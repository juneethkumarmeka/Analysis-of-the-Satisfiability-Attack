module basic_750_5000_1000_25_levels_5xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
xor U0 (N_0,In_570,In_545);
or U1 (N_1,In_392,In_483);
or U2 (N_2,In_472,In_144);
or U3 (N_3,In_663,In_51);
or U4 (N_4,In_717,In_83);
or U5 (N_5,In_65,In_679);
and U6 (N_6,In_420,In_373);
and U7 (N_7,In_77,In_452);
or U8 (N_8,In_26,In_199);
xnor U9 (N_9,In_149,In_290);
nor U10 (N_10,In_372,In_362);
nand U11 (N_11,In_422,In_682);
or U12 (N_12,In_175,In_361);
nor U13 (N_13,In_527,In_415);
nor U14 (N_14,In_88,In_720);
and U15 (N_15,In_329,In_419);
nand U16 (N_16,In_695,In_708);
or U17 (N_17,In_198,In_575);
or U18 (N_18,In_342,In_270);
xnor U19 (N_19,In_724,In_40);
nand U20 (N_20,In_384,In_439);
nand U21 (N_21,In_664,In_670);
and U22 (N_22,In_102,In_122);
nand U23 (N_23,In_359,In_580);
nand U24 (N_24,In_332,In_746);
and U25 (N_25,In_227,In_397);
nand U26 (N_26,In_311,In_601);
nand U27 (N_27,In_597,In_0);
and U28 (N_28,In_119,In_704);
and U29 (N_29,In_236,In_433);
and U30 (N_30,In_159,In_540);
xnor U31 (N_31,In_37,In_234);
or U32 (N_32,In_275,In_479);
nand U33 (N_33,In_310,In_85);
and U34 (N_34,In_230,In_209);
and U35 (N_35,In_696,In_716);
nand U36 (N_36,In_139,In_656);
nand U37 (N_37,In_453,In_201);
nand U38 (N_38,In_374,In_401);
nor U39 (N_39,In_733,In_331);
and U40 (N_40,In_147,In_685);
or U41 (N_41,In_661,In_448);
nor U42 (N_42,In_421,In_181);
or U43 (N_43,In_140,In_168);
nand U44 (N_44,In_418,In_87);
and U45 (N_45,In_30,In_585);
nor U46 (N_46,In_72,In_183);
nand U47 (N_47,In_727,In_5);
or U48 (N_48,In_531,In_743);
or U49 (N_49,In_606,In_210);
and U50 (N_50,In_651,In_650);
xor U51 (N_51,In_493,In_365);
nor U52 (N_52,In_609,In_615);
and U53 (N_53,In_607,In_382);
nor U54 (N_54,In_646,In_120);
or U55 (N_55,In_709,In_506);
xor U56 (N_56,In_42,In_348);
nor U57 (N_57,In_516,In_276);
and U58 (N_58,In_546,In_297);
or U59 (N_59,In_549,In_521);
nand U60 (N_60,In_610,In_619);
nor U61 (N_61,In_315,In_394);
or U62 (N_62,In_21,In_22);
nand U63 (N_63,In_689,In_426);
xnor U64 (N_64,In_490,In_671);
xnor U65 (N_65,In_279,In_553);
or U66 (N_66,In_283,In_599);
nand U67 (N_67,In_247,In_379);
nor U68 (N_68,In_626,In_518);
nand U69 (N_69,In_167,In_559);
or U70 (N_70,In_355,In_707);
nand U71 (N_71,In_10,In_195);
nor U72 (N_72,In_173,In_587);
nor U73 (N_73,In_114,In_80);
or U74 (N_74,In_36,In_1);
and U75 (N_75,In_665,In_13);
or U76 (N_76,In_742,In_454);
nor U77 (N_77,In_206,In_576);
nor U78 (N_78,In_445,In_202);
nor U79 (N_79,In_414,In_349);
or U80 (N_80,In_150,In_56);
nor U81 (N_81,In_410,In_244);
or U82 (N_82,In_133,In_556);
nor U83 (N_83,In_161,In_517);
nor U84 (N_84,In_522,In_125);
nor U85 (N_85,In_591,In_558);
nand U86 (N_86,In_388,In_738);
or U87 (N_87,In_267,In_14);
nand U88 (N_88,In_269,In_135);
nor U89 (N_89,In_151,In_478);
nand U90 (N_90,In_245,In_487);
nor U91 (N_91,In_327,In_293);
nand U92 (N_92,In_258,In_191);
nor U93 (N_93,In_308,In_101);
nor U94 (N_94,In_482,In_430);
nor U95 (N_95,In_259,In_203);
or U96 (N_96,In_237,In_456);
and U97 (N_97,In_171,In_480);
or U98 (N_98,In_450,In_215);
nand U99 (N_99,In_550,In_579);
and U100 (N_100,In_221,In_27);
nand U101 (N_101,In_712,In_255);
nand U102 (N_102,In_674,In_618);
nor U103 (N_103,In_376,In_443);
or U104 (N_104,In_152,In_312);
nor U105 (N_105,In_163,In_455);
nor U106 (N_106,In_188,In_288);
nand U107 (N_107,In_509,In_192);
xor U108 (N_108,In_100,In_132);
or U109 (N_109,In_701,In_251);
nor U110 (N_110,In_395,In_498);
and U111 (N_111,In_508,In_108);
nand U112 (N_112,In_338,In_596);
nor U113 (N_113,In_411,In_325);
and U114 (N_114,In_687,In_492);
or U115 (N_115,In_241,In_67);
nor U116 (N_116,In_555,In_145);
nor U117 (N_117,In_407,In_567);
or U118 (N_118,In_593,In_113);
or U119 (N_119,In_631,In_474);
or U120 (N_120,In_49,In_232);
nor U121 (N_121,In_475,In_340);
nor U122 (N_122,In_437,In_386);
xor U123 (N_123,In_95,In_638);
nand U124 (N_124,In_328,In_189);
xnor U125 (N_125,In_557,In_467);
or U126 (N_126,In_322,In_364);
nor U127 (N_127,In_569,In_383);
or U128 (N_128,In_284,In_260);
or U129 (N_129,In_605,In_718);
or U130 (N_130,In_337,In_371);
xor U131 (N_131,In_200,In_485);
nor U132 (N_132,In_621,In_252);
or U133 (N_133,In_360,In_86);
nand U134 (N_134,In_131,In_624);
nand U135 (N_135,In_18,In_653);
or U136 (N_136,In_45,In_633);
nand U137 (N_137,In_519,In_143);
nand U138 (N_138,In_600,In_463);
or U139 (N_139,In_64,In_317);
and U140 (N_140,In_250,In_398);
or U141 (N_141,In_729,In_197);
nor U142 (N_142,In_345,In_461);
and U143 (N_143,In_261,In_693);
xor U144 (N_144,In_124,In_481);
nor U145 (N_145,In_675,In_616);
and U146 (N_146,In_115,In_61);
nand U147 (N_147,In_226,In_686);
and U148 (N_148,In_705,In_416);
nor U149 (N_149,In_212,In_614);
and U150 (N_150,In_160,In_280);
xnor U151 (N_151,In_469,In_231);
and U152 (N_152,In_539,In_451);
and U153 (N_153,In_477,In_381);
xor U154 (N_154,In_354,In_229);
nand U155 (N_155,In_243,In_565);
nand U156 (N_156,In_417,In_399);
nand U157 (N_157,In_214,In_341);
nand U158 (N_158,In_58,In_528);
nand U159 (N_159,In_35,In_7);
nor U160 (N_160,In_166,In_494);
or U161 (N_161,In_59,In_378);
nand U162 (N_162,In_91,In_211);
or U163 (N_163,In_368,In_391);
nor U164 (N_164,In_654,In_655);
or U165 (N_165,In_678,In_387);
xor U166 (N_166,In_177,In_543);
nand U167 (N_167,In_172,In_714);
nor U168 (N_168,In_32,In_97);
nor U169 (N_169,In_105,In_488);
nor U170 (N_170,In_533,In_577);
nand U171 (N_171,In_79,In_8);
nand U172 (N_172,In_320,In_476);
and U173 (N_173,In_272,In_121);
nand U174 (N_174,In_684,In_425);
or U175 (N_175,In_564,In_586);
nor U176 (N_176,In_99,In_748);
or U177 (N_177,In_6,In_363);
or U178 (N_178,In_432,In_370);
nand U179 (N_179,In_639,In_41);
or U180 (N_180,In_323,In_734);
nor U181 (N_181,In_220,In_57);
or U182 (N_182,In_74,In_578);
or U183 (N_183,In_257,In_63);
and U184 (N_184,In_262,In_560);
or U185 (N_185,In_683,In_300);
nand U186 (N_186,In_566,In_627);
nand U187 (N_187,In_254,In_622);
and U188 (N_188,In_12,In_356);
and U189 (N_189,In_530,In_692);
xor U190 (N_190,In_179,In_289);
and U191 (N_191,In_389,In_643);
nor U192 (N_192,In_48,In_703);
and U193 (N_193,In_617,In_28);
xnor U194 (N_194,In_69,In_719);
and U195 (N_195,In_157,In_213);
nor U196 (N_196,In_38,In_691);
nand U197 (N_197,In_43,In_731);
or U198 (N_198,In_589,In_598);
nor U199 (N_199,In_17,In_604);
and U200 (N_200,In_103,In_351);
nor U201 (N_201,N_129,In_647);
and U202 (N_202,In_291,N_31);
and U203 (N_203,In_574,In_256);
and U204 (N_204,N_68,N_184);
or U205 (N_205,N_43,In_292);
nor U206 (N_206,N_82,In_645);
nor U207 (N_207,In_148,N_57);
xnor U208 (N_208,N_34,N_125);
and U209 (N_209,In_745,N_196);
or U210 (N_210,N_153,In_699);
and U211 (N_211,In_218,In_126);
or U212 (N_212,N_26,In_268);
or U213 (N_213,N_99,In_666);
and U214 (N_214,In_640,In_282);
or U215 (N_215,N_127,In_158);
and U216 (N_216,N_124,N_6);
and U217 (N_217,In_429,N_133);
nand U218 (N_218,In_138,In_644);
and U219 (N_219,In_129,In_515);
nand U220 (N_220,In_524,N_194);
nor U221 (N_221,In_669,In_46);
or U222 (N_222,In_73,N_131);
and U223 (N_223,In_694,In_563);
and U224 (N_224,In_673,N_114);
and U225 (N_225,N_186,N_126);
xor U226 (N_226,N_171,N_72);
or U227 (N_227,In_723,N_150);
nand U228 (N_228,In_286,In_235);
or U229 (N_229,In_590,In_471);
and U230 (N_230,In_611,In_130);
and U231 (N_231,In_608,In_740);
or U232 (N_232,N_66,In_304);
or U233 (N_233,In_681,In_702);
nand U234 (N_234,N_179,In_511);
nor U235 (N_235,In_154,N_49);
or U236 (N_236,In_613,N_143);
nor U237 (N_237,In_535,In_54);
nor U238 (N_238,In_174,In_296);
nor U239 (N_239,In_390,In_503);
nand U240 (N_240,In_39,In_440);
and U241 (N_241,N_54,In_544);
xnor U242 (N_242,In_238,In_82);
or U243 (N_243,In_406,In_541);
nor U244 (N_244,In_620,N_197);
nand U245 (N_245,N_178,In_110);
nand U246 (N_246,In_265,N_110);
nor U247 (N_247,In_648,N_132);
or U248 (N_248,In_588,N_12);
or U249 (N_249,In_697,In_281);
and U250 (N_250,N_155,N_44);
nand U251 (N_251,In_592,N_3);
and U252 (N_252,In_513,In_169);
nand U253 (N_253,In_441,In_2);
nor U254 (N_254,In_409,N_187);
nand U255 (N_255,In_294,N_45);
or U256 (N_256,In_193,In_228);
or U257 (N_257,In_510,In_552);
xnor U258 (N_258,N_8,N_139);
nand U259 (N_259,In_636,In_662);
nor U260 (N_260,In_75,In_500);
nor U261 (N_261,N_119,In_413);
nand U262 (N_262,N_91,In_134);
xor U263 (N_263,In_47,N_80);
and U264 (N_264,In_529,N_115);
or U265 (N_265,In_625,N_149);
or U266 (N_266,N_181,N_142);
and U267 (N_267,In_298,In_184);
nand U268 (N_268,In_305,In_403);
and U269 (N_269,In_525,In_412);
or U270 (N_270,N_67,In_343);
and U271 (N_271,N_16,N_159);
and U272 (N_272,N_93,In_90);
or U273 (N_273,N_63,In_538);
nand U274 (N_274,In_690,In_93);
and U275 (N_275,In_111,In_194);
nand U276 (N_276,In_29,N_33);
and U277 (N_277,In_358,In_715);
and U278 (N_278,N_168,N_135);
or U279 (N_279,In_584,In_208);
nor U280 (N_280,N_27,N_78);
nor U281 (N_281,N_199,In_107);
nand U282 (N_282,In_747,In_400);
or U283 (N_283,In_307,In_447);
nor U284 (N_284,N_50,In_190);
or U285 (N_285,In_271,In_464);
nand U286 (N_286,In_459,N_188);
or U287 (N_287,N_122,In_295);
and U288 (N_288,N_164,In_496);
or U289 (N_289,In_15,N_38);
or U290 (N_290,In_187,In_698);
nor U291 (N_291,In_680,N_18);
nand U292 (N_292,N_83,N_158);
nor U293 (N_293,N_151,N_148);
or U294 (N_294,N_48,N_73);
or U295 (N_295,In_635,In_562);
and U296 (N_296,In_19,N_166);
nand U297 (N_297,In_109,N_86);
nor U298 (N_298,In_335,In_710);
nand U299 (N_299,N_156,In_658);
and U300 (N_300,In_396,In_595);
nand U301 (N_301,In_219,In_20);
nand U302 (N_302,In_641,In_165);
and U303 (N_303,In_660,N_191);
or U304 (N_304,In_623,N_97);
nor U305 (N_305,N_74,In_319);
or U306 (N_306,In_507,In_242);
nand U307 (N_307,N_9,N_4);
nor U308 (N_308,N_162,In_23);
xnor U309 (N_309,In_16,In_652);
nand U310 (N_310,N_21,N_52);
nand U311 (N_311,N_163,In_239);
nor U312 (N_312,In_224,In_274);
nor U313 (N_313,N_193,In_749);
nor U314 (N_314,In_526,In_96);
and U315 (N_315,In_542,In_62);
nor U316 (N_316,In_405,In_112);
nor U317 (N_317,N_15,In_117);
and U318 (N_318,In_116,In_739);
nor U319 (N_319,N_130,N_109);
nor U320 (N_320,N_62,N_180);
nor U321 (N_321,N_42,N_89);
nor U322 (N_322,In_357,N_134);
and U323 (N_323,In_502,In_489);
or U324 (N_324,In_153,N_145);
nand U325 (N_325,In_466,N_157);
nand U326 (N_326,N_120,In_735);
or U327 (N_327,In_721,In_505);
xnor U328 (N_328,In_722,N_22);
or U329 (N_329,In_444,In_196);
nand U330 (N_330,N_76,In_726);
nand U331 (N_331,In_185,In_512);
xnor U332 (N_332,N_87,In_602);
nand U333 (N_333,In_4,N_173);
nor U334 (N_334,In_277,N_161);
nor U335 (N_335,In_287,N_28);
xor U336 (N_336,In_285,In_486);
xor U337 (N_337,N_195,In_78);
or U338 (N_338,In_668,In_71);
nand U339 (N_339,In_31,N_189);
nand U340 (N_340,In_98,N_198);
and U341 (N_341,N_136,In_302);
or U342 (N_342,In_728,In_347);
nor U343 (N_343,In_499,In_520);
and U344 (N_344,N_116,In_299);
and U345 (N_345,N_88,N_174);
or U346 (N_346,In_92,In_264);
or U347 (N_347,N_172,N_70);
and U348 (N_348,In_94,In_408);
xor U349 (N_349,In_657,In_55);
or U350 (N_350,N_90,In_630);
or U351 (N_351,In_568,N_7);
or U352 (N_352,In_222,N_2);
or U353 (N_353,In_318,In_225);
nor U354 (N_354,N_29,N_165);
and U355 (N_355,In_581,In_551);
nor U356 (N_356,In_632,N_182);
or U357 (N_357,N_128,N_94);
or U358 (N_358,In_446,In_324);
nor U359 (N_359,N_183,In_118);
nor U360 (N_360,N_19,In_460);
nor U361 (N_361,In_68,N_84);
or U362 (N_362,N_175,N_137);
and U363 (N_363,N_30,N_71);
nand U364 (N_364,In_423,In_182);
and U365 (N_365,N_5,In_66);
or U366 (N_366,In_316,In_501);
or U367 (N_367,In_442,In_273);
or U368 (N_368,In_402,In_491);
nor U369 (N_369,In_248,In_128);
nor U370 (N_370,N_58,In_217);
or U371 (N_371,In_34,In_170);
xnor U372 (N_372,In_534,N_23);
nor U373 (N_373,In_438,N_121);
xor U374 (N_374,In_301,In_572);
nand U375 (N_375,N_41,N_47);
nor U376 (N_376,In_249,N_113);
or U377 (N_377,N_141,N_177);
nand U378 (N_378,In_313,In_554);
nand U379 (N_379,N_51,N_1);
nand U380 (N_380,In_677,In_303);
nand U381 (N_381,In_207,N_95);
and U382 (N_382,N_100,In_730);
and U383 (N_383,N_20,In_367);
and U384 (N_384,In_583,In_84);
and U385 (N_385,N_170,In_688);
or U386 (N_386,In_350,In_186);
nand U387 (N_387,In_263,In_428);
nand U388 (N_388,N_152,In_431);
nand U389 (N_389,In_706,N_60);
nor U390 (N_390,In_336,In_333);
nand U391 (N_391,In_321,In_3);
or U392 (N_392,N_25,In_457);
or U393 (N_393,In_9,In_369);
or U394 (N_394,In_223,N_55);
and U395 (N_395,In_309,In_667);
and U396 (N_396,N_39,N_176);
nor U397 (N_397,N_185,In_278);
or U398 (N_398,In_741,N_154);
and U399 (N_399,In_123,In_136);
and U400 (N_400,N_311,In_104);
nand U401 (N_401,N_262,N_330);
nor U402 (N_402,In_637,N_256);
or U403 (N_403,N_75,N_358);
xor U404 (N_404,N_200,N_138);
xnor U405 (N_405,In_424,N_306);
and U406 (N_406,N_102,N_224);
and U407 (N_407,N_398,N_304);
and U408 (N_408,N_389,N_321);
or U409 (N_409,In_326,In_582);
nand U410 (N_410,N_322,In_629);
or U411 (N_411,N_140,In_127);
and U412 (N_412,N_327,In_523);
or U413 (N_413,N_59,N_104);
or U414 (N_414,N_264,N_323);
xnor U415 (N_415,N_147,N_277);
nor U416 (N_416,In_106,N_212);
xnor U417 (N_417,N_268,N_14);
or U418 (N_418,In_385,N_215);
and U419 (N_419,N_263,In_393);
or U420 (N_420,N_303,In_366);
nand U421 (N_421,N_231,N_288);
nand U422 (N_422,N_343,In_11);
or U423 (N_423,In_162,N_293);
and U424 (N_424,N_282,N_286);
xnor U425 (N_425,N_10,N_299);
and U426 (N_426,N_274,N_229);
nand U427 (N_427,N_365,In_404);
or U428 (N_428,N_247,In_33);
xnor U429 (N_429,N_337,N_363);
xor U430 (N_430,N_285,N_386);
xor U431 (N_431,In_634,N_237);
or U432 (N_432,N_56,In_137);
xnor U433 (N_433,In_50,N_316);
nand U434 (N_434,N_345,N_118);
xor U435 (N_435,In_548,N_0);
nand U436 (N_436,In_435,N_222);
nor U437 (N_437,In_330,N_313);
and U438 (N_438,N_112,N_387);
nor U439 (N_439,In_216,N_305);
and U440 (N_440,N_310,N_326);
nor U441 (N_441,In_700,N_220);
and U442 (N_442,N_317,N_244);
nor U443 (N_443,N_354,N_211);
nor U444 (N_444,N_240,N_85);
nand U445 (N_445,N_329,N_65);
or U446 (N_446,N_383,N_396);
nand U447 (N_447,N_361,In_353);
nand U448 (N_448,In_736,In_344);
xnor U449 (N_449,In_253,N_223);
or U450 (N_450,N_98,N_397);
xor U451 (N_451,In_178,N_290);
nor U452 (N_452,N_267,N_342);
or U453 (N_453,N_367,N_312);
nor U454 (N_454,N_101,N_210);
or U455 (N_455,N_366,N_69);
nor U456 (N_456,N_209,N_217);
nand U457 (N_457,N_292,In_352);
xnor U458 (N_458,N_160,N_40);
and U459 (N_459,N_214,In_76);
nor U460 (N_460,N_271,In_732);
and U461 (N_461,N_294,N_394);
nor U462 (N_462,N_123,N_279);
or U463 (N_463,N_275,N_207);
and U464 (N_464,In_205,N_333);
nor U465 (N_465,In_571,N_249);
nand U466 (N_466,In_676,N_364);
or U467 (N_467,N_258,N_379);
and U468 (N_468,N_225,N_340);
xor U469 (N_469,N_261,In_497);
nor U470 (N_470,N_332,In_547);
nand U471 (N_471,In_495,In_266);
and U472 (N_472,N_111,N_219);
nand U473 (N_473,N_314,N_350);
and U474 (N_474,N_190,N_339);
and U475 (N_475,N_106,N_360);
and U476 (N_476,In_659,N_24);
xor U477 (N_477,N_105,N_192);
and U478 (N_478,N_117,In_155);
and U479 (N_479,N_13,N_362);
nor U480 (N_480,In_146,N_205);
and U481 (N_481,N_260,N_353);
nor U482 (N_482,In_672,N_295);
and U483 (N_483,N_301,N_218);
nor U484 (N_484,In_484,N_169);
xor U485 (N_485,N_357,N_11);
and U486 (N_486,In_204,N_341);
xnor U487 (N_487,N_308,N_241);
xnor U488 (N_488,N_35,In_346);
nor U489 (N_489,N_349,N_399);
nor U490 (N_490,N_272,N_92);
or U491 (N_491,N_289,N_287);
nor U492 (N_492,N_108,N_372);
or U493 (N_493,N_36,N_320);
nor U494 (N_494,In_176,In_52);
xor U495 (N_495,N_255,N_17);
nor U496 (N_496,N_234,In_514);
and U497 (N_497,N_77,N_388);
xor U498 (N_498,In_380,In_713);
nor U499 (N_499,N_296,In_504);
and U500 (N_500,In_725,N_375);
nand U501 (N_501,In_314,N_368);
nand U502 (N_502,N_319,In_44);
or U503 (N_503,N_235,N_167);
or U504 (N_504,N_324,In_434);
nand U505 (N_505,N_226,N_238);
and U506 (N_506,N_391,N_242);
xor U507 (N_507,In_470,N_259);
nand U508 (N_508,N_307,N_257);
nor U509 (N_509,N_331,In_25);
and U510 (N_510,N_385,N_216);
and U511 (N_511,In_81,N_270);
nor U512 (N_512,N_278,N_273);
or U513 (N_513,N_79,In_339);
or U514 (N_514,N_309,In_306);
nand U515 (N_515,N_254,N_315);
or U516 (N_516,N_236,N_239);
or U517 (N_517,In_156,N_46);
nor U518 (N_518,N_233,N_248);
or U519 (N_519,N_377,N_359);
nor U520 (N_520,In_536,N_146);
and U521 (N_521,In_24,N_206);
xor U522 (N_522,In_164,In_458);
nor U523 (N_523,N_374,N_338);
and U524 (N_524,In_53,N_266);
nand U525 (N_525,N_221,N_53);
and U526 (N_526,N_103,In_711);
or U527 (N_527,N_61,N_201);
nor U528 (N_528,N_245,In_462);
and U529 (N_529,N_284,N_107);
xnor U530 (N_530,N_334,N_291);
nand U531 (N_531,In_737,N_395);
nand U532 (N_532,In_377,N_81);
and U533 (N_533,In_375,N_392);
nand U534 (N_534,N_346,In_240);
or U535 (N_535,N_378,N_32);
nor U536 (N_536,N_265,In_561);
xor U537 (N_537,In_744,N_228);
nand U538 (N_538,N_203,In_449);
nand U539 (N_539,N_227,N_280);
or U540 (N_540,N_96,N_204);
and U541 (N_541,N_328,In_642);
nand U542 (N_542,N_297,In_60);
or U543 (N_543,N_376,N_318);
and U544 (N_544,N_276,N_355);
nand U545 (N_545,In_628,N_302);
nand U546 (N_546,In_436,In_180);
nand U547 (N_547,N_352,N_381);
nor U548 (N_548,In_246,In_603);
nand U549 (N_549,N_230,In_473);
nor U550 (N_550,In_465,N_336);
nor U551 (N_551,In_468,N_253);
xor U552 (N_552,In_141,N_37);
or U553 (N_553,N_144,N_246);
or U554 (N_554,In_142,N_281);
or U555 (N_555,N_390,In_70);
nor U556 (N_556,N_393,N_269);
and U557 (N_557,N_232,In_334);
nand U558 (N_558,N_298,N_370);
and U559 (N_559,N_348,N_325);
and U560 (N_560,In_612,N_213);
nor U561 (N_561,In_594,N_335);
or U562 (N_562,N_202,N_351);
nor U563 (N_563,N_64,N_344);
and U564 (N_564,N_283,N_371);
nand U565 (N_565,In_573,N_252);
or U566 (N_566,N_356,In_89);
or U567 (N_567,N_382,N_384);
nor U568 (N_568,N_369,N_251);
nand U569 (N_569,N_347,N_373);
and U570 (N_570,In_532,N_300);
xnor U571 (N_571,In_427,N_380);
xnor U572 (N_572,N_243,N_250);
or U573 (N_573,In_233,In_537);
and U574 (N_574,N_208,In_649);
xor U575 (N_575,N_355,In_649);
and U576 (N_576,N_286,N_335);
nand U577 (N_577,N_242,N_209);
nand U578 (N_578,N_311,N_224);
or U579 (N_579,N_284,In_60);
nand U580 (N_580,In_634,N_32);
xnor U581 (N_581,In_246,In_504);
and U582 (N_582,N_350,N_385);
nor U583 (N_583,N_374,N_204);
nor U584 (N_584,N_144,In_142);
and U585 (N_585,In_377,N_104);
and U586 (N_586,N_294,N_329);
nand U587 (N_587,N_65,N_344);
nand U588 (N_588,N_282,N_366);
and U589 (N_589,N_392,N_105);
or U590 (N_590,N_235,N_317);
or U591 (N_591,N_219,N_206);
or U592 (N_592,N_235,N_190);
nand U593 (N_593,In_536,N_254);
xnor U594 (N_594,N_225,In_142);
nor U595 (N_595,N_318,N_265);
nand U596 (N_596,N_232,N_242);
nor U597 (N_597,N_246,In_523);
and U598 (N_598,N_221,N_291);
xnor U599 (N_599,In_44,N_207);
or U600 (N_600,N_562,N_541);
or U601 (N_601,N_534,N_445);
and U602 (N_602,N_429,N_455);
xor U603 (N_603,N_554,N_415);
or U604 (N_604,N_488,N_544);
and U605 (N_605,N_405,N_589);
or U606 (N_606,N_512,N_414);
or U607 (N_607,N_545,N_555);
xnor U608 (N_608,N_566,N_523);
xor U609 (N_609,N_474,N_542);
nand U610 (N_610,N_591,N_410);
nand U611 (N_611,N_597,N_568);
nor U612 (N_612,N_519,N_498);
or U613 (N_613,N_400,N_482);
nor U614 (N_614,N_434,N_437);
or U615 (N_615,N_490,N_501);
and U616 (N_616,N_463,N_470);
nand U617 (N_617,N_583,N_559);
or U618 (N_618,N_586,N_503);
xor U619 (N_619,N_409,N_528);
nand U620 (N_620,N_466,N_489);
nor U621 (N_621,N_502,N_428);
nor U622 (N_622,N_570,N_472);
nor U623 (N_623,N_522,N_465);
and U624 (N_624,N_438,N_550);
nand U625 (N_625,N_582,N_560);
or U626 (N_626,N_546,N_547);
nand U627 (N_627,N_483,N_468);
and U628 (N_628,N_495,N_442);
or U629 (N_629,N_510,N_593);
nand U630 (N_630,N_424,N_529);
nand U631 (N_631,N_416,N_491);
nor U632 (N_632,N_594,N_599);
and U633 (N_633,N_543,N_451);
xor U634 (N_634,N_408,N_581);
nand U635 (N_635,N_426,N_432);
nor U636 (N_636,N_453,N_507);
and U637 (N_637,N_595,N_475);
nand U638 (N_638,N_513,N_592);
nor U639 (N_639,N_494,N_580);
and U640 (N_640,N_412,N_462);
nor U641 (N_641,N_558,N_407);
nor U642 (N_642,N_485,N_471);
nor U643 (N_643,N_402,N_454);
xor U644 (N_644,N_446,N_441);
or U645 (N_645,N_535,N_436);
nand U646 (N_646,N_479,N_508);
nand U647 (N_647,N_443,N_458);
or U648 (N_648,N_499,N_506);
nand U649 (N_649,N_456,N_411);
or U650 (N_650,N_504,N_553);
or U651 (N_651,N_486,N_448);
and U652 (N_652,N_469,N_406);
or U653 (N_653,N_567,N_496);
and U654 (N_654,N_527,N_571);
xnor U655 (N_655,N_533,N_575);
nor U656 (N_656,N_588,N_435);
and U657 (N_657,N_572,N_477);
nand U658 (N_658,N_564,N_493);
or U659 (N_659,N_425,N_497);
nor U660 (N_660,N_505,N_526);
nand U661 (N_661,N_577,N_413);
nor U662 (N_662,N_450,N_473);
and U663 (N_663,N_430,N_515);
xor U664 (N_664,N_417,N_452);
or U665 (N_665,N_557,N_511);
nor U666 (N_666,N_532,N_585);
and U667 (N_667,N_478,N_537);
or U668 (N_668,N_584,N_587);
nor U669 (N_669,N_467,N_509);
xnor U670 (N_670,N_457,N_569);
nand U671 (N_671,N_464,N_403);
or U672 (N_672,N_573,N_563);
nand U673 (N_673,N_538,N_422);
or U674 (N_674,N_440,N_520);
or U675 (N_675,N_433,N_579);
xnor U676 (N_676,N_459,N_548);
xnor U677 (N_677,N_427,N_518);
or U678 (N_678,N_514,N_521);
and U679 (N_679,N_480,N_525);
nand U680 (N_680,N_476,N_574);
and U681 (N_681,N_549,N_552);
and U682 (N_682,N_431,N_460);
nor U683 (N_683,N_561,N_449);
nor U684 (N_684,N_419,N_461);
nand U685 (N_685,N_401,N_516);
or U686 (N_686,N_576,N_565);
or U687 (N_687,N_492,N_444);
nor U688 (N_688,N_536,N_596);
nand U689 (N_689,N_590,N_530);
and U690 (N_690,N_578,N_524);
and U691 (N_691,N_418,N_447);
and U692 (N_692,N_539,N_484);
nand U693 (N_693,N_556,N_500);
and U694 (N_694,N_517,N_439);
nand U695 (N_695,N_598,N_481);
or U696 (N_696,N_551,N_423);
or U697 (N_697,N_487,N_421);
or U698 (N_698,N_404,N_540);
nor U699 (N_699,N_531,N_420);
and U700 (N_700,N_539,N_593);
or U701 (N_701,N_491,N_516);
xnor U702 (N_702,N_561,N_439);
nor U703 (N_703,N_583,N_480);
nand U704 (N_704,N_505,N_587);
nand U705 (N_705,N_492,N_497);
or U706 (N_706,N_494,N_544);
nor U707 (N_707,N_408,N_446);
nor U708 (N_708,N_500,N_469);
or U709 (N_709,N_536,N_547);
and U710 (N_710,N_439,N_423);
nor U711 (N_711,N_498,N_531);
nor U712 (N_712,N_459,N_519);
nor U713 (N_713,N_586,N_524);
xor U714 (N_714,N_463,N_478);
xor U715 (N_715,N_426,N_541);
or U716 (N_716,N_573,N_518);
and U717 (N_717,N_515,N_590);
nor U718 (N_718,N_595,N_510);
and U719 (N_719,N_468,N_486);
or U720 (N_720,N_581,N_510);
nor U721 (N_721,N_462,N_431);
or U722 (N_722,N_507,N_485);
nor U723 (N_723,N_540,N_566);
nand U724 (N_724,N_545,N_443);
xnor U725 (N_725,N_462,N_512);
and U726 (N_726,N_521,N_414);
nand U727 (N_727,N_446,N_411);
or U728 (N_728,N_529,N_461);
and U729 (N_729,N_448,N_524);
nand U730 (N_730,N_506,N_418);
or U731 (N_731,N_433,N_475);
and U732 (N_732,N_505,N_460);
and U733 (N_733,N_587,N_438);
nor U734 (N_734,N_485,N_522);
nand U735 (N_735,N_450,N_557);
and U736 (N_736,N_460,N_500);
or U737 (N_737,N_455,N_584);
and U738 (N_738,N_579,N_403);
xor U739 (N_739,N_432,N_452);
nand U740 (N_740,N_473,N_523);
nand U741 (N_741,N_557,N_531);
nor U742 (N_742,N_405,N_409);
nor U743 (N_743,N_426,N_442);
xnor U744 (N_744,N_509,N_464);
and U745 (N_745,N_494,N_485);
and U746 (N_746,N_482,N_497);
xnor U747 (N_747,N_405,N_524);
and U748 (N_748,N_402,N_445);
or U749 (N_749,N_468,N_410);
nor U750 (N_750,N_446,N_431);
and U751 (N_751,N_540,N_488);
xnor U752 (N_752,N_566,N_539);
or U753 (N_753,N_596,N_562);
nor U754 (N_754,N_573,N_434);
nand U755 (N_755,N_599,N_415);
xnor U756 (N_756,N_551,N_429);
nor U757 (N_757,N_414,N_569);
and U758 (N_758,N_552,N_528);
and U759 (N_759,N_518,N_599);
nand U760 (N_760,N_445,N_555);
and U761 (N_761,N_583,N_426);
nand U762 (N_762,N_565,N_519);
xnor U763 (N_763,N_526,N_528);
nor U764 (N_764,N_545,N_482);
nand U765 (N_765,N_430,N_488);
nand U766 (N_766,N_510,N_596);
and U767 (N_767,N_560,N_496);
nand U768 (N_768,N_511,N_421);
xor U769 (N_769,N_589,N_452);
nor U770 (N_770,N_525,N_562);
nand U771 (N_771,N_516,N_469);
or U772 (N_772,N_410,N_544);
or U773 (N_773,N_402,N_450);
and U774 (N_774,N_469,N_529);
nor U775 (N_775,N_541,N_573);
nor U776 (N_776,N_484,N_493);
and U777 (N_777,N_416,N_402);
or U778 (N_778,N_445,N_552);
nor U779 (N_779,N_442,N_430);
nand U780 (N_780,N_599,N_595);
nand U781 (N_781,N_445,N_443);
xor U782 (N_782,N_544,N_403);
nand U783 (N_783,N_571,N_450);
or U784 (N_784,N_415,N_455);
and U785 (N_785,N_466,N_467);
nor U786 (N_786,N_409,N_475);
nand U787 (N_787,N_401,N_447);
nor U788 (N_788,N_546,N_597);
nand U789 (N_789,N_499,N_557);
nand U790 (N_790,N_468,N_470);
nor U791 (N_791,N_478,N_575);
nor U792 (N_792,N_453,N_597);
and U793 (N_793,N_456,N_409);
nor U794 (N_794,N_560,N_579);
nand U795 (N_795,N_577,N_423);
and U796 (N_796,N_544,N_516);
and U797 (N_797,N_597,N_413);
nand U798 (N_798,N_507,N_449);
nand U799 (N_799,N_477,N_488);
xnor U800 (N_800,N_734,N_649);
or U801 (N_801,N_779,N_638);
and U802 (N_802,N_786,N_747);
nor U803 (N_803,N_765,N_678);
nand U804 (N_804,N_735,N_651);
nand U805 (N_805,N_750,N_784);
nor U806 (N_806,N_761,N_719);
nand U807 (N_807,N_654,N_736);
nand U808 (N_808,N_668,N_661);
nand U809 (N_809,N_697,N_686);
and U810 (N_810,N_755,N_799);
and U811 (N_811,N_614,N_780);
and U812 (N_812,N_739,N_754);
and U813 (N_813,N_798,N_776);
and U814 (N_814,N_743,N_667);
nor U815 (N_815,N_647,N_698);
xor U816 (N_816,N_695,N_742);
xor U817 (N_817,N_669,N_774);
or U818 (N_818,N_716,N_636);
nand U819 (N_819,N_628,N_744);
nor U820 (N_820,N_660,N_673);
and U821 (N_821,N_741,N_642);
and U822 (N_822,N_637,N_748);
nand U823 (N_823,N_603,N_785);
and U824 (N_824,N_728,N_769);
xor U825 (N_825,N_778,N_757);
or U826 (N_826,N_763,N_718);
nand U827 (N_827,N_632,N_730);
xor U828 (N_828,N_713,N_665);
and U829 (N_829,N_620,N_662);
xor U830 (N_830,N_766,N_704);
nand U831 (N_831,N_625,N_705);
or U832 (N_832,N_733,N_717);
and U833 (N_833,N_737,N_659);
nand U834 (N_834,N_771,N_684);
nand U835 (N_835,N_723,N_756);
or U836 (N_836,N_663,N_680);
nand U837 (N_837,N_687,N_714);
nand U838 (N_838,N_773,N_609);
or U839 (N_839,N_781,N_611);
and U840 (N_840,N_615,N_711);
nor U841 (N_841,N_729,N_648);
or U842 (N_842,N_722,N_631);
or U843 (N_843,N_624,N_618);
xor U844 (N_844,N_789,N_783);
nor U845 (N_845,N_629,N_787);
and U846 (N_846,N_749,N_792);
nand U847 (N_847,N_788,N_664);
or U848 (N_848,N_708,N_682);
or U849 (N_849,N_709,N_655);
xor U850 (N_850,N_732,N_796);
nor U851 (N_851,N_703,N_623);
or U852 (N_852,N_639,N_634);
nor U853 (N_853,N_752,N_683);
nand U854 (N_854,N_710,N_726);
xor U855 (N_855,N_715,N_671);
nor U856 (N_856,N_681,N_644);
or U857 (N_857,N_791,N_653);
nand U858 (N_858,N_658,N_762);
or U859 (N_859,N_692,N_613);
nand U860 (N_860,N_617,N_690);
or U861 (N_861,N_707,N_760);
nor U862 (N_862,N_610,N_677);
or U863 (N_863,N_641,N_712);
and U864 (N_864,N_689,N_605);
or U865 (N_865,N_670,N_616);
nor U866 (N_866,N_652,N_626);
nand U867 (N_867,N_694,N_740);
nand U868 (N_868,N_674,N_643);
and U869 (N_869,N_797,N_640);
nor U870 (N_870,N_795,N_604);
nand U871 (N_871,N_608,N_635);
nor U872 (N_872,N_606,N_724);
nor U873 (N_873,N_633,N_793);
nor U874 (N_874,N_701,N_721);
nor U875 (N_875,N_645,N_772);
nor U876 (N_876,N_700,N_731);
nand U877 (N_877,N_702,N_746);
nand U878 (N_878,N_777,N_646);
and U879 (N_879,N_759,N_693);
or U880 (N_880,N_758,N_612);
or U881 (N_881,N_767,N_782);
nand U882 (N_882,N_672,N_790);
nand U883 (N_883,N_770,N_738);
and U884 (N_884,N_751,N_627);
and U885 (N_885,N_656,N_619);
nor U886 (N_886,N_602,N_691);
nand U887 (N_887,N_775,N_764);
nor U888 (N_888,N_650,N_622);
nand U889 (N_889,N_657,N_600);
nand U890 (N_890,N_607,N_696);
or U891 (N_891,N_621,N_745);
xnor U892 (N_892,N_666,N_676);
nor U893 (N_893,N_753,N_685);
and U894 (N_894,N_699,N_706);
nor U895 (N_895,N_720,N_794);
nor U896 (N_896,N_727,N_679);
xor U897 (N_897,N_675,N_725);
nand U898 (N_898,N_688,N_630);
and U899 (N_899,N_768,N_601);
nor U900 (N_900,N_733,N_619);
nor U901 (N_901,N_760,N_772);
nand U902 (N_902,N_788,N_707);
nand U903 (N_903,N_729,N_713);
or U904 (N_904,N_626,N_733);
nand U905 (N_905,N_678,N_738);
or U906 (N_906,N_735,N_728);
and U907 (N_907,N_736,N_745);
nor U908 (N_908,N_679,N_763);
nand U909 (N_909,N_799,N_739);
nor U910 (N_910,N_745,N_789);
and U911 (N_911,N_653,N_738);
and U912 (N_912,N_775,N_654);
xor U913 (N_913,N_757,N_624);
or U914 (N_914,N_671,N_660);
or U915 (N_915,N_772,N_723);
and U916 (N_916,N_722,N_748);
nand U917 (N_917,N_709,N_649);
nand U918 (N_918,N_637,N_777);
xor U919 (N_919,N_602,N_790);
nor U920 (N_920,N_734,N_629);
nand U921 (N_921,N_763,N_790);
nor U922 (N_922,N_685,N_778);
nand U923 (N_923,N_684,N_626);
nand U924 (N_924,N_691,N_797);
or U925 (N_925,N_626,N_728);
and U926 (N_926,N_711,N_670);
nand U927 (N_927,N_655,N_794);
nand U928 (N_928,N_721,N_696);
and U929 (N_929,N_728,N_779);
and U930 (N_930,N_778,N_756);
and U931 (N_931,N_727,N_696);
nand U932 (N_932,N_663,N_682);
nand U933 (N_933,N_671,N_664);
nand U934 (N_934,N_701,N_737);
xor U935 (N_935,N_671,N_708);
and U936 (N_936,N_789,N_660);
and U937 (N_937,N_781,N_627);
or U938 (N_938,N_788,N_789);
or U939 (N_939,N_614,N_651);
nor U940 (N_940,N_686,N_799);
nor U941 (N_941,N_669,N_650);
nor U942 (N_942,N_791,N_667);
nand U943 (N_943,N_637,N_715);
and U944 (N_944,N_601,N_772);
nor U945 (N_945,N_733,N_798);
nand U946 (N_946,N_689,N_779);
nand U947 (N_947,N_724,N_760);
nand U948 (N_948,N_731,N_778);
xnor U949 (N_949,N_633,N_687);
and U950 (N_950,N_739,N_678);
nor U951 (N_951,N_670,N_767);
nand U952 (N_952,N_770,N_774);
and U953 (N_953,N_719,N_603);
xor U954 (N_954,N_727,N_652);
or U955 (N_955,N_791,N_660);
or U956 (N_956,N_678,N_783);
xor U957 (N_957,N_630,N_734);
and U958 (N_958,N_734,N_635);
nor U959 (N_959,N_643,N_712);
nand U960 (N_960,N_709,N_684);
or U961 (N_961,N_792,N_652);
nand U962 (N_962,N_703,N_780);
nor U963 (N_963,N_687,N_659);
or U964 (N_964,N_752,N_695);
xnor U965 (N_965,N_777,N_766);
and U966 (N_966,N_632,N_683);
nand U967 (N_967,N_733,N_654);
nand U968 (N_968,N_763,N_663);
and U969 (N_969,N_640,N_769);
xnor U970 (N_970,N_739,N_716);
and U971 (N_971,N_749,N_682);
and U972 (N_972,N_760,N_731);
or U973 (N_973,N_735,N_726);
or U974 (N_974,N_777,N_731);
and U975 (N_975,N_720,N_766);
or U976 (N_976,N_600,N_783);
or U977 (N_977,N_746,N_736);
or U978 (N_978,N_712,N_789);
and U979 (N_979,N_611,N_782);
nor U980 (N_980,N_605,N_653);
nor U981 (N_981,N_622,N_725);
and U982 (N_982,N_665,N_739);
and U983 (N_983,N_657,N_768);
nor U984 (N_984,N_689,N_648);
or U985 (N_985,N_656,N_695);
and U986 (N_986,N_727,N_761);
nand U987 (N_987,N_788,N_616);
and U988 (N_988,N_744,N_785);
nand U989 (N_989,N_625,N_667);
and U990 (N_990,N_605,N_723);
xor U991 (N_991,N_634,N_638);
or U992 (N_992,N_777,N_636);
or U993 (N_993,N_767,N_691);
or U994 (N_994,N_648,N_753);
nand U995 (N_995,N_600,N_775);
and U996 (N_996,N_795,N_705);
and U997 (N_997,N_600,N_694);
xnor U998 (N_998,N_640,N_733);
and U999 (N_999,N_701,N_678);
nand U1000 (N_1000,N_960,N_940);
nand U1001 (N_1001,N_834,N_878);
or U1002 (N_1002,N_870,N_867);
nand U1003 (N_1003,N_836,N_843);
xor U1004 (N_1004,N_865,N_885);
nor U1005 (N_1005,N_970,N_888);
nand U1006 (N_1006,N_936,N_955);
nor U1007 (N_1007,N_835,N_900);
or U1008 (N_1008,N_829,N_875);
and U1009 (N_1009,N_999,N_945);
and U1010 (N_1010,N_896,N_930);
nand U1011 (N_1011,N_952,N_899);
and U1012 (N_1012,N_949,N_832);
and U1013 (N_1013,N_946,N_889);
or U1014 (N_1014,N_884,N_980);
nand U1015 (N_1015,N_909,N_969);
and U1016 (N_1016,N_987,N_830);
nor U1017 (N_1017,N_943,N_803);
nor U1018 (N_1018,N_931,N_887);
nand U1019 (N_1019,N_804,N_976);
and U1020 (N_1020,N_893,N_918);
or U1021 (N_1021,N_806,N_983);
nand U1022 (N_1022,N_845,N_932);
or U1023 (N_1023,N_805,N_905);
and U1024 (N_1024,N_965,N_817);
xnor U1025 (N_1025,N_935,N_881);
xor U1026 (N_1026,N_994,N_948);
or U1027 (N_1027,N_807,N_810);
xor U1028 (N_1028,N_852,N_974);
nor U1029 (N_1029,N_814,N_964);
or U1030 (N_1030,N_846,N_851);
nand U1031 (N_1031,N_892,N_847);
or U1032 (N_1032,N_876,N_860);
nor U1033 (N_1033,N_883,N_928);
nand U1034 (N_1034,N_841,N_819);
nand U1035 (N_1035,N_837,N_938);
nor U1036 (N_1036,N_990,N_833);
or U1037 (N_1037,N_890,N_947);
or U1038 (N_1038,N_861,N_951);
and U1039 (N_1039,N_920,N_842);
nand U1040 (N_1040,N_911,N_986);
or U1041 (N_1041,N_854,N_816);
xor U1042 (N_1042,N_917,N_815);
xnor U1043 (N_1043,N_996,N_992);
and U1044 (N_1044,N_995,N_823);
nand U1045 (N_1045,N_941,N_886);
or U1046 (N_1046,N_985,N_984);
nand U1047 (N_1047,N_978,N_997);
and U1048 (N_1048,N_981,N_916);
or U1049 (N_1049,N_959,N_801);
or U1050 (N_1050,N_988,N_894);
nor U1051 (N_1051,N_904,N_825);
nand U1052 (N_1052,N_872,N_827);
nor U1053 (N_1053,N_828,N_864);
xnor U1054 (N_1054,N_874,N_954);
or U1055 (N_1055,N_968,N_897);
nand U1056 (N_1056,N_868,N_973);
nand U1057 (N_1057,N_877,N_840);
nand U1058 (N_1058,N_822,N_812);
nor U1059 (N_1059,N_891,N_939);
nand U1060 (N_1060,N_901,N_913);
nor U1061 (N_1061,N_925,N_950);
or U1062 (N_1062,N_855,N_879);
nor U1063 (N_1063,N_907,N_922);
nand U1064 (N_1064,N_859,N_824);
nor U1065 (N_1065,N_929,N_991);
nor U1066 (N_1066,N_831,N_971);
nor U1067 (N_1067,N_937,N_979);
nor U1068 (N_1068,N_849,N_963);
nand U1069 (N_1069,N_802,N_921);
and U1070 (N_1070,N_906,N_998);
nand U1071 (N_1071,N_924,N_813);
nor U1072 (N_1072,N_914,N_848);
and U1073 (N_1073,N_957,N_956);
and U1074 (N_1074,N_934,N_800);
and U1075 (N_1075,N_869,N_944);
or U1076 (N_1076,N_838,N_821);
or U1077 (N_1077,N_923,N_880);
or U1078 (N_1078,N_912,N_818);
or U1079 (N_1079,N_982,N_871);
nor U1080 (N_1080,N_903,N_858);
nor U1081 (N_1081,N_808,N_942);
xor U1082 (N_1082,N_933,N_926);
and U1083 (N_1083,N_919,N_972);
and U1084 (N_1084,N_961,N_895);
and U1085 (N_1085,N_908,N_853);
nand U1086 (N_1086,N_993,N_910);
and U1087 (N_1087,N_977,N_902);
or U1088 (N_1088,N_866,N_967);
nand U1089 (N_1089,N_958,N_927);
nor U1090 (N_1090,N_873,N_856);
xor U1091 (N_1091,N_975,N_826);
nand U1092 (N_1092,N_839,N_882);
or U1093 (N_1093,N_857,N_962);
nand U1094 (N_1094,N_811,N_915);
xnor U1095 (N_1095,N_989,N_809);
xnor U1096 (N_1096,N_898,N_820);
nand U1097 (N_1097,N_953,N_844);
or U1098 (N_1098,N_966,N_862);
xor U1099 (N_1099,N_863,N_850);
xor U1100 (N_1100,N_956,N_813);
or U1101 (N_1101,N_949,N_945);
nand U1102 (N_1102,N_813,N_931);
or U1103 (N_1103,N_901,N_908);
nor U1104 (N_1104,N_800,N_947);
nand U1105 (N_1105,N_833,N_925);
nor U1106 (N_1106,N_956,N_883);
nor U1107 (N_1107,N_852,N_819);
nand U1108 (N_1108,N_905,N_923);
nand U1109 (N_1109,N_936,N_975);
or U1110 (N_1110,N_826,N_894);
or U1111 (N_1111,N_953,N_988);
and U1112 (N_1112,N_856,N_828);
nand U1113 (N_1113,N_964,N_919);
xnor U1114 (N_1114,N_921,N_863);
nand U1115 (N_1115,N_811,N_883);
or U1116 (N_1116,N_947,N_832);
nand U1117 (N_1117,N_873,N_881);
xnor U1118 (N_1118,N_927,N_974);
and U1119 (N_1119,N_948,N_987);
nand U1120 (N_1120,N_897,N_959);
or U1121 (N_1121,N_932,N_802);
nand U1122 (N_1122,N_911,N_808);
nor U1123 (N_1123,N_814,N_901);
nand U1124 (N_1124,N_853,N_972);
and U1125 (N_1125,N_982,N_877);
or U1126 (N_1126,N_965,N_959);
nand U1127 (N_1127,N_955,N_909);
xnor U1128 (N_1128,N_899,N_809);
nand U1129 (N_1129,N_856,N_972);
xor U1130 (N_1130,N_909,N_881);
and U1131 (N_1131,N_981,N_900);
or U1132 (N_1132,N_941,N_820);
and U1133 (N_1133,N_954,N_937);
nor U1134 (N_1134,N_887,N_890);
or U1135 (N_1135,N_815,N_887);
xnor U1136 (N_1136,N_923,N_979);
nand U1137 (N_1137,N_819,N_981);
or U1138 (N_1138,N_918,N_936);
nor U1139 (N_1139,N_806,N_909);
nand U1140 (N_1140,N_942,N_928);
nand U1141 (N_1141,N_830,N_984);
nand U1142 (N_1142,N_876,N_847);
or U1143 (N_1143,N_927,N_900);
and U1144 (N_1144,N_818,N_862);
and U1145 (N_1145,N_814,N_948);
nor U1146 (N_1146,N_997,N_936);
or U1147 (N_1147,N_885,N_936);
xor U1148 (N_1148,N_887,N_965);
or U1149 (N_1149,N_862,N_857);
or U1150 (N_1150,N_800,N_857);
xnor U1151 (N_1151,N_832,N_958);
xnor U1152 (N_1152,N_943,N_947);
and U1153 (N_1153,N_871,N_816);
nor U1154 (N_1154,N_895,N_969);
or U1155 (N_1155,N_952,N_945);
and U1156 (N_1156,N_875,N_938);
nor U1157 (N_1157,N_895,N_907);
or U1158 (N_1158,N_822,N_901);
or U1159 (N_1159,N_971,N_866);
and U1160 (N_1160,N_884,N_967);
or U1161 (N_1161,N_969,N_907);
nand U1162 (N_1162,N_848,N_954);
nand U1163 (N_1163,N_950,N_977);
or U1164 (N_1164,N_809,N_816);
or U1165 (N_1165,N_873,N_915);
nor U1166 (N_1166,N_840,N_924);
xnor U1167 (N_1167,N_903,N_874);
or U1168 (N_1168,N_906,N_982);
nand U1169 (N_1169,N_818,N_878);
or U1170 (N_1170,N_991,N_846);
and U1171 (N_1171,N_911,N_984);
and U1172 (N_1172,N_960,N_821);
or U1173 (N_1173,N_975,N_965);
or U1174 (N_1174,N_951,N_839);
nor U1175 (N_1175,N_947,N_956);
nor U1176 (N_1176,N_988,N_842);
or U1177 (N_1177,N_883,N_819);
nor U1178 (N_1178,N_831,N_868);
and U1179 (N_1179,N_929,N_949);
nor U1180 (N_1180,N_898,N_871);
nor U1181 (N_1181,N_998,N_981);
nand U1182 (N_1182,N_907,N_960);
nand U1183 (N_1183,N_919,N_904);
or U1184 (N_1184,N_822,N_855);
nand U1185 (N_1185,N_814,N_904);
nor U1186 (N_1186,N_816,N_934);
xor U1187 (N_1187,N_999,N_930);
or U1188 (N_1188,N_941,N_861);
and U1189 (N_1189,N_859,N_917);
nor U1190 (N_1190,N_859,N_902);
nor U1191 (N_1191,N_967,N_964);
nor U1192 (N_1192,N_854,N_917);
nand U1193 (N_1193,N_933,N_861);
nand U1194 (N_1194,N_924,N_871);
and U1195 (N_1195,N_872,N_869);
nor U1196 (N_1196,N_973,N_993);
nand U1197 (N_1197,N_856,N_979);
or U1198 (N_1198,N_963,N_972);
nand U1199 (N_1199,N_941,N_912);
nor U1200 (N_1200,N_1100,N_1190);
or U1201 (N_1201,N_1098,N_1104);
nor U1202 (N_1202,N_1080,N_1150);
or U1203 (N_1203,N_1056,N_1194);
nor U1204 (N_1204,N_1009,N_1182);
and U1205 (N_1205,N_1192,N_1055);
or U1206 (N_1206,N_1162,N_1160);
and U1207 (N_1207,N_1093,N_1019);
and U1208 (N_1208,N_1096,N_1095);
or U1209 (N_1209,N_1127,N_1085);
or U1210 (N_1210,N_1193,N_1136);
nor U1211 (N_1211,N_1010,N_1147);
or U1212 (N_1212,N_1121,N_1043);
nand U1213 (N_1213,N_1082,N_1024);
and U1214 (N_1214,N_1181,N_1040);
or U1215 (N_1215,N_1105,N_1003);
nand U1216 (N_1216,N_1196,N_1076);
and U1217 (N_1217,N_1044,N_1028);
and U1218 (N_1218,N_1049,N_1065);
or U1219 (N_1219,N_1186,N_1035);
and U1220 (N_1220,N_1144,N_1087);
nand U1221 (N_1221,N_1083,N_1107);
nor U1222 (N_1222,N_1119,N_1091);
or U1223 (N_1223,N_1166,N_1124);
nor U1224 (N_1224,N_1089,N_1026);
and U1225 (N_1225,N_1059,N_1167);
nand U1226 (N_1226,N_1061,N_1111);
nor U1227 (N_1227,N_1036,N_1139);
nor U1228 (N_1228,N_1140,N_1015);
or U1229 (N_1229,N_1081,N_1143);
nand U1230 (N_1230,N_1016,N_1042);
and U1231 (N_1231,N_1030,N_1070);
and U1232 (N_1232,N_1156,N_1165);
or U1233 (N_1233,N_1041,N_1155);
and U1234 (N_1234,N_1057,N_1051);
nor U1235 (N_1235,N_1185,N_1176);
and U1236 (N_1236,N_1067,N_1172);
nor U1237 (N_1237,N_1161,N_1189);
nand U1238 (N_1238,N_1000,N_1064);
and U1239 (N_1239,N_1106,N_1163);
and U1240 (N_1240,N_1005,N_1118);
and U1241 (N_1241,N_1017,N_1187);
nor U1242 (N_1242,N_1066,N_1123);
xor U1243 (N_1243,N_1075,N_1006);
nor U1244 (N_1244,N_1126,N_1099);
nand U1245 (N_1245,N_1008,N_1177);
nor U1246 (N_1246,N_1053,N_1020);
and U1247 (N_1247,N_1060,N_1045);
nor U1248 (N_1248,N_1063,N_1029);
nor U1249 (N_1249,N_1102,N_1062);
nor U1250 (N_1250,N_1046,N_1110);
xnor U1251 (N_1251,N_1004,N_1135);
or U1252 (N_1252,N_1047,N_1175);
or U1253 (N_1253,N_1039,N_1131);
nand U1254 (N_1254,N_1113,N_1115);
nor U1255 (N_1255,N_1138,N_1159);
nand U1256 (N_1256,N_1183,N_1178);
nand U1257 (N_1257,N_1050,N_1112);
nor U1258 (N_1258,N_1125,N_1074);
or U1259 (N_1259,N_1164,N_1197);
nand U1260 (N_1260,N_1184,N_1173);
or U1261 (N_1261,N_1191,N_1168);
xnor U1262 (N_1262,N_1097,N_1092);
and U1263 (N_1263,N_1086,N_1025);
or U1264 (N_1264,N_1179,N_1014);
nor U1265 (N_1265,N_1077,N_1058);
nand U1266 (N_1266,N_1145,N_1149);
or U1267 (N_1267,N_1120,N_1033);
and U1268 (N_1268,N_1108,N_1137);
nand U1269 (N_1269,N_1169,N_1171);
nor U1270 (N_1270,N_1130,N_1002);
nand U1271 (N_1271,N_1023,N_1148);
xor U1272 (N_1272,N_1001,N_1132);
nand U1273 (N_1273,N_1195,N_1038);
or U1274 (N_1274,N_1069,N_1198);
and U1275 (N_1275,N_1054,N_1084);
nor U1276 (N_1276,N_1117,N_1153);
or U1277 (N_1277,N_1079,N_1101);
and U1278 (N_1278,N_1007,N_1068);
nor U1279 (N_1279,N_1013,N_1031);
xnor U1280 (N_1280,N_1073,N_1078);
and U1281 (N_1281,N_1174,N_1180);
nor U1282 (N_1282,N_1021,N_1011);
nor U1283 (N_1283,N_1134,N_1037);
xor U1284 (N_1284,N_1052,N_1018);
and U1285 (N_1285,N_1199,N_1152);
or U1286 (N_1286,N_1034,N_1032);
nand U1287 (N_1287,N_1090,N_1071);
nand U1288 (N_1288,N_1154,N_1170);
or U1289 (N_1289,N_1116,N_1158);
nand U1290 (N_1290,N_1151,N_1122);
nor U1291 (N_1291,N_1146,N_1157);
nand U1292 (N_1292,N_1103,N_1072);
and U1293 (N_1293,N_1114,N_1109);
xnor U1294 (N_1294,N_1133,N_1027);
nand U1295 (N_1295,N_1048,N_1188);
or U1296 (N_1296,N_1129,N_1022);
nor U1297 (N_1297,N_1088,N_1141);
nand U1298 (N_1298,N_1128,N_1094);
nor U1299 (N_1299,N_1012,N_1142);
xnor U1300 (N_1300,N_1064,N_1078);
and U1301 (N_1301,N_1165,N_1163);
and U1302 (N_1302,N_1187,N_1024);
nor U1303 (N_1303,N_1119,N_1160);
or U1304 (N_1304,N_1137,N_1058);
nand U1305 (N_1305,N_1126,N_1198);
or U1306 (N_1306,N_1154,N_1153);
xnor U1307 (N_1307,N_1078,N_1173);
or U1308 (N_1308,N_1128,N_1134);
xnor U1309 (N_1309,N_1056,N_1042);
or U1310 (N_1310,N_1046,N_1060);
nor U1311 (N_1311,N_1123,N_1009);
nor U1312 (N_1312,N_1060,N_1197);
xnor U1313 (N_1313,N_1117,N_1173);
xor U1314 (N_1314,N_1178,N_1027);
nand U1315 (N_1315,N_1035,N_1166);
and U1316 (N_1316,N_1119,N_1162);
or U1317 (N_1317,N_1016,N_1081);
nand U1318 (N_1318,N_1046,N_1035);
nor U1319 (N_1319,N_1038,N_1036);
and U1320 (N_1320,N_1072,N_1166);
and U1321 (N_1321,N_1048,N_1032);
or U1322 (N_1322,N_1012,N_1125);
nor U1323 (N_1323,N_1026,N_1082);
or U1324 (N_1324,N_1149,N_1157);
nor U1325 (N_1325,N_1090,N_1197);
xor U1326 (N_1326,N_1091,N_1052);
and U1327 (N_1327,N_1084,N_1170);
or U1328 (N_1328,N_1032,N_1153);
nor U1329 (N_1329,N_1143,N_1014);
xor U1330 (N_1330,N_1017,N_1141);
and U1331 (N_1331,N_1039,N_1030);
nand U1332 (N_1332,N_1040,N_1139);
nor U1333 (N_1333,N_1116,N_1056);
or U1334 (N_1334,N_1087,N_1138);
nand U1335 (N_1335,N_1199,N_1082);
or U1336 (N_1336,N_1124,N_1034);
and U1337 (N_1337,N_1090,N_1181);
and U1338 (N_1338,N_1066,N_1016);
and U1339 (N_1339,N_1031,N_1195);
nand U1340 (N_1340,N_1198,N_1146);
nand U1341 (N_1341,N_1095,N_1058);
nand U1342 (N_1342,N_1173,N_1051);
nand U1343 (N_1343,N_1171,N_1107);
and U1344 (N_1344,N_1090,N_1180);
or U1345 (N_1345,N_1190,N_1008);
nand U1346 (N_1346,N_1107,N_1047);
and U1347 (N_1347,N_1093,N_1173);
nor U1348 (N_1348,N_1184,N_1047);
nor U1349 (N_1349,N_1147,N_1110);
or U1350 (N_1350,N_1134,N_1173);
or U1351 (N_1351,N_1056,N_1072);
nor U1352 (N_1352,N_1095,N_1112);
or U1353 (N_1353,N_1098,N_1015);
nor U1354 (N_1354,N_1176,N_1085);
and U1355 (N_1355,N_1117,N_1027);
and U1356 (N_1356,N_1196,N_1123);
nand U1357 (N_1357,N_1007,N_1017);
or U1358 (N_1358,N_1180,N_1199);
and U1359 (N_1359,N_1187,N_1075);
and U1360 (N_1360,N_1165,N_1104);
xnor U1361 (N_1361,N_1125,N_1030);
nor U1362 (N_1362,N_1199,N_1041);
nor U1363 (N_1363,N_1092,N_1063);
and U1364 (N_1364,N_1040,N_1052);
and U1365 (N_1365,N_1043,N_1124);
nand U1366 (N_1366,N_1192,N_1021);
nand U1367 (N_1367,N_1154,N_1150);
nand U1368 (N_1368,N_1121,N_1169);
and U1369 (N_1369,N_1073,N_1017);
or U1370 (N_1370,N_1053,N_1060);
nor U1371 (N_1371,N_1026,N_1180);
nor U1372 (N_1372,N_1039,N_1019);
xnor U1373 (N_1373,N_1167,N_1184);
and U1374 (N_1374,N_1195,N_1148);
nor U1375 (N_1375,N_1115,N_1100);
nor U1376 (N_1376,N_1160,N_1145);
and U1377 (N_1377,N_1169,N_1050);
nand U1378 (N_1378,N_1117,N_1141);
nor U1379 (N_1379,N_1047,N_1105);
xnor U1380 (N_1380,N_1055,N_1029);
and U1381 (N_1381,N_1001,N_1081);
and U1382 (N_1382,N_1146,N_1192);
or U1383 (N_1383,N_1124,N_1038);
and U1384 (N_1384,N_1074,N_1191);
nand U1385 (N_1385,N_1190,N_1120);
or U1386 (N_1386,N_1165,N_1067);
or U1387 (N_1387,N_1096,N_1116);
nor U1388 (N_1388,N_1094,N_1188);
and U1389 (N_1389,N_1072,N_1088);
and U1390 (N_1390,N_1156,N_1012);
nor U1391 (N_1391,N_1076,N_1003);
and U1392 (N_1392,N_1076,N_1005);
xnor U1393 (N_1393,N_1015,N_1139);
nor U1394 (N_1394,N_1029,N_1048);
or U1395 (N_1395,N_1082,N_1036);
nor U1396 (N_1396,N_1091,N_1135);
and U1397 (N_1397,N_1145,N_1060);
or U1398 (N_1398,N_1114,N_1159);
xor U1399 (N_1399,N_1078,N_1139);
nor U1400 (N_1400,N_1237,N_1318);
nor U1401 (N_1401,N_1337,N_1308);
xor U1402 (N_1402,N_1234,N_1369);
nor U1403 (N_1403,N_1288,N_1353);
xor U1404 (N_1404,N_1329,N_1378);
xor U1405 (N_1405,N_1219,N_1304);
nand U1406 (N_1406,N_1356,N_1231);
and U1407 (N_1407,N_1362,N_1306);
and U1408 (N_1408,N_1317,N_1243);
nor U1409 (N_1409,N_1289,N_1343);
xnor U1410 (N_1410,N_1293,N_1204);
or U1411 (N_1411,N_1344,N_1380);
xor U1412 (N_1412,N_1280,N_1364);
or U1413 (N_1413,N_1248,N_1349);
or U1414 (N_1414,N_1253,N_1225);
nor U1415 (N_1415,N_1249,N_1257);
or U1416 (N_1416,N_1340,N_1292);
nand U1417 (N_1417,N_1295,N_1279);
or U1418 (N_1418,N_1213,N_1205);
or U1419 (N_1419,N_1332,N_1223);
nor U1420 (N_1420,N_1321,N_1247);
or U1421 (N_1421,N_1323,N_1284);
and U1422 (N_1422,N_1316,N_1265);
nor U1423 (N_1423,N_1324,N_1297);
or U1424 (N_1424,N_1250,N_1387);
nand U1425 (N_1425,N_1375,N_1334);
and U1426 (N_1426,N_1273,N_1202);
and U1427 (N_1427,N_1258,N_1326);
or U1428 (N_1428,N_1281,N_1392);
nand U1429 (N_1429,N_1301,N_1307);
and U1430 (N_1430,N_1294,N_1239);
xnor U1431 (N_1431,N_1212,N_1328);
nor U1432 (N_1432,N_1261,N_1252);
or U1433 (N_1433,N_1347,N_1310);
or U1434 (N_1434,N_1256,N_1206);
nor U1435 (N_1435,N_1263,N_1389);
and U1436 (N_1436,N_1386,N_1331);
nor U1437 (N_1437,N_1207,N_1325);
nor U1438 (N_1438,N_1214,N_1246);
or U1439 (N_1439,N_1228,N_1235);
nor U1440 (N_1440,N_1300,N_1285);
nand U1441 (N_1441,N_1287,N_1391);
nand U1442 (N_1442,N_1299,N_1309);
nand U1443 (N_1443,N_1278,N_1314);
and U1444 (N_1444,N_1365,N_1333);
xor U1445 (N_1445,N_1381,N_1264);
nand U1446 (N_1446,N_1254,N_1335);
nand U1447 (N_1447,N_1251,N_1315);
and U1448 (N_1448,N_1377,N_1218);
nor U1449 (N_1449,N_1255,N_1360);
nand U1450 (N_1450,N_1373,N_1245);
or U1451 (N_1451,N_1348,N_1221);
xor U1452 (N_1452,N_1296,N_1262);
or U1453 (N_1453,N_1211,N_1275);
or U1454 (N_1454,N_1398,N_1216);
nor U1455 (N_1455,N_1371,N_1282);
and U1456 (N_1456,N_1269,N_1267);
and U1457 (N_1457,N_1266,N_1209);
or U1458 (N_1458,N_1270,N_1240);
nor U1459 (N_1459,N_1286,N_1390);
nand U1460 (N_1460,N_1352,N_1217);
nor U1461 (N_1461,N_1220,N_1305);
nand U1462 (N_1462,N_1203,N_1394);
nand U1463 (N_1463,N_1260,N_1372);
nand U1464 (N_1464,N_1366,N_1388);
nand U1465 (N_1465,N_1383,N_1367);
and U1466 (N_1466,N_1290,N_1313);
nor U1467 (N_1467,N_1342,N_1302);
or U1468 (N_1468,N_1238,N_1396);
nand U1469 (N_1469,N_1227,N_1276);
and U1470 (N_1470,N_1271,N_1355);
or U1471 (N_1471,N_1230,N_1229);
or U1472 (N_1472,N_1222,N_1345);
or U1473 (N_1473,N_1330,N_1376);
and U1474 (N_1474,N_1320,N_1298);
nor U1475 (N_1475,N_1354,N_1339);
and U1476 (N_1476,N_1233,N_1395);
xnor U1477 (N_1477,N_1399,N_1200);
and U1478 (N_1478,N_1338,N_1379);
xnor U1479 (N_1479,N_1359,N_1312);
nand U1480 (N_1480,N_1368,N_1201);
or U1481 (N_1481,N_1327,N_1272);
nor U1482 (N_1482,N_1241,N_1336);
nor U1483 (N_1483,N_1351,N_1277);
and U1484 (N_1484,N_1397,N_1370);
nor U1485 (N_1485,N_1346,N_1341);
and U1486 (N_1486,N_1259,N_1303);
xnor U1487 (N_1487,N_1384,N_1210);
xnor U1488 (N_1488,N_1232,N_1226);
nand U1489 (N_1489,N_1244,N_1224);
and U1490 (N_1490,N_1358,N_1357);
and U1491 (N_1491,N_1385,N_1350);
nand U1492 (N_1492,N_1274,N_1311);
nand U1493 (N_1493,N_1236,N_1208);
nor U1494 (N_1494,N_1393,N_1268);
nand U1495 (N_1495,N_1283,N_1319);
and U1496 (N_1496,N_1291,N_1382);
and U1497 (N_1497,N_1374,N_1363);
nand U1498 (N_1498,N_1215,N_1322);
or U1499 (N_1499,N_1361,N_1242);
and U1500 (N_1500,N_1371,N_1354);
nand U1501 (N_1501,N_1239,N_1243);
or U1502 (N_1502,N_1235,N_1308);
and U1503 (N_1503,N_1365,N_1315);
nand U1504 (N_1504,N_1340,N_1314);
and U1505 (N_1505,N_1340,N_1389);
or U1506 (N_1506,N_1285,N_1345);
xnor U1507 (N_1507,N_1362,N_1254);
nor U1508 (N_1508,N_1247,N_1204);
or U1509 (N_1509,N_1208,N_1264);
and U1510 (N_1510,N_1320,N_1358);
nor U1511 (N_1511,N_1357,N_1345);
or U1512 (N_1512,N_1375,N_1356);
nor U1513 (N_1513,N_1380,N_1219);
nor U1514 (N_1514,N_1230,N_1244);
nand U1515 (N_1515,N_1227,N_1349);
nor U1516 (N_1516,N_1208,N_1274);
or U1517 (N_1517,N_1270,N_1383);
and U1518 (N_1518,N_1287,N_1397);
nand U1519 (N_1519,N_1229,N_1269);
nor U1520 (N_1520,N_1398,N_1318);
and U1521 (N_1521,N_1389,N_1264);
nor U1522 (N_1522,N_1303,N_1288);
nor U1523 (N_1523,N_1333,N_1254);
and U1524 (N_1524,N_1250,N_1324);
and U1525 (N_1525,N_1358,N_1242);
and U1526 (N_1526,N_1230,N_1321);
or U1527 (N_1527,N_1242,N_1376);
nor U1528 (N_1528,N_1260,N_1395);
or U1529 (N_1529,N_1207,N_1285);
or U1530 (N_1530,N_1398,N_1242);
and U1531 (N_1531,N_1304,N_1267);
nor U1532 (N_1532,N_1302,N_1357);
and U1533 (N_1533,N_1240,N_1238);
and U1534 (N_1534,N_1372,N_1399);
or U1535 (N_1535,N_1244,N_1354);
and U1536 (N_1536,N_1233,N_1391);
nor U1537 (N_1537,N_1297,N_1223);
and U1538 (N_1538,N_1295,N_1352);
nand U1539 (N_1539,N_1287,N_1293);
and U1540 (N_1540,N_1304,N_1388);
and U1541 (N_1541,N_1396,N_1252);
or U1542 (N_1542,N_1233,N_1344);
xnor U1543 (N_1543,N_1398,N_1282);
nand U1544 (N_1544,N_1250,N_1319);
xor U1545 (N_1545,N_1246,N_1238);
nand U1546 (N_1546,N_1358,N_1307);
nor U1547 (N_1547,N_1395,N_1373);
or U1548 (N_1548,N_1226,N_1201);
or U1549 (N_1549,N_1249,N_1236);
or U1550 (N_1550,N_1380,N_1281);
nand U1551 (N_1551,N_1307,N_1208);
nor U1552 (N_1552,N_1262,N_1341);
and U1553 (N_1553,N_1369,N_1322);
nor U1554 (N_1554,N_1224,N_1207);
and U1555 (N_1555,N_1388,N_1290);
nand U1556 (N_1556,N_1293,N_1300);
nand U1557 (N_1557,N_1362,N_1282);
or U1558 (N_1558,N_1386,N_1359);
and U1559 (N_1559,N_1331,N_1210);
nand U1560 (N_1560,N_1257,N_1255);
nor U1561 (N_1561,N_1248,N_1224);
or U1562 (N_1562,N_1297,N_1367);
nand U1563 (N_1563,N_1318,N_1302);
or U1564 (N_1564,N_1382,N_1342);
and U1565 (N_1565,N_1233,N_1288);
and U1566 (N_1566,N_1346,N_1393);
xnor U1567 (N_1567,N_1233,N_1206);
and U1568 (N_1568,N_1352,N_1202);
or U1569 (N_1569,N_1353,N_1293);
and U1570 (N_1570,N_1292,N_1373);
and U1571 (N_1571,N_1314,N_1359);
or U1572 (N_1572,N_1363,N_1235);
or U1573 (N_1573,N_1276,N_1245);
or U1574 (N_1574,N_1242,N_1324);
xor U1575 (N_1575,N_1255,N_1325);
or U1576 (N_1576,N_1356,N_1398);
or U1577 (N_1577,N_1324,N_1235);
or U1578 (N_1578,N_1248,N_1358);
or U1579 (N_1579,N_1255,N_1247);
and U1580 (N_1580,N_1344,N_1376);
and U1581 (N_1581,N_1381,N_1377);
or U1582 (N_1582,N_1299,N_1241);
nor U1583 (N_1583,N_1301,N_1240);
nand U1584 (N_1584,N_1240,N_1219);
nor U1585 (N_1585,N_1224,N_1218);
nand U1586 (N_1586,N_1397,N_1226);
xor U1587 (N_1587,N_1222,N_1318);
and U1588 (N_1588,N_1239,N_1330);
and U1589 (N_1589,N_1319,N_1379);
nand U1590 (N_1590,N_1292,N_1298);
nand U1591 (N_1591,N_1235,N_1305);
nand U1592 (N_1592,N_1381,N_1314);
nand U1593 (N_1593,N_1382,N_1229);
and U1594 (N_1594,N_1316,N_1324);
nor U1595 (N_1595,N_1269,N_1203);
or U1596 (N_1596,N_1324,N_1360);
nand U1597 (N_1597,N_1261,N_1250);
nor U1598 (N_1598,N_1329,N_1240);
nor U1599 (N_1599,N_1259,N_1214);
nor U1600 (N_1600,N_1512,N_1413);
nand U1601 (N_1601,N_1555,N_1505);
or U1602 (N_1602,N_1401,N_1547);
or U1603 (N_1603,N_1490,N_1501);
nor U1604 (N_1604,N_1408,N_1492);
and U1605 (N_1605,N_1587,N_1471);
and U1606 (N_1606,N_1565,N_1524);
or U1607 (N_1607,N_1446,N_1405);
nand U1608 (N_1608,N_1516,N_1462);
xor U1609 (N_1609,N_1450,N_1518);
nand U1610 (N_1610,N_1478,N_1507);
or U1611 (N_1611,N_1578,N_1564);
xor U1612 (N_1612,N_1553,N_1498);
nor U1613 (N_1613,N_1530,N_1540);
and U1614 (N_1614,N_1593,N_1489);
nor U1615 (N_1615,N_1594,N_1487);
or U1616 (N_1616,N_1491,N_1438);
nand U1617 (N_1617,N_1580,N_1416);
or U1618 (N_1618,N_1430,N_1597);
nor U1619 (N_1619,N_1543,N_1452);
and U1620 (N_1620,N_1417,N_1402);
xor U1621 (N_1621,N_1460,N_1411);
nor U1622 (N_1622,N_1421,N_1534);
and U1623 (N_1623,N_1483,N_1585);
nand U1624 (N_1624,N_1464,N_1445);
and U1625 (N_1625,N_1476,N_1549);
nor U1626 (N_1626,N_1496,N_1493);
nand U1627 (N_1627,N_1560,N_1531);
nand U1628 (N_1628,N_1463,N_1538);
nand U1629 (N_1629,N_1584,N_1514);
and U1630 (N_1630,N_1554,N_1466);
nand U1631 (N_1631,N_1432,N_1403);
and U1632 (N_1632,N_1522,N_1418);
xnor U1633 (N_1633,N_1599,N_1509);
or U1634 (N_1634,N_1448,N_1563);
or U1635 (N_1635,N_1495,N_1423);
nand U1636 (N_1636,N_1519,N_1447);
nor U1637 (N_1637,N_1488,N_1459);
nor U1638 (N_1638,N_1535,N_1461);
or U1639 (N_1639,N_1470,N_1588);
nand U1640 (N_1640,N_1454,N_1542);
nand U1641 (N_1641,N_1465,N_1412);
and U1642 (N_1642,N_1410,N_1548);
nor U1643 (N_1643,N_1520,N_1550);
xor U1644 (N_1644,N_1526,N_1596);
nand U1645 (N_1645,N_1428,N_1433);
nand U1646 (N_1646,N_1467,N_1582);
or U1647 (N_1647,N_1562,N_1575);
xor U1648 (N_1648,N_1482,N_1533);
and U1649 (N_1649,N_1571,N_1529);
and U1650 (N_1650,N_1474,N_1473);
xor U1651 (N_1651,N_1427,N_1545);
nand U1652 (N_1652,N_1481,N_1424);
nand U1653 (N_1653,N_1472,N_1544);
nand U1654 (N_1654,N_1570,N_1523);
nand U1655 (N_1655,N_1579,N_1451);
nand U1656 (N_1656,N_1400,N_1532);
or U1657 (N_1657,N_1485,N_1415);
and U1658 (N_1658,N_1572,N_1589);
nand U1659 (N_1659,N_1458,N_1431);
nor U1660 (N_1660,N_1442,N_1573);
or U1661 (N_1661,N_1577,N_1528);
and U1662 (N_1662,N_1502,N_1497);
or U1663 (N_1663,N_1557,N_1499);
and U1664 (N_1664,N_1574,N_1590);
and U1665 (N_1665,N_1419,N_1515);
nor U1666 (N_1666,N_1468,N_1444);
and U1667 (N_1667,N_1581,N_1443);
nor U1668 (N_1668,N_1511,N_1494);
nor U1669 (N_1669,N_1404,N_1434);
or U1670 (N_1670,N_1521,N_1552);
xnor U1671 (N_1671,N_1500,N_1569);
nor U1672 (N_1672,N_1551,N_1475);
nand U1673 (N_1673,N_1561,N_1504);
nor U1674 (N_1674,N_1539,N_1536);
nor U1675 (N_1675,N_1559,N_1592);
or U1676 (N_1676,N_1591,N_1558);
or U1677 (N_1677,N_1414,N_1429);
nand U1678 (N_1678,N_1527,N_1409);
or U1679 (N_1679,N_1513,N_1510);
and U1680 (N_1680,N_1541,N_1508);
or U1681 (N_1681,N_1598,N_1435);
nand U1682 (N_1682,N_1583,N_1469);
or U1683 (N_1683,N_1586,N_1546);
nor U1684 (N_1684,N_1420,N_1426);
nand U1685 (N_1685,N_1595,N_1455);
or U1686 (N_1686,N_1456,N_1506);
nand U1687 (N_1687,N_1436,N_1525);
nand U1688 (N_1688,N_1479,N_1567);
nor U1689 (N_1689,N_1425,N_1440);
and U1690 (N_1690,N_1449,N_1406);
and U1691 (N_1691,N_1439,N_1407);
nand U1692 (N_1692,N_1453,N_1484);
and U1693 (N_1693,N_1441,N_1537);
nor U1694 (N_1694,N_1517,N_1556);
xnor U1695 (N_1695,N_1437,N_1568);
or U1696 (N_1696,N_1566,N_1503);
nor U1697 (N_1697,N_1576,N_1480);
and U1698 (N_1698,N_1486,N_1422);
and U1699 (N_1699,N_1477,N_1457);
or U1700 (N_1700,N_1592,N_1471);
xor U1701 (N_1701,N_1458,N_1558);
nor U1702 (N_1702,N_1524,N_1571);
nand U1703 (N_1703,N_1484,N_1401);
nand U1704 (N_1704,N_1486,N_1460);
or U1705 (N_1705,N_1592,N_1585);
nand U1706 (N_1706,N_1526,N_1588);
and U1707 (N_1707,N_1437,N_1515);
or U1708 (N_1708,N_1596,N_1557);
and U1709 (N_1709,N_1433,N_1506);
nor U1710 (N_1710,N_1558,N_1454);
or U1711 (N_1711,N_1521,N_1598);
or U1712 (N_1712,N_1562,N_1494);
nor U1713 (N_1713,N_1586,N_1587);
and U1714 (N_1714,N_1431,N_1436);
nor U1715 (N_1715,N_1510,N_1452);
or U1716 (N_1716,N_1450,N_1551);
nand U1717 (N_1717,N_1472,N_1414);
xor U1718 (N_1718,N_1407,N_1571);
and U1719 (N_1719,N_1571,N_1430);
nor U1720 (N_1720,N_1402,N_1547);
or U1721 (N_1721,N_1462,N_1405);
nand U1722 (N_1722,N_1474,N_1468);
and U1723 (N_1723,N_1458,N_1471);
and U1724 (N_1724,N_1449,N_1579);
nand U1725 (N_1725,N_1409,N_1519);
or U1726 (N_1726,N_1541,N_1490);
nor U1727 (N_1727,N_1546,N_1409);
or U1728 (N_1728,N_1426,N_1514);
nand U1729 (N_1729,N_1542,N_1502);
and U1730 (N_1730,N_1510,N_1461);
nand U1731 (N_1731,N_1527,N_1444);
and U1732 (N_1732,N_1462,N_1422);
nor U1733 (N_1733,N_1584,N_1561);
or U1734 (N_1734,N_1414,N_1559);
nand U1735 (N_1735,N_1425,N_1492);
nor U1736 (N_1736,N_1445,N_1510);
and U1737 (N_1737,N_1503,N_1454);
nand U1738 (N_1738,N_1452,N_1496);
xor U1739 (N_1739,N_1438,N_1474);
and U1740 (N_1740,N_1497,N_1551);
or U1741 (N_1741,N_1479,N_1497);
and U1742 (N_1742,N_1569,N_1477);
nor U1743 (N_1743,N_1562,N_1404);
nor U1744 (N_1744,N_1471,N_1552);
and U1745 (N_1745,N_1501,N_1531);
nor U1746 (N_1746,N_1431,N_1481);
nor U1747 (N_1747,N_1468,N_1441);
nor U1748 (N_1748,N_1511,N_1480);
and U1749 (N_1749,N_1452,N_1421);
nand U1750 (N_1750,N_1556,N_1430);
or U1751 (N_1751,N_1451,N_1588);
and U1752 (N_1752,N_1596,N_1552);
nor U1753 (N_1753,N_1570,N_1481);
nor U1754 (N_1754,N_1504,N_1566);
or U1755 (N_1755,N_1519,N_1404);
or U1756 (N_1756,N_1546,N_1427);
and U1757 (N_1757,N_1444,N_1488);
and U1758 (N_1758,N_1537,N_1545);
and U1759 (N_1759,N_1496,N_1518);
or U1760 (N_1760,N_1568,N_1510);
xnor U1761 (N_1761,N_1520,N_1495);
or U1762 (N_1762,N_1548,N_1423);
nand U1763 (N_1763,N_1498,N_1509);
nand U1764 (N_1764,N_1568,N_1522);
and U1765 (N_1765,N_1590,N_1556);
and U1766 (N_1766,N_1438,N_1430);
and U1767 (N_1767,N_1543,N_1438);
nor U1768 (N_1768,N_1425,N_1566);
and U1769 (N_1769,N_1449,N_1550);
and U1770 (N_1770,N_1472,N_1477);
nor U1771 (N_1771,N_1533,N_1562);
xor U1772 (N_1772,N_1472,N_1574);
and U1773 (N_1773,N_1573,N_1490);
nand U1774 (N_1774,N_1585,N_1594);
nor U1775 (N_1775,N_1559,N_1505);
and U1776 (N_1776,N_1493,N_1429);
and U1777 (N_1777,N_1532,N_1441);
or U1778 (N_1778,N_1470,N_1586);
nor U1779 (N_1779,N_1498,N_1421);
nor U1780 (N_1780,N_1481,N_1437);
or U1781 (N_1781,N_1454,N_1473);
nand U1782 (N_1782,N_1539,N_1407);
xnor U1783 (N_1783,N_1577,N_1553);
and U1784 (N_1784,N_1596,N_1525);
nor U1785 (N_1785,N_1412,N_1501);
and U1786 (N_1786,N_1500,N_1552);
and U1787 (N_1787,N_1504,N_1533);
and U1788 (N_1788,N_1541,N_1503);
and U1789 (N_1789,N_1533,N_1571);
nand U1790 (N_1790,N_1401,N_1430);
nand U1791 (N_1791,N_1591,N_1457);
and U1792 (N_1792,N_1536,N_1523);
nor U1793 (N_1793,N_1564,N_1503);
or U1794 (N_1794,N_1444,N_1548);
and U1795 (N_1795,N_1474,N_1553);
or U1796 (N_1796,N_1443,N_1573);
nor U1797 (N_1797,N_1580,N_1492);
nand U1798 (N_1798,N_1543,N_1518);
nor U1799 (N_1799,N_1480,N_1562);
nor U1800 (N_1800,N_1718,N_1693);
nand U1801 (N_1801,N_1613,N_1759);
and U1802 (N_1802,N_1659,N_1711);
nor U1803 (N_1803,N_1676,N_1608);
or U1804 (N_1804,N_1771,N_1698);
nor U1805 (N_1805,N_1794,N_1627);
and U1806 (N_1806,N_1722,N_1728);
and U1807 (N_1807,N_1607,N_1615);
or U1808 (N_1808,N_1609,N_1719);
nor U1809 (N_1809,N_1733,N_1618);
nand U1810 (N_1810,N_1656,N_1649);
and U1811 (N_1811,N_1604,N_1663);
or U1812 (N_1812,N_1681,N_1764);
xor U1813 (N_1813,N_1601,N_1738);
nand U1814 (N_1814,N_1640,N_1625);
xor U1815 (N_1815,N_1798,N_1763);
or U1816 (N_1816,N_1780,N_1707);
or U1817 (N_1817,N_1743,N_1732);
nor U1818 (N_1818,N_1713,N_1611);
xor U1819 (N_1819,N_1778,N_1682);
nand U1820 (N_1820,N_1715,N_1716);
nand U1821 (N_1821,N_1773,N_1660);
nand U1822 (N_1822,N_1644,N_1740);
nor U1823 (N_1823,N_1638,N_1623);
or U1824 (N_1824,N_1662,N_1650);
or U1825 (N_1825,N_1755,N_1674);
nand U1826 (N_1826,N_1709,N_1683);
nor U1827 (N_1827,N_1687,N_1782);
and U1828 (N_1828,N_1767,N_1741);
nand U1829 (N_1829,N_1726,N_1749);
nand U1830 (N_1830,N_1723,N_1757);
xor U1831 (N_1831,N_1793,N_1702);
nand U1832 (N_1832,N_1747,N_1641);
nand U1833 (N_1833,N_1686,N_1622);
nand U1834 (N_1834,N_1671,N_1721);
nand U1835 (N_1835,N_1751,N_1673);
and U1836 (N_1836,N_1626,N_1768);
nor U1837 (N_1837,N_1787,N_1727);
nor U1838 (N_1838,N_1679,N_1642);
nand U1839 (N_1839,N_1668,N_1678);
xor U1840 (N_1840,N_1729,N_1691);
xor U1841 (N_1841,N_1756,N_1672);
nand U1842 (N_1842,N_1720,N_1704);
and U1843 (N_1843,N_1788,N_1688);
nor U1844 (N_1844,N_1657,N_1648);
xnor U1845 (N_1845,N_1635,N_1708);
and U1846 (N_1846,N_1646,N_1637);
and U1847 (N_1847,N_1760,N_1700);
or U1848 (N_1848,N_1724,N_1603);
nand U1849 (N_1849,N_1610,N_1765);
nor U1850 (N_1850,N_1776,N_1617);
or U1851 (N_1851,N_1777,N_1664);
nand U1852 (N_1852,N_1792,N_1620);
and U1853 (N_1853,N_1670,N_1628);
nor U1854 (N_1854,N_1789,N_1614);
nand U1855 (N_1855,N_1624,N_1612);
or U1856 (N_1856,N_1631,N_1616);
nor U1857 (N_1857,N_1653,N_1643);
nand U1858 (N_1858,N_1761,N_1742);
and U1859 (N_1859,N_1621,N_1651);
and U1860 (N_1860,N_1694,N_1697);
or U1861 (N_1861,N_1665,N_1745);
nor U1862 (N_1862,N_1645,N_1606);
xor U1863 (N_1863,N_1696,N_1796);
or U1864 (N_1864,N_1797,N_1762);
xnor U1865 (N_1865,N_1735,N_1705);
nor U1866 (N_1866,N_1689,N_1712);
nand U1867 (N_1867,N_1717,N_1669);
and U1868 (N_1868,N_1690,N_1731);
nor U1869 (N_1869,N_1750,N_1799);
nor U1870 (N_1870,N_1632,N_1739);
nand U1871 (N_1871,N_1675,N_1725);
nand U1872 (N_1872,N_1661,N_1752);
and U1873 (N_1873,N_1685,N_1647);
xnor U1874 (N_1874,N_1658,N_1680);
nand U1875 (N_1875,N_1695,N_1706);
and U1876 (N_1876,N_1786,N_1744);
xnor U1877 (N_1877,N_1766,N_1667);
nand U1878 (N_1878,N_1710,N_1795);
or U1879 (N_1879,N_1783,N_1774);
nand U1880 (N_1880,N_1701,N_1779);
or U1881 (N_1881,N_1605,N_1684);
or U1882 (N_1882,N_1703,N_1746);
nand U1883 (N_1883,N_1734,N_1775);
and U1884 (N_1884,N_1619,N_1666);
xnor U1885 (N_1885,N_1677,N_1748);
nand U1886 (N_1886,N_1600,N_1770);
nor U1887 (N_1887,N_1753,N_1790);
nand U1888 (N_1888,N_1772,N_1754);
nand U1889 (N_1889,N_1781,N_1655);
and U1890 (N_1890,N_1636,N_1629);
or U1891 (N_1891,N_1699,N_1639);
and U1892 (N_1892,N_1633,N_1791);
nand U1893 (N_1893,N_1652,N_1730);
nor U1894 (N_1894,N_1736,N_1714);
nand U1895 (N_1895,N_1784,N_1630);
and U1896 (N_1896,N_1602,N_1634);
nor U1897 (N_1897,N_1785,N_1758);
nor U1898 (N_1898,N_1769,N_1737);
nand U1899 (N_1899,N_1692,N_1654);
xor U1900 (N_1900,N_1743,N_1660);
nand U1901 (N_1901,N_1793,N_1651);
and U1902 (N_1902,N_1704,N_1776);
nand U1903 (N_1903,N_1692,N_1663);
and U1904 (N_1904,N_1603,N_1715);
or U1905 (N_1905,N_1629,N_1752);
nor U1906 (N_1906,N_1715,N_1769);
nand U1907 (N_1907,N_1751,N_1780);
nand U1908 (N_1908,N_1796,N_1652);
nand U1909 (N_1909,N_1634,N_1720);
or U1910 (N_1910,N_1796,N_1750);
or U1911 (N_1911,N_1729,N_1741);
nand U1912 (N_1912,N_1764,N_1771);
and U1913 (N_1913,N_1714,N_1698);
nand U1914 (N_1914,N_1752,N_1721);
and U1915 (N_1915,N_1745,N_1751);
nand U1916 (N_1916,N_1659,N_1778);
nor U1917 (N_1917,N_1672,N_1779);
or U1918 (N_1918,N_1714,N_1631);
or U1919 (N_1919,N_1738,N_1610);
and U1920 (N_1920,N_1659,N_1751);
xor U1921 (N_1921,N_1752,N_1706);
and U1922 (N_1922,N_1765,N_1625);
xnor U1923 (N_1923,N_1650,N_1698);
nor U1924 (N_1924,N_1691,N_1795);
or U1925 (N_1925,N_1648,N_1612);
and U1926 (N_1926,N_1732,N_1794);
or U1927 (N_1927,N_1620,N_1615);
and U1928 (N_1928,N_1786,N_1765);
nand U1929 (N_1929,N_1726,N_1761);
and U1930 (N_1930,N_1646,N_1713);
nand U1931 (N_1931,N_1614,N_1778);
xnor U1932 (N_1932,N_1730,N_1733);
nand U1933 (N_1933,N_1688,N_1630);
nor U1934 (N_1934,N_1788,N_1757);
nor U1935 (N_1935,N_1776,N_1649);
or U1936 (N_1936,N_1604,N_1638);
and U1937 (N_1937,N_1736,N_1757);
nand U1938 (N_1938,N_1792,N_1756);
or U1939 (N_1939,N_1702,N_1663);
nor U1940 (N_1940,N_1796,N_1721);
or U1941 (N_1941,N_1624,N_1673);
nor U1942 (N_1942,N_1629,N_1698);
nand U1943 (N_1943,N_1636,N_1791);
or U1944 (N_1944,N_1780,N_1726);
nor U1945 (N_1945,N_1743,N_1650);
nand U1946 (N_1946,N_1766,N_1723);
nor U1947 (N_1947,N_1731,N_1668);
nor U1948 (N_1948,N_1716,N_1691);
nor U1949 (N_1949,N_1663,N_1738);
nor U1950 (N_1950,N_1615,N_1702);
or U1951 (N_1951,N_1634,N_1726);
and U1952 (N_1952,N_1751,N_1775);
nand U1953 (N_1953,N_1644,N_1605);
and U1954 (N_1954,N_1649,N_1668);
and U1955 (N_1955,N_1766,N_1765);
nor U1956 (N_1956,N_1760,N_1775);
or U1957 (N_1957,N_1773,N_1797);
nand U1958 (N_1958,N_1785,N_1791);
and U1959 (N_1959,N_1794,N_1662);
nor U1960 (N_1960,N_1679,N_1750);
nand U1961 (N_1961,N_1784,N_1603);
and U1962 (N_1962,N_1751,N_1664);
nor U1963 (N_1963,N_1738,N_1697);
nor U1964 (N_1964,N_1615,N_1732);
nor U1965 (N_1965,N_1602,N_1799);
nand U1966 (N_1966,N_1656,N_1624);
nand U1967 (N_1967,N_1618,N_1677);
or U1968 (N_1968,N_1748,N_1757);
and U1969 (N_1969,N_1624,N_1683);
or U1970 (N_1970,N_1699,N_1625);
nor U1971 (N_1971,N_1745,N_1686);
and U1972 (N_1972,N_1604,N_1736);
or U1973 (N_1973,N_1764,N_1685);
nand U1974 (N_1974,N_1750,N_1698);
or U1975 (N_1975,N_1607,N_1630);
nand U1976 (N_1976,N_1701,N_1724);
nand U1977 (N_1977,N_1697,N_1754);
xnor U1978 (N_1978,N_1651,N_1697);
nor U1979 (N_1979,N_1730,N_1667);
nand U1980 (N_1980,N_1769,N_1773);
and U1981 (N_1981,N_1674,N_1628);
nand U1982 (N_1982,N_1704,N_1742);
or U1983 (N_1983,N_1690,N_1753);
xnor U1984 (N_1984,N_1689,N_1796);
nor U1985 (N_1985,N_1731,N_1781);
and U1986 (N_1986,N_1754,N_1654);
nor U1987 (N_1987,N_1782,N_1715);
nand U1988 (N_1988,N_1639,N_1772);
or U1989 (N_1989,N_1774,N_1661);
nor U1990 (N_1990,N_1781,N_1620);
or U1991 (N_1991,N_1606,N_1613);
or U1992 (N_1992,N_1704,N_1604);
nand U1993 (N_1993,N_1743,N_1684);
and U1994 (N_1994,N_1750,N_1646);
or U1995 (N_1995,N_1706,N_1624);
and U1996 (N_1996,N_1684,N_1736);
or U1997 (N_1997,N_1614,N_1708);
or U1998 (N_1998,N_1757,N_1733);
or U1999 (N_1999,N_1601,N_1685);
nand U2000 (N_2000,N_1910,N_1926);
nor U2001 (N_2001,N_1946,N_1955);
nand U2002 (N_2002,N_1824,N_1947);
nor U2003 (N_2003,N_1873,N_1945);
or U2004 (N_2004,N_1819,N_1999);
xnor U2005 (N_2005,N_1986,N_1997);
and U2006 (N_2006,N_1922,N_1932);
nand U2007 (N_2007,N_1982,N_1889);
or U2008 (N_2008,N_1826,N_1830);
nor U2009 (N_2009,N_1851,N_1940);
nand U2010 (N_2010,N_1992,N_1958);
and U2011 (N_2011,N_1886,N_1924);
nor U2012 (N_2012,N_1832,N_1879);
nand U2013 (N_2013,N_1857,N_1899);
nand U2014 (N_2014,N_1988,N_1833);
or U2015 (N_2015,N_1961,N_1934);
nand U2016 (N_2016,N_1964,N_1822);
nor U2017 (N_2017,N_1878,N_1952);
nand U2018 (N_2018,N_1845,N_1810);
and U2019 (N_2019,N_1925,N_1912);
nor U2020 (N_2020,N_1954,N_1908);
and U2021 (N_2021,N_1866,N_1990);
or U2022 (N_2022,N_1973,N_1820);
xnor U2023 (N_2023,N_1861,N_1981);
nand U2024 (N_2024,N_1842,N_1980);
and U2025 (N_2025,N_1882,N_1966);
or U2026 (N_2026,N_1829,N_1801);
nand U2027 (N_2027,N_1978,N_1813);
and U2028 (N_2028,N_1812,N_1840);
nor U2029 (N_2029,N_1859,N_1962);
nand U2030 (N_2030,N_1898,N_1894);
xnor U2031 (N_2031,N_1960,N_1855);
nor U2032 (N_2032,N_1809,N_1904);
and U2033 (N_2033,N_1849,N_1805);
nand U2034 (N_2034,N_1834,N_1807);
or U2035 (N_2035,N_1970,N_1967);
nor U2036 (N_2036,N_1837,N_1868);
nand U2037 (N_2037,N_1874,N_1974);
nand U2038 (N_2038,N_1883,N_1825);
xor U2039 (N_2039,N_1872,N_1880);
or U2040 (N_2040,N_1907,N_1891);
nor U2041 (N_2041,N_1987,N_1916);
or U2042 (N_2042,N_1817,N_1993);
and U2043 (N_2043,N_1839,N_1877);
nand U2044 (N_2044,N_1802,N_1864);
xnor U2045 (N_2045,N_1835,N_1911);
and U2046 (N_2046,N_1957,N_1887);
and U2047 (N_2047,N_1959,N_1863);
or U2048 (N_2048,N_1943,N_1989);
nand U2049 (N_2049,N_1804,N_1821);
and U2050 (N_2050,N_1928,N_1975);
and U2051 (N_2051,N_1923,N_1929);
or U2052 (N_2052,N_1838,N_1853);
or U2053 (N_2053,N_1930,N_1848);
and U2054 (N_2054,N_1843,N_1800);
and U2055 (N_2055,N_1884,N_1858);
nand U2056 (N_2056,N_1998,N_1870);
or U2057 (N_2057,N_1939,N_1875);
nand U2058 (N_2058,N_1921,N_1920);
nand U2059 (N_2059,N_1919,N_1950);
xor U2060 (N_2060,N_1915,N_1971);
nand U2061 (N_2061,N_1867,N_1996);
or U2062 (N_2062,N_1828,N_1948);
xor U2063 (N_2063,N_1977,N_1965);
or U2064 (N_2064,N_1953,N_1896);
nand U2065 (N_2065,N_1869,N_1936);
or U2066 (N_2066,N_1933,N_1914);
nand U2067 (N_2067,N_1900,N_1836);
or U2068 (N_2068,N_1856,N_1860);
nor U2069 (N_2069,N_1865,N_1902);
and U2070 (N_2070,N_1892,N_1942);
nor U2071 (N_2071,N_1979,N_1917);
or U2072 (N_2072,N_1803,N_1905);
nand U2073 (N_2073,N_1818,N_1888);
nor U2074 (N_2074,N_1956,N_1850);
nor U2075 (N_2075,N_1949,N_1854);
or U2076 (N_2076,N_1852,N_1984);
xor U2077 (N_2077,N_1806,N_1876);
nand U2078 (N_2078,N_1808,N_1951);
nand U2079 (N_2079,N_1871,N_1938);
or U2080 (N_2080,N_1969,N_1831);
nor U2081 (N_2081,N_1903,N_1963);
nand U2082 (N_2082,N_1895,N_1811);
and U2083 (N_2083,N_1816,N_1968);
and U2084 (N_2084,N_1944,N_1823);
xnor U2085 (N_2085,N_1881,N_1991);
nor U2086 (N_2086,N_1983,N_1994);
xor U2087 (N_2087,N_1901,N_1815);
and U2088 (N_2088,N_1847,N_1985);
and U2089 (N_2089,N_1918,N_1941);
nand U2090 (N_2090,N_1841,N_1893);
or U2091 (N_2091,N_1927,N_1885);
nor U2092 (N_2092,N_1897,N_1890);
nand U2093 (N_2093,N_1995,N_1935);
or U2094 (N_2094,N_1862,N_1937);
or U2095 (N_2095,N_1909,N_1972);
nand U2096 (N_2096,N_1814,N_1827);
nand U2097 (N_2097,N_1913,N_1844);
and U2098 (N_2098,N_1846,N_1976);
and U2099 (N_2099,N_1906,N_1931);
or U2100 (N_2100,N_1956,N_1885);
or U2101 (N_2101,N_1852,N_1938);
nand U2102 (N_2102,N_1982,N_1925);
and U2103 (N_2103,N_1976,N_1998);
and U2104 (N_2104,N_1854,N_1999);
xnor U2105 (N_2105,N_1878,N_1946);
and U2106 (N_2106,N_1980,N_1859);
and U2107 (N_2107,N_1819,N_1989);
and U2108 (N_2108,N_1976,N_1950);
nor U2109 (N_2109,N_1803,N_1832);
nand U2110 (N_2110,N_1892,N_1943);
nor U2111 (N_2111,N_1855,N_1822);
nor U2112 (N_2112,N_1811,N_1889);
nor U2113 (N_2113,N_1909,N_1921);
nor U2114 (N_2114,N_1948,N_1998);
nand U2115 (N_2115,N_1802,N_1806);
nand U2116 (N_2116,N_1933,N_1938);
nand U2117 (N_2117,N_1908,N_1838);
xor U2118 (N_2118,N_1958,N_1971);
nand U2119 (N_2119,N_1971,N_1881);
or U2120 (N_2120,N_1975,N_1823);
and U2121 (N_2121,N_1806,N_1917);
nand U2122 (N_2122,N_1934,N_1811);
nand U2123 (N_2123,N_1845,N_1916);
nand U2124 (N_2124,N_1964,N_1888);
or U2125 (N_2125,N_1882,N_1919);
nand U2126 (N_2126,N_1840,N_1940);
or U2127 (N_2127,N_1907,N_1952);
or U2128 (N_2128,N_1867,N_1809);
and U2129 (N_2129,N_1912,N_1988);
nor U2130 (N_2130,N_1866,N_1852);
or U2131 (N_2131,N_1852,N_1838);
nor U2132 (N_2132,N_1934,N_1815);
nand U2133 (N_2133,N_1848,N_1850);
or U2134 (N_2134,N_1960,N_1965);
nand U2135 (N_2135,N_1939,N_1883);
and U2136 (N_2136,N_1923,N_1903);
nor U2137 (N_2137,N_1859,N_1868);
or U2138 (N_2138,N_1925,N_1963);
and U2139 (N_2139,N_1974,N_1976);
and U2140 (N_2140,N_1900,N_1977);
nor U2141 (N_2141,N_1812,N_1829);
nand U2142 (N_2142,N_1956,N_1800);
and U2143 (N_2143,N_1999,N_1978);
and U2144 (N_2144,N_1870,N_1838);
and U2145 (N_2145,N_1852,N_1839);
nor U2146 (N_2146,N_1951,N_1911);
or U2147 (N_2147,N_1965,N_1819);
nand U2148 (N_2148,N_1831,N_1874);
nor U2149 (N_2149,N_1987,N_1802);
and U2150 (N_2150,N_1827,N_1854);
nand U2151 (N_2151,N_1825,N_1882);
or U2152 (N_2152,N_1948,N_1887);
nand U2153 (N_2153,N_1966,N_1876);
nand U2154 (N_2154,N_1956,N_1977);
nand U2155 (N_2155,N_1915,N_1977);
or U2156 (N_2156,N_1940,N_1981);
nor U2157 (N_2157,N_1830,N_1940);
nor U2158 (N_2158,N_1817,N_1896);
and U2159 (N_2159,N_1917,N_1805);
nor U2160 (N_2160,N_1988,N_1855);
xor U2161 (N_2161,N_1897,N_1836);
xor U2162 (N_2162,N_1940,N_1955);
and U2163 (N_2163,N_1917,N_1983);
nand U2164 (N_2164,N_1886,N_1997);
nor U2165 (N_2165,N_1816,N_1891);
or U2166 (N_2166,N_1821,N_1911);
or U2167 (N_2167,N_1940,N_1934);
nor U2168 (N_2168,N_1865,N_1810);
and U2169 (N_2169,N_1986,N_1879);
nor U2170 (N_2170,N_1873,N_1977);
nand U2171 (N_2171,N_1859,N_1902);
nor U2172 (N_2172,N_1981,N_1872);
nor U2173 (N_2173,N_1847,N_1895);
nor U2174 (N_2174,N_1943,N_1947);
and U2175 (N_2175,N_1827,N_1965);
xnor U2176 (N_2176,N_1807,N_1959);
nand U2177 (N_2177,N_1904,N_1846);
nand U2178 (N_2178,N_1831,N_1859);
nand U2179 (N_2179,N_1893,N_1952);
and U2180 (N_2180,N_1815,N_1971);
or U2181 (N_2181,N_1810,N_1944);
nor U2182 (N_2182,N_1871,N_1875);
and U2183 (N_2183,N_1879,N_1971);
nor U2184 (N_2184,N_1824,N_1856);
and U2185 (N_2185,N_1939,N_1843);
and U2186 (N_2186,N_1919,N_1842);
xnor U2187 (N_2187,N_1837,N_1908);
or U2188 (N_2188,N_1870,N_1949);
or U2189 (N_2189,N_1878,N_1965);
or U2190 (N_2190,N_1937,N_1986);
and U2191 (N_2191,N_1916,N_1908);
nor U2192 (N_2192,N_1936,N_1865);
and U2193 (N_2193,N_1987,N_1899);
xnor U2194 (N_2194,N_1867,N_1889);
nor U2195 (N_2195,N_1861,N_1894);
and U2196 (N_2196,N_1978,N_1835);
nor U2197 (N_2197,N_1962,N_1954);
nor U2198 (N_2198,N_1912,N_1856);
or U2199 (N_2199,N_1835,N_1876);
and U2200 (N_2200,N_2139,N_2194);
nor U2201 (N_2201,N_2089,N_2025);
and U2202 (N_2202,N_2122,N_2173);
xnor U2203 (N_2203,N_2027,N_2063);
nor U2204 (N_2204,N_2034,N_2151);
nand U2205 (N_2205,N_2073,N_2159);
and U2206 (N_2206,N_2044,N_2129);
and U2207 (N_2207,N_2060,N_2024);
nor U2208 (N_2208,N_2006,N_2142);
and U2209 (N_2209,N_2187,N_2178);
nor U2210 (N_2210,N_2056,N_2076);
nand U2211 (N_2211,N_2085,N_2175);
or U2212 (N_2212,N_2161,N_2118);
xor U2213 (N_2213,N_2057,N_2133);
nor U2214 (N_2214,N_2047,N_2052);
or U2215 (N_2215,N_2198,N_2048);
xor U2216 (N_2216,N_2032,N_2018);
or U2217 (N_2217,N_2120,N_2136);
nor U2218 (N_2218,N_2038,N_2112);
nand U2219 (N_2219,N_2177,N_2017);
xnor U2220 (N_2220,N_2072,N_2082);
nand U2221 (N_2221,N_2147,N_2163);
nand U2222 (N_2222,N_2043,N_2121);
nor U2223 (N_2223,N_2169,N_2108);
and U2224 (N_2224,N_2170,N_2003);
nand U2225 (N_2225,N_2126,N_2093);
nor U2226 (N_2226,N_2167,N_2095);
or U2227 (N_2227,N_2158,N_2176);
or U2228 (N_2228,N_2011,N_2004);
and U2229 (N_2229,N_2045,N_2081);
or U2230 (N_2230,N_2109,N_2131);
or U2231 (N_2231,N_2141,N_2197);
nor U2232 (N_2232,N_2116,N_2182);
and U2233 (N_2233,N_2171,N_2042);
nand U2234 (N_2234,N_2154,N_2155);
nor U2235 (N_2235,N_2101,N_2067);
or U2236 (N_2236,N_2033,N_2180);
xor U2237 (N_2237,N_2053,N_2021);
and U2238 (N_2238,N_2064,N_2168);
nand U2239 (N_2239,N_2022,N_2166);
and U2240 (N_2240,N_2041,N_2099);
or U2241 (N_2241,N_2137,N_2192);
nand U2242 (N_2242,N_2104,N_2014);
and U2243 (N_2243,N_2113,N_2146);
nand U2244 (N_2244,N_2068,N_2054);
and U2245 (N_2245,N_2156,N_2026);
nor U2246 (N_2246,N_2123,N_2020);
nor U2247 (N_2247,N_2111,N_2196);
and U2248 (N_2248,N_2102,N_2119);
nor U2249 (N_2249,N_2097,N_2075);
nor U2250 (N_2250,N_2181,N_2035);
nor U2251 (N_2251,N_2190,N_2199);
nor U2252 (N_2252,N_2023,N_2002);
nor U2253 (N_2253,N_2059,N_2144);
nand U2254 (N_2254,N_2110,N_2103);
and U2255 (N_2255,N_2050,N_2008);
or U2256 (N_2256,N_2174,N_2183);
nand U2257 (N_2257,N_2055,N_2028);
or U2258 (N_2258,N_2062,N_2149);
nor U2259 (N_2259,N_2090,N_2127);
xnor U2260 (N_2260,N_2077,N_2005);
xor U2261 (N_2261,N_2152,N_2193);
and U2262 (N_2262,N_2130,N_2049);
and U2263 (N_2263,N_2040,N_2009);
nand U2264 (N_2264,N_2153,N_2150);
nor U2265 (N_2265,N_2019,N_2036);
nand U2266 (N_2266,N_2013,N_2143);
nor U2267 (N_2267,N_2058,N_2069);
nor U2268 (N_2268,N_2189,N_2012);
nor U2269 (N_2269,N_2105,N_2071);
nor U2270 (N_2270,N_2132,N_2185);
nor U2271 (N_2271,N_2083,N_2046);
nand U2272 (N_2272,N_2065,N_2078);
nand U2273 (N_2273,N_2195,N_2179);
nand U2274 (N_2274,N_2117,N_2100);
nand U2275 (N_2275,N_2079,N_2066);
nand U2276 (N_2276,N_2070,N_2094);
or U2277 (N_2277,N_2162,N_2107);
or U2278 (N_2278,N_2114,N_2138);
nand U2279 (N_2279,N_2088,N_2039);
or U2280 (N_2280,N_2091,N_2031);
or U2281 (N_2281,N_2092,N_2080);
and U2282 (N_2282,N_2051,N_2087);
nor U2283 (N_2283,N_2184,N_2001);
or U2284 (N_2284,N_2188,N_2016);
or U2285 (N_2285,N_2164,N_2172);
nand U2286 (N_2286,N_2106,N_2128);
nor U2287 (N_2287,N_2096,N_2186);
or U2288 (N_2288,N_2115,N_2124);
xor U2289 (N_2289,N_2148,N_2140);
and U2290 (N_2290,N_2157,N_2145);
nand U2291 (N_2291,N_2061,N_2029);
nand U2292 (N_2292,N_2030,N_2125);
xnor U2293 (N_2293,N_2007,N_2165);
or U2294 (N_2294,N_2135,N_2000);
nand U2295 (N_2295,N_2134,N_2191);
nor U2296 (N_2296,N_2037,N_2098);
nor U2297 (N_2297,N_2010,N_2074);
nand U2298 (N_2298,N_2086,N_2084);
xnor U2299 (N_2299,N_2160,N_2015);
xnor U2300 (N_2300,N_2126,N_2014);
nand U2301 (N_2301,N_2118,N_2044);
nand U2302 (N_2302,N_2165,N_2120);
and U2303 (N_2303,N_2043,N_2143);
or U2304 (N_2304,N_2051,N_2160);
nand U2305 (N_2305,N_2149,N_2120);
and U2306 (N_2306,N_2006,N_2163);
nor U2307 (N_2307,N_2057,N_2022);
nor U2308 (N_2308,N_2073,N_2024);
or U2309 (N_2309,N_2024,N_2096);
and U2310 (N_2310,N_2191,N_2172);
nand U2311 (N_2311,N_2146,N_2167);
or U2312 (N_2312,N_2038,N_2110);
nand U2313 (N_2313,N_2058,N_2167);
nand U2314 (N_2314,N_2134,N_2118);
nand U2315 (N_2315,N_2160,N_2119);
or U2316 (N_2316,N_2044,N_2080);
and U2317 (N_2317,N_2178,N_2090);
and U2318 (N_2318,N_2039,N_2069);
or U2319 (N_2319,N_2128,N_2060);
nor U2320 (N_2320,N_2091,N_2076);
or U2321 (N_2321,N_2023,N_2176);
or U2322 (N_2322,N_2077,N_2034);
nor U2323 (N_2323,N_2036,N_2152);
nand U2324 (N_2324,N_2180,N_2041);
xnor U2325 (N_2325,N_2158,N_2076);
and U2326 (N_2326,N_2012,N_2114);
or U2327 (N_2327,N_2083,N_2017);
and U2328 (N_2328,N_2056,N_2020);
nor U2329 (N_2329,N_2141,N_2030);
or U2330 (N_2330,N_2063,N_2145);
xnor U2331 (N_2331,N_2099,N_2085);
nand U2332 (N_2332,N_2101,N_2002);
and U2333 (N_2333,N_2081,N_2160);
or U2334 (N_2334,N_2192,N_2123);
nor U2335 (N_2335,N_2089,N_2046);
xor U2336 (N_2336,N_2065,N_2075);
nand U2337 (N_2337,N_2089,N_2095);
nand U2338 (N_2338,N_2113,N_2086);
xnor U2339 (N_2339,N_2168,N_2076);
or U2340 (N_2340,N_2003,N_2156);
nand U2341 (N_2341,N_2195,N_2015);
nor U2342 (N_2342,N_2120,N_2037);
nor U2343 (N_2343,N_2031,N_2123);
and U2344 (N_2344,N_2025,N_2127);
and U2345 (N_2345,N_2117,N_2038);
and U2346 (N_2346,N_2122,N_2145);
or U2347 (N_2347,N_2011,N_2140);
and U2348 (N_2348,N_2195,N_2055);
nor U2349 (N_2349,N_2098,N_2001);
and U2350 (N_2350,N_2171,N_2166);
or U2351 (N_2351,N_2067,N_2111);
nand U2352 (N_2352,N_2016,N_2137);
nand U2353 (N_2353,N_2154,N_2099);
nand U2354 (N_2354,N_2123,N_2147);
or U2355 (N_2355,N_2168,N_2126);
xor U2356 (N_2356,N_2001,N_2129);
and U2357 (N_2357,N_2052,N_2080);
and U2358 (N_2358,N_2074,N_2085);
nand U2359 (N_2359,N_2181,N_2152);
nor U2360 (N_2360,N_2017,N_2060);
or U2361 (N_2361,N_2066,N_2014);
or U2362 (N_2362,N_2005,N_2093);
nor U2363 (N_2363,N_2109,N_2051);
or U2364 (N_2364,N_2103,N_2035);
nor U2365 (N_2365,N_2015,N_2106);
and U2366 (N_2366,N_2133,N_2131);
nor U2367 (N_2367,N_2186,N_2194);
and U2368 (N_2368,N_2172,N_2002);
nand U2369 (N_2369,N_2099,N_2059);
nor U2370 (N_2370,N_2048,N_2053);
nor U2371 (N_2371,N_2197,N_2111);
nand U2372 (N_2372,N_2093,N_2083);
nor U2373 (N_2373,N_2027,N_2156);
and U2374 (N_2374,N_2182,N_2079);
nor U2375 (N_2375,N_2126,N_2146);
xnor U2376 (N_2376,N_2011,N_2072);
and U2377 (N_2377,N_2058,N_2107);
and U2378 (N_2378,N_2013,N_2198);
xnor U2379 (N_2379,N_2176,N_2178);
nand U2380 (N_2380,N_2099,N_2172);
nor U2381 (N_2381,N_2017,N_2184);
or U2382 (N_2382,N_2022,N_2134);
or U2383 (N_2383,N_2093,N_2047);
xnor U2384 (N_2384,N_2000,N_2184);
or U2385 (N_2385,N_2163,N_2016);
and U2386 (N_2386,N_2136,N_2105);
nor U2387 (N_2387,N_2196,N_2138);
nand U2388 (N_2388,N_2133,N_2013);
nor U2389 (N_2389,N_2148,N_2052);
nand U2390 (N_2390,N_2181,N_2112);
nand U2391 (N_2391,N_2087,N_2187);
and U2392 (N_2392,N_2198,N_2130);
or U2393 (N_2393,N_2195,N_2005);
or U2394 (N_2394,N_2172,N_2032);
nor U2395 (N_2395,N_2101,N_2001);
or U2396 (N_2396,N_2002,N_2069);
and U2397 (N_2397,N_2038,N_2068);
and U2398 (N_2398,N_2183,N_2041);
or U2399 (N_2399,N_2165,N_2057);
nand U2400 (N_2400,N_2283,N_2309);
nor U2401 (N_2401,N_2333,N_2384);
nand U2402 (N_2402,N_2232,N_2281);
nand U2403 (N_2403,N_2397,N_2342);
nand U2404 (N_2404,N_2340,N_2211);
or U2405 (N_2405,N_2396,N_2362);
and U2406 (N_2406,N_2318,N_2288);
and U2407 (N_2407,N_2261,N_2260);
nor U2408 (N_2408,N_2364,N_2291);
nand U2409 (N_2409,N_2382,N_2371);
and U2410 (N_2410,N_2373,N_2344);
xnor U2411 (N_2411,N_2392,N_2264);
nor U2412 (N_2412,N_2311,N_2323);
nor U2413 (N_2413,N_2259,N_2295);
xnor U2414 (N_2414,N_2269,N_2247);
nor U2415 (N_2415,N_2312,N_2315);
nand U2416 (N_2416,N_2374,N_2367);
or U2417 (N_2417,N_2271,N_2262);
nor U2418 (N_2418,N_2387,N_2265);
nand U2419 (N_2419,N_2248,N_2388);
and U2420 (N_2420,N_2357,N_2368);
nand U2421 (N_2421,N_2365,N_2219);
nand U2422 (N_2422,N_2251,N_2274);
nand U2423 (N_2423,N_2363,N_2358);
xor U2424 (N_2424,N_2266,N_2205);
and U2425 (N_2425,N_2341,N_2328);
and U2426 (N_2426,N_2221,N_2237);
and U2427 (N_2427,N_2238,N_2338);
nor U2428 (N_2428,N_2310,N_2393);
nor U2429 (N_2429,N_2343,N_2245);
or U2430 (N_2430,N_2216,N_2249);
and U2431 (N_2431,N_2280,N_2337);
and U2432 (N_2432,N_2324,N_2330);
nor U2433 (N_2433,N_2297,N_2256);
and U2434 (N_2434,N_2218,N_2376);
nor U2435 (N_2435,N_2317,N_2234);
nand U2436 (N_2436,N_2307,N_2300);
or U2437 (N_2437,N_2206,N_2361);
or U2438 (N_2438,N_2395,N_2278);
nand U2439 (N_2439,N_2349,N_2226);
nand U2440 (N_2440,N_2224,N_2285);
or U2441 (N_2441,N_2352,N_2359);
nand U2442 (N_2442,N_2389,N_2293);
nand U2443 (N_2443,N_2214,N_2209);
nand U2444 (N_2444,N_2294,N_2306);
nand U2445 (N_2445,N_2304,N_2277);
or U2446 (N_2446,N_2217,N_2326);
or U2447 (N_2447,N_2284,N_2275);
and U2448 (N_2448,N_2331,N_2203);
or U2449 (N_2449,N_2231,N_2287);
nand U2450 (N_2450,N_2336,N_2270);
and U2451 (N_2451,N_2394,N_2204);
or U2452 (N_2452,N_2235,N_2348);
nand U2453 (N_2453,N_2222,N_2273);
nor U2454 (N_2454,N_2268,N_2254);
xnor U2455 (N_2455,N_2350,N_2355);
nand U2456 (N_2456,N_2215,N_2213);
and U2457 (N_2457,N_2244,N_2228);
nor U2458 (N_2458,N_2339,N_2366);
nor U2459 (N_2459,N_2313,N_2332);
nor U2460 (N_2460,N_2298,N_2282);
nor U2461 (N_2461,N_2272,N_2267);
nor U2462 (N_2462,N_2370,N_2289);
or U2463 (N_2463,N_2223,N_2225);
xor U2464 (N_2464,N_2386,N_2303);
xor U2465 (N_2465,N_2353,N_2200);
or U2466 (N_2466,N_2286,N_2372);
or U2467 (N_2467,N_2202,N_2229);
nor U2468 (N_2468,N_2210,N_2314);
xor U2469 (N_2469,N_2322,N_2241);
nand U2470 (N_2470,N_2335,N_2279);
nand U2471 (N_2471,N_2201,N_2346);
and U2472 (N_2472,N_2255,N_2383);
nand U2473 (N_2473,N_2236,N_2220);
nand U2474 (N_2474,N_2212,N_2239);
or U2475 (N_2475,N_2246,N_2305);
nor U2476 (N_2476,N_2399,N_2351);
nand U2477 (N_2477,N_2381,N_2321);
xnor U2478 (N_2478,N_2390,N_2380);
nand U2479 (N_2479,N_2360,N_2252);
nor U2480 (N_2480,N_2258,N_2378);
and U2481 (N_2481,N_2243,N_2230);
or U2482 (N_2482,N_2233,N_2379);
nand U2483 (N_2483,N_2377,N_2325);
or U2484 (N_2484,N_2302,N_2290);
xnor U2485 (N_2485,N_2354,N_2276);
nand U2486 (N_2486,N_2227,N_2345);
and U2487 (N_2487,N_2250,N_2316);
or U2488 (N_2488,N_2253,N_2320);
and U2489 (N_2489,N_2356,N_2208);
nand U2490 (N_2490,N_2369,N_2329);
nor U2491 (N_2491,N_2347,N_2391);
nor U2492 (N_2492,N_2299,N_2385);
or U2493 (N_2493,N_2308,N_2334);
nand U2494 (N_2494,N_2257,N_2375);
nand U2495 (N_2495,N_2292,N_2398);
nor U2496 (N_2496,N_2319,N_2296);
or U2497 (N_2497,N_2207,N_2327);
xnor U2498 (N_2498,N_2263,N_2242);
xor U2499 (N_2499,N_2240,N_2301);
xor U2500 (N_2500,N_2322,N_2311);
nor U2501 (N_2501,N_2319,N_2212);
nor U2502 (N_2502,N_2363,N_2308);
nand U2503 (N_2503,N_2311,N_2364);
and U2504 (N_2504,N_2383,N_2245);
or U2505 (N_2505,N_2332,N_2317);
and U2506 (N_2506,N_2235,N_2247);
or U2507 (N_2507,N_2375,N_2283);
nand U2508 (N_2508,N_2201,N_2312);
nor U2509 (N_2509,N_2253,N_2263);
or U2510 (N_2510,N_2200,N_2397);
or U2511 (N_2511,N_2278,N_2307);
and U2512 (N_2512,N_2369,N_2367);
or U2513 (N_2513,N_2270,N_2322);
and U2514 (N_2514,N_2381,N_2208);
nor U2515 (N_2515,N_2303,N_2308);
nor U2516 (N_2516,N_2313,N_2235);
nand U2517 (N_2517,N_2357,N_2353);
and U2518 (N_2518,N_2392,N_2282);
and U2519 (N_2519,N_2318,N_2314);
or U2520 (N_2520,N_2228,N_2393);
and U2521 (N_2521,N_2292,N_2351);
and U2522 (N_2522,N_2285,N_2373);
and U2523 (N_2523,N_2348,N_2221);
and U2524 (N_2524,N_2224,N_2376);
and U2525 (N_2525,N_2397,N_2396);
nand U2526 (N_2526,N_2258,N_2240);
nor U2527 (N_2527,N_2276,N_2272);
and U2528 (N_2528,N_2357,N_2376);
or U2529 (N_2529,N_2314,N_2396);
nor U2530 (N_2530,N_2339,N_2227);
nand U2531 (N_2531,N_2276,N_2348);
and U2532 (N_2532,N_2367,N_2395);
nor U2533 (N_2533,N_2365,N_2341);
and U2534 (N_2534,N_2395,N_2244);
nand U2535 (N_2535,N_2234,N_2262);
nand U2536 (N_2536,N_2308,N_2274);
or U2537 (N_2537,N_2272,N_2379);
nor U2538 (N_2538,N_2221,N_2336);
nand U2539 (N_2539,N_2220,N_2361);
xor U2540 (N_2540,N_2268,N_2235);
nor U2541 (N_2541,N_2305,N_2243);
and U2542 (N_2542,N_2317,N_2249);
and U2543 (N_2543,N_2375,N_2390);
nor U2544 (N_2544,N_2311,N_2388);
nand U2545 (N_2545,N_2379,N_2257);
nor U2546 (N_2546,N_2324,N_2200);
and U2547 (N_2547,N_2271,N_2322);
and U2548 (N_2548,N_2350,N_2397);
nor U2549 (N_2549,N_2266,N_2373);
or U2550 (N_2550,N_2319,N_2308);
nand U2551 (N_2551,N_2210,N_2206);
nor U2552 (N_2552,N_2352,N_2309);
nor U2553 (N_2553,N_2265,N_2333);
or U2554 (N_2554,N_2395,N_2327);
nor U2555 (N_2555,N_2373,N_2361);
nor U2556 (N_2556,N_2204,N_2343);
nor U2557 (N_2557,N_2265,N_2345);
and U2558 (N_2558,N_2359,N_2205);
nand U2559 (N_2559,N_2360,N_2385);
nand U2560 (N_2560,N_2265,N_2381);
xnor U2561 (N_2561,N_2360,N_2287);
xnor U2562 (N_2562,N_2338,N_2321);
nand U2563 (N_2563,N_2361,N_2269);
and U2564 (N_2564,N_2279,N_2291);
nand U2565 (N_2565,N_2248,N_2241);
nand U2566 (N_2566,N_2343,N_2354);
xnor U2567 (N_2567,N_2397,N_2331);
or U2568 (N_2568,N_2378,N_2208);
nor U2569 (N_2569,N_2316,N_2252);
and U2570 (N_2570,N_2268,N_2351);
and U2571 (N_2571,N_2281,N_2392);
or U2572 (N_2572,N_2231,N_2212);
and U2573 (N_2573,N_2363,N_2313);
and U2574 (N_2574,N_2274,N_2385);
or U2575 (N_2575,N_2352,N_2362);
or U2576 (N_2576,N_2268,N_2373);
nand U2577 (N_2577,N_2283,N_2254);
nor U2578 (N_2578,N_2224,N_2239);
xnor U2579 (N_2579,N_2264,N_2304);
or U2580 (N_2580,N_2336,N_2340);
nor U2581 (N_2581,N_2382,N_2297);
nor U2582 (N_2582,N_2306,N_2223);
xor U2583 (N_2583,N_2358,N_2289);
nand U2584 (N_2584,N_2318,N_2273);
or U2585 (N_2585,N_2304,N_2379);
and U2586 (N_2586,N_2340,N_2380);
nand U2587 (N_2587,N_2209,N_2262);
xnor U2588 (N_2588,N_2211,N_2247);
and U2589 (N_2589,N_2315,N_2251);
and U2590 (N_2590,N_2330,N_2294);
or U2591 (N_2591,N_2200,N_2310);
nand U2592 (N_2592,N_2211,N_2351);
nand U2593 (N_2593,N_2382,N_2201);
nand U2594 (N_2594,N_2201,N_2217);
nor U2595 (N_2595,N_2334,N_2342);
or U2596 (N_2596,N_2397,N_2223);
or U2597 (N_2597,N_2285,N_2303);
nor U2598 (N_2598,N_2269,N_2305);
and U2599 (N_2599,N_2253,N_2377);
and U2600 (N_2600,N_2519,N_2411);
nand U2601 (N_2601,N_2484,N_2569);
nor U2602 (N_2602,N_2420,N_2444);
or U2603 (N_2603,N_2560,N_2403);
and U2604 (N_2604,N_2416,N_2417);
nor U2605 (N_2605,N_2460,N_2504);
nor U2606 (N_2606,N_2478,N_2424);
nand U2607 (N_2607,N_2529,N_2441);
and U2608 (N_2608,N_2584,N_2563);
or U2609 (N_2609,N_2485,N_2454);
and U2610 (N_2610,N_2525,N_2581);
nor U2611 (N_2611,N_2461,N_2443);
and U2612 (N_2612,N_2524,N_2538);
nand U2613 (N_2613,N_2566,N_2542);
nand U2614 (N_2614,N_2415,N_2430);
nor U2615 (N_2615,N_2533,N_2477);
or U2616 (N_2616,N_2404,N_2541);
nor U2617 (N_2617,N_2448,N_2419);
nor U2618 (N_2618,N_2570,N_2435);
nor U2619 (N_2619,N_2423,N_2549);
and U2620 (N_2620,N_2599,N_2571);
nor U2621 (N_2621,N_2580,N_2465);
xnor U2622 (N_2622,N_2530,N_2586);
nand U2623 (N_2623,N_2493,N_2589);
nand U2624 (N_2624,N_2507,N_2467);
or U2625 (N_2625,N_2442,N_2528);
nand U2626 (N_2626,N_2418,N_2475);
or U2627 (N_2627,N_2592,N_2481);
or U2628 (N_2628,N_2596,N_2518);
and U2629 (N_2629,N_2591,N_2577);
or U2630 (N_2630,N_2585,N_2550);
nand U2631 (N_2631,N_2429,N_2492);
xor U2632 (N_2632,N_2401,N_2597);
or U2633 (N_2633,N_2576,N_2422);
or U2634 (N_2634,N_2554,N_2489);
or U2635 (N_2635,N_2520,N_2509);
nand U2636 (N_2636,N_2474,N_2548);
nor U2637 (N_2637,N_2498,N_2438);
nor U2638 (N_2638,N_2532,N_2428);
or U2639 (N_2639,N_2426,N_2412);
nor U2640 (N_2640,N_2501,N_2436);
nand U2641 (N_2641,N_2425,N_2526);
nand U2642 (N_2642,N_2405,N_2557);
and U2643 (N_2643,N_2497,N_2480);
and U2644 (N_2644,N_2536,N_2495);
xor U2645 (N_2645,N_2567,N_2445);
or U2646 (N_2646,N_2552,N_2470);
or U2647 (N_2647,N_2510,N_2464);
nor U2648 (N_2648,N_2521,N_2402);
and U2649 (N_2649,N_2453,N_2583);
nor U2650 (N_2650,N_2506,N_2468);
or U2651 (N_2651,N_2575,N_2434);
nand U2652 (N_2652,N_2499,N_2527);
nor U2653 (N_2653,N_2496,N_2494);
or U2654 (N_2654,N_2523,N_2451);
nand U2655 (N_2655,N_2573,N_2457);
or U2656 (N_2656,N_2503,N_2466);
nand U2657 (N_2657,N_2482,N_2512);
or U2658 (N_2658,N_2439,N_2410);
or U2659 (N_2659,N_2508,N_2488);
nand U2660 (N_2660,N_2455,N_2514);
or U2661 (N_2661,N_2409,N_2537);
and U2662 (N_2662,N_2561,N_2515);
nor U2663 (N_2663,N_2491,N_2421);
and U2664 (N_2664,N_2505,N_2551);
nand U2665 (N_2665,N_2593,N_2598);
nor U2666 (N_2666,N_2547,N_2456);
and U2667 (N_2667,N_2534,N_2446);
nor U2668 (N_2668,N_2539,N_2463);
nor U2669 (N_2669,N_2502,N_2559);
nand U2670 (N_2670,N_2458,N_2452);
and U2671 (N_2671,N_2433,N_2522);
nand U2672 (N_2672,N_2511,N_2572);
and U2673 (N_2673,N_2486,N_2431);
or U2674 (N_2674,N_2535,N_2587);
nand U2675 (N_2675,N_2483,N_2479);
and U2676 (N_2676,N_2574,N_2565);
or U2677 (N_2677,N_2544,N_2449);
nand U2678 (N_2678,N_2517,N_2447);
or U2679 (N_2679,N_2462,N_2490);
nand U2680 (N_2680,N_2595,N_2414);
or U2681 (N_2681,N_2546,N_2437);
and U2682 (N_2682,N_2471,N_2487);
nand U2683 (N_2683,N_2568,N_2553);
nor U2684 (N_2684,N_2588,N_2558);
nor U2685 (N_2685,N_2579,N_2543);
nand U2686 (N_2686,N_2594,N_2516);
nor U2687 (N_2687,N_2432,N_2555);
or U2688 (N_2688,N_2562,N_2540);
xor U2689 (N_2689,N_2564,N_2413);
or U2690 (N_2690,N_2582,N_2473);
and U2691 (N_2691,N_2531,N_2513);
nand U2692 (N_2692,N_2556,N_2406);
nand U2693 (N_2693,N_2476,N_2408);
and U2694 (N_2694,N_2400,N_2459);
and U2695 (N_2695,N_2450,N_2427);
nand U2696 (N_2696,N_2407,N_2472);
nor U2697 (N_2697,N_2500,N_2578);
or U2698 (N_2698,N_2545,N_2469);
and U2699 (N_2699,N_2590,N_2440);
and U2700 (N_2700,N_2521,N_2554);
nor U2701 (N_2701,N_2578,N_2457);
xnor U2702 (N_2702,N_2560,N_2577);
or U2703 (N_2703,N_2541,N_2594);
and U2704 (N_2704,N_2554,N_2459);
xnor U2705 (N_2705,N_2430,N_2478);
and U2706 (N_2706,N_2574,N_2573);
nor U2707 (N_2707,N_2464,N_2433);
nor U2708 (N_2708,N_2546,N_2463);
nor U2709 (N_2709,N_2582,N_2497);
xor U2710 (N_2710,N_2519,N_2402);
or U2711 (N_2711,N_2548,N_2450);
nand U2712 (N_2712,N_2508,N_2466);
nand U2713 (N_2713,N_2547,N_2495);
or U2714 (N_2714,N_2517,N_2560);
nor U2715 (N_2715,N_2589,N_2547);
or U2716 (N_2716,N_2421,N_2479);
nor U2717 (N_2717,N_2422,N_2556);
nor U2718 (N_2718,N_2489,N_2421);
xnor U2719 (N_2719,N_2432,N_2417);
xor U2720 (N_2720,N_2436,N_2595);
or U2721 (N_2721,N_2443,N_2467);
nor U2722 (N_2722,N_2594,N_2442);
nand U2723 (N_2723,N_2414,N_2409);
nand U2724 (N_2724,N_2452,N_2560);
or U2725 (N_2725,N_2435,N_2415);
and U2726 (N_2726,N_2468,N_2576);
nand U2727 (N_2727,N_2532,N_2553);
nand U2728 (N_2728,N_2551,N_2502);
or U2729 (N_2729,N_2533,N_2579);
and U2730 (N_2730,N_2506,N_2419);
xnor U2731 (N_2731,N_2545,N_2589);
or U2732 (N_2732,N_2485,N_2549);
or U2733 (N_2733,N_2478,N_2440);
and U2734 (N_2734,N_2498,N_2570);
nor U2735 (N_2735,N_2542,N_2562);
nor U2736 (N_2736,N_2574,N_2521);
nor U2737 (N_2737,N_2497,N_2413);
nand U2738 (N_2738,N_2569,N_2506);
and U2739 (N_2739,N_2518,N_2536);
or U2740 (N_2740,N_2536,N_2421);
nand U2741 (N_2741,N_2535,N_2538);
nand U2742 (N_2742,N_2562,N_2524);
nor U2743 (N_2743,N_2462,N_2494);
nand U2744 (N_2744,N_2411,N_2482);
xor U2745 (N_2745,N_2495,N_2573);
or U2746 (N_2746,N_2508,N_2478);
nand U2747 (N_2747,N_2516,N_2546);
xnor U2748 (N_2748,N_2450,N_2558);
or U2749 (N_2749,N_2527,N_2579);
and U2750 (N_2750,N_2586,N_2589);
nor U2751 (N_2751,N_2510,N_2591);
xnor U2752 (N_2752,N_2419,N_2433);
nand U2753 (N_2753,N_2577,N_2575);
or U2754 (N_2754,N_2412,N_2575);
or U2755 (N_2755,N_2401,N_2563);
nand U2756 (N_2756,N_2466,N_2481);
and U2757 (N_2757,N_2547,N_2446);
or U2758 (N_2758,N_2463,N_2510);
and U2759 (N_2759,N_2528,N_2596);
or U2760 (N_2760,N_2466,N_2446);
nand U2761 (N_2761,N_2562,N_2412);
nor U2762 (N_2762,N_2531,N_2440);
and U2763 (N_2763,N_2585,N_2464);
nand U2764 (N_2764,N_2412,N_2431);
nand U2765 (N_2765,N_2523,N_2478);
and U2766 (N_2766,N_2501,N_2522);
and U2767 (N_2767,N_2415,N_2481);
nor U2768 (N_2768,N_2426,N_2591);
nor U2769 (N_2769,N_2569,N_2406);
and U2770 (N_2770,N_2418,N_2517);
nor U2771 (N_2771,N_2511,N_2544);
nand U2772 (N_2772,N_2490,N_2400);
nor U2773 (N_2773,N_2521,N_2481);
or U2774 (N_2774,N_2510,N_2580);
and U2775 (N_2775,N_2551,N_2521);
nor U2776 (N_2776,N_2541,N_2552);
and U2777 (N_2777,N_2555,N_2428);
or U2778 (N_2778,N_2584,N_2555);
nand U2779 (N_2779,N_2509,N_2510);
and U2780 (N_2780,N_2489,N_2474);
nand U2781 (N_2781,N_2494,N_2457);
or U2782 (N_2782,N_2450,N_2547);
and U2783 (N_2783,N_2453,N_2472);
nor U2784 (N_2784,N_2489,N_2452);
nand U2785 (N_2785,N_2593,N_2471);
nor U2786 (N_2786,N_2469,N_2461);
and U2787 (N_2787,N_2592,N_2447);
or U2788 (N_2788,N_2408,N_2422);
nand U2789 (N_2789,N_2599,N_2414);
nor U2790 (N_2790,N_2548,N_2549);
nor U2791 (N_2791,N_2546,N_2432);
or U2792 (N_2792,N_2589,N_2417);
nand U2793 (N_2793,N_2593,N_2457);
nand U2794 (N_2794,N_2489,N_2504);
or U2795 (N_2795,N_2576,N_2535);
xnor U2796 (N_2796,N_2439,N_2573);
and U2797 (N_2797,N_2531,N_2426);
nand U2798 (N_2798,N_2484,N_2583);
and U2799 (N_2799,N_2514,N_2446);
nand U2800 (N_2800,N_2778,N_2648);
nand U2801 (N_2801,N_2767,N_2738);
or U2802 (N_2802,N_2706,N_2600);
nor U2803 (N_2803,N_2664,N_2676);
or U2804 (N_2804,N_2724,N_2729);
nor U2805 (N_2805,N_2726,N_2709);
nand U2806 (N_2806,N_2675,N_2783);
or U2807 (N_2807,N_2785,N_2772);
nor U2808 (N_2808,N_2768,N_2680);
nor U2809 (N_2809,N_2736,N_2735);
xor U2810 (N_2810,N_2687,N_2752);
and U2811 (N_2811,N_2635,N_2702);
xnor U2812 (N_2812,N_2793,N_2650);
nand U2813 (N_2813,N_2669,N_2603);
nor U2814 (N_2814,N_2712,N_2643);
nor U2815 (N_2815,N_2660,N_2761);
nor U2816 (N_2816,N_2796,N_2705);
nor U2817 (N_2817,N_2758,N_2777);
nor U2818 (N_2818,N_2682,N_2641);
nand U2819 (N_2819,N_2638,N_2794);
or U2820 (N_2820,N_2658,N_2618);
and U2821 (N_2821,N_2751,N_2708);
nor U2822 (N_2822,N_2710,N_2619);
and U2823 (N_2823,N_2734,N_2616);
or U2824 (N_2824,N_2779,N_2757);
or U2825 (N_2825,N_2646,N_2681);
and U2826 (N_2826,N_2694,N_2728);
nand U2827 (N_2827,N_2717,N_2642);
and U2828 (N_2828,N_2713,N_2606);
nand U2829 (N_2829,N_2731,N_2602);
and U2830 (N_2830,N_2659,N_2652);
and U2831 (N_2831,N_2756,N_2698);
and U2832 (N_2832,N_2733,N_2656);
nand U2833 (N_2833,N_2673,N_2700);
nand U2834 (N_2834,N_2649,N_2748);
and U2835 (N_2835,N_2770,N_2604);
or U2836 (N_2836,N_2701,N_2787);
nand U2837 (N_2837,N_2674,N_2615);
or U2838 (N_2838,N_2759,N_2760);
nor U2839 (N_2839,N_2684,N_2666);
nor U2840 (N_2840,N_2750,N_2632);
xnor U2841 (N_2841,N_2747,N_2620);
or U2842 (N_2842,N_2639,N_2753);
nor U2843 (N_2843,N_2695,N_2626);
nor U2844 (N_2844,N_2628,N_2630);
nor U2845 (N_2845,N_2697,N_2730);
nand U2846 (N_2846,N_2611,N_2746);
and U2847 (N_2847,N_2634,N_2773);
or U2848 (N_2848,N_2786,N_2671);
or U2849 (N_2849,N_2774,N_2790);
and U2850 (N_2850,N_2755,N_2633);
and U2851 (N_2851,N_2686,N_2601);
or U2852 (N_2852,N_2624,N_2792);
or U2853 (N_2853,N_2683,N_2692);
nor U2854 (N_2854,N_2764,N_2754);
nor U2855 (N_2855,N_2678,N_2769);
nor U2856 (N_2856,N_2645,N_2742);
nor U2857 (N_2857,N_2791,N_2623);
nand U2858 (N_2858,N_2690,N_2627);
and U2859 (N_2859,N_2636,N_2667);
xor U2860 (N_2860,N_2795,N_2799);
xnor U2861 (N_2861,N_2703,N_2727);
nor U2862 (N_2862,N_2797,N_2661);
or U2863 (N_2863,N_2655,N_2637);
or U2864 (N_2864,N_2607,N_2605);
nand U2865 (N_2865,N_2718,N_2775);
nand U2866 (N_2866,N_2691,N_2631);
nor U2867 (N_2867,N_2610,N_2771);
nor U2868 (N_2868,N_2629,N_2621);
nand U2869 (N_2869,N_2739,N_2654);
nand U2870 (N_2870,N_2725,N_2720);
and U2871 (N_2871,N_2716,N_2653);
or U2872 (N_2872,N_2640,N_2613);
xnor U2873 (N_2873,N_2665,N_2696);
nor U2874 (N_2874,N_2693,N_2685);
or U2875 (N_2875,N_2744,N_2788);
nand U2876 (N_2876,N_2765,N_2644);
or U2877 (N_2877,N_2688,N_2781);
xnor U2878 (N_2878,N_2743,N_2776);
nor U2879 (N_2879,N_2740,N_2657);
and U2880 (N_2880,N_2798,N_2714);
nand U2881 (N_2881,N_2719,N_2647);
or U2882 (N_2882,N_2651,N_2745);
nand U2883 (N_2883,N_2715,N_2612);
and U2884 (N_2884,N_2784,N_2625);
nor U2885 (N_2885,N_2677,N_2608);
or U2886 (N_2886,N_2668,N_2609);
nor U2887 (N_2887,N_2617,N_2782);
and U2888 (N_2888,N_2689,N_2780);
and U2889 (N_2889,N_2672,N_2679);
nand U2890 (N_2890,N_2723,N_2663);
and U2891 (N_2891,N_2707,N_2741);
nor U2892 (N_2892,N_2670,N_2622);
nand U2893 (N_2893,N_2614,N_2732);
xnor U2894 (N_2894,N_2763,N_2766);
and U2895 (N_2895,N_2722,N_2704);
nand U2896 (N_2896,N_2762,N_2789);
or U2897 (N_2897,N_2721,N_2699);
nand U2898 (N_2898,N_2737,N_2749);
nor U2899 (N_2899,N_2662,N_2711);
nor U2900 (N_2900,N_2610,N_2699);
and U2901 (N_2901,N_2672,N_2782);
or U2902 (N_2902,N_2693,N_2710);
and U2903 (N_2903,N_2624,N_2784);
and U2904 (N_2904,N_2789,N_2697);
nor U2905 (N_2905,N_2602,N_2748);
or U2906 (N_2906,N_2651,N_2778);
nor U2907 (N_2907,N_2726,N_2725);
xnor U2908 (N_2908,N_2642,N_2633);
nand U2909 (N_2909,N_2660,N_2632);
nor U2910 (N_2910,N_2604,N_2715);
nor U2911 (N_2911,N_2714,N_2729);
or U2912 (N_2912,N_2774,N_2727);
or U2913 (N_2913,N_2761,N_2690);
nor U2914 (N_2914,N_2706,N_2734);
and U2915 (N_2915,N_2726,N_2702);
and U2916 (N_2916,N_2763,N_2728);
nand U2917 (N_2917,N_2791,N_2787);
nand U2918 (N_2918,N_2637,N_2794);
xnor U2919 (N_2919,N_2605,N_2749);
nand U2920 (N_2920,N_2760,N_2719);
nand U2921 (N_2921,N_2774,N_2791);
nor U2922 (N_2922,N_2608,N_2655);
or U2923 (N_2923,N_2685,N_2716);
nor U2924 (N_2924,N_2733,N_2718);
nand U2925 (N_2925,N_2651,N_2672);
nor U2926 (N_2926,N_2634,N_2781);
and U2927 (N_2927,N_2752,N_2650);
nor U2928 (N_2928,N_2757,N_2773);
or U2929 (N_2929,N_2642,N_2791);
or U2930 (N_2930,N_2763,N_2778);
and U2931 (N_2931,N_2742,N_2747);
nor U2932 (N_2932,N_2761,N_2680);
nand U2933 (N_2933,N_2718,N_2711);
or U2934 (N_2934,N_2669,N_2768);
or U2935 (N_2935,N_2710,N_2659);
xnor U2936 (N_2936,N_2623,N_2733);
or U2937 (N_2937,N_2639,N_2730);
nand U2938 (N_2938,N_2694,N_2657);
and U2939 (N_2939,N_2682,N_2757);
and U2940 (N_2940,N_2697,N_2644);
or U2941 (N_2941,N_2702,N_2742);
nand U2942 (N_2942,N_2796,N_2626);
and U2943 (N_2943,N_2758,N_2642);
nor U2944 (N_2944,N_2759,N_2695);
xor U2945 (N_2945,N_2751,N_2741);
nand U2946 (N_2946,N_2601,N_2732);
or U2947 (N_2947,N_2762,N_2711);
nand U2948 (N_2948,N_2659,N_2668);
or U2949 (N_2949,N_2627,N_2783);
or U2950 (N_2950,N_2721,N_2612);
xor U2951 (N_2951,N_2789,N_2613);
and U2952 (N_2952,N_2606,N_2681);
nor U2953 (N_2953,N_2766,N_2685);
or U2954 (N_2954,N_2624,N_2740);
and U2955 (N_2955,N_2797,N_2731);
and U2956 (N_2956,N_2656,N_2771);
and U2957 (N_2957,N_2780,N_2657);
and U2958 (N_2958,N_2761,N_2644);
nand U2959 (N_2959,N_2623,N_2650);
nand U2960 (N_2960,N_2725,N_2650);
and U2961 (N_2961,N_2777,N_2681);
or U2962 (N_2962,N_2698,N_2630);
and U2963 (N_2963,N_2608,N_2741);
and U2964 (N_2964,N_2667,N_2755);
nor U2965 (N_2965,N_2667,N_2768);
nand U2966 (N_2966,N_2627,N_2619);
or U2967 (N_2967,N_2747,N_2762);
nor U2968 (N_2968,N_2740,N_2794);
or U2969 (N_2969,N_2654,N_2642);
and U2970 (N_2970,N_2703,N_2649);
nand U2971 (N_2971,N_2625,N_2743);
and U2972 (N_2972,N_2699,N_2684);
and U2973 (N_2973,N_2620,N_2680);
nand U2974 (N_2974,N_2618,N_2613);
and U2975 (N_2975,N_2708,N_2697);
or U2976 (N_2976,N_2683,N_2785);
or U2977 (N_2977,N_2748,N_2705);
and U2978 (N_2978,N_2705,N_2755);
and U2979 (N_2979,N_2734,N_2778);
nand U2980 (N_2980,N_2754,N_2638);
nand U2981 (N_2981,N_2622,N_2716);
nor U2982 (N_2982,N_2626,N_2744);
or U2983 (N_2983,N_2666,N_2775);
or U2984 (N_2984,N_2781,N_2692);
nor U2985 (N_2985,N_2771,N_2753);
xnor U2986 (N_2986,N_2768,N_2774);
or U2987 (N_2987,N_2661,N_2622);
nand U2988 (N_2988,N_2702,N_2637);
or U2989 (N_2989,N_2699,N_2659);
xnor U2990 (N_2990,N_2610,N_2799);
nand U2991 (N_2991,N_2785,N_2645);
and U2992 (N_2992,N_2670,N_2728);
nor U2993 (N_2993,N_2624,N_2654);
and U2994 (N_2994,N_2737,N_2746);
or U2995 (N_2995,N_2620,N_2618);
and U2996 (N_2996,N_2644,N_2623);
and U2997 (N_2997,N_2750,N_2780);
nor U2998 (N_2998,N_2624,N_2611);
nor U2999 (N_2999,N_2760,N_2735);
and U3000 (N_3000,N_2952,N_2942);
and U3001 (N_3001,N_2903,N_2977);
and U3002 (N_3002,N_2959,N_2895);
nor U3003 (N_3003,N_2946,N_2823);
and U3004 (N_3004,N_2811,N_2933);
or U3005 (N_3005,N_2882,N_2804);
nor U3006 (N_3006,N_2867,N_2824);
nand U3007 (N_3007,N_2845,N_2944);
nand U3008 (N_3008,N_2938,N_2885);
xor U3009 (N_3009,N_2857,N_2881);
xnor U3010 (N_3010,N_2987,N_2925);
nor U3011 (N_3011,N_2991,N_2806);
or U3012 (N_3012,N_2931,N_2874);
xor U3013 (N_3013,N_2937,N_2920);
nand U3014 (N_3014,N_2837,N_2955);
nor U3015 (N_3015,N_2922,N_2829);
and U3016 (N_3016,N_2973,N_2868);
or U3017 (N_3017,N_2919,N_2914);
nand U3018 (N_3018,N_2932,N_2842);
xnor U3019 (N_3019,N_2865,N_2912);
or U3020 (N_3020,N_2956,N_2815);
nand U3021 (N_3021,N_2966,N_2856);
and U3022 (N_3022,N_2838,N_2821);
xor U3023 (N_3023,N_2846,N_2855);
and U3024 (N_3024,N_2849,N_2820);
or U3025 (N_3025,N_2911,N_2992);
and U3026 (N_3026,N_2803,N_2915);
nand U3027 (N_3027,N_2801,N_2904);
nor U3028 (N_3028,N_2861,N_2945);
nand U3029 (N_3029,N_2962,N_2948);
and U3030 (N_3030,N_2957,N_2941);
or U3031 (N_3031,N_2984,N_2917);
or U3032 (N_3032,N_2918,N_2809);
nand U3033 (N_3033,N_2864,N_2875);
nand U3034 (N_3034,N_2817,N_2923);
nand U3035 (N_3035,N_2884,N_2947);
or U3036 (N_3036,N_2900,N_2808);
or U3037 (N_3037,N_2913,N_2985);
and U3038 (N_3038,N_2847,N_2862);
and U3039 (N_3039,N_2907,N_2814);
or U3040 (N_3040,N_2971,N_2830);
nand U3041 (N_3041,N_2954,N_2980);
nor U3042 (N_3042,N_2958,N_2975);
and U3043 (N_3043,N_2848,N_2894);
nand U3044 (N_3044,N_2889,N_2807);
nand U3045 (N_3045,N_2892,N_2939);
nand U3046 (N_3046,N_2998,N_2990);
nand U3047 (N_3047,N_2978,N_2982);
and U3048 (N_3048,N_2983,N_2981);
nor U3049 (N_3049,N_2877,N_2970);
and U3050 (N_3050,N_2963,N_2924);
nor U3051 (N_3051,N_2886,N_2943);
or U3052 (N_3052,N_2831,N_2967);
or U3053 (N_3053,N_2995,N_2835);
and U3054 (N_3054,N_2974,N_2960);
and U3055 (N_3055,N_2896,N_2927);
nor U3056 (N_3056,N_2964,N_2839);
and U3057 (N_3057,N_2841,N_2993);
nand U3058 (N_3058,N_2879,N_2816);
nand U3059 (N_3059,N_2910,N_2908);
xor U3060 (N_3060,N_2986,N_2812);
and U3061 (N_3061,N_2870,N_2972);
nor U3062 (N_3062,N_2836,N_2961);
nand U3063 (N_3063,N_2872,N_2826);
nor U3064 (N_3064,N_2858,N_2949);
or U3065 (N_3065,N_2888,N_2953);
nand U3066 (N_3066,N_2905,N_2869);
or U3067 (N_3067,N_2880,N_2822);
and U3068 (N_3068,N_2940,N_2936);
nand U3069 (N_3069,N_2828,N_2883);
nor U3070 (N_3070,N_2916,N_2832);
and U3071 (N_3071,N_2988,N_2890);
or U3072 (N_3072,N_2851,N_2802);
or U3073 (N_3073,N_2813,N_2928);
nor U3074 (N_3074,N_2929,N_2897);
nor U3075 (N_3075,N_2901,N_2976);
and U3076 (N_3076,N_2860,N_2989);
or U3077 (N_3077,N_2852,N_2997);
xor U3078 (N_3078,N_2853,N_2891);
nand U3079 (N_3079,N_2921,N_2878);
xor U3080 (N_3080,N_2930,N_2844);
nand U3081 (N_3081,N_2909,N_2935);
nor U3082 (N_3082,N_2873,N_2906);
and U3083 (N_3083,N_2876,N_2850);
xor U3084 (N_3084,N_2833,N_2840);
and U3085 (N_3085,N_2994,N_2968);
xor U3086 (N_3086,N_2859,N_2996);
xnor U3087 (N_3087,N_2887,N_2819);
and U3088 (N_3088,N_2893,N_2871);
nand U3089 (N_3089,N_2934,N_2866);
or U3090 (N_3090,N_2825,N_2854);
nand U3091 (N_3091,N_2898,N_2965);
nor U3092 (N_3092,N_2999,N_2950);
and U3093 (N_3093,N_2899,N_2843);
nor U3094 (N_3094,N_2827,N_2979);
or U3095 (N_3095,N_2926,N_2800);
nand U3096 (N_3096,N_2805,N_2863);
and U3097 (N_3097,N_2818,N_2969);
and U3098 (N_3098,N_2810,N_2951);
nand U3099 (N_3099,N_2834,N_2902);
xor U3100 (N_3100,N_2889,N_2979);
nand U3101 (N_3101,N_2937,N_2869);
or U3102 (N_3102,N_2810,N_2839);
and U3103 (N_3103,N_2845,N_2989);
nor U3104 (N_3104,N_2979,N_2881);
or U3105 (N_3105,N_2953,N_2923);
nand U3106 (N_3106,N_2998,N_2942);
nor U3107 (N_3107,N_2831,N_2981);
or U3108 (N_3108,N_2955,N_2919);
and U3109 (N_3109,N_2933,N_2971);
nand U3110 (N_3110,N_2828,N_2933);
nor U3111 (N_3111,N_2847,N_2826);
or U3112 (N_3112,N_2805,N_2992);
or U3113 (N_3113,N_2897,N_2954);
nor U3114 (N_3114,N_2806,N_2938);
nor U3115 (N_3115,N_2891,N_2955);
nor U3116 (N_3116,N_2868,N_2845);
nand U3117 (N_3117,N_2840,N_2955);
nand U3118 (N_3118,N_2969,N_2864);
and U3119 (N_3119,N_2948,N_2826);
and U3120 (N_3120,N_2959,N_2956);
nor U3121 (N_3121,N_2801,N_2828);
and U3122 (N_3122,N_2993,N_2859);
and U3123 (N_3123,N_2806,N_2868);
nor U3124 (N_3124,N_2821,N_2905);
and U3125 (N_3125,N_2992,N_2800);
or U3126 (N_3126,N_2908,N_2899);
or U3127 (N_3127,N_2958,N_2890);
nand U3128 (N_3128,N_2850,N_2918);
and U3129 (N_3129,N_2995,N_2917);
nor U3130 (N_3130,N_2939,N_2990);
nand U3131 (N_3131,N_2865,N_2896);
and U3132 (N_3132,N_2979,N_2896);
nand U3133 (N_3133,N_2963,N_2939);
nor U3134 (N_3134,N_2899,N_2956);
nand U3135 (N_3135,N_2830,N_2835);
nand U3136 (N_3136,N_2970,N_2988);
or U3137 (N_3137,N_2909,N_2835);
and U3138 (N_3138,N_2985,N_2982);
nand U3139 (N_3139,N_2837,N_2804);
nand U3140 (N_3140,N_2967,N_2839);
and U3141 (N_3141,N_2910,N_2938);
and U3142 (N_3142,N_2979,N_2992);
or U3143 (N_3143,N_2876,N_2912);
xor U3144 (N_3144,N_2804,N_2898);
nand U3145 (N_3145,N_2990,N_2820);
nor U3146 (N_3146,N_2892,N_2860);
or U3147 (N_3147,N_2929,N_2942);
or U3148 (N_3148,N_2862,N_2957);
nand U3149 (N_3149,N_2811,N_2958);
nor U3150 (N_3150,N_2889,N_2901);
nand U3151 (N_3151,N_2969,N_2873);
nand U3152 (N_3152,N_2871,N_2874);
and U3153 (N_3153,N_2952,N_2924);
nor U3154 (N_3154,N_2941,N_2869);
nor U3155 (N_3155,N_2945,N_2914);
and U3156 (N_3156,N_2854,N_2956);
and U3157 (N_3157,N_2818,N_2813);
and U3158 (N_3158,N_2915,N_2817);
and U3159 (N_3159,N_2842,N_2876);
or U3160 (N_3160,N_2884,N_2861);
or U3161 (N_3161,N_2928,N_2939);
or U3162 (N_3162,N_2949,N_2904);
nor U3163 (N_3163,N_2893,N_2950);
nand U3164 (N_3164,N_2855,N_2978);
nand U3165 (N_3165,N_2964,N_2931);
and U3166 (N_3166,N_2934,N_2992);
and U3167 (N_3167,N_2934,N_2922);
nor U3168 (N_3168,N_2853,N_2883);
nor U3169 (N_3169,N_2823,N_2933);
or U3170 (N_3170,N_2806,N_2839);
or U3171 (N_3171,N_2967,N_2923);
or U3172 (N_3172,N_2829,N_2972);
nor U3173 (N_3173,N_2898,N_2867);
or U3174 (N_3174,N_2834,N_2959);
nor U3175 (N_3175,N_2929,N_2902);
xnor U3176 (N_3176,N_2840,N_2903);
or U3177 (N_3177,N_2853,N_2893);
nor U3178 (N_3178,N_2965,N_2909);
nand U3179 (N_3179,N_2891,N_2824);
nand U3180 (N_3180,N_2802,N_2858);
and U3181 (N_3181,N_2843,N_2878);
nor U3182 (N_3182,N_2857,N_2959);
and U3183 (N_3183,N_2815,N_2804);
nor U3184 (N_3184,N_2844,N_2972);
nor U3185 (N_3185,N_2862,N_2899);
and U3186 (N_3186,N_2838,N_2954);
or U3187 (N_3187,N_2882,N_2841);
nor U3188 (N_3188,N_2898,N_2842);
nor U3189 (N_3189,N_2929,N_2826);
or U3190 (N_3190,N_2962,N_2857);
nor U3191 (N_3191,N_2935,N_2804);
and U3192 (N_3192,N_2905,N_2894);
and U3193 (N_3193,N_2857,N_2804);
nand U3194 (N_3194,N_2895,N_2813);
xor U3195 (N_3195,N_2863,N_2829);
nor U3196 (N_3196,N_2921,N_2853);
nor U3197 (N_3197,N_2818,N_2871);
or U3198 (N_3198,N_2802,N_2899);
and U3199 (N_3199,N_2948,N_2895);
or U3200 (N_3200,N_3070,N_3005);
and U3201 (N_3201,N_3098,N_3068);
nor U3202 (N_3202,N_3161,N_3185);
xnor U3203 (N_3203,N_3197,N_3053);
or U3204 (N_3204,N_3015,N_3082);
or U3205 (N_3205,N_3138,N_3007);
and U3206 (N_3206,N_3170,N_3013);
and U3207 (N_3207,N_3081,N_3093);
and U3208 (N_3208,N_3184,N_3104);
or U3209 (N_3209,N_3164,N_3146);
or U3210 (N_3210,N_3171,N_3177);
and U3211 (N_3211,N_3190,N_3012);
xor U3212 (N_3212,N_3024,N_3017);
and U3213 (N_3213,N_3144,N_3052);
and U3214 (N_3214,N_3096,N_3191);
nor U3215 (N_3215,N_3108,N_3189);
nor U3216 (N_3216,N_3183,N_3139);
nor U3217 (N_3217,N_3182,N_3167);
nand U3218 (N_3218,N_3100,N_3030);
nand U3219 (N_3219,N_3141,N_3049);
and U3220 (N_3220,N_3157,N_3174);
or U3221 (N_3221,N_3113,N_3175);
or U3222 (N_3222,N_3143,N_3055);
nor U3223 (N_3223,N_3045,N_3065);
nor U3224 (N_3224,N_3173,N_3048);
or U3225 (N_3225,N_3155,N_3033);
nor U3226 (N_3226,N_3066,N_3057);
nor U3227 (N_3227,N_3089,N_3014);
or U3228 (N_3228,N_3000,N_3072);
or U3229 (N_3229,N_3136,N_3036);
or U3230 (N_3230,N_3181,N_3067);
and U3231 (N_3231,N_3169,N_3087);
nor U3232 (N_3232,N_3004,N_3102);
or U3233 (N_3233,N_3010,N_3140);
nand U3234 (N_3234,N_3129,N_3124);
xor U3235 (N_3235,N_3097,N_3076);
nand U3236 (N_3236,N_3160,N_3121);
nand U3237 (N_3237,N_3162,N_3147);
or U3238 (N_3238,N_3018,N_3195);
or U3239 (N_3239,N_3071,N_3176);
nand U3240 (N_3240,N_3056,N_3064);
or U3241 (N_3241,N_3074,N_3073);
xnor U3242 (N_3242,N_3192,N_3040);
nor U3243 (N_3243,N_3106,N_3092);
or U3244 (N_3244,N_3101,N_3103);
nand U3245 (N_3245,N_3107,N_3084);
nor U3246 (N_3246,N_3080,N_3026);
or U3247 (N_3247,N_3008,N_3047);
or U3248 (N_3248,N_3088,N_3193);
nand U3249 (N_3249,N_3148,N_3196);
and U3250 (N_3250,N_3091,N_3060);
and U3251 (N_3251,N_3038,N_3127);
nand U3252 (N_3252,N_3044,N_3166);
nor U3253 (N_3253,N_3020,N_3165);
nand U3254 (N_3254,N_3151,N_3125);
nand U3255 (N_3255,N_3051,N_3130);
nand U3256 (N_3256,N_3134,N_3094);
or U3257 (N_3257,N_3043,N_3194);
nand U3258 (N_3258,N_3159,N_3090);
or U3259 (N_3259,N_3180,N_3118);
or U3260 (N_3260,N_3077,N_3109);
and U3261 (N_3261,N_3079,N_3062);
or U3262 (N_3262,N_3027,N_3172);
and U3263 (N_3263,N_3150,N_3086);
nor U3264 (N_3264,N_3003,N_3059);
and U3265 (N_3265,N_3023,N_3112);
xnor U3266 (N_3266,N_3119,N_3085);
nor U3267 (N_3267,N_3163,N_3039);
xnor U3268 (N_3268,N_3032,N_3029);
or U3269 (N_3269,N_3002,N_3132);
nor U3270 (N_3270,N_3135,N_3016);
nand U3271 (N_3271,N_3123,N_3110);
nand U3272 (N_3272,N_3154,N_3061);
or U3273 (N_3273,N_3105,N_3041);
and U3274 (N_3274,N_3006,N_3050);
nor U3275 (N_3275,N_3042,N_3156);
nor U3276 (N_3276,N_3011,N_3178);
xor U3277 (N_3277,N_3021,N_3019);
and U3278 (N_3278,N_3054,N_3199);
nor U3279 (N_3279,N_3037,N_3025);
nor U3280 (N_3280,N_3187,N_3149);
nand U3281 (N_3281,N_3001,N_3046);
nand U3282 (N_3282,N_3153,N_3133);
nor U3283 (N_3283,N_3095,N_3117);
and U3284 (N_3284,N_3145,N_3126);
xor U3285 (N_3285,N_3028,N_3111);
and U3286 (N_3286,N_3131,N_3075);
xnor U3287 (N_3287,N_3122,N_3069);
or U3288 (N_3288,N_3114,N_3009);
or U3289 (N_3289,N_3022,N_3142);
nand U3290 (N_3290,N_3179,N_3128);
xor U3291 (N_3291,N_3034,N_3137);
nand U3292 (N_3292,N_3120,N_3083);
nor U3293 (N_3293,N_3188,N_3078);
nand U3294 (N_3294,N_3035,N_3099);
and U3295 (N_3295,N_3058,N_3152);
or U3296 (N_3296,N_3186,N_3168);
and U3297 (N_3297,N_3063,N_3031);
and U3298 (N_3298,N_3158,N_3115);
nand U3299 (N_3299,N_3198,N_3116);
nand U3300 (N_3300,N_3003,N_3136);
xnor U3301 (N_3301,N_3010,N_3106);
nor U3302 (N_3302,N_3081,N_3043);
nor U3303 (N_3303,N_3169,N_3043);
and U3304 (N_3304,N_3097,N_3176);
or U3305 (N_3305,N_3158,N_3191);
xor U3306 (N_3306,N_3063,N_3141);
and U3307 (N_3307,N_3042,N_3102);
or U3308 (N_3308,N_3014,N_3150);
nor U3309 (N_3309,N_3174,N_3197);
or U3310 (N_3310,N_3177,N_3043);
nor U3311 (N_3311,N_3073,N_3063);
or U3312 (N_3312,N_3185,N_3074);
nand U3313 (N_3313,N_3085,N_3136);
and U3314 (N_3314,N_3007,N_3124);
and U3315 (N_3315,N_3006,N_3111);
and U3316 (N_3316,N_3161,N_3162);
or U3317 (N_3317,N_3009,N_3035);
xor U3318 (N_3318,N_3003,N_3176);
nor U3319 (N_3319,N_3002,N_3031);
nor U3320 (N_3320,N_3061,N_3003);
nor U3321 (N_3321,N_3011,N_3175);
nand U3322 (N_3322,N_3017,N_3089);
nand U3323 (N_3323,N_3156,N_3198);
nor U3324 (N_3324,N_3002,N_3152);
nor U3325 (N_3325,N_3124,N_3020);
xor U3326 (N_3326,N_3062,N_3021);
nand U3327 (N_3327,N_3007,N_3101);
nor U3328 (N_3328,N_3010,N_3024);
nand U3329 (N_3329,N_3173,N_3049);
or U3330 (N_3330,N_3138,N_3139);
or U3331 (N_3331,N_3070,N_3094);
nor U3332 (N_3332,N_3164,N_3049);
or U3333 (N_3333,N_3103,N_3162);
or U3334 (N_3334,N_3036,N_3052);
nor U3335 (N_3335,N_3070,N_3096);
nor U3336 (N_3336,N_3161,N_3044);
or U3337 (N_3337,N_3020,N_3000);
or U3338 (N_3338,N_3164,N_3044);
and U3339 (N_3339,N_3015,N_3025);
xor U3340 (N_3340,N_3049,N_3152);
nand U3341 (N_3341,N_3072,N_3134);
or U3342 (N_3342,N_3099,N_3009);
or U3343 (N_3343,N_3001,N_3007);
and U3344 (N_3344,N_3188,N_3147);
nor U3345 (N_3345,N_3084,N_3097);
nand U3346 (N_3346,N_3118,N_3032);
and U3347 (N_3347,N_3101,N_3160);
nand U3348 (N_3348,N_3049,N_3193);
nor U3349 (N_3349,N_3081,N_3180);
or U3350 (N_3350,N_3102,N_3087);
or U3351 (N_3351,N_3063,N_3169);
nor U3352 (N_3352,N_3089,N_3035);
nand U3353 (N_3353,N_3044,N_3152);
or U3354 (N_3354,N_3036,N_3133);
and U3355 (N_3355,N_3181,N_3084);
nor U3356 (N_3356,N_3095,N_3032);
nand U3357 (N_3357,N_3108,N_3169);
or U3358 (N_3358,N_3003,N_3149);
and U3359 (N_3359,N_3173,N_3046);
and U3360 (N_3360,N_3107,N_3117);
nor U3361 (N_3361,N_3080,N_3100);
nand U3362 (N_3362,N_3066,N_3087);
xor U3363 (N_3363,N_3012,N_3195);
nor U3364 (N_3364,N_3188,N_3193);
nor U3365 (N_3365,N_3046,N_3181);
nand U3366 (N_3366,N_3096,N_3123);
and U3367 (N_3367,N_3193,N_3184);
and U3368 (N_3368,N_3131,N_3195);
nand U3369 (N_3369,N_3176,N_3140);
or U3370 (N_3370,N_3100,N_3040);
or U3371 (N_3371,N_3029,N_3051);
nand U3372 (N_3372,N_3184,N_3091);
nand U3373 (N_3373,N_3178,N_3092);
or U3374 (N_3374,N_3077,N_3007);
or U3375 (N_3375,N_3100,N_3138);
nor U3376 (N_3376,N_3132,N_3102);
xor U3377 (N_3377,N_3188,N_3050);
nand U3378 (N_3378,N_3127,N_3067);
or U3379 (N_3379,N_3018,N_3193);
or U3380 (N_3380,N_3049,N_3085);
or U3381 (N_3381,N_3157,N_3068);
nand U3382 (N_3382,N_3118,N_3092);
nor U3383 (N_3383,N_3163,N_3121);
nor U3384 (N_3384,N_3146,N_3125);
and U3385 (N_3385,N_3006,N_3046);
nand U3386 (N_3386,N_3129,N_3125);
nand U3387 (N_3387,N_3139,N_3105);
nor U3388 (N_3388,N_3040,N_3008);
xor U3389 (N_3389,N_3156,N_3087);
or U3390 (N_3390,N_3157,N_3171);
nor U3391 (N_3391,N_3002,N_3189);
xor U3392 (N_3392,N_3078,N_3095);
and U3393 (N_3393,N_3194,N_3135);
nand U3394 (N_3394,N_3106,N_3111);
or U3395 (N_3395,N_3126,N_3182);
nand U3396 (N_3396,N_3010,N_3134);
and U3397 (N_3397,N_3090,N_3126);
nor U3398 (N_3398,N_3139,N_3001);
nor U3399 (N_3399,N_3114,N_3157);
nor U3400 (N_3400,N_3270,N_3218);
nor U3401 (N_3401,N_3343,N_3209);
nor U3402 (N_3402,N_3210,N_3333);
nand U3403 (N_3403,N_3264,N_3371);
and U3404 (N_3404,N_3356,N_3368);
xnor U3405 (N_3405,N_3211,N_3361);
or U3406 (N_3406,N_3373,N_3257);
xnor U3407 (N_3407,N_3310,N_3359);
nor U3408 (N_3408,N_3347,N_3362);
or U3409 (N_3409,N_3379,N_3224);
nand U3410 (N_3410,N_3354,N_3344);
nand U3411 (N_3411,N_3364,N_3208);
nand U3412 (N_3412,N_3340,N_3276);
nand U3413 (N_3413,N_3203,N_3274);
xnor U3414 (N_3414,N_3200,N_3380);
nand U3415 (N_3415,N_3350,N_3248);
nand U3416 (N_3416,N_3281,N_3271);
or U3417 (N_3417,N_3235,N_3267);
nand U3418 (N_3418,N_3346,N_3323);
or U3419 (N_3419,N_3345,N_3374);
or U3420 (N_3420,N_3355,N_3278);
and U3421 (N_3421,N_3334,N_3256);
nor U3422 (N_3422,N_3395,N_3304);
xnor U3423 (N_3423,N_3279,N_3324);
and U3424 (N_3424,N_3313,N_3341);
or U3425 (N_3425,N_3298,N_3321);
or U3426 (N_3426,N_3363,N_3201);
or U3427 (N_3427,N_3352,N_3383);
xor U3428 (N_3428,N_3392,N_3282);
nand U3429 (N_3429,N_3360,N_3311);
nand U3430 (N_3430,N_3222,N_3295);
nand U3431 (N_3431,N_3205,N_3296);
or U3432 (N_3432,N_3314,N_3332);
or U3433 (N_3433,N_3221,N_3250);
and U3434 (N_3434,N_3317,N_3348);
nor U3435 (N_3435,N_3391,N_3312);
or U3436 (N_3436,N_3377,N_3214);
or U3437 (N_3437,N_3398,N_3286);
nor U3438 (N_3438,N_3358,N_3397);
xnor U3439 (N_3439,N_3337,N_3249);
xnor U3440 (N_3440,N_3285,N_3236);
xor U3441 (N_3441,N_3389,N_3390);
nand U3442 (N_3442,N_3247,N_3303);
nand U3443 (N_3443,N_3302,N_3294);
xnor U3444 (N_3444,N_3233,N_3231);
or U3445 (N_3445,N_3386,N_3255);
nand U3446 (N_3446,N_3382,N_3365);
nand U3447 (N_3447,N_3297,N_3225);
and U3448 (N_3448,N_3378,N_3385);
and U3449 (N_3449,N_3399,N_3384);
or U3450 (N_3450,N_3239,N_3237);
nand U3451 (N_3451,N_3353,N_3393);
or U3452 (N_3452,N_3202,N_3308);
and U3453 (N_3453,N_3326,N_3375);
nor U3454 (N_3454,N_3357,N_3316);
nor U3455 (N_3455,N_3288,N_3215);
or U3456 (N_3456,N_3251,N_3227);
or U3457 (N_3457,N_3206,N_3226);
xor U3458 (N_3458,N_3238,N_3372);
or U3459 (N_3459,N_3260,N_3289);
or U3460 (N_3460,N_3263,N_3292);
nor U3461 (N_3461,N_3217,N_3376);
nor U3462 (N_3462,N_3327,N_3299);
nand U3463 (N_3463,N_3280,N_3325);
and U3464 (N_3464,N_3309,N_3212);
nor U3465 (N_3465,N_3349,N_3219);
nor U3466 (N_3466,N_3351,N_3223);
xor U3467 (N_3467,N_3213,N_3388);
nor U3468 (N_3468,N_3265,N_3240);
or U3469 (N_3469,N_3381,N_3246);
and U3470 (N_3470,N_3262,N_3230);
xor U3471 (N_3471,N_3319,N_3272);
or U3472 (N_3472,N_3300,N_3291);
or U3473 (N_3473,N_3336,N_3284);
nand U3474 (N_3474,N_3320,N_3366);
nand U3475 (N_3475,N_3305,N_3234);
or U3476 (N_3476,N_3396,N_3245);
and U3477 (N_3477,N_3273,N_3287);
nand U3478 (N_3478,N_3301,N_3318);
nand U3479 (N_3479,N_3329,N_3266);
nand U3480 (N_3480,N_3322,N_3220);
xnor U3481 (N_3481,N_3232,N_3290);
or U3482 (N_3482,N_3369,N_3242);
xnor U3483 (N_3483,N_3307,N_3204);
xnor U3484 (N_3484,N_3228,N_3253);
or U3485 (N_3485,N_3342,N_3261);
nor U3486 (N_3486,N_3306,N_3370);
xnor U3487 (N_3487,N_3269,N_3339);
nor U3488 (N_3488,N_3243,N_3338);
or U3489 (N_3489,N_3254,N_3328);
xor U3490 (N_3490,N_3330,N_3252);
nor U3491 (N_3491,N_3293,N_3229);
nand U3492 (N_3492,N_3241,N_3331);
or U3493 (N_3493,N_3258,N_3275);
or U3494 (N_3494,N_3367,N_3207);
and U3495 (N_3495,N_3259,N_3283);
or U3496 (N_3496,N_3335,N_3387);
and U3497 (N_3497,N_3394,N_3277);
nor U3498 (N_3498,N_3315,N_3244);
nor U3499 (N_3499,N_3216,N_3268);
xnor U3500 (N_3500,N_3371,N_3346);
and U3501 (N_3501,N_3374,N_3382);
nor U3502 (N_3502,N_3389,N_3365);
or U3503 (N_3503,N_3320,N_3243);
nor U3504 (N_3504,N_3226,N_3212);
or U3505 (N_3505,N_3380,N_3259);
nor U3506 (N_3506,N_3287,N_3297);
nand U3507 (N_3507,N_3276,N_3244);
nand U3508 (N_3508,N_3304,N_3268);
nor U3509 (N_3509,N_3359,N_3366);
or U3510 (N_3510,N_3214,N_3351);
nor U3511 (N_3511,N_3249,N_3362);
or U3512 (N_3512,N_3309,N_3369);
xor U3513 (N_3513,N_3309,N_3297);
or U3514 (N_3514,N_3394,N_3339);
or U3515 (N_3515,N_3220,N_3246);
and U3516 (N_3516,N_3293,N_3322);
xor U3517 (N_3517,N_3332,N_3289);
or U3518 (N_3518,N_3268,N_3309);
nand U3519 (N_3519,N_3350,N_3283);
and U3520 (N_3520,N_3245,N_3368);
nand U3521 (N_3521,N_3215,N_3347);
and U3522 (N_3522,N_3240,N_3263);
and U3523 (N_3523,N_3279,N_3398);
and U3524 (N_3524,N_3208,N_3299);
nand U3525 (N_3525,N_3303,N_3364);
or U3526 (N_3526,N_3320,N_3331);
nor U3527 (N_3527,N_3218,N_3395);
and U3528 (N_3528,N_3309,N_3366);
nor U3529 (N_3529,N_3204,N_3336);
or U3530 (N_3530,N_3319,N_3389);
or U3531 (N_3531,N_3283,N_3210);
nor U3532 (N_3532,N_3336,N_3387);
nand U3533 (N_3533,N_3244,N_3234);
nor U3534 (N_3534,N_3383,N_3272);
or U3535 (N_3535,N_3349,N_3304);
xor U3536 (N_3536,N_3368,N_3369);
nand U3537 (N_3537,N_3241,N_3297);
nor U3538 (N_3538,N_3356,N_3398);
and U3539 (N_3539,N_3285,N_3251);
xnor U3540 (N_3540,N_3218,N_3340);
or U3541 (N_3541,N_3259,N_3267);
and U3542 (N_3542,N_3303,N_3322);
and U3543 (N_3543,N_3264,N_3347);
and U3544 (N_3544,N_3333,N_3389);
nand U3545 (N_3545,N_3320,N_3299);
nand U3546 (N_3546,N_3393,N_3269);
and U3547 (N_3547,N_3309,N_3279);
nor U3548 (N_3548,N_3321,N_3286);
nor U3549 (N_3549,N_3300,N_3286);
and U3550 (N_3550,N_3295,N_3255);
nand U3551 (N_3551,N_3367,N_3357);
xor U3552 (N_3552,N_3294,N_3337);
nor U3553 (N_3553,N_3270,N_3220);
nand U3554 (N_3554,N_3318,N_3285);
nor U3555 (N_3555,N_3275,N_3351);
nand U3556 (N_3556,N_3339,N_3369);
nor U3557 (N_3557,N_3393,N_3289);
xnor U3558 (N_3558,N_3273,N_3327);
xor U3559 (N_3559,N_3287,N_3362);
nor U3560 (N_3560,N_3298,N_3354);
nor U3561 (N_3561,N_3376,N_3277);
and U3562 (N_3562,N_3205,N_3303);
nand U3563 (N_3563,N_3240,N_3343);
nand U3564 (N_3564,N_3311,N_3238);
and U3565 (N_3565,N_3319,N_3294);
xnor U3566 (N_3566,N_3239,N_3343);
nor U3567 (N_3567,N_3289,N_3361);
nor U3568 (N_3568,N_3335,N_3380);
and U3569 (N_3569,N_3314,N_3371);
nand U3570 (N_3570,N_3289,N_3239);
nand U3571 (N_3571,N_3285,N_3322);
nand U3572 (N_3572,N_3263,N_3297);
nor U3573 (N_3573,N_3256,N_3222);
and U3574 (N_3574,N_3303,N_3356);
or U3575 (N_3575,N_3317,N_3292);
nor U3576 (N_3576,N_3208,N_3282);
or U3577 (N_3577,N_3389,N_3305);
xor U3578 (N_3578,N_3321,N_3210);
xor U3579 (N_3579,N_3358,N_3388);
nor U3580 (N_3580,N_3355,N_3272);
nand U3581 (N_3581,N_3217,N_3341);
nand U3582 (N_3582,N_3331,N_3364);
xor U3583 (N_3583,N_3291,N_3323);
or U3584 (N_3584,N_3205,N_3311);
xnor U3585 (N_3585,N_3220,N_3217);
or U3586 (N_3586,N_3374,N_3245);
and U3587 (N_3587,N_3383,N_3348);
nor U3588 (N_3588,N_3395,N_3266);
nand U3589 (N_3589,N_3315,N_3258);
nor U3590 (N_3590,N_3288,N_3330);
or U3591 (N_3591,N_3320,N_3279);
or U3592 (N_3592,N_3361,N_3326);
or U3593 (N_3593,N_3254,N_3296);
or U3594 (N_3594,N_3388,N_3272);
nand U3595 (N_3595,N_3392,N_3215);
nand U3596 (N_3596,N_3210,N_3290);
nor U3597 (N_3597,N_3278,N_3240);
nor U3598 (N_3598,N_3243,N_3389);
or U3599 (N_3599,N_3332,N_3202);
and U3600 (N_3600,N_3482,N_3528);
nand U3601 (N_3601,N_3530,N_3485);
xnor U3602 (N_3602,N_3568,N_3555);
or U3603 (N_3603,N_3510,N_3554);
nand U3604 (N_3604,N_3419,N_3472);
xor U3605 (N_3605,N_3424,N_3545);
and U3606 (N_3606,N_3592,N_3417);
nand U3607 (N_3607,N_3562,N_3446);
nor U3608 (N_3608,N_3567,N_3453);
and U3609 (N_3609,N_3527,N_3549);
or U3610 (N_3610,N_3401,N_3440);
and U3611 (N_3611,N_3473,N_3563);
nand U3612 (N_3612,N_3483,N_3544);
xnor U3613 (N_3613,N_3529,N_3422);
xnor U3614 (N_3614,N_3409,N_3503);
nand U3615 (N_3615,N_3523,N_3546);
and U3616 (N_3616,N_3493,N_3556);
nand U3617 (N_3617,N_3414,N_3452);
nor U3618 (N_3618,N_3467,N_3486);
and U3619 (N_3619,N_3531,N_3437);
nor U3620 (N_3620,N_3598,N_3463);
and U3621 (N_3621,N_3465,N_3464);
nor U3622 (N_3622,N_3559,N_3584);
nor U3623 (N_3623,N_3541,N_3586);
and U3624 (N_3624,N_3405,N_3588);
or U3625 (N_3625,N_3438,N_3434);
xnor U3626 (N_3626,N_3479,N_3495);
nand U3627 (N_3627,N_3404,N_3475);
or U3628 (N_3628,N_3526,N_3560);
nor U3629 (N_3629,N_3427,N_3469);
nor U3630 (N_3630,N_3439,N_3577);
and U3631 (N_3631,N_3547,N_3597);
nor U3632 (N_3632,N_3506,N_3447);
nor U3633 (N_3633,N_3594,N_3599);
nand U3634 (N_3634,N_3566,N_3431);
or U3635 (N_3635,N_3569,N_3537);
nand U3636 (N_3636,N_3502,N_3575);
nor U3637 (N_3637,N_3536,N_3400);
and U3638 (N_3638,N_3406,N_3423);
nor U3639 (N_3639,N_3513,N_3505);
and U3640 (N_3640,N_3494,N_3497);
or U3641 (N_3641,N_3425,N_3455);
xnor U3642 (N_3642,N_3416,N_3520);
nand U3643 (N_3643,N_3471,N_3461);
and U3644 (N_3644,N_3490,N_3581);
nand U3645 (N_3645,N_3535,N_3408);
or U3646 (N_3646,N_3442,N_3420);
xor U3647 (N_3647,N_3524,N_3593);
and U3648 (N_3648,N_3543,N_3565);
xnor U3649 (N_3649,N_3553,N_3552);
and U3650 (N_3650,N_3561,N_3551);
or U3651 (N_3651,N_3507,N_3457);
or U3652 (N_3652,N_3449,N_3407);
nor U3653 (N_3653,N_3433,N_3430);
nand U3654 (N_3654,N_3432,N_3578);
or U3655 (N_3655,N_3585,N_3573);
nand U3656 (N_3656,N_3542,N_3410);
or U3657 (N_3657,N_3538,N_3571);
and U3658 (N_3658,N_3477,N_3454);
xor U3659 (N_3659,N_3525,N_3583);
xnor U3660 (N_3660,N_3444,N_3484);
or U3661 (N_3661,N_3451,N_3436);
and U3662 (N_3662,N_3415,N_3499);
xnor U3663 (N_3663,N_3492,N_3458);
nor U3664 (N_3664,N_3480,N_3496);
or U3665 (N_3665,N_3403,N_3596);
nand U3666 (N_3666,N_3421,N_3476);
nor U3667 (N_3667,N_3521,N_3550);
nor U3668 (N_3668,N_3540,N_3501);
nand U3669 (N_3669,N_3570,N_3532);
nor U3670 (N_3670,N_3448,N_3591);
nor U3671 (N_3671,N_3411,N_3489);
nand U3672 (N_3672,N_3487,N_3435);
or U3673 (N_3673,N_3441,N_3548);
nor U3674 (N_3674,N_3518,N_3558);
nand U3675 (N_3675,N_3481,N_3580);
or U3676 (N_3676,N_3519,N_3564);
xnor U3677 (N_3677,N_3429,N_3462);
nor U3678 (N_3678,N_3504,N_3508);
xnor U3679 (N_3679,N_3515,N_3402);
nor U3680 (N_3680,N_3478,N_3500);
xnor U3681 (N_3681,N_3474,N_3512);
and U3682 (N_3682,N_3533,N_3514);
nand U3683 (N_3683,N_3445,N_3579);
and U3684 (N_3684,N_3468,N_3456);
and U3685 (N_3685,N_3443,N_3517);
or U3686 (N_3686,N_3498,N_3516);
or U3687 (N_3687,N_3412,N_3589);
xnor U3688 (N_3688,N_3470,N_3491);
or U3689 (N_3689,N_3509,N_3534);
nand U3690 (N_3690,N_3488,N_3413);
and U3691 (N_3691,N_3428,N_3595);
and U3692 (N_3692,N_3539,N_3522);
xnor U3693 (N_3693,N_3460,N_3466);
and U3694 (N_3694,N_3582,N_3426);
or U3695 (N_3695,N_3572,N_3557);
nand U3696 (N_3696,N_3418,N_3590);
nor U3697 (N_3697,N_3587,N_3511);
and U3698 (N_3698,N_3574,N_3576);
and U3699 (N_3699,N_3450,N_3459);
or U3700 (N_3700,N_3475,N_3523);
and U3701 (N_3701,N_3452,N_3427);
nor U3702 (N_3702,N_3583,N_3581);
nand U3703 (N_3703,N_3530,N_3570);
xor U3704 (N_3704,N_3593,N_3531);
xnor U3705 (N_3705,N_3587,N_3460);
and U3706 (N_3706,N_3568,N_3418);
xnor U3707 (N_3707,N_3472,N_3490);
nor U3708 (N_3708,N_3443,N_3421);
or U3709 (N_3709,N_3464,N_3584);
and U3710 (N_3710,N_3584,N_3440);
nor U3711 (N_3711,N_3478,N_3502);
and U3712 (N_3712,N_3497,N_3409);
xor U3713 (N_3713,N_3483,N_3404);
and U3714 (N_3714,N_3520,N_3490);
or U3715 (N_3715,N_3598,N_3535);
nand U3716 (N_3716,N_3480,N_3547);
xnor U3717 (N_3717,N_3468,N_3432);
or U3718 (N_3718,N_3575,N_3457);
nor U3719 (N_3719,N_3552,N_3487);
and U3720 (N_3720,N_3597,N_3591);
or U3721 (N_3721,N_3531,N_3503);
and U3722 (N_3722,N_3419,N_3493);
and U3723 (N_3723,N_3535,N_3437);
nor U3724 (N_3724,N_3556,N_3466);
and U3725 (N_3725,N_3589,N_3423);
and U3726 (N_3726,N_3421,N_3536);
nor U3727 (N_3727,N_3453,N_3436);
nor U3728 (N_3728,N_3523,N_3457);
or U3729 (N_3729,N_3432,N_3532);
nand U3730 (N_3730,N_3586,N_3432);
nand U3731 (N_3731,N_3403,N_3416);
nand U3732 (N_3732,N_3449,N_3593);
xnor U3733 (N_3733,N_3501,N_3548);
nor U3734 (N_3734,N_3495,N_3583);
or U3735 (N_3735,N_3476,N_3498);
nand U3736 (N_3736,N_3551,N_3441);
and U3737 (N_3737,N_3579,N_3449);
or U3738 (N_3738,N_3504,N_3594);
nand U3739 (N_3739,N_3509,N_3501);
or U3740 (N_3740,N_3442,N_3596);
nor U3741 (N_3741,N_3503,N_3538);
and U3742 (N_3742,N_3583,N_3474);
and U3743 (N_3743,N_3432,N_3595);
xor U3744 (N_3744,N_3441,N_3570);
nor U3745 (N_3745,N_3471,N_3589);
or U3746 (N_3746,N_3574,N_3599);
nand U3747 (N_3747,N_3501,N_3574);
nor U3748 (N_3748,N_3441,N_3561);
and U3749 (N_3749,N_3583,N_3506);
nand U3750 (N_3750,N_3409,N_3465);
or U3751 (N_3751,N_3551,N_3424);
nand U3752 (N_3752,N_3544,N_3449);
nor U3753 (N_3753,N_3444,N_3415);
and U3754 (N_3754,N_3511,N_3576);
nand U3755 (N_3755,N_3539,N_3575);
and U3756 (N_3756,N_3578,N_3400);
nor U3757 (N_3757,N_3467,N_3534);
or U3758 (N_3758,N_3437,N_3511);
nor U3759 (N_3759,N_3454,N_3474);
and U3760 (N_3760,N_3478,N_3564);
nand U3761 (N_3761,N_3517,N_3449);
nor U3762 (N_3762,N_3407,N_3493);
or U3763 (N_3763,N_3441,N_3506);
and U3764 (N_3764,N_3416,N_3537);
nor U3765 (N_3765,N_3441,N_3494);
or U3766 (N_3766,N_3447,N_3539);
and U3767 (N_3767,N_3598,N_3546);
xor U3768 (N_3768,N_3421,N_3438);
nand U3769 (N_3769,N_3587,N_3412);
and U3770 (N_3770,N_3588,N_3552);
or U3771 (N_3771,N_3458,N_3535);
nand U3772 (N_3772,N_3402,N_3548);
nand U3773 (N_3773,N_3553,N_3452);
and U3774 (N_3774,N_3413,N_3496);
nand U3775 (N_3775,N_3442,N_3449);
and U3776 (N_3776,N_3433,N_3536);
nor U3777 (N_3777,N_3437,N_3597);
and U3778 (N_3778,N_3582,N_3533);
xor U3779 (N_3779,N_3523,N_3594);
nand U3780 (N_3780,N_3519,N_3547);
nand U3781 (N_3781,N_3402,N_3407);
nor U3782 (N_3782,N_3557,N_3530);
nor U3783 (N_3783,N_3505,N_3497);
xor U3784 (N_3784,N_3520,N_3420);
nor U3785 (N_3785,N_3411,N_3530);
nand U3786 (N_3786,N_3497,N_3487);
nand U3787 (N_3787,N_3453,N_3464);
nand U3788 (N_3788,N_3441,N_3580);
and U3789 (N_3789,N_3454,N_3429);
nand U3790 (N_3790,N_3542,N_3569);
nand U3791 (N_3791,N_3563,N_3536);
and U3792 (N_3792,N_3423,N_3485);
xor U3793 (N_3793,N_3408,N_3568);
xor U3794 (N_3794,N_3551,N_3435);
and U3795 (N_3795,N_3471,N_3533);
nand U3796 (N_3796,N_3576,N_3425);
and U3797 (N_3797,N_3593,N_3540);
or U3798 (N_3798,N_3479,N_3484);
and U3799 (N_3799,N_3498,N_3518);
nor U3800 (N_3800,N_3726,N_3797);
and U3801 (N_3801,N_3616,N_3682);
xor U3802 (N_3802,N_3735,N_3652);
nand U3803 (N_3803,N_3645,N_3796);
or U3804 (N_3804,N_3621,N_3600);
nor U3805 (N_3805,N_3658,N_3603);
nor U3806 (N_3806,N_3665,N_3715);
and U3807 (N_3807,N_3632,N_3692);
nor U3808 (N_3808,N_3719,N_3608);
xnor U3809 (N_3809,N_3684,N_3623);
and U3810 (N_3810,N_3663,N_3650);
xor U3811 (N_3811,N_3664,N_3694);
nand U3812 (N_3812,N_3611,N_3745);
nand U3813 (N_3813,N_3732,N_3761);
xnor U3814 (N_3814,N_3673,N_3606);
nand U3815 (N_3815,N_3791,N_3751);
xor U3816 (N_3816,N_3773,N_3693);
nand U3817 (N_3817,N_3769,N_3641);
nor U3818 (N_3818,N_3794,N_3772);
and U3819 (N_3819,N_3776,N_3727);
xnor U3820 (N_3820,N_3753,N_3638);
and U3821 (N_3821,N_3625,N_3701);
nand U3822 (N_3822,N_3672,N_3618);
and U3823 (N_3823,N_3774,N_3728);
nor U3824 (N_3824,N_3669,N_3661);
nor U3825 (N_3825,N_3768,N_3764);
nor U3826 (N_3826,N_3782,N_3709);
nor U3827 (N_3827,N_3722,N_3636);
xnor U3828 (N_3828,N_3703,N_3690);
or U3829 (N_3829,N_3646,N_3688);
nand U3830 (N_3830,N_3757,N_3786);
nor U3831 (N_3831,N_3729,N_3799);
and U3832 (N_3832,N_3642,N_3734);
or U3833 (N_3833,N_3754,N_3619);
and U3834 (N_3834,N_3676,N_3689);
and U3835 (N_3835,N_3717,N_3679);
xor U3836 (N_3836,N_3651,N_3724);
or U3837 (N_3837,N_3637,N_3617);
nor U3838 (N_3838,N_3749,N_3639);
nand U3839 (N_3839,N_3765,N_3696);
nand U3840 (N_3840,N_3718,N_3777);
and U3841 (N_3841,N_3737,N_3654);
nor U3842 (N_3842,N_3779,N_3771);
nor U3843 (N_3843,N_3612,N_3738);
or U3844 (N_3844,N_3667,N_3793);
nand U3845 (N_3845,N_3685,N_3741);
xor U3846 (N_3846,N_3788,N_3756);
nand U3847 (N_3847,N_3628,N_3748);
and U3848 (N_3848,N_3613,N_3784);
or U3849 (N_3849,N_3708,N_3666);
or U3850 (N_3850,N_3721,N_3712);
and U3851 (N_3851,N_3795,N_3674);
nor U3852 (N_3852,N_3624,N_3755);
nor U3853 (N_3853,N_3750,N_3675);
xor U3854 (N_3854,N_3716,N_3766);
xnor U3855 (N_3855,N_3775,N_3798);
nor U3856 (N_3856,N_3730,N_3605);
nand U3857 (N_3857,N_3622,N_3720);
nor U3858 (N_3858,N_3760,N_3648);
nand U3859 (N_3859,N_3683,N_3697);
or U3860 (N_3860,N_3781,N_3739);
and U3861 (N_3861,N_3759,N_3604);
and U3862 (N_3862,N_3691,N_3758);
or U3863 (N_3863,N_3762,N_3670);
nor U3864 (N_3864,N_3660,N_3662);
nor U3865 (N_3865,N_3677,N_3725);
or U3866 (N_3866,N_3742,N_3681);
nand U3867 (N_3867,N_3644,N_3713);
nand U3868 (N_3868,N_3671,N_3614);
and U3869 (N_3869,N_3680,N_3678);
nand U3870 (N_3870,N_3626,N_3746);
xor U3871 (N_3871,N_3783,N_3634);
and U3872 (N_3872,N_3607,N_3789);
and U3873 (N_3873,N_3640,N_3711);
or U3874 (N_3874,N_3744,N_3747);
or U3875 (N_3875,N_3695,N_3643);
nor U3876 (N_3876,N_3647,N_3687);
nor U3877 (N_3877,N_3723,N_3792);
and U3878 (N_3878,N_3627,N_3706);
nor U3879 (N_3879,N_3705,N_3610);
or U3880 (N_3880,N_3767,N_3710);
or U3881 (N_3881,N_3699,N_3707);
nor U3882 (N_3882,N_3700,N_3630);
nand U3883 (N_3883,N_3657,N_3714);
nor U3884 (N_3884,N_3733,N_3736);
or U3885 (N_3885,N_3602,N_3790);
or U3886 (N_3886,N_3780,N_3743);
nand U3887 (N_3887,N_3763,N_3609);
nand U3888 (N_3888,N_3655,N_3698);
and U3889 (N_3889,N_3702,N_3633);
or U3890 (N_3890,N_3653,N_3601);
and U3891 (N_3891,N_3740,N_3686);
and U3892 (N_3892,N_3787,N_3785);
nand U3893 (N_3893,N_3731,N_3615);
nand U3894 (N_3894,N_3631,N_3659);
and U3895 (N_3895,N_3635,N_3704);
and U3896 (N_3896,N_3668,N_3649);
or U3897 (N_3897,N_3770,N_3629);
and U3898 (N_3898,N_3656,N_3752);
or U3899 (N_3899,N_3778,N_3620);
nand U3900 (N_3900,N_3709,N_3641);
nand U3901 (N_3901,N_3755,N_3687);
or U3902 (N_3902,N_3678,N_3724);
nand U3903 (N_3903,N_3704,N_3711);
nor U3904 (N_3904,N_3784,N_3695);
nand U3905 (N_3905,N_3699,N_3691);
or U3906 (N_3906,N_3788,N_3649);
and U3907 (N_3907,N_3678,N_3623);
nor U3908 (N_3908,N_3663,N_3748);
nand U3909 (N_3909,N_3777,N_3656);
or U3910 (N_3910,N_3699,N_3740);
nand U3911 (N_3911,N_3663,N_3683);
nand U3912 (N_3912,N_3741,N_3612);
nand U3913 (N_3913,N_3701,N_3631);
or U3914 (N_3914,N_3653,N_3755);
and U3915 (N_3915,N_3749,N_3732);
nand U3916 (N_3916,N_3698,N_3696);
nor U3917 (N_3917,N_3686,N_3664);
and U3918 (N_3918,N_3655,N_3601);
xor U3919 (N_3919,N_3691,N_3667);
or U3920 (N_3920,N_3728,N_3753);
and U3921 (N_3921,N_3615,N_3711);
nor U3922 (N_3922,N_3761,N_3606);
nand U3923 (N_3923,N_3710,N_3634);
nor U3924 (N_3924,N_3612,N_3680);
nor U3925 (N_3925,N_3720,N_3607);
nand U3926 (N_3926,N_3697,N_3646);
nor U3927 (N_3927,N_3660,N_3718);
xnor U3928 (N_3928,N_3690,N_3689);
xor U3929 (N_3929,N_3645,N_3798);
nor U3930 (N_3930,N_3672,N_3755);
nand U3931 (N_3931,N_3650,N_3746);
nand U3932 (N_3932,N_3671,N_3620);
nor U3933 (N_3933,N_3633,N_3693);
or U3934 (N_3934,N_3694,N_3792);
xor U3935 (N_3935,N_3729,N_3756);
and U3936 (N_3936,N_3691,N_3752);
nand U3937 (N_3937,N_3613,N_3677);
and U3938 (N_3938,N_3718,N_3608);
nand U3939 (N_3939,N_3727,N_3636);
nand U3940 (N_3940,N_3636,N_3609);
nor U3941 (N_3941,N_3687,N_3639);
and U3942 (N_3942,N_3682,N_3653);
and U3943 (N_3943,N_3764,N_3747);
nand U3944 (N_3944,N_3674,N_3770);
nor U3945 (N_3945,N_3671,N_3667);
or U3946 (N_3946,N_3725,N_3631);
or U3947 (N_3947,N_3635,N_3681);
nand U3948 (N_3948,N_3785,N_3604);
nand U3949 (N_3949,N_3601,N_3774);
or U3950 (N_3950,N_3728,N_3742);
nor U3951 (N_3951,N_3635,N_3712);
and U3952 (N_3952,N_3761,N_3617);
and U3953 (N_3953,N_3716,N_3726);
nor U3954 (N_3954,N_3686,N_3657);
and U3955 (N_3955,N_3755,N_3657);
nand U3956 (N_3956,N_3681,N_3753);
or U3957 (N_3957,N_3629,N_3663);
nand U3958 (N_3958,N_3699,N_3779);
or U3959 (N_3959,N_3603,N_3647);
nand U3960 (N_3960,N_3749,N_3604);
nor U3961 (N_3961,N_3610,N_3671);
nand U3962 (N_3962,N_3767,N_3690);
nor U3963 (N_3963,N_3652,N_3710);
or U3964 (N_3964,N_3725,N_3621);
nor U3965 (N_3965,N_3712,N_3777);
and U3966 (N_3966,N_3672,N_3645);
or U3967 (N_3967,N_3643,N_3766);
nand U3968 (N_3968,N_3672,N_3752);
nand U3969 (N_3969,N_3623,N_3657);
nor U3970 (N_3970,N_3746,N_3756);
xnor U3971 (N_3971,N_3687,N_3785);
and U3972 (N_3972,N_3709,N_3793);
xnor U3973 (N_3973,N_3620,N_3696);
or U3974 (N_3974,N_3797,N_3724);
or U3975 (N_3975,N_3725,N_3732);
nor U3976 (N_3976,N_3726,N_3715);
nand U3977 (N_3977,N_3617,N_3608);
or U3978 (N_3978,N_3794,N_3736);
nor U3979 (N_3979,N_3621,N_3767);
nand U3980 (N_3980,N_3609,N_3628);
and U3981 (N_3981,N_3772,N_3787);
and U3982 (N_3982,N_3783,N_3680);
xor U3983 (N_3983,N_3738,N_3633);
nor U3984 (N_3984,N_3778,N_3794);
nand U3985 (N_3985,N_3612,N_3644);
or U3986 (N_3986,N_3706,N_3622);
nand U3987 (N_3987,N_3679,N_3612);
or U3988 (N_3988,N_3754,N_3677);
and U3989 (N_3989,N_3736,N_3637);
nand U3990 (N_3990,N_3759,N_3736);
nor U3991 (N_3991,N_3707,N_3632);
nor U3992 (N_3992,N_3789,N_3692);
nand U3993 (N_3993,N_3645,N_3649);
nor U3994 (N_3994,N_3605,N_3674);
nor U3995 (N_3995,N_3676,N_3600);
and U3996 (N_3996,N_3634,N_3670);
or U3997 (N_3997,N_3710,N_3782);
or U3998 (N_3998,N_3643,N_3717);
and U3999 (N_3999,N_3775,N_3652);
nand U4000 (N_4000,N_3871,N_3922);
and U4001 (N_4001,N_3901,N_3807);
or U4002 (N_4002,N_3878,N_3904);
nand U4003 (N_4003,N_3903,N_3961);
or U4004 (N_4004,N_3847,N_3941);
or U4005 (N_4005,N_3802,N_3953);
nor U4006 (N_4006,N_3841,N_3945);
nand U4007 (N_4007,N_3869,N_3921);
and U4008 (N_4008,N_3943,N_3894);
xnor U4009 (N_4009,N_3818,N_3984);
or U4010 (N_4010,N_3990,N_3987);
nor U4011 (N_4011,N_3825,N_3932);
xor U4012 (N_4012,N_3929,N_3914);
and U4013 (N_4013,N_3811,N_3843);
nand U4014 (N_4014,N_3872,N_3832);
nor U4015 (N_4015,N_3853,N_3973);
nor U4016 (N_4016,N_3955,N_3977);
or U4017 (N_4017,N_3909,N_3979);
nor U4018 (N_4018,N_3900,N_3873);
and U4019 (N_4019,N_3851,N_3927);
or U4020 (N_4020,N_3924,N_3888);
and U4021 (N_4021,N_3960,N_3854);
nor U4022 (N_4022,N_3896,N_3947);
nand U4023 (N_4023,N_3857,N_3980);
xor U4024 (N_4024,N_3966,N_3835);
nand U4025 (N_4025,N_3848,N_3938);
nand U4026 (N_4026,N_3908,N_3877);
xor U4027 (N_4027,N_3928,N_3856);
nor U4028 (N_4028,N_3940,N_3994);
nand U4029 (N_4029,N_3817,N_3936);
nand U4030 (N_4030,N_3864,N_3920);
or U4031 (N_4031,N_3972,N_3923);
xor U4032 (N_4032,N_3992,N_3944);
nor U4033 (N_4033,N_3804,N_3842);
or U4034 (N_4034,N_3988,N_3800);
and U4035 (N_4035,N_3998,N_3897);
or U4036 (N_4036,N_3926,N_3812);
and U4037 (N_4037,N_3912,N_3892);
nor U4038 (N_4038,N_3859,N_3836);
or U4039 (N_4039,N_3917,N_3883);
xnor U4040 (N_4040,N_3957,N_3861);
or U4041 (N_4041,N_3821,N_3946);
xor U4042 (N_4042,N_3951,N_3891);
nand U4043 (N_4043,N_3875,N_3833);
or U4044 (N_4044,N_3815,N_3886);
xor U4045 (N_4045,N_3898,N_3975);
xnor U4046 (N_4046,N_3824,N_3814);
nor U4047 (N_4047,N_3813,N_3999);
or U4048 (N_4048,N_3959,N_3884);
or U4049 (N_4049,N_3838,N_3822);
or U4050 (N_4050,N_3865,N_3970);
nor U4051 (N_4051,N_3965,N_3952);
xor U4052 (N_4052,N_3902,N_3808);
nand U4053 (N_4053,N_3880,N_3950);
or U4054 (N_4054,N_3963,N_3976);
nor U4055 (N_4055,N_3868,N_3849);
xnor U4056 (N_4056,N_3906,N_3937);
or U4057 (N_4057,N_3819,N_3925);
nor U4058 (N_4058,N_3930,N_3840);
nand U4059 (N_4059,N_3964,N_3866);
or U4060 (N_4060,N_3845,N_3863);
xnor U4061 (N_4061,N_3968,N_3874);
nor U4062 (N_4062,N_3803,N_3887);
and U4063 (N_4063,N_3971,N_3837);
nor U4064 (N_4064,N_3809,N_3962);
or U4065 (N_4065,N_3935,N_3991);
and U4066 (N_4066,N_3844,N_3983);
nor U4067 (N_4067,N_3846,N_3805);
nor U4068 (N_4068,N_3893,N_3997);
or U4069 (N_4069,N_3890,N_3995);
nand U4070 (N_4070,N_3850,N_3934);
and U4071 (N_4071,N_3905,N_3867);
and U4072 (N_4072,N_3830,N_3823);
xnor U4073 (N_4073,N_3870,N_3834);
and U4074 (N_4074,N_3852,N_3942);
or U4075 (N_4075,N_3882,N_3860);
nor U4076 (N_4076,N_3820,N_3829);
nor U4077 (N_4077,N_3967,N_3801);
nor U4078 (N_4078,N_3981,N_3985);
or U4079 (N_4079,N_3978,N_3956);
xnor U4080 (N_4080,N_3939,N_3996);
or U4081 (N_4081,N_3858,N_3974);
nor U4082 (N_4082,N_3933,N_3911);
or U4083 (N_4083,N_3918,N_3958);
nand U4084 (N_4084,N_3895,N_3862);
nor U4085 (N_4085,N_3910,N_3881);
or U4086 (N_4086,N_3919,N_3806);
or U4087 (N_4087,N_3931,N_3949);
nor U4088 (N_4088,N_3831,N_3828);
and U4089 (N_4089,N_3993,N_3839);
nand U4090 (N_4090,N_3826,N_3885);
or U4091 (N_4091,N_3969,N_3889);
nor U4092 (N_4092,N_3855,N_3907);
nor U4093 (N_4093,N_3954,N_3913);
nand U4094 (N_4094,N_3810,N_3916);
nand U4095 (N_4095,N_3989,N_3827);
and U4096 (N_4096,N_3816,N_3986);
nor U4097 (N_4097,N_3915,N_3876);
nand U4098 (N_4098,N_3899,N_3982);
xnor U4099 (N_4099,N_3879,N_3948);
and U4100 (N_4100,N_3805,N_3872);
xor U4101 (N_4101,N_3821,N_3966);
or U4102 (N_4102,N_3847,N_3875);
nor U4103 (N_4103,N_3973,N_3878);
nor U4104 (N_4104,N_3948,N_3966);
nor U4105 (N_4105,N_3844,N_3989);
nand U4106 (N_4106,N_3917,N_3964);
nand U4107 (N_4107,N_3804,N_3874);
and U4108 (N_4108,N_3877,N_3960);
nor U4109 (N_4109,N_3819,N_3982);
nand U4110 (N_4110,N_3908,N_3899);
or U4111 (N_4111,N_3955,N_3974);
nand U4112 (N_4112,N_3844,N_3881);
and U4113 (N_4113,N_3958,N_3804);
and U4114 (N_4114,N_3894,N_3891);
or U4115 (N_4115,N_3973,N_3962);
nand U4116 (N_4116,N_3973,N_3877);
or U4117 (N_4117,N_3998,N_3962);
xor U4118 (N_4118,N_3979,N_3883);
nand U4119 (N_4119,N_3921,N_3909);
nand U4120 (N_4120,N_3931,N_3886);
nor U4121 (N_4121,N_3844,N_3859);
nor U4122 (N_4122,N_3941,N_3923);
xor U4123 (N_4123,N_3975,N_3871);
nor U4124 (N_4124,N_3898,N_3845);
nor U4125 (N_4125,N_3897,N_3934);
xor U4126 (N_4126,N_3941,N_3857);
nor U4127 (N_4127,N_3845,N_3884);
or U4128 (N_4128,N_3870,N_3958);
nor U4129 (N_4129,N_3810,N_3848);
xor U4130 (N_4130,N_3811,N_3820);
and U4131 (N_4131,N_3928,N_3910);
nand U4132 (N_4132,N_3873,N_3996);
nor U4133 (N_4133,N_3959,N_3880);
or U4134 (N_4134,N_3832,N_3983);
nor U4135 (N_4135,N_3828,N_3945);
nor U4136 (N_4136,N_3907,N_3874);
and U4137 (N_4137,N_3880,N_3961);
nand U4138 (N_4138,N_3871,N_3935);
and U4139 (N_4139,N_3860,N_3896);
nand U4140 (N_4140,N_3835,N_3822);
and U4141 (N_4141,N_3835,N_3996);
nand U4142 (N_4142,N_3936,N_3969);
xnor U4143 (N_4143,N_3883,N_3873);
nand U4144 (N_4144,N_3826,N_3835);
nor U4145 (N_4145,N_3954,N_3896);
xnor U4146 (N_4146,N_3905,N_3859);
nand U4147 (N_4147,N_3952,N_3961);
xor U4148 (N_4148,N_3906,N_3994);
xor U4149 (N_4149,N_3816,N_3929);
xor U4150 (N_4150,N_3811,N_3806);
nand U4151 (N_4151,N_3875,N_3858);
or U4152 (N_4152,N_3807,N_3885);
or U4153 (N_4153,N_3979,N_3859);
nand U4154 (N_4154,N_3805,N_3862);
and U4155 (N_4155,N_3895,N_3916);
and U4156 (N_4156,N_3846,N_3979);
xnor U4157 (N_4157,N_3849,N_3906);
and U4158 (N_4158,N_3841,N_3988);
nor U4159 (N_4159,N_3988,N_3809);
and U4160 (N_4160,N_3805,N_3857);
nor U4161 (N_4161,N_3856,N_3847);
or U4162 (N_4162,N_3948,N_3946);
nor U4163 (N_4163,N_3891,N_3980);
nor U4164 (N_4164,N_3910,N_3819);
or U4165 (N_4165,N_3883,N_3877);
nand U4166 (N_4166,N_3839,N_3822);
nor U4167 (N_4167,N_3820,N_3944);
nor U4168 (N_4168,N_3822,N_3894);
nand U4169 (N_4169,N_3999,N_3916);
nor U4170 (N_4170,N_3853,N_3890);
nor U4171 (N_4171,N_3922,N_3977);
nor U4172 (N_4172,N_3983,N_3836);
nand U4173 (N_4173,N_3995,N_3975);
xor U4174 (N_4174,N_3909,N_3874);
nor U4175 (N_4175,N_3868,N_3957);
nand U4176 (N_4176,N_3975,N_3805);
nor U4177 (N_4177,N_3891,N_3846);
and U4178 (N_4178,N_3903,N_3921);
xnor U4179 (N_4179,N_3969,N_3880);
and U4180 (N_4180,N_3971,N_3883);
nor U4181 (N_4181,N_3963,N_3827);
and U4182 (N_4182,N_3876,N_3904);
and U4183 (N_4183,N_3931,N_3902);
nor U4184 (N_4184,N_3935,N_3984);
or U4185 (N_4185,N_3844,N_3848);
nor U4186 (N_4186,N_3948,N_3864);
and U4187 (N_4187,N_3845,N_3896);
or U4188 (N_4188,N_3881,N_3973);
or U4189 (N_4189,N_3993,N_3960);
nand U4190 (N_4190,N_3812,N_3898);
nor U4191 (N_4191,N_3945,N_3966);
and U4192 (N_4192,N_3951,N_3923);
nor U4193 (N_4193,N_3818,N_3841);
or U4194 (N_4194,N_3818,N_3971);
or U4195 (N_4195,N_3910,N_3800);
or U4196 (N_4196,N_3963,N_3966);
or U4197 (N_4197,N_3861,N_3935);
or U4198 (N_4198,N_3909,N_3983);
and U4199 (N_4199,N_3800,N_3998);
nor U4200 (N_4200,N_4127,N_4192);
nand U4201 (N_4201,N_4072,N_4083);
and U4202 (N_4202,N_4197,N_4071);
or U4203 (N_4203,N_4195,N_4092);
and U4204 (N_4204,N_4185,N_4038);
nor U4205 (N_4205,N_4084,N_4052);
nand U4206 (N_4206,N_4015,N_4163);
or U4207 (N_4207,N_4187,N_4147);
and U4208 (N_4208,N_4130,N_4003);
nor U4209 (N_4209,N_4004,N_4011);
xor U4210 (N_4210,N_4090,N_4077);
xnor U4211 (N_4211,N_4001,N_4093);
or U4212 (N_4212,N_4022,N_4153);
nand U4213 (N_4213,N_4044,N_4189);
nor U4214 (N_4214,N_4050,N_4021);
nor U4215 (N_4215,N_4150,N_4199);
nor U4216 (N_4216,N_4117,N_4188);
nor U4217 (N_4217,N_4014,N_4110);
nor U4218 (N_4218,N_4159,N_4142);
nand U4219 (N_4219,N_4023,N_4157);
nand U4220 (N_4220,N_4193,N_4113);
nand U4221 (N_4221,N_4190,N_4032);
or U4222 (N_4222,N_4122,N_4134);
nand U4223 (N_4223,N_4051,N_4094);
nand U4224 (N_4224,N_4140,N_4065);
nand U4225 (N_4225,N_4174,N_4115);
nor U4226 (N_4226,N_4136,N_4098);
and U4227 (N_4227,N_4025,N_4133);
xor U4228 (N_4228,N_4165,N_4036);
nor U4229 (N_4229,N_4000,N_4102);
nor U4230 (N_4230,N_4103,N_4074);
or U4231 (N_4231,N_4033,N_4068);
nand U4232 (N_4232,N_4069,N_4131);
or U4233 (N_4233,N_4108,N_4176);
nor U4234 (N_4234,N_4008,N_4137);
or U4235 (N_4235,N_4064,N_4018);
nor U4236 (N_4236,N_4155,N_4081);
or U4237 (N_4237,N_4141,N_4107);
or U4238 (N_4238,N_4059,N_4027);
or U4239 (N_4239,N_4168,N_4112);
nor U4240 (N_4240,N_4184,N_4170);
and U4241 (N_4241,N_4191,N_4013);
nor U4242 (N_4242,N_4166,N_4161);
or U4243 (N_4243,N_4078,N_4118);
and U4244 (N_4244,N_4009,N_4047);
and U4245 (N_4245,N_4086,N_4178);
and U4246 (N_4246,N_4172,N_4125);
nor U4247 (N_4247,N_4097,N_4030);
nand U4248 (N_4248,N_4063,N_4148);
nand U4249 (N_4249,N_4169,N_4160);
nor U4250 (N_4250,N_4180,N_4196);
nor U4251 (N_4251,N_4056,N_4143);
and U4252 (N_4252,N_4067,N_4075);
and U4253 (N_4253,N_4046,N_4173);
or U4254 (N_4254,N_4167,N_4091);
or U4255 (N_4255,N_4181,N_4010);
xnor U4256 (N_4256,N_4007,N_4151);
and U4257 (N_4257,N_4149,N_4177);
nor U4258 (N_4258,N_4182,N_4126);
and U4259 (N_4259,N_4034,N_4154);
or U4260 (N_4260,N_4058,N_4061);
and U4261 (N_4261,N_4146,N_4162);
and U4262 (N_4262,N_4128,N_4198);
xor U4263 (N_4263,N_4152,N_4079);
nor U4264 (N_4264,N_4049,N_4116);
xnor U4265 (N_4265,N_4085,N_4089);
xnor U4266 (N_4266,N_4119,N_4144);
or U4267 (N_4267,N_4186,N_4179);
or U4268 (N_4268,N_4017,N_4120);
nand U4269 (N_4269,N_4145,N_4053);
nand U4270 (N_4270,N_4055,N_4037);
or U4271 (N_4271,N_4080,N_4002);
and U4272 (N_4272,N_4100,N_4139);
and U4273 (N_4273,N_4066,N_4024);
or U4274 (N_4274,N_4121,N_4158);
nor U4275 (N_4275,N_4028,N_4073);
nor U4276 (N_4276,N_4114,N_4026);
nand U4277 (N_4277,N_4076,N_4135);
nor U4278 (N_4278,N_4104,N_4109);
xnor U4279 (N_4279,N_4138,N_4096);
and U4280 (N_4280,N_4175,N_4020);
or U4281 (N_4281,N_4087,N_4048);
and U4282 (N_4282,N_4054,N_4043);
xor U4283 (N_4283,N_4099,N_4060);
and U4284 (N_4284,N_4040,N_4057);
and U4285 (N_4285,N_4132,N_4012);
or U4286 (N_4286,N_4183,N_4111);
nand U4287 (N_4287,N_4129,N_4123);
nand U4288 (N_4288,N_4016,N_4171);
nand U4289 (N_4289,N_4070,N_4194);
nand U4290 (N_4290,N_4105,N_4062);
nor U4291 (N_4291,N_4005,N_4045);
nor U4292 (N_4292,N_4124,N_4095);
and U4293 (N_4293,N_4042,N_4082);
or U4294 (N_4294,N_4106,N_4164);
and U4295 (N_4295,N_4029,N_4031);
and U4296 (N_4296,N_4006,N_4019);
nand U4297 (N_4297,N_4156,N_4039);
and U4298 (N_4298,N_4088,N_4101);
and U4299 (N_4299,N_4041,N_4035);
and U4300 (N_4300,N_4118,N_4079);
or U4301 (N_4301,N_4027,N_4007);
and U4302 (N_4302,N_4069,N_4019);
nand U4303 (N_4303,N_4124,N_4180);
or U4304 (N_4304,N_4040,N_4070);
nor U4305 (N_4305,N_4089,N_4170);
xor U4306 (N_4306,N_4021,N_4107);
or U4307 (N_4307,N_4110,N_4022);
or U4308 (N_4308,N_4191,N_4046);
nand U4309 (N_4309,N_4043,N_4062);
or U4310 (N_4310,N_4081,N_4025);
nand U4311 (N_4311,N_4133,N_4183);
or U4312 (N_4312,N_4156,N_4174);
nor U4313 (N_4313,N_4196,N_4190);
or U4314 (N_4314,N_4117,N_4186);
and U4315 (N_4315,N_4029,N_4145);
nand U4316 (N_4316,N_4178,N_4128);
nand U4317 (N_4317,N_4180,N_4183);
and U4318 (N_4318,N_4127,N_4035);
and U4319 (N_4319,N_4149,N_4008);
nor U4320 (N_4320,N_4120,N_4085);
or U4321 (N_4321,N_4116,N_4156);
nand U4322 (N_4322,N_4093,N_4139);
nand U4323 (N_4323,N_4126,N_4017);
and U4324 (N_4324,N_4185,N_4031);
nor U4325 (N_4325,N_4137,N_4047);
xnor U4326 (N_4326,N_4159,N_4046);
or U4327 (N_4327,N_4118,N_4181);
xnor U4328 (N_4328,N_4082,N_4024);
nor U4329 (N_4329,N_4189,N_4100);
nand U4330 (N_4330,N_4001,N_4062);
nor U4331 (N_4331,N_4047,N_4156);
nor U4332 (N_4332,N_4076,N_4107);
nor U4333 (N_4333,N_4169,N_4054);
or U4334 (N_4334,N_4035,N_4116);
nor U4335 (N_4335,N_4149,N_4145);
nand U4336 (N_4336,N_4052,N_4069);
nor U4337 (N_4337,N_4189,N_4003);
and U4338 (N_4338,N_4105,N_4051);
nor U4339 (N_4339,N_4079,N_4065);
xor U4340 (N_4340,N_4197,N_4015);
nor U4341 (N_4341,N_4132,N_4160);
nand U4342 (N_4342,N_4138,N_4012);
or U4343 (N_4343,N_4098,N_4051);
or U4344 (N_4344,N_4022,N_4067);
or U4345 (N_4345,N_4116,N_4071);
nor U4346 (N_4346,N_4102,N_4152);
xnor U4347 (N_4347,N_4145,N_4017);
and U4348 (N_4348,N_4154,N_4026);
nor U4349 (N_4349,N_4066,N_4112);
nand U4350 (N_4350,N_4146,N_4062);
or U4351 (N_4351,N_4086,N_4144);
and U4352 (N_4352,N_4155,N_4156);
nand U4353 (N_4353,N_4129,N_4148);
and U4354 (N_4354,N_4178,N_4020);
nor U4355 (N_4355,N_4160,N_4141);
or U4356 (N_4356,N_4162,N_4153);
nor U4357 (N_4357,N_4138,N_4065);
and U4358 (N_4358,N_4008,N_4148);
and U4359 (N_4359,N_4068,N_4098);
and U4360 (N_4360,N_4181,N_4182);
nor U4361 (N_4361,N_4056,N_4090);
or U4362 (N_4362,N_4045,N_4012);
nand U4363 (N_4363,N_4025,N_4046);
nor U4364 (N_4364,N_4175,N_4120);
and U4365 (N_4365,N_4124,N_4158);
nor U4366 (N_4366,N_4018,N_4181);
and U4367 (N_4367,N_4035,N_4160);
and U4368 (N_4368,N_4035,N_4197);
xnor U4369 (N_4369,N_4169,N_4050);
and U4370 (N_4370,N_4054,N_4078);
nand U4371 (N_4371,N_4037,N_4092);
or U4372 (N_4372,N_4047,N_4159);
xnor U4373 (N_4373,N_4040,N_4161);
or U4374 (N_4374,N_4093,N_4174);
nand U4375 (N_4375,N_4103,N_4147);
nor U4376 (N_4376,N_4095,N_4184);
nand U4377 (N_4377,N_4177,N_4104);
and U4378 (N_4378,N_4165,N_4172);
nand U4379 (N_4379,N_4035,N_4130);
and U4380 (N_4380,N_4052,N_4040);
nand U4381 (N_4381,N_4027,N_4089);
or U4382 (N_4382,N_4131,N_4119);
and U4383 (N_4383,N_4018,N_4057);
and U4384 (N_4384,N_4083,N_4017);
and U4385 (N_4385,N_4049,N_4147);
nand U4386 (N_4386,N_4010,N_4018);
and U4387 (N_4387,N_4082,N_4038);
and U4388 (N_4388,N_4179,N_4075);
nand U4389 (N_4389,N_4045,N_4009);
nand U4390 (N_4390,N_4068,N_4159);
nand U4391 (N_4391,N_4097,N_4122);
nor U4392 (N_4392,N_4121,N_4166);
nand U4393 (N_4393,N_4012,N_4141);
nand U4394 (N_4394,N_4033,N_4036);
or U4395 (N_4395,N_4003,N_4111);
or U4396 (N_4396,N_4181,N_4009);
or U4397 (N_4397,N_4171,N_4191);
and U4398 (N_4398,N_4154,N_4120);
nor U4399 (N_4399,N_4095,N_4017);
or U4400 (N_4400,N_4209,N_4291);
xnor U4401 (N_4401,N_4312,N_4363);
and U4402 (N_4402,N_4304,N_4210);
and U4403 (N_4403,N_4317,N_4337);
nor U4404 (N_4404,N_4314,N_4333);
and U4405 (N_4405,N_4229,N_4364);
nand U4406 (N_4406,N_4388,N_4372);
and U4407 (N_4407,N_4336,N_4306);
xnor U4408 (N_4408,N_4320,N_4362);
nor U4409 (N_4409,N_4370,N_4201);
nor U4410 (N_4410,N_4350,N_4261);
and U4411 (N_4411,N_4205,N_4380);
nand U4412 (N_4412,N_4325,N_4351);
and U4413 (N_4413,N_4385,N_4219);
nand U4414 (N_4414,N_4313,N_4202);
and U4415 (N_4415,N_4376,N_4398);
and U4416 (N_4416,N_4305,N_4311);
or U4417 (N_4417,N_4259,N_4238);
nor U4418 (N_4418,N_4399,N_4240);
and U4419 (N_4419,N_4348,N_4239);
and U4420 (N_4420,N_4371,N_4278);
xnor U4421 (N_4421,N_4224,N_4270);
and U4422 (N_4422,N_4373,N_4241);
nand U4423 (N_4423,N_4288,N_4206);
xor U4424 (N_4424,N_4384,N_4332);
and U4425 (N_4425,N_4299,N_4282);
nand U4426 (N_4426,N_4297,N_4386);
or U4427 (N_4427,N_4276,N_4272);
or U4428 (N_4428,N_4242,N_4281);
nand U4429 (N_4429,N_4267,N_4343);
or U4430 (N_4430,N_4285,N_4392);
nor U4431 (N_4431,N_4319,N_4322);
nor U4432 (N_4432,N_4323,N_4216);
nor U4433 (N_4433,N_4356,N_4228);
xnor U4434 (N_4434,N_4315,N_4328);
or U4435 (N_4435,N_4353,N_4243);
nor U4436 (N_4436,N_4381,N_4221);
nor U4437 (N_4437,N_4227,N_4212);
nand U4438 (N_4438,N_4302,N_4346);
or U4439 (N_4439,N_4361,N_4266);
nand U4440 (N_4440,N_4377,N_4258);
nand U4441 (N_4441,N_4389,N_4365);
and U4442 (N_4442,N_4391,N_4340);
nor U4443 (N_4443,N_4215,N_4283);
or U4444 (N_4444,N_4349,N_4339);
nor U4445 (N_4445,N_4247,N_4220);
or U4446 (N_4446,N_4244,N_4255);
nor U4447 (N_4447,N_4289,N_4301);
nor U4448 (N_4448,N_4357,N_4300);
nand U4449 (N_4449,N_4284,N_4369);
xnor U4450 (N_4450,N_4207,N_4366);
or U4451 (N_4451,N_4321,N_4214);
or U4452 (N_4452,N_4268,N_4257);
or U4453 (N_4453,N_4355,N_4232);
nor U4454 (N_4454,N_4360,N_4251);
nor U4455 (N_4455,N_4330,N_4287);
and U4456 (N_4456,N_4230,N_4290);
xor U4457 (N_4457,N_4263,N_4393);
or U4458 (N_4458,N_4326,N_4245);
nand U4459 (N_4459,N_4310,N_4235);
and U4460 (N_4460,N_4303,N_4277);
or U4461 (N_4461,N_4234,N_4274);
or U4462 (N_4462,N_4262,N_4286);
and U4463 (N_4463,N_4390,N_4249);
xor U4464 (N_4464,N_4252,N_4331);
nor U4465 (N_4465,N_4378,N_4307);
nand U4466 (N_4466,N_4352,N_4279);
nor U4467 (N_4467,N_4273,N_4256);
and U4468 (N_4468,N_4396,N_4327);
nand U4469 (N_4469,N_4231,N_4233);
xor U4470 (N_4470,N_4395,N_4260);
or U4471 (N_4471,N_4397,N_4211);
nor U4472 (N_4472,N_4318,N_4367);
nor U4473 (N_4473,N_4264,N_4265);
and U4474 (N_4474,N_4254,N_4204);
xnor U4475 (N_4475,N_4250,N_4294);
or U4476 (N_4476,N_4218,N_4383);
nand U4477 (N_4477,N_4342,N_4298);
or U4478 (N_4478,N_4271,N_4293);
or U4479 (N_4479,N_4246,N_4347);
nor U4480 (N_4480,N_4394,N_4358);
nor U4481 (N_4481,N_4359,N_4225);
xor U4482 (N_4482,N_4253,N_4375);
nand U4483 (N_4483,N_4237,N_4354);
nand U4484 (N_4484,N_4226,N_4248);
and U4485 (N_4485,N_4208,N_4345);
or U4486 (N_4486,N_4309,N_4203);
and U4487 (N_4487,N_4368,N_4329);
nor U4488 (N_4488,N_4379,N_4223);
nand U4489 (N_4489,N_4269,N_4338);
and U4490 (N_4490,N_4213,N_4222);
or U4491 (N_4491,N_4308,N_4324);
xor U4492 (N_4492,N_4374,N_4344);
nor U4493 (N_4493,N_4280,N_4334);
nand U4494 (N_4494,N_4316,N_4296);
and U4495 (N_4495,N_4341,N_4200);
nor U4496 (N_4496,N_4382,N_4335);
or U4497 (N_4497,N_4292,N_4295);
and U4498 (N_4498,N_4387,N_4217);
and U4499 (N_4499,N_4236,N_4275);
nor U4500 (N_4500,N_4248,N_4241);
and U4501 (N_4501,N_4206,N_4379);
or U4502 (N_4502,N_4377,N_4349);
and U4503 (N_4503,N_4333,N_4355);
nor U4504 (N_4504,N_4234,N_4391);
or U4505 (N_4505,N_4236,N_4210);
nor U4506 (N_4506,N_4291,N_4387);
nand U4507 (N_4507,N_4355,N_4276);
nand U4508 (N_4508,N_4252,N_4302);
xnor U4509 (N_4509,N_4306,N_4328);
or U4510 (N_4510,N_4287,N_4345);
or U4511 (N_4511,N_4392,N_4229);
nor U4512 (N_4512,N_4279,N_4330);
nand U4513 (N_4513,N_4309,N_4389);
and U4514 (N_4514,N_4264,N_4305);
and U4515 (N_4515,N_4333,N_4301);
or U4516 (N_4516,N_4387,N_4313);
or U4517 (N_4517,N_4371,N_4217);
or U4518 (N_4518,N_4289,N_4320);
nor U4519 (N_4519,N_4230,N_4398);
nor U4520 (N_4520,N_4200,N_4384);
nand U4521 (N_4521,N_4325,N_4291);
and U4522 (N_4522,N_4332,N_4248);
or U4523 (N_4523,N_4342,N_4245);
nand U4524 (N_4524,N_4214,N_4296);
or U4525 (N_4525,N_4310,N_4353);
and U4526 (N_4526,N_4290,N_4359);
nand U4527 (N_4527,N_4339,N_4242);
nor U4528 (N_4528,N_4297,N_4395);
nor U4529 (N_4529,N_4305,N_4296);
nor U4530 (N_4530,N_4286,N_4292);
or U4531 (N_4531,N_4305,N_4219);
or U4532 (N_4532,N_4399,N_4223);
and U4533 (N_4533,N_4271,N_4397);
nand U4534 (N_4534,N_4385,N_4237);
or U4535 (N_4535,N_4272,N_4264);
nand U4536 (N_4536,N_4352,N_4262);
and U4537 (N_4537,N_4273,N_4205);
nor U4538 (N_4538,N_4387,N_4326);
xnor U4539 (N_4539,N_4252,N_4311);
xnor U4540 (N_4540,N_4322,N_4375);
and U4541 (N_4541,N_4238,N_4340);
and U4542 (N_4542,N_4274,N_4362);
nand U4543 (N_4543,N_4224,N_4353);
and U4544 (N_4544,N_4228,N_4244);
nor U4545 (N_4545,N_4215,N_4242);
and U4546 (N_4546,N_4223,N_4299);
and U4547 (N_4547,N_4288,N_4290);
nand U4548 (N_4548,N_4357,N_4222);
or U4549 (N_4549,N_4333,N_4305);
or U4550 (N_4550,N_4350,N_4317);
nor U4551 (N_4551,N_4259,N_4343);
nor U4552 (N_4552,N_4330,N_4291);
nand U4553 (N_4553,N_4365,N_4216);
or U4554 (N_4554,N_4397,N_4223);
xnor U4555 (N_4555,N_4298,N_4345);
nand U4556 (N_4556,N_4294,N_4263);
nand U4557 (N_4557,N_4256,N_4242);
nand U4558 (N_4558,N_4273,N_4222);
and U4559 (N_4559,N_4337,N_4282);
nand U4560 (N_4560,N_4200,N_4328);
or U4561 (N_4561,N_4399,N_4276);
nor U4562 (N_4562,N_4222,N_4399);
nand U4563 (N_4563,N_4203,N_4274);
and U4564 (N_4564,N_4350,N_4361);
or U4565 (N_4565,N_4299,N_4305);
and U4566 (N_4566,N_4289,N_4347);
nor U4567 (N_4567,N_4264,N_4329);
or U4568 (N_4568,N_4210,N_4375);
and U4569 (N_4569,N_4323,N_4338);
nand U4570 (N_4570,N_4278,N_4348);
or U4571 (N_4571,N_4202,N_4336);
or U4572 (N_4572,N_4372,N_4394);
nand U4573 (N_4573,N_4298,N_4313);
nand U4574 (N_4574,N_4260,N_4399);
nor U4575 (N_4575,N_4325,N_4320);
or U4576 (N_4576,N_4233,N_4371);
and U4577 (N_4577,N_4345,N_4277);
nand U4578 (N_4578,N_4391,N_4399);
nand U4579 (N_4579,N_4286,N_4347);
nor U4580 (N_4580,N_4224,N_4231);
nand U4581 (N_4581,N_4359,N_4304);
and U4582 (N_4582,N_4394,N_4325);
or U4583 (N_4583,N_4394,N_4242);
or U4584 (N_4584,N_4357,N_4251);
nand U4585 (N_4585,N_4215,N_4286);
and U4586 (N_4586,N_4305,N_4351);
nor U4587 (N_4587,N_4214,N_4245);
or U4588 (N_4588,N_4303,N_4345);
nand U4589 (N_4589,N_4356,N_4202);
nand U4590 (N_4590,N_4362,N_4367);
or U4591 (N_4591,N_4383,N_4267);
nand U4592 (N_4592,N_4241,N_4210);
or U4593 (N_4593,N_4334,N_4222);
nand U4594 (N_4594,N_4294,N_4303);
and U4595 (N_4595,N_4374,N_4234);
and U4596 (N_4596,N_4376,N_4314);
or U4597 (N_4597,N_4282,N_4228);
nand U4598 (N_4598,N_4241,N_4359);
or U4599 (N_4599,N_4204,N_4222);
nor U4600 (N_4600,N_4555,N_4522);
or U4601 (N_4601,N_4543,N_4423);
nor U4602 (N_4602,N_4521,N_4575);
nor U4603 (N_4603,N_4517,N_4402);
nor U4604 (N_4604,N_4540,N_4421);
nand U4605 (N_4605,N_4530,N_4587);
xnor U4606 (N_4606,N_4579,N_4584);
and U4607 (N_4607,N_4478,N_4409);
and U4608 (N_4608,N_4593,N_4516);
and U4609 (N_4609,N_4531,N_4470);
or U4610 (N_4610,N_4519,N_4414);
nand U4611 (N_4611,N_4556,N_4568);
nand U4612 (N_4612,N_4498,N_4407);
nor U4613 (N_4613,N_4432,N_4411);
xor U4614 (N_4614,N_4529,N_4582);
or U4615 (N_4615,N_4412,N_4471);
nor U4616 (N_4616,N_4477,N_4580);
nand U4617 (N_4617,N_4511,N_4461);
nand U4618 (N_4618,N_4501,N_4401);
and U4619 (N_4619,N_4539,N_4462);
and U4620 (N_4620,N_4417,N_4437);
or U4621 (N_4621,N_4436,N_4541);
xnor U4622 (N_4622,N_4496,N_4561);
or U4623 (N_4623,N_4586,N_4528);
or U4624 (N_4624,N_4583,N_4549);
nor U4625 (N_4625,N_4419,N_4502);
or U4626 (N_4626,N_4524,N_4546);
and U4627 (N_4627,N_4597,N_4483);
xor U4628 (N_4628,N_4426,N_4591);
or U4629 (N_4629,N_4515,N_4576);
nand U4630 (N_4630,N_4420,N_4507);
and U4631 (N_4631,N_4504,N_4469);
nand U4632 (N_4632,N_4512,N_4443);
nor U4633 (N_4633,N_4525,N_4481);
nor U4634 (N_4634,N_4454,N_4486);
xor U4635 (N_4635,N_4594,N_4503);
or U4636 (N_4636,N_4588,N_4415);
and U4637 (N_4637,N_4434,N_4431);
nor U4638 (N_4638,N_4554,N_4413);
nor U4639 (N_4639,N_4505,N_4596);
and U4640 (N_4640,N_4405,N_4571);
nand U4641 (N_4641,N_4425,N_4450);
or U4642 (N_4642,N_4466,N_4557);
and U4643 (N_4643,N_4495,N_4572);
and U4644 (N_4644,N_4534,N_4564);
nor U4645 (N_4645,N_4533,N_4445);
nor U4646 (N_4646,N_4416,N_4562);
nand U4647 (N_4647,N_4422,N_4492);
nand U4648 (N_4648,N_4491,N_4453);
and U4649 (N_4649,N_4460,N_4508);
and U4650 (N_4650,N_4433,N_4509);
nand U4651 (N_4651,N_4551,N_4590);
nor U4652 (N_4652,N_4544,N_4464);
xor U4653 (N_4653,N_4410,N_4441);
or U4654 (N_4654,N_4552,N_4500);
nand U4655 (N_4655,N_4468,N_4446);
and U4656 (N_4656,N_4456,N_4518);
or U4657 (N_4657,N_4506,N_4573);
nand U4658 (N_4658,N_4536,N_4489);
and U4659 (N_4659,N_4459,N_4463);
xor U4660 (N_4660,N_4563,N_4400);
nor U4661 (N_4661,N_4570,N_4484);
xnor U4662 (N_4662,N_4542,N_4550);
and U4663 (N_4663,N_4472,N_4592);
nand U4664 (N_4664,N_4424,N_4581);
and U4665 (N_4665,N_4473,N_4440);
nor U4666 (N_4666,N_4532,N_4520);
nor U4667 (N_4667,N_4558,N_4435);
or U4668 (N_4668,N_4490,N_4577);
and U4669 (N_4669,N_4447,N_4428);
nand U4670 (N_4670,N_4574,N_4452);
nand U4671 (N_4671,N_4449,N_4438);
xnor U4672 (N_4672,N_4480,N_4439);
nor U4673 (N_4673,N_4510,N_4487);
or U4674 (N_4674,N_4514,N_4427);
nor U4675 (N_4675,N_4595,N_4406);
nand U4676 (N_4676,N_4526,N_4589);
and U4677 (N_4677,N_4479,N_4567);
nor U4678 (N_4678,N_4451,N_4547);
or U4679 (N_4679,N_4523,N_4457);
or U4680 (N_4680,N_4408,N_4527);
nor U4681 (N_4681,N_4559,N_4538);
or U4682 (N_4682,N_4497,N_4545);
nand U4683 (N_4683,N_4494,N_4535);
and U4684 (N_4684,N_4429,N_4598);
and U4685 (N_4685,N_4403,N_4578);
and U4686 (N_4686,N_4474,N_4499);
or U4687 (N_4687,N_4548,N_4430);
xor U4688 (N_4688,N_4442,N_4513);
or U4689 (N_4689,N_4485,N_4560);
xnor U4690 (N_4690,N_4444,N_4553);
and U4691 (N_4691,N_4482,N_4455);
nor U4692 (N_4692,N_4493,N_4599);
nand U4693 (N_4693,N_4537,N_4569);
or U4694 (N_4694,N_4448,N_4418);
nor U4695 (N_4695,N_4465,N_4467);
or U4696 (N_4696,N_4458,N_4475);
nand U4697 (N_4697,N_4585,N_4488);
or U4698 (N_4698,N_4476,N_4404);
nand U4699 (N_4699,N_4565,N_4566);
nand U4700 (N_4700,N_4567,N_4402);
or U4701 (N_4701,N_4539,N_4452);
nand U4702 (N_4702,N_4548,N_4561);
nand U4703 (N_4703,N_4501,N_4583);
nor U4704 (N_4704,N_4506,N_4545);
or U4705 (N_4705,N_4558,N_4492);
or U4706 (N_4706,N_4502,N_4570);
nor U4707 (N_4707,N_4459,N_4464);
nor U4708 (N_4708,N_4468,N_4493);
and U4709 (N_4709,N_4434,N_4457);
or U4710 (N_4710,N_4503,N_4483);
nand U4711 (N_4711,N_4529,N_4574);
xnor U4712 (N_4712,N_4438,N_4431);
nor U4713 (N_4713,N_4519,N_4421);
nor U4714 (N_4714,N_4410,N_4462);
nand U4715 (N_4715,N_4564,N_4529);
nand U4716 (N_4716,N_4443,N_4586);
xnor U4717 (N_4717,N_4427,N_4490);
and U4718 (N_4718,N_4431,N_4562);
nand U4719 (N_4719,N_4462,N_4593);
nor U4720 (N_4720,N_4552,N_4539);
nand U4721 (N_4721,N_4437,N_4442);
nand U4722 (N_4722,N_4403,N_4570);
xor U4723 (N_4723,N_4430,N_4495);
or U4724 (N_4724,N_4474,N_4514);
nand U4725 (N_4725,N_4488,N_4468);
nand U4726 (N_4726,N_4405,N_4504);
and U4727 (N_4727,N_4489,N_4517);
nor U4728 (N_4728,N_4571,N_4517);
and U4729 (N_4729,N_4435,N_4500);
or U4730 (N_4730,N_4574,N_4429);
nor U4731 (N_4731,N_4408,N_4594);
nor U4732 (N_4732,N_4453,N_4556);
nor U4733 (N_4733,N_4431,N_4566);
and U4734 (N_4734,N_4528,N_4505);
and U4735 (N_4735,N_4416,N_4457);
or U4736 (N_4736,N_4455,N_4479);
and U4737 (N_4737,N_4520,N_4465);
nor U4738 (N_4738,N_4575,N_4578);
nand U4739 (N_4739,N_4491,N_4570);
and U4740 (N_4740,N_4403,N_4550);
nor U4741 (N_4741,N_4564,N_4467);
or U4742 (N_4742,N_4453,N_4551);
and U4743 (N_4743,N_4549,N_4586);
and U4744 (N_4744,N_4496,N_4409);
or U4745 (N_4745,N_4535,N_4519);
nand U4746 (N_4746,N_4592,N_4537);
or U4747 (N_4747,N_4411,N_4515);
nand U4748 (N_4748,N_4462,N_4492);
nor U4749 (N_4749,N_4453,N_4481);
and U4750 (N_4750,N_4448,N_4458);
and U4751 (N_4751,N_4494,N_4461);
and U4752 (N_4752,N_4528,N_4560);
nor U4753 (N_4753,N_4527,N_4540);
xor U4754 (N_4754,N_4400,N_4401);
or U4755 (N_4755,N_4564,N_4500);
and U4756 (N_4756,N_4581,N_4526);
nand U4757 (N_4757,N_4400,N_4509);
xor U4758 (N_4758,N_4510,N_4466);
nor U4759 (N_4759,N_4452,N_4486);
or U4760 (N_4760,N_4473,N_4547);
nand U4761 (N_4761,N_4547,N_4514);
nor U4762 (N_4762,N_4421,N_4582);
nand U4763 (N_4763,N_4581,N_4552);
or U4764 (N_4764,N_4418,N_4532);
xor U4765 (N_4765,N_4499,N_4475);
xor U4766 (N_4766,N_4466,N_4560);
nor U4767 (N_4767,N_4544,N_4542);
nand U4768 (N_4768,N_4460,N_4400);
or U4769 (N_4769,N_4511,N_4455);
and U4770 (N_4770,N_4598,N_4587);
and U4771 (N_4771,N_4509,N_4455);
nor U4772 (N_4772,N_4588,N_4414);
nand U4773 (N_4773,N_4418,N_4587);
xor U4774 (N_4774,N_4492,N_4474);
and U4775 (N_4775,N_4473,N_4588);
xor U4776 (N_4776,N_4415,N_4507);
nor U4777 (N_4777,N_4478,N_4534);
nand U4778 (N_4778,N_4444,N_4523);
xnor U4779 (N_4779,N_4458,N_4469);
or U4780 (N_4780,N_4553,N_4475);
and U4781 (N_4781,N_4433,N_4404);
or U4782 (N_4782,N_4514,N_4401);
and U4783 (N_4783,N_4561,N_4545);
and U4784 (N_4784,N_4542,N_4566);
nand U4785 (N_4785,N_4465,N_4416);
nor U4786 (N_4786,N_4577,N_4593);
nand U4787 (N_4787,N_4576,N_4561);
nor U4788 (N_4788,N_4588,N_4488);
nor U4789 (N_4789,N_4494,N_4508);
or U4790 (N_4790,N_4564,N_4456);
and U4791 (N_4791,N_4425,N_4451);
nor U4792 (N_4792,N_4531,N_4407);
nor U4793 (N_4793,N_4594,N_4425);
xor U4794 (N_4794,N_4468,N_4542);
nand U4795 (N_4795,N_4519,N_4465);
and U4796 (N_4796,N_4462,N_4568);
or U4797 (N_4797,N_4588,N_4460);
nand U4798 (N_4798,N_4519,N_4500);
nor U4799 (N_4799,N_4506,N_4510);
nand U4800 (N_4800,N_4725,N_4677);
xor U4801 (N_4801,N_4692,N_4676);
nand U4802 (N_4802,N_4628,N_4738);
xnor U4803 (N_4803,N_4616,N_4795);
nand U4804 (N_4804,N_4771,N_4758);
or U4805 (N_4805,N_4757,N_4642);
xnor U4806 (N_4806,N_4624,N_4764);
or U4807 (N_4807,N_4675,N_4635);
and U4808 (N_4808,N_4629,N_4678);
nand U4809 (N_4809,N_4690,N_4761);
or U4810 (N_4810,N_4740,N_4664);
or U4811 (N_4811,N_4620,N_4696);
and U4812 (N_4812,N_4614,N_4734);
nand U4813 (N_4813,N_4760,N_4631);
nand U4814 (N_4814,N_4778,N_4777);
xnor U4815 (N_4815,N_4663,N_4657);
xor U4816 (N_4816,N_4712,N_4794);
nor U4817 (N_4817,N_4773,N_4708);
xnor U4818 (N_4818,N_4759,N_4766);
nor U4819 (N_4819,N_4662,N_4775);
nand U4820 (N_4820,N_4653,N_4736);
and U4821 (N_4821,N_4729,N_4717);
or U4822 (N_4822,N_4674,N_4721);
or U4823 (N_4823,N_4601,N_4711);
and U4824 (N_4824,N_4680,N_4672);
and U4825 (N_4825,N_4750,N_4641);
nor U4826 (N_4826,N_4748,N_4713);
nand U4827 (N_4827,N_4656,N_4707);
nor U4828 (N_4828,N_4646,N_4667);
and U4829 (N_4829,N_4787,N_4726);
and U4830 (N_4830,N_4767,N_4751);
nor U4831 (N_4831,N_4654,N_4798);
and U4832 (N_4832,N_4665,N_4689);
or U4833 (N_4833,N_4705,N_4763);
and U4834 (N_4834,N_4745,N_4791);
nor U4835 (N_4835,N_4617,N_4682);
or U4836 (N_4836,N_4639,N_4783);
xor U4837 (N_4837,N_4686,N_4782);
nand U4838 (N_4838,N_4733,N_4737);
nor U4839 (N_4839,N_4785,N_4718);
and U4840 (N_4840,N_4703,N_4735);
and U4841 (N_4841,N_4730,N_4604);
nand U4842 (N_4842,N_4799,N_4790);
nor U4843 (N_4843,N_4609,N_4784);
xnor U4844 (N_4844,N_4728,N_4753);
or U4845 (N_4845,N_4781,N_4636);
nor U4846 (N_4846,N_4659,N_4684);
or U4847 (N_4847,N_4621,N_4739);
and U4848 (N_4848,N_4688,N_4797);
and U4849 (N_4849,N_4752,N_4666);
nand U4850 (N_4850,N_4608,N_4619);
and U4851 (N_4851,N_4694,N_4744);
nor U4852 (N_4852,N_4727,N_4647);
or U4853 (N_4853,N_4710,N_4632);
xor U4854 (N_4854,N_4695,N_4706);
or U4855 (N_4855,N_4768,N_4731);
and U4856 (N_4856,N_4792,N_4716);
or U4857 (N_4857,N_4762,N_4774);
nor U4858 (N_4858,N_4698,N_4671);
nand U4859 (N_4859,N_4613,N_4724);
and U4860 (N_4860,N_4786,N_4651);
nand U4861 (N_4861,N_4650,N_4648);
or U4862 (N_4862,N_4749,N_4723);
xor U4863 (N_4863,N_4746,N_4637);
nor U4864 (N_4864,N_4779,N_4722);
nand U4865 (N_4865,N_4670,N_4643);
or U4866 (N_4866,N_4742,N_4719);
nand U4867 (N_4867,N_4605,N_4600);
and U4868 (N_4868,N_4640,N_4715);
and U4869 (N_4869,N_4693,N_4615);
xor U4870 (N_4870,N_4658,N_4732);
nor U4871 (N_4871,N_4679,N_4660);
and U4872 (N_4872,N_4612,N_4687);
nand U4873 (N_4873,N_4630,N_4625);
nor U4874 (N_4874,N_4691,N_4606);
nand U4875 (N_4875,N_4638,N_4623);
and U4876 (N_4876,N_4627,N_4607);
xor U4877 (N_4877,N_4714,N_4789);
and U4878 (N_4878,N_4754,N_4673);
xor U4879 (N_4879,N_4634,N_4741);
nor U4880 (N_4880,N_4683,N_4776);
nor U4881 (N_4881,N_4743,N_4769);
nor U4882 (N_4882,N_4793,N_4649);
or U4883 (N_4883,N_4747,N_4644);
nor U4884 (N_4884,N_4645,N_4704);
and U4885 (N_4885,N_4701,N_4622);
and U4886 (N_4886,N_4626,N_4765);
nand U4887 (N_4887,N_4655,N_4681);
nor U4888 (N_4888,N_4668,N_4699);
xnor U4889 (N_4889,N_4697,N_4661);
and U4890 (N_4890,N_4772,N_4610);
xor U4891 (N_4891,N_4602,N_4669);
or U4892 (N_4892,N_4780,N_4755);
or U4893 (N_4893,N_4611,N_4770);
nor U4894 (N_4894,N_4603,N_4633);
nand U4895 (N_4895,N_4756,N_4652);
nor U4896 (N_4896,N_4720,N_4618);
nand U4897 (N_4897,N_4796,N_4709);
and U4898 (N_4898,N_4788,N_4700);
or U4899 (N_4899,N_4702,N_4685);
xor U4900 (N_4900,N_4733,N_4632);
nor U4901 (N_4901,N_4684,N_4643);
xnor U4902 (N_4902,N_4610,N_4684);
and U4903 (N_4903,N_4753,N_4674);
nand U4904 (N_4904,N_4708,N_4629);
nor U4905 (N_4905,N_4795,N_4719);
and U4906 (N_4906,N_4622,N_4717);
or U4907 (N_4907,N_4722,N_4678);
nor U4908 (N_4908,N_4708,N_4706);
nor U4909 (N_4909,N_4624,N_4714);
or U4910 (N_4910,N_4628,N_4618);
and U4911 (N_4911,N_4733,N_4762);
and U4912 (N_4912,N_4768,N_4611);
nand U4913 (N_4913,N_4732,N_4718);
nand U4914 (N_4914,N_4799,N_4776);
nand U4915 (N_4915,N_4799,N_4740);
nand U4916 (N_4916,N_4660,N_4651);
nor U4917 (N_4917,N_4669,N_4651);
nor U4918 (N_4918,N_4777,N_4792);
nor U4919 (N_4919,N_4735,N_4640);
nor U4920 (N_4920,N_4600,N_4761);
or U4921 (N_4921,N_4722,N_4683);
nor U4922 (N_4922,N_4677,N_4765);
nor U4923 (N_4923,N_4765,N_4699);
nor U4924 (N_4924,N_4629,N_4649);
xnor U4925 (N_4925,N_4644,N_4711);
and U4926 (N_4926,N_4700,N_4793);
and U4927 (N_4927,N_4702,N_4692);
and U4928 (N_4928,N_4687,N_4713);
or U4929 (N_4929,N_4794,N_4792);
nand U4930 (N_4930,N_4702,N_4785);
or U4931 (N_4931,N_4755,N_4620);
or U4932 (N_4932,N_4793,N_4772);
nand U4933 (N_4933,N_4779,N_4643);
nor U4934 (N_4934,N_4624,N_4611);
nor U4935 (N_4935,N_4737,N_4610);
nor U4936 (N_4936,N_4626,N_4753);
and U4937 (N_4937,N_4791,N_4723);
nand U4938 (N_4938,N_4740,N_4745);
or U4939 (N_4939,N_4779,N_4765);
xor U4940 (N_4940,N_4670,N_4731);
or U4941 (N_4941,N_4623,N_4783);
or U4942 (N_4942,N_4631,N_4751);
or U4943 (N_4943,N_4711,N_4635);
nand U4944 (N_4944,N_4665,N_4603);
nand U4945 (N_4945,N_4613,N_4760);
nand U4946 (N_4946,N_4680,N_4646);
nor U4947 (N_4947,N_4620,N_4677);
xor U4948 (N_4948,N_4669,N_4680);
and U4949 (N_4949,N_4764,N_4696);
or U4950 (N_4950,N_4658,N_4646);
or U4951 (N_4951,N_4757,N_4622);
nand U4952 (N_4952,N_4703,N_4684);
and U4953 (N_4953,N_4721,N_4739);
and U4954 (N_4954,N_4716,N_4666);
nor U4955 (N_4955,N_4660,N_4716);
or U4956 (N_4956,N_4718,N_4742);
nand U4957 (N_4957,N_4666,N_4625);
nor U4958 (N_4958,N_4686,N_4790);
nor U4959 (N_4959,N_4790,N_4754);
or U4960 (N_4960,N_4666,N_4657);
or U4961 (N_4961,N_4784,N_4603);
nor U4962 (N_4962,N_4688,N_4746);
or U4963 (N_4963,N_4778,N_4767);
nand U4964 (N_4964,N_4725,N_4767);
nor U4965 (N_4965,N_4789,N_4604);
and U4966 (N_4966,N_4724,N_4764);
nand U4967 (N_4967,N_4797,N_4628);
or U4968 (N_4968,N_4779,N_4731);
or U4969 (N_4969,N_4602,N_4769);
nand U4970 (N_4970,N_4798,N_4748);
nor U4971 (N_4971,N_4764,N_4645);
or U4972 (N_4972,N_4727,N_4638);
and U4973 (N_4973,N_4774,N_4678);
nand U4974 (N_4974,N_4603,N_4664);
or U4975 (N_4975,N_4626,N_4787);
nor U4976 (N_4976,N_4634,N_4747);
nand U4977 (N_4977,N_4604,N_4620);
nand U4978 (N_4978,N_4645,N_4652);
nor U4979 (N_4979,N_4796,N_4739);
xnor U4980 (N_4980,N_4664,N_4769);
and U4981 (N_4981,N_4754,N_4640);
nand U4982 (N_4982,N_4647,N_4640);
or U4983 (N_4983,N_4756,N_4605);
or U4984 (N_4984,N_4682,N_4658);
nor U4985 (N_4985,N_4794,N_4719);
or U4986 (N_4986,N_4709,N_4725);
and U4987 (N_4987,N_4755,N_4630);
or U4988 (N_4988,N_4730,N_4692);
and U4989 (N_4989,N_4690,N_4767);
or U4990 (N_4990,N_4647,N_4659);
nor U4991 (N_4991,N_4610,N_4649);
and U4992 (N_4992,N_4687,N_4702);
nand U4993 (N_4993,N_4786,N_4772);
and U4994 (N_4994,N_4621,N_4674);
and U4995 (N_4995,N_4622,N_4697);
or U4996 (N_4996,N_4678,N_4641);
nor U4997 (N_4997,N_4665,N_4680);
xnor U4998 (N_4998,N_4640,N_4714);
and U4999 (N_4999,N_4644,N_4640);
xor UO_0 (O_0,N_4967,N_4943);
nor UO_1 (O_1,N_4824,N_4997);
and UO_2 (O_2,N_4843,N_4882);
and UO_3 (O_3,N_4945,N_4984);
or UO_4 (O_4,N_4926,N_4925);
nand UO_5 (O_5,N_4807,N_4937);
or UO_6 (O_6,N_4877,N_4863);
xnor UO_7 (O_7,N_4973,N_4914);
nand UO_8 (O_8,N_4846,N_4944);
nor UO_9 (O_9,N_4961,N_4855);
and UO_10 (O_10,N_4930,N_4959);
nor UO_11 (O_11,N_4848,N_4902);
nor UO_12 (O_12,N_4886,N_4871);
and UO_13 (O_13,N_4983,N_4819);
and UO_14 (O_14,N_4890,N_4918);
nor UO_15 (O_15,N_4903,N_4999);
nand UO_16 (O_16,N_4935,N_4951);
nand UO_17 (O_17,N_4936,N_4852);
nand UO_18 (O_18,N_4904,N_4895);
nor UO_19 (O_19,N_4899,N_4847);
nand UO_20 (O_20,N_4979,N_4956);
nor UO_21 (O_21,N_4885,N_4911);
and UO_22 (O_22,N_4953,N_4927);
or UO_23 (O_23,N_4928,N_4978);
nand UO_24 (O_24,N_4864,N_4804);
nand UO_25 (O_25,N_4907,N_4962);
xnor UO_26 (O_26,N_4866,N_4809);
and UO_27 (O_27,N_4958,N_4888);
and UO_28 (O_28,N_4872,N_4805);
nor UO_29 (O_29,N_4988,N_4875);
xor UO_30 (O_30,N_4938,N_4917);
or UO_31 (O_31,N_4876,N_4830);
and UO_32 (O_32,N_4870,N_4835);
and UO_33 (O_33,N_4832,N_4822);
nand UO_34 (O_34,N_4892,N_4836);
nand UO_35 (O_35,N_4932,N_4933);
xor UO_36 (O_36,N_4985,N_4839);
nor UO_37 (O_37,N_4982,N_4976);
and UO_38 (O_38,N_4874,N_4996);
nor UO_39 (O_39,N_4901,N_4981);
nor UO_40 (O_40,N_4906,N_4849);
nand UO_41 (O_41,N_4919,N_4905);
and UO_42 (O_42,N_4861,N_4912);
nand UO_43 (O_43,N_4869,N_4811);
xor UO_44 (O_44,N_4854,N_4980);
and UO_45 (O_45,N_4820,N_4994);
and UO_46 (O_46,N_4970,N_4896);
nor UO_47 (O_47,N_4841,N_4858);
nor UO_48 (O_48,N_4884,N_4845);
or UO_49 (O_49,N_4891,N_4887);
and UO_50 (O_50,N_4987,N_4860);
or UO_51 (O_51,N_4881,N_4964);
or UO_52 (O_52,N_4800,N_4837);
nor UO_53 (O_53,N_4810,N_4920);
nor UO_54 (O_54,N_4900,N_4816);
nor UO_55 (O_55,N_4868,N_4921);
and UO_56 (O_56,N_4878,N_4865);
or UO_57 (O_57,N_4812,N_4850);
nor UO_58 (O_58,N_4889,N_4802);
or UO_59 (O_59,N_4814,N_4828);
or UO_60 (O_60,N_4898,N_4826);
or UO_61 (O_61,N_4894,N_4965);
and UO_62 (O_62,N_4989,N_4946);
and UO_63 (O_63,N_4853,N_4813);
nand UO_64 (O_64,N_4977,N_4823);
xor UO_65 (O_65,N_4992,N_4833);
nand UO_66 (O_66,N_4924,N_4908);
and UO_67 (O_67,N_4842,N_4838);
or UO_68 (O_68,N_4829,N_4954);
nor UO_69 (O_69,N_4806,N_4840);
nor UO_70 (O_70,N_4952,N_4949);
or UO_71 (O_71,N_4915,N_4880);
nand UO_72 (O_72,N_4960,N_4942);
nand UO_73 (O_73,N_4986,N_4897);
nor UO_74 (O_74,N_4966,N_4883);
nor UO_75 (O_75,N_4859,N_4940);
or UO_76 (O_76,N_4939,N_4815);
nor UO_77 (O_77,N_4975,N_4818);
xor UO_78 (O_78,N_4947,N_4929);
and UO_79 (O_79,N_4963,N_4873);
or UO_80 (O_80,N_4856,N_4957);
nand UO_81 (O_81,N_4827,N_4893);
and UO_82 (O_82,N_4916,N_4834);
nand UO_83 (O_83,N_4851,N_4968);
or UO_84 (O_84,N_4879,N_4995);
nor UO_85 (O_85,N_4910,N_4990);
and UO_86 (O_86,N_4998,N_4934);
and UO_87 (O_87,N_4825,N_4801);
and UO_88 (O_88,N_4972,N_4913);
nor UO_89 (O_89,N_4971,N_4931);
nor UO_90 (O_90,N_4991,N_4922);
nor UO_91 (O_91,N_4974,N_4948);
or UO_92 (O_92,N_4844,N_4862);
xnor UO_93 (O_93,N_4831,N_4857);
nor UO_94 (O_94,N_4969,N_4803);
nor UO_95 (O_95,N_4941,N_4923);
xor UO_96 (O_96,N_4955,N_4821);
or UO_97 (O_97,N_4867,N_4950);
nand UO_98 (O_98,N_4993,N_4909);
and UO_99 (O_99,N_4808,N_4817);
or UO_100 (O_100,N_4909,N_4834);
nor UO_101 (O_101,N_4873,N_4976);
and UO_102 (O_102,N_4815,N_4857);
xnor UO_103 (O_103,N_4952,N_4808);
nand UO_104 (O_104,N_4994,N_4812);
nor UO_105 (O_105,N_4968,N_4913);
and UO_106 (O_106,N_4866,N_4974);
nand UO_107 (O_107,N_4907,N_4845);
or UO_108 (O_108,N_4923,N_4860);
nor UO_109 (O_109,N_4821,N_4891);
and UO_110 (O_110,N_4852,N_4820);
and UO_111 (O_111,N_4966,N_4928);
and UO_112 (O_112,N_4955,N_4888);
nand UO_113 (O_113,N_4997,N_4899);
nor UO_114 (O_114,N_4855,N_4809);
nand UO_115 (O_115,N_4842,N_4856);
or UO_116 (O_116,N_4887,N_4883);
nand UO_117 (O_117,N_4938,N_4965);
nand UO_118 (O_118,N_4864,N_4961);
nand UO_119 (O_119,N_4851,N_4974);
nand UO_120 (O_120,N_4931,N_4870);
nand UO_121 (O_121,N_4995,N_4965);
and UO_122 (O_122,N_4847,N_4967);
nand UO_123 (O_123,N_4921,N_4950);
nand UO_124 (O_124,N_4891,N_4858);
or UO_125 (O_125,N_4968,N_4856);
and UO_126 (O_126,N_4824,N_4863);
xor UO_127 (O_127,N_4875,N_4879);
nor UO_128 (O_128,N_4965,N_4823);
or UO_129 (O_129,N_4969,N_4962);
or UO_130 (O_130,N_4976,N_4838);
or UO_131 (O_131,N_4833,N_4814);
and UO_132 (O_132,N_4963,N_4879);
nand UO_133 (O_133,N_4974,N_4847);
and UO_134 (O_134,N_4927,N_4923);
nor UO_135 (O_135,N_4803,N_4936);
or UO_136 (O_136,N_4962,N_4924);
nand UO_137 (O_137,N_4911,N_4877);
nor UO_138 (O_138,N_4986,N_4858);
nor UO_139 (O_139,N_4874,N_4901);
nor UO_140 (O_140,N_4986,N_4971);
and UO_141 (O_141,N_4964,N_4996);
and UO_142 (O_142,N_4917,N_4811);
nor UO_143 (O_143,N_4806,N_4926);
nand UO_144 (O_144,N_4903,N_4927);
xor UO_145 (O_145,N_4864,N_4955);
and UO_146 (O_146,N_4814,N_4870);
nand UO_147 (O_147,N_4815,N_4810);
xnor UO_148 (O_148,N_4989,N_4970);
xor UO_149 (O_149,N_4980,N_4816);
or UO_150 (O_150,N_4837,N_4982);
nand UO_151 (O_151,N_4941,N_4979);
nor UO_152 (O_152,N_4809,N_4946);
and UO_153 (O_153,N_4995,N_4888);
xnor UO_154 (O_154,N_4895,N_4805);
or UO_155 (O_155,N_4849,N_4925);
nor UO_156 (O_156,N_4970,N_4890);
or UO_157 (O_157,N_4893,N_4803);
and UO_158 (O_158,N_4853,N_4931);
or UO_159 (O_159,N_4830,N_4833);
nor UO_160 (O_160,N_4886,N_4957);
xor UO_161 (O_161,N_4809,N_4898);
and UO_162 (O_162,N_4891,N_4915);
xnor UO_163 (O_163,N_4916,N_4838);
and UO_164 (O_164,N_4823,N_4839);
nor UO_165 (O_165,N_4883,N_4825);
nor UO_166 (O_166,N_4998,N_4844);
nor UO_167 (O_167,N_4810,N_4936);
nand UO_168 (O_168,N_4903,N_4936);
nand UO_169 (O_169,N_4963,N_4938);
nor UO_170 (O_170,N_4870,N_4810);
and UO_171 (O_171,N_4862,N_4951);
nor UO_172 (O_172,N_4824,N_4994);
and UO_173 (O_173,N_4947,N_4996);
xnor UO_174 (O_174,N_4922,N_4846);
nand UO_175 (O_175,N_4900,N_4832);
nand UO_176 (O_176,N_4901,N_4974);
nor UO_177 (O_177,N_4846,N_4984);
nor UO_178 (O_178,N_4909,N_4817);
and UO_179 (O_179,N_4984,N_4832);
xnor UO_180 (O_180,N_4860,N_4916);
or UO_181 (O_181,N_4808,N_4970);
nor UO_182 (O_182,N_4842,N_4972);
nand UO_183 (O_183,N_4886,N_4863);
and UO_184 (O_184,N_4897,N_4805);
nor UO_185 (O_185,N_4948,N_4916);
and UO_186 (O_186,N_4998,N_4856);
or UO_187 (O_187,N_4882,N_4903);
nand UO_188 (O_188,N_4934,N_4875);
nor UO_189 (O_189,N_4984,N_4861);
nor UO_190 (O_190,N_4957,N_4942);
or UO_191 (O_191,N_4897,N_4987);
nor UO_192 (O_192,N_4842,N_4872);
nor UO_193 (O_193,N_4971,N_4845);
xnor UO_194 (O_194,N_4903,N_4833);
and UO_195 (O_195,N_4968,N_4843);
nand UO_196 (O_196,N_4904,N_4983);
nor UO_197 (O_197,N_4886,N_4937);
nor UO_198 (O_198,N_4810,N_4833);
or UO_199 (O_199,N_4811,N_4882);
xnor UO_200 (O_200,N_4899,N_4817);
or UO_201 (O_201,N_4995,N_4822);
or UO_202 (O_202,N_4837,N_4971);
or UO_203 (O_203,N_4930,N_4944);
xnor UO_204 (O_204,N_4800,N_4977);
nand UO_205 (O_205,N_4841,N_4979);
nor UO_206 (O_206,N_4867,N_4804);
or UO_207 (O_207,N_4879,N_4870);
nor UO_208 (O_208,N_4998,N_4897);
nand UO_209 (O_209,N_4820,N_4807);
xor UO_210 (O_210,N_4863,N_4888);
nor UO_211 (O_211,N_4897,N_4965);
and UO_212 (O_212,N_4904,N_4951);
nand UO_213 (O_213,N_4867,N_4872);
xor UO_214 (O_214,N_4823,N_4858);
nor UO_215 (O_215,N_4907,N_4975);
and UO_216 (O_216,N_4903,N_4830);
nor UO_217 (O_217,N_4830,N_4806);
nor UO_218 (O_218,N_4933,N_4858);
nand UO_219 (O_219,N_4876,N_4838);
and UO_220 (O_220,N_4883,N_4913);
xnor UO_221 (O_221,N_4962,N_4954);
and UO_222 (O_222,N_4835,N_4810);
and UO_223 (O_223,N_4861,N_4948);
xnor UO_224 (O_224,N_4986,N_4956);
or UO_225 (O_225,N_4865,N_4805);
nor UO_226 (O_226,N_4894,N_4930);
or UO_227 (O_227,N_4988,N_4940);
nor UO_228 (O_228,N_4802,N_4946);
and UO_229 (O_229,N_4823,N_4828);
nor UO_230 (O_230,N_4888,N_4933);
or UO_231 (O_231,N_4935,N_4854);
nor UO_232 (O_232,N_4964,N_4814);
and UO_233 (O_233,N_4826,N_4922);
nand UO_234 (O_234,N_4893,N_4906);
and UO_235 (O_235,N_4985,N_4901);
and UO_236 (O_236,N_4839,N_4931);
and UO_237 (O_237,N_4872,N_4917);
or UO_238 (O_238,N_4901,N_4890);
nor UO_239 (O_239,N_4826,N_4841);
and UO_240 (O_240,N_4961,N_4993);
and UO_241 (O_241,N_4967,N_4834);
and UO_242 (O_242,N_4800,N_4852);
or UO_243 (O_243,N_4965,N_4943);
and UO_244 (O_244,N_4926,N_4939);
nand UO_245 (O_245,N_4871,N_4926);
or UO_246 (O_246,N_4853,N_4997);
xnor UO_247 (O_247,N_4900,N_4888);
nor UO_248 (O_248,N_4981,N_4894);
and UO_249 (O_249,N_4992,N_4960);
or UO_250 (O_250,N_4854,N_4890);
or UO_251 (O_251,N_4900,N_4826);
and UO_252 (O_252,N_4997,N_4925);
nand UO_253 (O_253,N_4936,N_4854);
nand UO_254 (O_254,N_4976,N_4912);
or UO_255 (O_255,N_4855,N_4861);
nor UO_256 (O_256,N_4820,N_4822);
nand UO_257 (O_257,N_4872,N_4839);
nor UO_258 (O_258,N_4813,N_4807);
xor UO_259 (O_259,N_4811,N_4876);
and UO_260 (O_260,N_4891,N_4810);
and UO_261 (O_261,N_4849,N_4911);
or UO_262 (O_262,N_4922,N_4880);
nor UO_263 (O_263,N_4970,N_4957);
nor UO_264 (O_264,N_4890,N_4947);
and UO_265 (O_265,N_4813,N_4859);
or UO_266 (O_266,N_4892,N_4923);
nor UO_267 (O_267,N_4843,N_4899);
nand UO_268 (O_268,N_4962,N_4930);
nor UO_269 (O_269,N_4830,N_4993);
nand UO_270 (O_270,N_4906,N_4978);
and UO_271 (O_271,N_4875,N_4999);
or UO_272 (O_272,N_4859,N_4983);
and UO_273 (O_273,N_4943,N_4955);
nand UO_274 (O_274,N_4989,N_4969);
and UO_275 (O_275,N_4992,N_4834);
or UO_276 (O_276,N_4832,N_4853);
and UO_277 (O_277,N_4974,N_4919);
and UO_278 (O_278,N_4928,N_4991);
nor UO_279 (O_279,N_4800,N_4897);
nor UO_280 (O_280,N_4962,N_4856);
xnor UO_281 (O_281,N_4895,N_4994);
nand UO_282 (O_282,N_4949,N_4946);
nand UO_283 (O_283,N_4872,N_4968);
or UO_284 (O_284,N_4840,N_4990);
nand UO_285 (O_285,N_4809,N_4863);
nand UO_286 (O_286,N_4832,N_4978);
nor UO_287 (O_287,N_4974,N_4909);
nor UO_288 (O_288,N_4923,N_4969);
nand UO_289 (O_289,N_4937,N_4890);
nand UO_290 (O_290,N_4961,N_4962);
or UO_291 (O_291,N_4860,N_4935);
nand UO_292 (O_292,N_4876,N_4849);
nand UO_293 (O_293,N_4875,N_4994);
nor UO_294 (O_294,N_4955,N_4930);
nand UO_295 (O_295,N_4945,N_4859);
and UO_296 (O_296,N_4992,N_4874);
and UO_297 (O_297,N_4801,N_4836);
nor UO_298 (O_298,N_4802,N_4920);
and UO_299 (O_299,N_4979,N_4900);
nand UO_300 (O_300,N_4987,N_4979);
nor UO_301 (O_301,N_4958,N_4858);
or UO_302 (O_302,N_4952,N_4855);
or UO_303 (O_303,N_4825,N_4925);
nand UO_304 (O_304,N_4900,N_4848);
and UO_305 (O_305,N_4995,N_4932);
and UO_306 (O_306,N_4930,N_4983);
nor UO_307 (O_307,N_4982,N_4862);
and UO_308 (O_308,N_4963,N_4916);
or UO_309 (O_309,N_4804,N_4933);
and UO_310 (O_310,N_4895,N_4970);
and UO_311 (O_311,N_4806,N_4894);
xor UO_312 (O_312,N_4959,N_4859);
and UO_313 (O_313,N_4972,N_4814);
nor UO_314 (O_314,N_4877,N_4997);
and UO_315 (O_315,N_4864,N_4968);
and UO_316 (O_316,N_4844,N_4996);
nor UO_317 (O_317,N_4946,N_4863);
nand UO_318 (O_318,N_4978,N_4877);
nor UO_319 (O_319,N_4960,N_4905);
nand UO_320 (O_320,N_4825,N_4870);
xor UO_321 (O_321,N_4859,N_4846);
or UO_322 (O_322,N_4942,N_4883);
xor UO_323 (O_323,N_4874,N_4938);
or UO_324 (O_324,N_4930,N_4829);
nand UO_325 (O_325,N_4978,N_4887);
nand UO_326 (O_326,N_4909,N_4803);
and UO_327 (O_327,N_4987,N_4831);
nor UO_328 (O_328,N_4925,N_4842);
nand UO_329 (O_329,N_4894,N_4922);
nand UO_330 (O_330,N_4849,N_4963);
nand UO_331 (O_331,N_4849,N_4856);
and UO_332 (O_332,N_4838,N_4975);
or UO_333 (O_333,N_4981,N_4861);
nor UO_334 (O_334,N_4803,N_4821);
or UO_335 (O_335,N_4823,N_4833);
nand UO_336 (O_336,N_4979,N_4869);
nor UO_337 (O_337,N_4958,N_4980);
and UO_338 (O_338,N_4962,N_4863);
and UO_339 (O_339,N_4940,N_4854);
or UO_340 (O_340,N_4842,N_4991);
nor UO_341 (O_341,N_4979,N_4920);
or UO_342 (O_342,N_4871,N_4969);
or UO_343 (O_343,N_4899,N_4928);
nand UO_344 (O_344,N_4814,N_4861);
xnor UO_345 (O_345,N_4873,N_4821);
nor UO_346 (O_346,N_4983,N_4801);
and UO_347 (O_347,N_4826,N_4849);
and UO_348 (O_348,N_4891,N_4888);
xnor UO_349 (O_349,N_4942,N_4866);
and UO_350 (O_350,N_4926,N_4969);
and UO_351 (O_351,N_4812,N_4857);
nand UO_352 (O_352,N_4945,N_4822);
or UO_353 (O_353,N_4802,N_4854);
nand UO_354 (O_354,N_4919,N_4941);
nand UO_355 (O_355,N_4803,N_4884);
and UO_356 (O_356,N_4937,N_4875);
nor UO_357 (O_357,N_4881,N_4907);
or UO_358 (O_358,N_4830,N_4842);
or UO_359 (O_359,N_4837,N_4929);
and UO_360 (O_360,N_4919,N_4928);
nand UO_361 (O_361,N_4884,N_4949);
nand UO_362 (O_362,N_4862,N_4899);
and UO_363 (O_363,N_4830,N_4868);
or UO_364 (O_364,N_4864,N_4869);
nor UO_365 (O_365,N_4915,N_4916);
nor UO_366 (O_366,N_4922,N_4924);
or UO_367 (O_367,N_4978,N_4837);
and UO_368 (O_368,N_4807,N_4837);
xnor UO_369 (O_369,N_4818,N_4991);
nand UO_370 (O_370,N_4938,N_4823);
nor UO_371 (O_371,N_4949,N_4983);
nor UO_372 (O_372,N_4882,N_4961);
and UO_373 (O_373,N_4991,N_4921);
nor UO_374 (O_374,N_4850,N_4918);
or UO_375 (O_375,N_4979,N_4977);
nand UO_376 (O_376,N_4804,N_4848);
nor UO_377 (O_377,N_4972,N_4937);
xor UO_378 (O_378,N_4956,N_4910);
nor UO_379 (O_379,N_4938,N_4831);
nand UO_380 (O_380,N_4913,N_4805);
nor UO_381 (O_381,N_4953,N_4919);
nand UO_382 (O_382,N_4920,N_4847);
nand UO_383 (O_383,N_4960,N_4943);
or UO_384 (O_384,N_4856,N_4971);
nand UO_385 (O_385,N_4945,N_4957);
or UO_386 (O_386,N_4890,N_4823);
nand UO_387 (O_387,N_4958,N_4931);
xnor UO_388 (O_388,N_4812,N_4879);
nor UO_389 (O_389,N_4913,N_4956);
nor UO_390 (O_390,N_4935,N_4912);
and UO_391 (O_391,N_4924,N_4875);
or UO_392 (O_392,N_4815,N_4968);
and UO_393 (O_393,N_4897,N_4990);
nor UO_394 (O_394,N_4976,N_4833);
and UO_395 (O_395,N_4891,N_4959);
and UO_396 (O_396,N_4814,N_4869);
or UO_397 (O_397,N_4851,N_4915);
nand UO_398 (O_398,N_4862,N_4969);
nand UO_399 (O_399,N_4870,N_4846);
nand UO_400 (O_400,N_4861,N_4980);
and UO_401 (O_401,N_4966,N_4821);
or UO_402 (O_402,N_4947,N_4927);
nor UO_403 (O_403,N_4912,N_4872);
nand UO_404 (O_404,N_4813,N_4842);
or UO_405 (O_405,N_4850,N_4974);
xor UO_406 (O_406,N_4856,N_4834);
and UO_407 (O_407,N_4939,N_4992);
and UO_408 (O_408,N_4821,N_4836);
or UO_409 (O_409,N_4906,N_4819);
or UO_410 (O_410,N_4895,N_4984);
and UO_411 (O_411,N_4856,N_4843);
or UO_412 (O_412,N_4991,N_4876);
and UO_413 (O_413,N_4881,N_4805);
or UO_414 (O_414,N_4995,N_4952);
nor UO_415 (O_415,N_4865,N_4942);
nor UO_416 (O_416,N_4828,N_4839);
xnor UO_417 (O_417,N_4823,N_4816);
or UO_418 (O_418,N_4844,N_4854);
xnor UO_419 (O_419,N_4973,N_4870);
nor UO_420 (O_420,N_4987,N_4810);
nor UO_421 (O_421,N_4856,N_4930);
or UO_422 (O_422,N_4950,N_4808);
nand UO_423 (O_423,N_4805,N_4894);
nand UO_424 (O_424,N_4995,N_4999);
xor UO_425 (O_425,N_4820,N_4984);
nand UO_426 (O_426,N_4968,N_4966);
nand UO_427 (O_427,N_4849,N_4894);
or UO_428 (O_428,N_4821,N_4972);
and UO_429 (O_429,N_4817,N_4923);
and UO_430 (O_430,N_4991,N_4838);
and UO_431 (O_431,N_4978,N_4854);
xor UO_432 (O_432,N_4908,N_4934);
or UO_433 (O_433,N_4955,N_4896);
nor UO_434 (O_434,N_4831,N_4825);
or UO_435 (O_435,N_4813,N_4829);
nor UO_436 (O_436,N_4988,N_4841);
or UO_437 (O_437,N_4939,N_4906);
nand UO_438 (O_438,N_4935,N_4888);
or UO_439 (O_439,N_4951,N_4873);
xnor UO_440 (O_440,N_4861,N_4830);
nand UO_441 (O_441,N_4834,N_4948);
nor UO_442 (O_442,N_4987,N_4963);
nand UO_443 (O_443,N_4984,N_4998);
nor UO_444 (O_444,N_4974,N_4913);
nand UO_445 (O_445,N_4866,N_4963);
or UO_446 (O_446,N_4925,N_4906);
or UO_447 (O_447,N_4861,N_4964);
or UO_448 (O_448,N_4813,N_4993);
xor UO_449 (O_449,N_4948,N_4901);
nor UO_450 (O_450,N_4870,N_4889);
or UO_451 (O_451,N_4819,N_4982);
nor UO_452 (O_452,N_4811,N_4814);
or UO_453 (O_453,N_4928,N_4874);
nand UO_454 (O_454,N_4912,N_4822);
nand UO_455 (O_455,N_4995,N_4982);
xor UO_456 (O_456,N_4868,N_4904);
nor UO_457 (O_457,N_4871,N_4991);
and UO_458 (O_458,N_4910,N_4906);
nor UO_459 (O_459,N_4943,N_4818);
or UO_460 (O_460,N_4874,N_4998);
or UO_461 (O_461,N_4857,N_4892);
xnor UO_462 (O_462,N_4866,N_4957);
or UO_463 (O_463,N_4818,N_4928);
or UO_464 (O_464,N_4993,N_4846);
and UO_465 (O_465,N_4939,N_4919);
and UO_466 (O_466,N_4923,N_4862);
or UO_467 (O_467,N_4992,N_4843);
and UO_468 (O_468,N_4874,N_4840);
nor UO_469 (O_469,N_4989,N_4959);
or UO_470 (O_470,N_4891,N_4843);
or UO_471 (O_471,N_4964,N_4813);
xnor UO_472 (O_472,N_4897,N_4924);
and UO_473 (O_473,N_4966,N_4960);
or UO_474 (O_474,N_4986,N_4952);
or UO_475 (O_475,N_4927,N_4875);
nand UO_476 (O_476,N_4860,N_4848);
nand UO_477 (O_477,N_4827,N_4881);
nor UO_478 (O_478,N_4842,N_4877);
nor UO_479 (O_479,N_4936,N_4818);
and UO_480 (O_480,N_4844,N_4926);
or UO_481 (O_481,N_4904,N_4806);
nor UO_482 (O_482,N_4815,N_4825);
and UO_483 (O_483,N_4914,N_4830);
nor UO_484 (O_484,N_4942,N_4982);
or UO_485 (O_485,N_4813,N_4987);
nor UO_486 (O_486,N_4809,N_4864);
xnor UO_487 (O_487,N_4864,N_4997);
nor UO_488 (O_488,N_4800,N_4956);
nor UO_489 (O_489,N_4920,N_4874);
or UO_490 (O_490,N_4996,N_4925);
nand UO_491 (O_491,N_4941,N_4930);
nor UO_492 (O_492,N_4924,N_4991);
nand UO_493 (O_493,N_4813,N_4906);
and UO_494 (O_494,N_4842,N_4839);
nor UO_495 (O_495,N_4935,N_4954);
nand UO_496 (O_496,N_4853,N_4968);
or UO_497 (O_497,N_4923,N_4844);
or UO_498 (O_498,N_4851,N_4864);
or UO_499 (O_499,N_4869,N_4809);
or UO_500 (O_500,N_4813,N_4983);
nor UO_501 (O_501,N_4857,N_4969);
nor UO_502 (O_502,N_4835,N_4965);
or UO_503 (O_503,N_4955,N_4945);
nand UO_504 (O_504,N_4834,N_4924);
nor UO_505 (O_505,N_4860,N_4823);
and UO_506 (O_506,N_4921,N_4941);
nor UO_507 (O_507,N_4845,N_4978);
and UO_508 (O_508,N_4975,N_4895);
and UO_509 (O_509,N_4823,N_4966);
or UO_510 (O_510,N_4898,N_4862);
nor UO_511 (O_511,N_4857,N_4961);
nor UO_512 (O_512,N_4863,N_4844);
nand UO_513 (O_513,N_4908,N_4916);
nor UO_514 (O_514,N_4836,N_4904);
and UO_515 (O_515,N_4863,N_4949);
nand UO_516 (O_516,N_4967,N_4878);
and UO_517 (O_517,N_4882,N_4973);
nor UO_518 (O_518,N_4859,N_4982);
nand UO_519 (O_519,N_4803,N_4840);
or UO_520 (O_520,N_4824,N_4920);
or UO_521 (O_521,N_4993,N_4900);
nor UO_522 (O_522,N_4883,N_4837);
or UO_523 (O_523,N_4990,N_4944);
nor UO_524 (O_524,N_4918,N_4971);
and UO_525 (O_525,N_4879,N_4933);
or UO_526 (O_526,N_4870,N_4878);
and UO_527 (O_527,N_4919,N_4891);
nand UO_528 (O_528,N_4819,N_4813);
or UO_529 (O_529,N_4977,N_4860);
nand UO_530 (O_530,N_4800,N_4935);
nand UO_531 (O_531,N_4972,N_4859);
nand UO_532 (O_532,N_4938,N_4934);
or UO_533 (O_533,N_4923,N_4830);
nand UO_534 (O_534,N_4935,N_4891);
nor UO_535 (O_535,N_4820,N_4800);
or UO_536 (O_536,N_4942,N_4886);
nand UO_537 (O_537,N_4803,N_4812);
and UO_538 (O_538,N_4840,N_4932);
nand UO_539 (O_539,N_4940,N_4862);
nor UO_540 (O_540,N_4915,N_4976);
and UO_541 (O_541,N_4957,N_4824);
nand UO_542 (O_542,N_4942,N_4933);
nor UO_543 (O_543,N_4935,N_4852);
and UO_544 (O_544,N_4889,N_4916);
and UO_545 (O_545,N_4922,N_4942);
and UO_546 (O_546,N_4967,N_4970);
and UO_547 (O_547,N_4852,N_4905);
nand UO_548 (O_548,N_4848,N_4820);
and UO_549 (O_549,N_4863,N_4994);
nand UO_550 (O_550,N_4856,N_4950);
and UO_551 (O_551,N_4845,N_4901);
nor UO_552 (O_552,N_4963,N_4966);
xnor UO_553 (O_553,N_4891,N_4809);
or UO_554 (O_554,N_4849,N_4863);
or UO_555 (O_555,N_4849,N_4824);
nor UO_556 (O_556,N_4961,N_4833);
nor UO_557 (O_557,N_4888,N_4823);
or UO_558 (O_558,N_4882,N_4850);
nand UO_559 (O_559,N_4937,N_4936);
nor UO_560 (O_560,N_4997,N_4866);
and UO_561 (O_561,N_4870,N_4983);
or UO_562 (O_562,N_4878,N_4855);
nand UO_563 (O_563,N_4959,N_4988);
or UO_564 (O_564,N_4984,N_4880);
or UO_565 (O_565,N_4818,N_4821);
or UO_566 (O_566,N_4866,N_4972);
nand UO_567 (O_567,N_4926,N_4991);
nand UO_568 (O_568,N_4914,N_4979);
nor UO_569 (O_569,N_4844,N_4879);
and UO_570 (O_570,N_4884,N_4915);
and UO_571 (O_571,N_4925,N_4937);
nand UO_572 (O_572,N_4966,N_4930);
nand UO_573 (O_573,N_4870,N_4996);
and UO_574 (O_574,N_4861,N_4946);
xor UO_575 (O_575,N_4842,N_4814);
nor UO_576 (O_576,N_4966,N_4965);
or UO_577 (O_577,N_4828,N_4816);
or UO_578 (O_578,N_4980,N_4948);
nand UO_579 (O_579,N_4907,N_4949);
or UO_580 (O_580,N_4889,N_4906);
and UO_581 (O_581,N_4980,N_4928);
or UO_582 (O_582,N_4970,N_4899);
or UO_583 (O_583,N_4923,N_4963);
and UO_584 (O_584,N_4882,N_4813);
or UO_585 (O_585,N_4979,N_4846);
nor UO_586 (O_586,N_4807,N_4847);
nand UO_587 (O_587,N_4912,N_4962);
or UO_588 (O_588,N_4838,N_4852);
and UO_589 (O_589,N_4990,N_4992);
nor UO_590 (O_590,N_4986,N_4816);
xor UO_591 (O_591,N_4820,N_4929);
and UO_592 (O_592,N_4921,N_4879);
or UO_593 (O_593,N_4987,N_4967);
and UO_594 (O_594,N_4827,N_4957);
xnor UO_595 (O_595,N_4822,N_4990);
nor UO_596 (O_596,N_4970,N_4994);
nor UO_597 (O_597,N_4967,N_4806);
and UO_598 (O_598,N_4994,N_4835);
nor UO_599 (O_599,N_4945,N_4968);
nand UO_600 (O_600,N_4923,N_4899);
or UO_601 (O_601,N_4956,N_4886);
nand UO_602 (O_602,N_4892,N_4835);
xor UO_603 (O_603,N_4857,N_4856);
and UO_604 (O_604,N_4972,N_4905);
or UO_605 (O_605,N_4859,N_4864);
xnor UO_606 (O_606,N_4866,N_4919);
and UO_607 (O_607,N_4942,N_4912);
or UO_608 (O_608,N_4916,N_4815);
xor UO_609 (O_609,N_4894,N_4832);
nand UO_610 (O_610,N_4972,N_4989);
nand UO_611 (O_611,N_4945,N_4922);
nand UO_612 (O_612,N_4966,N_4851);
nor UO_613 (O_613,N_4824,N_4944);
or UO_614 (O_614,N_4930,N_4854);
and UO_615 (O_615,N_4913,N_4840);
and UO_616 (O_616,N_4923,N_4935);
nor UO_617 (O_617,N_4840,N_4823);
nand UO_618 (O_618,N_4966,N_4879);
and UO_619 (O_619,N_4837,N_4834);
and UO_620 (O_620,N_4957,N_4816);
nand UO_621 (O_621,N_4801,N_4969);
nor UO_622 (O_622,N_4977,N_4987);
or UO_623 (O_623,N_4820,N_4942);
nand UO_624 (O_624,N_4846,N_4836);
nand UO_625 (O_625,N_4862,N_4856);
nor UO_626 (O_626,N_4873,N_4945);
nor UO_627 (O_627,N_4907,N_4854);
xnor UO_628 (O_628,N_4997,N_4990);
nor UO_629 (O_629,N_4835,N_4847);
xor UO_630 (O_630,N_4903,N_4923);
or UO_631 (O_631,N_4998,N_4931);
nand UO_632 (O_632,N_4851,N_4804);
nor UO_633 (O_633,N_4844,N_4987);
and UO_634 (O_634,N_4985,N_4861);
nor UO_635 (O_635,N_4932,N_4953);
nand UO_636 (O_636,N_4995,N_4854);
xnor UO_637 (O_637,N_4982,N_4992);
and UO_638 (O_638,N_4834,N_4805);
or UO_639 (O_639,N_4946,N_4817);
and UO_640 (O_640,N_4990,N_4964);
and UO_641 (O_641,N_4962,N_4919);
nand UO_642 (O_642,N_4900,N_4837);
nand UO_643 (O_643,N_4872,N_4851);
or UO_644 (O_644,N_4847,N_4906);
xor UO_645 (O_645,N_4927,N_4868);
and UO_646 (O_646,N_4889,N_4846);
nor UO_647 (O_647,N_4880,N_4841);
nor UO_648 (O_648,N_4802,N_4848);
xor UO_649 (O_649,N_4876,N_4824);
nand UO_650 (O_650,N_4836,N_4845);
or UO_651 (O_651,N_4984,N_4890);
nand UO_652 (O_652,N_4809,N_4931);
or UO_653 (O_653,N_4841,N_4820);
nor UO_654 (O_654,N_4897,N_4890);
and UO_655 (O_655,N_4822,N_4874);
xor UO_656 (O_656,N_4881,N_4935);
nor UO_657 (O_657,N_4966,N_4972);
xor UO_658 (O_658,N_4985,N_4884);
nor UO_659 (O_659,N_4969,N_4869);
nand UO_660 (O_660,N_4866,N_4826);
nor UO_661 (O_661,N_4987,N_4972);
xor UO_662 (O_662,N_4832,N_4995);
and UO_663 (O_663,N_4916,N_4906);
nor UO_664 (O_664,N_4839,N_4990);
nand UO_665 (O_665,N_4977,N_4968);
nor UO_666 (O_666,N_4866,N_4895);
nand UO_667 (O_667,N_4881,N_4977);
nor UO_668 (O_668,N_4923,N_4884);
or UO_669 (O_669,N_4962,N_4854);
xnor UO_670 (O_670,N_4989,N_4859);
and UO_671 (O_671,N_4986,N_4917);
or UO_672 (O_672,N_4981,N_4938);
nand UO_673 (O_673,N_4859,N_4865);
and UO_674 (O_674,N_4923,N_4824);
nand UO_675 (O_675,N_4936,N_4994);
nor UO_676 (O_676,N_4994,N_4974);
xor UO_677 (O_677,N_4831,N_4884);
or UO_678 (O_678,N_4994,N_4952);
nand UO_679 (O_679,N_4833,N_4840);
nand UO_680 (O_680,N_4903,N_4931);
and UO_681 (O_681,N_4815,N_4921);
and UO_682 (O_682,N_4940,N_4899);
and UO_683 (O_683,N_4890,N_4842);
nand UO_684 (O_684,N_4975,N_4954);
nand UO_685 (O_685,N_4977,N_4826);
xnor UO_686 (O_686,N_4833,N_4996);
nor UO_687 (O_687,N_4817,N_4872);
nor UO_688 (O_688,N_4970,N_4852);
and UO_689 (O_689,N_4859,N_4857);
or UO_690 (O_690,N_4943,N_4904);
nor UO_691 (O_691,N_4914,N_4992);
nand UO_692 (O_692,N_4814,N_4841);
xnor UO_693 (O_693,N_4887,N_4969);
and UO_694 (O_694,N_4977,N_4971);
nand UO_695 (O_695,N_4849,N_4895);
and UO_696 (O_696,N_4946,N_4947);
nor UO_697 (O_697,N_4970,N_4873);
nand UO_698 (O_698,N_4859,N_4887);
nor UO_699 (O_699,N_4948,N_4915);
nand UO_700 (O_700,N_4990,N_4830);
nand UO_701 (O_701,N_4817,N_4950);
nor UO_702 (O_702,N_4954,N_4972);
nor UO_703 (O_703,N_4865,N_4876);
xor UO_704 (O_704,N_4800,N_4995);
nand UO_705 (O_705,N_4898,N_4995);
and UO_706 (O_706,N_4884,N_4812);
or UO_707 (O_707,N_4947,N_4933);
nor UO_708 (O_708,N_4872,N_4860);
or UO_709 (O_709,N_4959,N_4805);
and UO_710 (O_710,N_4875,N_4860);
nand UO_711 (O_711,N_4858,N_4916);
or UO_712 (O_712,N_4915,N_4892);
nor UO_713 (O_713,N_4890,N_4973);
and UO_714 (O_714,N_4982,N_4963);
or UO_715 (O_715,N_4946,N_4834);
or UO_716 (O_716,N_4905,N_4848);
nor UO_717 (O_717,N_4924,N_4894);
nor UO_718 (O_718,N_4877,N_4952);
and UO_719 (O_719,N_4845,N_4841);
or UO_720 (O_720,N_4821,N_4940);
nand UO_721 (O_721,N_4830,N_4875);
or UO_722 (O_722,N_4942,N_4835);
and UO_723 (O_723,N_4986,N_4817);
and UO_724 (O_724,N_4849,N_4973);
and UO_725 (O_725,N_4853,N_4877);
and UO_726 (O_726,N_4886,N_4809);
or UO_727 (O_727,N_4811,N_4985);
or UO_728 (O_728,N_4860,N_4955);
or UO_729 (O_729,N_4868,N_4882);
and UO_730 (O_730,N_4947,N_4935);
or UO_731 (O_731,N_4970,N_4990);
xor UO_732 (O_732,N_4993,N_4907);
and UO_733 (O_733,N_4934,N_4853);
and UO_734 (O_734,N_4831,N_4948);
and UO_735 (O_735,N_4823,N_4972);
and UO_736 (O_736,N_4937,N_4888);
nor UO_737 (O_737,N_4966,N_4991);
and UO_738 (O_738,N_4964,N_4801);
nand UO_739 (O_739,N_4884,N_4956);
or UO_740 (O_740,N_4899,N_4931);
xor UO_741 (O_741,N_4858,N_4844);
or UO_742 (O_742,N_4814,N_4989);
and UO_743 (O_743,N_4831,N_4872);
nand UO_744 (O_744,N_4919,N_4938);
or UO_745 (O_745,N_4993,N_4977);
nor UO_746 (O_746,N_4807,N_4963);
nand UO_747 (O_747,N_4944,N_4901);
and UO_748 (O_748,N_4992,N_4929);
and UO_749 (O_749,N_4948,N_4975);
nand UO_750 (O_750,N_4824,N_4979);
xor UO_751 (O_751,N_4857,N_4862);
or UO_752 (O_752,N_4941,N_4926);
and UO_753 (O_753,N_4825,N_4992);
or UO_754 (O_754,N_4825,N_4881);
nor UO_755 (O_755,N_4825,N_4844);
nand UO_756 (O_756,N_4994,N_4965);
or UO_757 (O_757,N_4989,N_4993);
nor UO_758 (O_758,N_4902,N_4926);
nor UO_759 (O_759,N_4981,N_4930);
or UO_760 (O_760,N_4881,N_4937);
nand UO_761 (O_761,N_4850,N_4898);
and UO_762 (O_762,N_4914,N_4968);
or UO_763 (O_763,N_4870,N_4851);
nand UO_764 (O_764,N_4981,N_4805);
nor UO_765 (O_765,N_4995,N_4825);
nor UO_766 (O_766,N_4911,N_4808);
or UO_767 (O_767,N_4878,N_4871);
and UO_768 (O_768,N_4961,N_4899);
and UO_769 (O_769,N_4928,N_4886);
and UO_770 (O_770,N_4996,N_4913);
nand UO_771 (O_771,N_4913,N_4835);
or UO_772 (O_772,N_4819,N_4889);
and UO_773 (O_773,N_4845,N_4840);
or UO_774 (O_774,N_4977,N_4943);
or UO_775 (O_775,N_4888,N_4875);
nor UO_776 (O_776,N_4995,N_4820);
or UO_777 (O_777,N_4926,N_4965);
or UO_778 (O_778,N_4857,N_4983);
and UO_779 (O_779,N_4985,N_4887);
nand UO_780 (O_780,N_4900,N_4857);
nor UO_781 (O_781,N_4848,N_4984);
nand UO_782 (O_782,N_4914,N_4827);
xor UO_783 (O_783,N_4800,N_4829);
nand UO_784 (O_784,N_4891,N_4844);
or UO_785 (O_785,N_4884,N_4963);
nor UO_786 (O_786,N_4802,N_4835);
nor UO_787 (O_787,N_4888,N_4818);
and UO_788 (O_788,N_4916,N_4930);
nor UO_789 (O_789,N_4891,N_4823);
nand UO_790 (O_790,N_4837,N_4843);
and UO_791 (O_791,N_4958,N_4915);
and UO_792 (O_792,N_4951,N_4852);
or UO_793 (O_793,N_4894,N_4900);
and UO_794 (O_794,N_4955,N_4933);
or UO_795 (O_795,N_4830,N_4949);
and UO_796 (O_796,N_4964,N_4981);
nor UO_797 (O_797,N_4870,N_4856);
or UO_798 (O_798,N_4827,N_4854);
xor UO_799 (O_799,N_4917,N_4976);
nand UO_800 (O_800,N_4951,N_4833);
nor UO_801 (O_801,N_4855,N_4931);
xnor UO_802 (O_802,N_4910,N_4813);
nor UO_803 (O_803,N_4902,N_4991);
or UO_804 (O_804,N_4891,N_4923);
or UO_805 (O_805,N_4998,N_4880);
and UO_806 (O_806,N_4951,N_4914);
and UO_807 (O_807,N_4996,N_4930);
nor UO_808 (O_808,N_4824,N_4961);
or UO_809 (O_809,N_4906,N_4935);
nor UO_810 (O_810,N_4971,N_4821);
and UO_811 (O_811,N_4845,N_4843);
xnor UO_812 (O_812,N_4906,N_4818);
or UO_813 (O_813,N_4905,N_4955);
nor UO_814 (O_814,N_4830,N_4819);
xnor UO_815 (O_815,N_4923,N_4956);
xnor UO_816 (O_816,N_4991,N_4885);
or UO_817 (O_817,N_4895,N_4882);
nand UO_818 (O_818,N_4834,N_4943);
or UO_819 (O_819,N_4825,N_4924);
or UO_820 (O_820,N_4836,N_4810);
or UO_821 (O_821,N_4869,N_4802);
and UO_822 (O_822,N_4822,N_4985);
and UO_823 (O_823,N_4999,N_4973);
nor UO_824 (O_824,N_4999,N_4824);
xnor UO_825 (O_825,N_4856,N_4881);
xnor UO_826 (O_826,N_4962,N_4917);
and UO_827 (O_827,N_4907,N_4825);
and UO_828 (O_828,N_4920,N_4883);
or UO_829 (O_829,N_4932,N_4873);
and UO_830 (O_830,N_4871,N_4977);
nand UO_831 (O_831,N_4922,N_4908);
nand UO_832 (O_832,N_4857,N_4945);
nand UO_833 (O_833,N_4904,N_4808);
and UO_834 (O_834,N_4831,N_4975);
nand UO_835 (O_835,N_4820,N_4876);
or UO_836 (O_836,N_4800,N_4874);
nand UO_837 (O_837,N_4903,N_4981);
or UO_838 (O_838,N_4914,N_4811);
or UO_839 (O_839,N_4823,N_4933);
or UO_840 (O_840,N_4829,N_4907);
nor UO_841 (O_841,N_4866,N_4987);
or UO_842 (O_842,N_4864,N_4974);
nor UO_843 (O_843,N_4856,N_4853);
and UO_844 (O_844,N_4941,N_4933);
nand UO_845 (O_845,N_4897,N_4961);
or UO_846 (O_846,N_4951,N_4851);
nor UO_847 (O_847,N_4940,N_4852);
and UO_848 (O_848,N_4828,N_4937);
and UO_849 (O_849,N_4884,N_4837);
xnor UO_850 (O_850,N_4959,N_4905);
and UO_851 (O_851,N_4879,N_4989);
nand UO_852 (O_852,N_4938,N_4943);
xor UO_853 (O_853,N_4966,N_4911);
xor UO_854 (O_854,N_4846,N_4891);
and UO_855 (O_855,N_4802,N_4880);
nand UO_856 (O_856,N_4896,N_4821);
nand UO_857 (O_857,N_4979,N_4973);
nand UO_858 (O_858,N_4926,N_4961);
nand UO_859 (O_859,N_4979,N_4945);
nor UO_860 (O_860,N_4913,N_4963);
or UO_861 (O_861,N_4827,N_4892);
or UO_862 (O_862,N_4860,N_4954);
or UO_863 (O_863,N_4869,N_4944);
or UO_864 (O_864,N_4960,N_4932);
or UO_865 (O_865,N_4900,N_4919);
or UO_866 (O_866,N_4808,N_4919);
nand UO_867 (O_867,N_4821,N_4980);
nand UO_868 (O_868,N_4994,N_4964);
and UO_869 (O_869,N_4915,N_4905);
and UO_870 (O_870,N_4993,N_4802);
or UO_871 (O_871,N_4982,N_4950);
and UO_872 (O_872,N_4949,N_4879);
nand UO_873 (O_873,N_4837,N_4926);
and UO_874 (O_874,N_4812,N_4887);
nor UO_875 (O_875,N_4944,N_4904);
or UO_876 (O_876,N_4940,N_4989);
or UO_877 (O_877,N_4984,N_4816);
or UO_878 (O_878,N_4868,N_4841);
or UO_879 (O_879,N_4872,N_4907);
nand UO_880 (O_880,N_4844,N_4977);
and UO_881 (O_881,N_4938,N_4928);
nand UO_882 (O_882,N_4888,N_4805);
and UO_883 (O_883,N_4903,N_4845);
xor UO_884 (O_884,N_4854,N_4808);
nand UO_885 (O_885,N_4888,N_4956);
nand UO_886 (O_886,N_4880,N_4865);
nand UO_887 (O_887,N_4825,N_4889);
or UO_888 (O_888,N_4828,N_4896);
nand UO_889 (O_889,N_4820,N_4868);
or UO_890 (O_890,N_4885,N_4941);
or UO_891 (O_891,N_4840,N_4926);
or UO_892 (O_892,N_4846,N_4848);
nor UO_893 (O_893,N_4805,N_4873);
nand UO_894 (O_894,N_4821,N_4992);
nand UO_895 (O_895,N_4912,N_4915);
xnor UO_896 (O_896,N_4910,N_4836);
or UO_897 (O_897,N_4900,N_4814);
nor UO_898 (O_898,N_4853,N_4849);
or UO_899 (O_899,N_4866,N_4915);
nand UO_900 (O_900,N_4837,N_4961);
nor UO_901 (O_901,N_4861,N_4974);
nor UO_902 (O_902,N_4973,N_4827);
nand UO_903 (O_903,N_4999,N_4813);
or UO_904 (O_904,N_4904,N_4989);
xor UO_905 (O_905,N_4968,N_4832);
nand UO_906 (O_906,N_4922,N_4870);
and UO_907 (O_907,N_4853,N_4905);
or UO_908 (O_908,N_4868,N_4854);
nand UO_909 (O_909,N_4917,N_4885);
or UO_910 (O_910,N_4909,N_4911);
xor UO_911 (O_911,N_4811,N_4898);
nand UO_912 (O_912,N_4993,N_4962);
nand UO_913 (O_913,N_4876,N_4993);
nand UO_914 (O_914,N_4848,N_4840);
nand UO_915 (O_915,N_4912,N_4991);
xnor UO_916 (O_916,N_4849,N_4952);
and UO_917 (O_917,N_4927,N_4881);
nor UO_918 (O_918,N_4842,N_4969);
xnor UO_919 (O_919,N_4802,N_4827);
nor UO_920 (O_920,N_4897,N_4929);
and UO_921 (O_921,N_4939,N_4851);
or UO_922 (O_922,N_4947,N_4882);
nor UO_923 (O_923,N_4961,N_4800);
nor UO_924 (O_924,N_4996,N_4867);
or UO_925 (O_925,N_4846,N_4845);
nand UO_926 (O_926,N_4910,N_4821);
and UO_927 (O_927,N_4825,N_4856);
nor UO_928 (O_928,N_4951,N_4837);
nor UO_929 (O_929,N_4920,N_4913);
and UO_930 (O_930,N_4823,N_4880);
or UO_931 (O_931,N_4960,N_4939);
or UO_932 (O_932,N_4916,N_4909);
nand UO_933 (O_933,N_4954,N_4976);
nor UO_934 (O_934,N_4845,N_4999);
nand UO_935 (O_935,N_4859,N_4936);
and UO_936 (O_936,N_4977,N_4877);
and UO_937 (O_937,N_4953,N_4807);
xnor UO_938 (O_938,N_4866,N_4894);
and UO_939 (O_939,N_4979,N_4955);
and UO_940 (O_940,N_4976,N_4959);
xor UO_941 (O_941,N_4849,N_4949);
nand UO_942 (O_942,N_4811,N_4845);
or UO_943 (O_943,N_4817,N_4953);
xor UO_944 (O_944,N_4932,N_4998);
or UO_945 (O_945,N_4836,N_4973);
nand UO_946 (O_946,N_4978,N_4885);
or UO_947 (O_947,N_4827,N_4834);
xnor UO_948 (O_948,N_4817,N_4830);
xnor UO_949 (O_949,N_4868,N_4825);
nor UO_950 (O_950,N_4953,N_4813);
or UO_951 (O_951,N_4916,N_4882);
or UO_952 (O_952,N_4807,N_4877);
nor UO_953 (O_953,N_4814,N_4981);
and UO_954 (O_954,N_4850,N_4901);
and UO_955 (O_955,N_4842,N_4845);
and UO_956 (O_956,N_4896,N_4814);
and UO_957 (O_957,N_4912,N_4849);
and UO_958 (O_958,N_4987,N_4927);
nand UO_959 (O_959,N_4887,N_4822);
nor UO_960 (O_960,N_4887,N_4929);
nand UO_961 (O_961,N_4971,N_4804);
or UO_962 (O_962,N_4818,N_4948);
and UO_963 (O_963,N_4908,N_4878);
nand UO_964 (O_964,N_4827,N_4868);
nor UO_965 (O_965,N_4975,N_4870);
nor UO_966 (O_966,N_4889,N_4873);
or UO_967 (O_967,N_4954,N_4970);
or UO_968 (O_968,N_4865,N_4932);
or UO_969 (O_969,N_4943,N_4833);
or UO_970 (O_970,N_4972,N_4863);
nor UO_971 (O_971,N_4999,N_4867);
or UO_972 (O_972,N_4932,N_4824);
and UO_973 (O_973,N_4836,N_4952);
nor UO_974 (O_974,N_4834,N_4970);
or UO_975 (O_975,N_4898,N_4998);
and UO_976 (O_976,N_4906,N_4806);
xnor UO_977 (O_977,N_4942,N_4927);
and UO_978 (O_978,N_4908,N_4925);
nor UO_979 (O_979,N_4918,N_4959);
and UO_980 (O_980,N_4901,N_4843);
nor UO_981 (O_981,N_4841,N_4964);
xnor UO_982 (O_982,N_4847,N_4983);
nor UO_983 (O_983,N_4860,N_4869);
or UO_984 (O_984,N_4973,N_4984);
nor UO_985 (O_985,N_4965,N_4960);
xor UO_986 (O_986,N_4835,N_4841);
and UO_987 (O_987,N_4842,N_4894);
and UO_988 (O_988,N_4861,N_4929);
and UO_989 (O_989,N_4920,N_4936);
nand UO_990 (O_990,N_4969,N_4984);
nor UO_991 (O_991,N_4805,N_4800);
or UO_992 (O_992,N_4952,N_4859);
or UO_993 (O_993,N_4807,N_4909);
or UO_994 (O_994,N_4952,N_4804);
nand UO_995 (O_995,N_4924,N_4822);
or UO_996 (O_996,N_4871,N_4978);
nand UO_997 (O_997,N_4804,N_4849);
nor UO_998 (O_998,N_4923,N_4917);
and UO_999 (O_999,N_4829,N_4871);
endmodule