module basic_500_3000_500_50_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_341,In_247);
nor U1 (N_1,In_115,In_429);
nor U2 (N_2,In_428,In_281);
nor U3 (N_3,In_352,In_482);
nand U4 (N_4,In_43,In_13);
and U5 (N_5,In_160,In_147);
and U6 (N_6,In_280,In_381);
nor U7 (N_7,In_212,In_228);
or U8 (N_8,In_211,In_473);
nand U9 (N_9,In_274,In_277);
and U10 (N_10,In_32,In_146);
nand U11 (N_11,In_89,In_271);
and U12 (N_12,In_229,In_472);
nor U13 (N_13,In_99,In_11);
nand U14 (N_14,In_359,In_363);
nand U15 (N_15,In_193,In_67);
nand U16 (N_16,In_322,In_476);
nand U17 (N_17,In_114,In_225);
nor U18 (N_18,In_12,In_201);
xor U19 (N_19,In_188,In_80);
nand U20 (N_20,In_199,In_182);
xor U21 (N_21,In_218,In_110);
or U22 (N_22,In_435,In_289);
and U23 (N_23,In_483,In_446);
xnor U24 (N_24,In_36,In_244);
and U25 (N_25,In_220,In_190);
or U26 (N_26,In_22,In_31);
and U27 (N_27,In_408,In_140);
and U28 (N_28,In_245,In_465);
xnor U29 (N_29,In_168,In_109);
nor U30 (N_30,In_276,In_16);
xnor U31 (N_31,In_368,In_165);
or U32 (N_32,In_18,In_139);
and U33 (N_33,In_237,In_296);
nor U34 (N_34,In_5,In_197);
nand U35 (N_35,In_65,In_464);
xnor U36 (N_36,In_495,In_486);
xnor U37 (N_37,In_377,In_273);
nor U38 (N_38,In_198,In_332);
or U39 (N_39,In_493,In_66);
xor U40 (N_40,In_174,In_24);
nand U41 (N_41,In_10,In_158);
or U42 (N_42,In_407,In_378);
and U43 (N_43,In_291,In_216);
nor U44 (N_44,In_223,In_309);
or U45 (N_45,In_152,In_58);
or U46 (N_46,In_369,In_302);
nand U47 (N_47,In_306,In_55);
xor U48 (N_48,In_163,In_29);
xor U49 (N_49,In_479,In_59);
or U50 (N_50,In_189,In_124);
nand U51 (N_51,In_343,In_321);
or U52 (N_52,In_414,In_405);
nand U53 (N_53,In_126,In_463);
xnor U54 (N_54,In_437,In_365);
nor U55 (N_55,In_349,In_316);
and U56 (N_56,In_45,In_200);
xnor U57 (N_57,In_346,In_286);
xnor U58 (N_58,In_362,In_42);
nand U59 (N_59,In_275,In_235);
nor U60 (N_60,N_51,In_459);
or U61 (N_61,N_28,In_287);
nand U62 (N_62,In_379,In_130);
nand U63 (N_63,In_143,N_27);
xor U64 (N_64,In_56,In_87);
or U65 (N_65,In_373,In_0);
xnor U66 (N_66,In_283,In_471);
nand U67 (N_67,In_453,In_14);
nor U68 (N_68,In_419,In_269);
nor U69 (N_69,In_44,N_14);
xor U70 (N_70,In_107,In_261);
nand U71 (N_71,N_26,In_221);
xnor U72 (N_72,In_490,In_250);
nor U73 (N_73,In_398,In_427);
nand U74 (N_74,In_454,In_30);
nor U75 (N_75,In_496,In_164);
or U76 (N_76,In_335,In_249);
nor U77 (N_77,In_451,In_345);
xor U78 (N_78,In_297,In_394);
nand U79 (N_79,In_272,In_450);
nand U80 (N_80,In_412,In_185);
nor U81 (N_81,In_366,In_4);
nand U82 (N_82,In_304,N_19);
nor U83 (N_83,In_62,N_42);
nor U84 (N_84,In_468,In_171);
and U85 (N_85,N_15,In_334);
xnor U86 (N_86,In_120,In_434);
nand U87 (N_87,In_238,In_466);
nor U88 (N_88,In_48,In_191);
or U89 (N_89,In_416,N_30);
xnor U90 (N_90,In_155,In_353);
or U91 (N_91,In_392,In_396);
nand U92 (N_92,In_118,N_40);
xnor U93 (N_93,In_282,In_461);
and U94 (N_94,In_433,In_457);
or U95 (N_95,N_17,In_447);
nor U96 (N_96,In_327,In_324);
and U97 (N_97,N_48,In_263);
and U98 (N_98,In_95,In_195);
and U99 (N_99,In_76,In_90);
and U100 (N_100,In_47,In_358);
nor U101 (N_101,In_279,N_52);
and U102 (N_102,In_367,In_492);
and U103 (N_103,In_315,In_129);
xnor U104 (N_104,In_77,In_208);
nand U105 (N_105,In_41,In_336);
and U106 (N_106,In_2,In_3);
and U107 (N_107,In_86,In_127);
nor U108 (N_108,In_219,In_179);
xnor U109 (N_109,In_106,In_243);
and U110 (N_110,In_293,In_424);
nor U111 (N_111,N_31,In_79);
and U112 (N_112,N_37,In_299);
xor U113 (N_113,In_49,In_415);
xor U114 (N_114,In_300,In_173);
and U115 (N_115,In_204,In_402);
or U116 (N_116,In_399,N_53);
xor U117 (N_117,N_16,In_338);
nor U118 (N_118,In_456,N_55);
and U119 (N_119,In_142,In_93);
and U120 (N_120,In_432,In_194);
nand U121 (N_121,In_102,In_330);
nand U122 (N_122,In_411,In_119);
nand U123 (N_123,In_175,N_90);
or U124 (N_124,N_110,In_387);
nand U125 (N_125,In_475,In_138);
xor U126 (N_126,N_6,In_497);
nor U127 (N_127,N_73,In_176);
and U128 (N_128,In_389,In_101);
nor U129 (N_129,N_104,In_21);
xor U130 (N_130,In_105,In_375);
nor U131 (N_131,In_170,In_131);
and U132 (N_132,N_18,In_210);
or U133 (N_133,In_372,In_395);
xor U134 (N_134,In_159,In_469);
and U135 (N_135,In_136,N_108);
xor U136 (N_136,N_7,In_292);
xnor U137 (N_137,In_391,In_117);
or U138 (N_138,In_357,In_157);
nor U139 (N_139,In_254,N_119);
nor U140 (N_140,In_9,In_294);
and U141 (N_141,N_72,N_97);
nor U142 (N_142,N_92,In_54);
nor U143 (N_143,In_374,N_32);
nand U144 (N_144,N_103,In_448);
nor U145 (N_145,In_312,In_488);
and U146 (N_146,In_307,In_78);
and U147 (N_147,In_376,In_401);
or U148 (N_148,In_187,In_305);
nand U149 (N_149,In_236,In_478);
or U150 (N_150,N_57,In_35);
xnor U151 (N_151,N_91,N_65);
xor U152 (N_152,In_270,In_224);
and U153 (N_153,In_60,In_183);
xnor U154 (N_154,In_442,In_134);
and U155 (N_155,In_319,In_284);
nor U156 (N_156,In_20,In_73);
or U157 (N_157,In_148,In_241);
nor U158 (N_158,N_106,N_105);
nor U159 (N_159,N_56,In_121);
or U160 (N_160,In_268,In_441);
nor U161 (N_161,In_104,In_103);
and U162 (N_162,In_356,In_423);
and U163 (N_163,In_206,In_149);
xnor U164 (N_164,N_100,In_361);
and U165 (N_165,N_38,In_213);
nor U166 (N_166,N_39,In_410);
nor U167 (N_167,In_85,In_278);
nand U168 (N_168,In_354,N_12);
xnor U169 (N_169,In_258,In_84);
or U170 (N_170,In_491,In_400);
xnor U171 (N_171,In_452,In_123);
xor U172 (N_172,In_474,In_351);
nor U173 (N_173,In_470,N_115);
nor U174 (N_174,In_253,In_371);
or U175 (N_175,In_494,N_69);
and U176 (N_176,In_128,In_458);
xor U177 (N_177,N_34,N_41);
and U178 (N_178,N_68,N_0);
nor U179 (N_179,In_37,In_82);
nand U180 (N_180,N_83,In_51);
nor U181 (N_181,N_130,N_62);
nor U182 (N_182,In_156,In_72);
or U183 (N_183,N_168,In_460);
nand U184 (N_184,In_234,In_57);
xnor U185 (N_185,In_205,In_81);
nand U186 (N_186,In_313,In_167);
and U187 (N_187,In_413,In_422);
and U188 (N_188,N_82,In_53);
and U189 (N_189,In_83,N_123);
nand U190 (N_190,N_46,In_111);
nor U191 (N_191,N_161,N_175);
nand U192 (N_192,N_134,In_339);
and U193 (N_193,N_145,N_144);
and U194 (N_194,N_84,In_257);
or U195 (N_195,N_75,In_137);
nand U196 (N_196,In_132,N_157);
xnor U197 (N_197,In_7,N_74);
nand U198 (N_198,In_40,In_467);
and U199 (N_199,N_177,In_100);
and U200 (N_200,N_80,In_325);
or U201 (N_201,N_129,In_240);
nand U202 (N_202,N_63,In_355);
nor U203 (N_203,N_60,In_285);
and U204 (N_204,In_231,In_184);
xor U205 (N_205,In_38,N_150);
and U206 (N_206,N_10,In_487);
nor U207 (N_207,In_153,In_317);
nor U208 (N_208,N_1,N_22);
and U209 (N_209,N_36,N_178);
and U210 (N_210,In_295,N_76);
xor U211 (N_211,In_262,In_1);
nand U212 (N_212,In_484,N_137);
and U213 (N_213,In_17,N_77);
xor U214 (N_214,N_87,In_438);
nor U215 (N_215,In_260,N_85);
nor U216 (N_216,N_24,N_33);
and U217 (N_217,In_88,In_485);
xnor U218 (N_218,In_154,N_45);
nor U219 (N_219,In_248,In_264);
and U220 (N_220,In_288,In_267);
or U221 (N_221,In_462,In_333);
nor U222 (N_222,In_25,N_166);
nand U223 (N_223,N_102,N_136);
or U224 (N_224,N_8,In_203);
nand U225 (N_225,In_337,N_169);
and U226 (N_226,In_230,In_112);
nand U227 (N_227,N_162,N_79);
nor U228 (N_228,N_152,In_348);
or U229 (N_229,In_310,In_323);
nand U230 (N_230,N_107,In_209);
nor U231 (N_231,In_409,N_101);
nor U232 (N_232,N_111,N_59);
or U233 (N_233,In_196,In_151);
xor U234 (N_234,In_96,N_160);
or U235 (N_235,In_39,In_145);
nor U236 (N_236,N_9,N_89);
nor U237 (N_237,N_127,N_148);
or U238 (N_238,In_251,In_144);
nor U239 (N_239,N_173,In_350);
or U240 (N_240,In_439,N_229);
nor U241 (N_241,In_420,In_311);
xnor U242 (N_242,N_95,N_176);
and U243 (N_243,N_143,N_214);
or U244 (N_244,N_182,In_498);
xnor U245 (N_245,N_142,N_50);
or U246 (N_246,N_122,In_180);
or U247 (N_247,N_186,N_133);
and U248 (N_248,In_233,N_86);
and U249 (N_249,N_158,N_140);
or U250 (N_250,In_445,In_181);
nand U251 (N_251,In_383,N_138);
xnor U252 (N_252,In_386,N_70);
and U253 (N_253,In_207,N_199);
nand U254 (N_254,In_426,N_155);
nand U255 (N_255,N_174,In_217);
nor U256 (N_256,N_125,N_121);
nand U257 (N_257,N_197,In_232);
nor U258 (N_258,In_318,N_235);
nand U259 (N_259,In_202,N_209);
and U260 (N_260,In_364,N_222);
or U261 (N_261,N_44,In_290);
nand U262 (N_262,In_265,N_2);
nor U263 (N_263,In_444,N_98);
xor U264 (N_264,In_64,N_189);
nor U265 (N_265,In_440,N_151);
or U266 (N_266,In_342,N_192);
or U267 (N_267,In_252,In_166);
xor U268 (N_268,N_219,N_179);
and U269 (N_269,N_35,N_211);
or U270 (N_270,In_403,N_96);
or U271 (N_271,In_50,N_208);
nor U272 (N_272,N_183,In_393);
and U273 (N_273,N_218,N_188);
and U274 (N_274,In_314,N_228);
or U275 (N_275,N_20,In_26);
and U276 (N_276,N_147,In_308);
and U277 (N_277,In_98,N_181);
or U278 (N_278,N_233,In_92);
nor U279 (N_279,In_303,In_34);
xnor U280 (N_280,In_404,In_390);
nand U281 (N_281,N_54,N_180);
and U282 (N_282,N_81,In_91);
or U283 (N_283,N_191,In_384);
nand U284 (N_284,In_430,In_449);
nand U285 (N_285,In_186,N_210);
xnor U286 (N_286,N_61,In_256);
xnor U287 (N_287,N_230,N_88);
xnor U288 (N_288,N_220,N_149);
or U289 (N_289,N_207,N_116);
and U290 (N_290,N_156,N_94);
nand U291 (N_291,In_239,In_481);
nor U292 (N_292,In_227,In_71);
or U293 (N_293,N_167,N_238);
nand U294 (N_294,In_116,In_380);
or U295 (N_295,N_205,In_222);
xnor U296 (N_296,N_190,N_67);
nand U297 (N_297,N_43,N_13);
nor U298 (N_298,N_217,N_216);
xnor U299 (N_299,In_19,N_120);
nor U300 (N_300,N_124,N_289);
xor U301 (N_301,In_52,In_421);
or U302 (N_302,N_285,N_267);
xor U303 (N_303,In_6,N_296);
nand U304 (N_304,In_33,N_258);
xnor U305 (N_305,In_489,N_5);
nand U306 (N_306,N_295,In_108);
xor U307 (N_307,N_198,N_283);
and U308 (N_308,N_170,In_214);
or U309 (N_309,N_294,N_268);
xnor U310 (N_310,In_326,In_266);
or U311 (N_311,In_455,N_244);
or U312 (N_312,N_250,N_251);
nand U313 (N_313,In_28,N_221);
xor U314 (N_314,In_75,In_499);
and U315 (N_315,In_141,In_417);
and U316 (N_316,N_227,In_242);
nor U317 (N_317,N_117,In_370);
xnor U318 (N_318,N_113,N_47);
nor U319 (N_319,N_249,N_212);
and U320 (N_320,In_226,In_68);
xor U321 (N_321,N_231,N_281);
nor U322 (N_322,N_21,N_275);
xnor U323 (N_323,In_169,N_262);
nand U324 (N_324,In_133,N_277);
nand U325 (N_325,In_480,N_195);
nor U326 (N_326,N_223,N_126);
or U327 (N_327,In_397,N_71);
or U328 (N_328,In_125,N_118);
and U329 (N_329,N_287,In_23);
or U330 (N_330,In_388,In_113);
or U331 (N_331,In_477,N_232);
nor U332 (N_332,N_257,N_135);
nand U333 (N_333,In_8,N_224);
nand U334 (N_334,N_242,N_291);
nand U335 (N_335,N_226,N_298);
and U336 (N_336,In_172,N_292);
or U337 (N_337,N_193,N_252);
and U338 (N_338,In_329,N_29);
xor U339 (N_339,N_297,In_443);
nor U340 (N_340,N_184,In_27);
nand U341 (N_341,N_256,N_164);
and U342 (N_342,In_135,N_202);
xnor U343 (N_343,N_154,N_128);
and U344 (N_344,N_23,N_248);
or U345 (N_345,N_172,N_288);
xor U346 (N_346,N_265,In_177);
or U347 (N_347,N_201,N_247);
nor U348 (N_348,N_163,N_78);
nor U349 (N_349,N_270,In_425);
or U350 (N_350,In_97,N_225);
xnor U351 (N_351,In_259,N_25);
nand U352 (N_352,In_122,N_284);
nand U353 (N_353,In_301,N_112);
xor U354 (N_354,N_11,In_418);
and U355 (N_355,In_347,In_406);
or U356 (N_356,N_215,In_382);
xnor U357 (N_357,In_162,N_264);
xor U358 (N_358,N_271,N_200);
nor U359 (N_359,In_344,N_273);
or U360 (N_360,N_354,N_260);
nor U361 (N_361,N_236,N_213);
or U362 (N_362,N_253,N_346);
nor U363 (N_363,N_318,In_320);
nand U364 (N_364,N_315,N_309);
nor U365 (N_365,N_259,N_301);
xor U366 (N_366,N_316,N_327);
nand U367 (N_367,N_356,N_317);
and U368 (N_368,N_109,N_357);
or U369 (N_369,In_15,N_355);
nand U370 (N_370,N_330,N_49);
nor U371 (N_371,N_302,In_69);
xnor U372 (N_372,N_245,N_328);
xor U373 (N_373,N_325,N_329);
or U374 (N_374,In_385,In_298);
or U375 (N_375,N_93,N_338);
xnor U376 (N_376,In_431,N_261);
nand U377 (N_377,N_353,In_150);
xnor U378 (N_378,N_299,In_328);
nor U379 (N_379,N_286,In_255);
and U380 (N_380,N_254,N_359);
or U381 (N_381,N_240,N_114);
xor U382 (N_382,N_324,N_332);
xor U383 (N_383,In_246,N_196);
nand U384 (N_384,N_185,N_351);
nor U385 (N_385,In_360,N_334);
nand U386 (N_386,N_349,N_3);
and U387 (N_387,N_340,N_352);
xor U388 (N_388,N_323,N_278);
and U389 (N_389,N_336,N_345);
nand U390 (N_390,N_99,N_206);
nand U391 (N_391,N_313,N_279);
nand U392 (N_392,N_326,N_331);
nand U393 (N_393,N_241,N_319);
xor U394 (N_394,In_61,In_192);
nor U395 (N_395,N_303,N_237);
xor U396 (N_396,In_161,N_333);
nor U397 (N_397,N_344,N_165);
and U398 (N_398,N_312,N_321);
nor U399 (N_399,N_304,N_266);
or U400 (N_400,N_243,N_171);
nor U401 (N_401,N_139,In_215);
nor U402 (N_402,In_46,N_339);
nor U403 (N_403,N_269,N_280);
or U404 (N_404,N_306,N_153);
and U405 (N_405,N_204,N_64);
or U406 (N_406,N_308,N_234);
and U407 (N_407,N_255,N_58);
or U408 (N_408,N_290,N_337);
nand U409 (N_409,N_159,N_314);
nor U410 (N_410,N_274,N_300);
or U411 (N_411,N_66,N_187);
nand U412 (N_412,In_63,N_348);
or U413 (N_413,In_178,N_263);
and U414 (N_414,N_141,N_307);
nand U415 (N_415,In_331,N_239);
and U416 (N_416,N_4,N_132);
and U417 (N_417,N_282,N_146);
nor U418 (N_418,N_310,In_74);
nand U419 (N_419,In_94,N_311);
xnor U420 (N_420,N_341,N_370);
and U421 (N_421,N_246,N_414);
nor U422 (N_422,N_377,N_374);
and U423 (N_423,N_403,N_413);
nand U424 (N_424,N_322,N_373);
nor U425 (N_425,N_358,N_397);
and U426 (N_426,N_203,N_379);
xnor U427 (N_427,N_361,N_396);
nand U428 (N_428,N_390,N_395);
xnor U429 (N_429,N_350,N_398);
nand U430 (N_430,N_388,N_386);
or U431 (N_431,N_418,N_385);
nand U432 (N_432,N_276,N_367);
or U433 (N_433,N_378,N_369);
nor U434 (N_434,N_381,N_363);
or U435 (N_435,In_340,N_392);
xor U436 (N_436,N_412,N_375);
nand U437 (N_437,N_411,N_305);
or U438 (N_438,N_399,N_409);
nor U439 (N_439,N_405,N_380);
xor U440 (N_440,N_371,N_419);
xor U441 (N_441,N_410,In_70);
and U442 (N_442,N_384,In_436);
nand U443 (N_443,N_362,N_364);
nor U444 (N_444,N_400,N_335);
nor U445 (N_445,N_365,N_293);
and U446 (N_446,N_366,N_415);
and U447 (N_447,N_347,N_417);
and U448 (N_448,N_383,N_320);
xnor U449 (N_449,N_272,N_360);
or U450 (N_450,N_389,N_407);
nor U451 (N_451,N_416,N_394);
xor U452 (N_452,N_393,N_391);
xor U453 (N_453,N_404,N_376);
nor U454 (N_454,N_194,N_387);
nor U455 (N_455,N_401,N_408);
nand U456 (N_456,N_406,N_402);
nor U457 (N_457,N_372,N_342);
xnor U458 (N_458,N_131,N_382);
or U459 (N_459,N_368,N_343);
nand U460 (N_460,N_379,N_411);
and U461 (N_461,N_390,N_372);
and U462 (N_462,N_401,N_402);
or U463 (N_463,N_380,N_409);
nor U464 (N_464,N_396,N_387);
or U465 (N_465,N_391,N_399);
or U466 (N_466,N_272,N_342);
nor U467 (N_467,N_341,N_360);
and U468 (N_468,N_406,N_408);
nand U469 (N_469,In_340,In_436);
nor U470 (N_470,N_415,N_131);
xnor U471 (N_471,N_362,N_400);
nor U472 (N_472,N_415,N_203);
xnor U473 (N_473,N_377,In_70);
and U474 (N_474,In_340,N_416);
and U475 (N_475,N_373,In_340);
xor U476 (N_476,N_361,N_366);
nor U477 (N_477,N_335,N_402);
and U478 (N_478,N_402,N_390);
and U479 (N_479,N_418,N_246);
nand U480 (N_480,N_423,N_478);
and U481 (N_481,N_442,N_477);
xor U482 (N_482,N_473,N_453);
or U483 (N_483,N_472,N_475);
or U484 (N_484,N_435,N_466);
and U485 (N_485,N_432,N_426);
nand U486 (N_486,N_448,N_433);
nand U487 (N_487,N_464,N_468);
nand U488 (N_488,N_471,N_467);
and U489 (N_489,N_422,N_447);
xor U490 (N_490,N_476,N_470);
xnor U491 (N_491,N_469,N_455);
or U492 (N_492,N_465,N_437);
or U493 (N_493,N_429,N_427);
xor U494 (N_494,N_431,N_446);
nor U495 (N_495,N_445,N_439);
nand U496 (N_496,N_459,N_451);
xnor U497 (N_497,N_454,N_449);
or U498 (N_498,N_436,N_456);
nor U499 (N_499,N_458,N_428);
or U500 (N_500,N_438,N_461);
nor U501 (N_501,N_421,N_425);
xor U502 (N_502,N_420,N_443);
or U503 (N_503,N_430,N_460);
and U504 (N_504,N_479,N_450);
nor U505 (N_505,N_463,N_434);
xnor U506 (N_506,N_462,N_440);
xnor U507 (N_507,N_444,N_424);
and U508 (N_508,N_441,N_457);
or U509 (N_509,N_474,N_452);
or U510 (N_510,N_424,N_428);
nor U511 (N_511,N_449,N_470);
or U512 (N_512,N_435,N_439);
or U513 (N_513,N_437,N_475);
or U514 (N_514,N_433,N_423);
and U515 (N_515,N_474,N_439);
nor U516 (N_516,N_458,N_456);
nor U517 (N_517,N_421,N_478);
xnor U518 (N_518,N_469,N_451);
xor U519 (N_519,N_447,N_465);
nor U520 (N_520,N_459,N_471);
nand U521 (N_521,N_434,N_457);
or U522 (N_522,N_456,N_447);
xnor U523 (N_523,N_466,N_447);
nor U524 (N_524,N_467,N_465);
or U525 (N_525,N_438,N_440);
and U526 (N_526,N_473,N_454);
or U527 (N_527,N_456,N_431);
nand U528 (N_528,N_438,N_460);
nand U529 (N_529,N_462,N_461);
xor U530 (N_530,N_450,N_463);
or U531 (N_531,N_454,N_434);
or U532 (N_532,N_433,N_458);
or U533 (N_533,N_447,N_441);
and U534 (N_534,N_463,N_424);
nand U535 (N_535,N_429,N_425);
or U536 (N_536,N_430,N_441);
nand U537 (N_537,N_452,N_424);
xor U538 (N_538,N_443,N_460);
nor U539 (N_539,N_430,N_452);
and U540 (N_540,N_520,N_481);
nor U541 (N_541,N_504,N_530);
or U542 (N_542,N_498,N_491);
nor U543 (N_543,N_523,N_485);
and U544 (N_544,N_517,N_509);
nand U545 (N_545,N_536,N_516);
and U546 (N_546,N_539,N_519);
nor U547 (N_547,N_528,N_511);
or U548 (N_548,N_488,N_533);
nand U549 (N_549,N_521,N_492);
nor U550 (N_550,N_487,N_518);
nor U551 (N_551,N_538,N_496);
nand U552 (N_552,N_515,N_506);
nand U553 (N_553,N_537,N_507);
nand U554 (N_554,N_529,N_514);
nor U555 (N_555,N_525,N_482);
xor U556 (N_556,N_494,N_527);
nor U557 (N_557,N_512,N_534);
and U558 (N_558,N_480,N_524);
xnor U559 (N_559,N_483,N_526);
or U560 (N_560,N_531,N_489);
xnor U561 (N_561,N_505,N_495);
and U562 (N_562,N_490,N_503);
xor U563 (N_563,N_510,N_486);
xnor U564 (N_564,N_497,N_499);
and U565 (N_565,N_493,N_484);
xnor U566 (N_566,N_501,N_502);
or U567 (N_567,N_532,N_522);
xnor U568 (N_568,N_508,N_500);
or U569 (N_569,N_535,N_513);
and U570 (N_570,N_522,N_521);
nand U571 (N_571,N_509,N_528);
or U572 (N_572,N_480,N_508);
xnor U573 (N_573,N_496,N_514);
and U574 (N_574,N_529,N_510);
and U575 (N_575,N_522,N_508);
xor U576 (N_576,N_512,N_539);
nand U577 (N_577,N_528,N_482);
xnor U578 (N_578,N_484,N_501);
xor U579 (N_579,N_498,N_514);
nor U580 (N_580,N_526,N_539);
xor U581 (N_581,N_488,N_481);
xnor U582 (N_582,N_518,N_523);
or U583 (N_583,N_532,N_495);
nand U584 (N_584,N_490,N_513);
nand U585 (N_585,N_500,N_482);
and U586 (N_586,N_501,N_516);
nor U587 (N_587,N_531,N_504);
or U588 (N_588,N_487,N_504);
nand U589 (N_589,N_512,N_491);
xnor U590 (N_590,N_509,N_499);
and U591 (N_591,N_522,N_534);
or U592 (N_592,N_535,N_512);
nor U593 (N_593,N_529,N_480);
nor U594 (N_594,N_483,N_515);
xnor U595 (N_595,N_519,N_508);
nand U596 (N_596,N_501,N_532);
and U597 (N_597,N_516,N_481);
nor U598 (N_598,N_512,N_480);
xor U599 (N_599,N_482,N_504);
nand U600 (N_600,N_586,N_569);
xor U601 (N_601,N_573,N_570);
nand U602 (N_602,N_592,N_568);
nand U603 (N_603,N_566,N_584);
and U604 (N_604,N_577,N_594);
xnor U605 (N_605,N_576,N_572);
nor U606 (N_606,N_547,N_558);
xnor U607 (N_607,N_587,N_578);
or U608 (N_608,N_562,N_559);
nand U609 (N_609,N_540,N_567);
nor U610 (N_610,N_557,N_597);
and U611 (N_611,N_596,N_548);
and U612 (N_612,N_589,N_595);
nand U613 (N_613,N_588,N_560);
or U614 (N_614,N_590,N_585);
or U615 (N_615,N_571,N_583);
nor U616 (N_616,N_555,N_549);
and U617 (N_617,N_598,N_563);
xnor U618 (N_618,N_582,N_553);
xnor U619 (N_619,N_580,N_543);
or U620 (N_620,N_591,N_564);
and U621 (N_621,N_574,N_542);
nand U622 (N_622,N_544,N_561);
or U623 (N_623,N_554,N_550);
and U624 (N_624,N_551,N_556);
xor U625 (N_625,N_579,N_545);
nand U626 (N_626,N_575,N_599);
nor U627 (N_627,N_581,N_593);
nand U628 (N_628,N_541,N_565);
nand U629 (N_629,N_552,N_546);
nand U630 (N_630,N_545,N_596);
or U631 (N_631,N_568,N_562);
or U632 (N_632,N_549,N_580);
nand U633 (N_633,N_577,N_562);
nor U634 (N_634,N_568,N_565);
or U635 (N_635,N_581,N_564);
nand U636 (N_636,N_579,N_570);
and U637 (N_637,N_577,N_552);
or U638 (N_638,N_550,N_577);
and U639 (N_639,N_548,N_550);
nor U640 (N_640,N_576,N_574);
and U641 (N_641,N_578,N_548);
nand U642 (N_642,N_544,N_570);
nand U643 (N_643,N_567,N_578);
and U644 (N_644,N_561,N_572);
nand U645 (N_645,N_594,N_551);
xnor U646 (N_646,N_545,N_576);
and U647 (N_647,N_591,N_542);
nand U648 (N_648,N_595,N_568);
xor U649 (N_649,N_574,N_558);
nand U650 (N_650,N_568,N_583);
nor U651 (N_651,N_598,N_596);
and U652 (N_652,N_541,N_584);
xnor U653 (N_653,N_582,N_594);
nor U654 (N_654,N_585,N_584);
nand U655 (N_655,N_599,N_598);
and U656 (N_656,N_592,N_559);
or U657 (N_657,N_585,N_555);
nand U658 (N_658,N_553,N_585);
nor U659 (N_659,N_541,N_563);
nand U660 (N_660,N_640,N_609);
nor U661 (N_661,N_604,N_607);
and U662 (N_662,N_625,N_644);
nor U663 (N_663,N_631,N_620);
and U664 (N_664,N_623,N_622);
or U665 (N_665,N_642,N_646);
and U666 (N_666,N_655,N_653);
nand U667 (N_667,N_654,N_610);
and U668 (N_668,N_641,N_616);
xor U669 (N_669,N_658,N_647);
nand U670 (N_670,N_639,N_638);
and U671 (N_671,N_606,N_656);
nand U672 (N_672,N_635,N_630);
or U673 (N_673,N_615,N_614);
nor U674 (N_674,N_636,N_649);
and U675 (N_675,N_650,N_652);
nand U676 (N_676,N_648,N_613);
and U677 (N_677,N_602,N_612);
xor U678 (N_678,N_617,N_628);
or U679 (N_679,N_618,N_632);
or U680 (N_680,N_601,N_624);
xor U681 (N_681,N_627,N_608);
xor U682 (N_682,N_634,N_603);
nand U683 (N_683,N_657,N_645);
nor U684 (N_684,N_651,N_605);
or U685 (N_685,N_633,N_600);
xor U686 (N_686,N_629,N_619);
nand U687 (N_687,N_659,N_643);
nand U688 (N_688,N_621,N_626);
nor U689 (N_689,N_637,N_611);
nor U690 (N_690,N_641,N_624);
nor U691 (N_691,N_623,N_649);
nor U692 (N_692,N_631,N_621);
or U693 (N_693,N_631,N_624);
nand U694 (N_694,N_610,N_620);
or U695 (N_695,N_635,N_606);
or U696 (N_696,N_608,N_650);
xor U697 (N_697,N_642,N_626);
xor U698 (N_698,N_629,N_627);
nand U699 (N_699,N_611,N_627);
xnor U700 (N_700,N_622,N_635);
xnor U701 (N_701,N_641,N_611);
xnor U702 (N_702,N_645,N_651);
nor U703 (N_703,N_641,N_607);
or U704 (N_704,N_610,N_650);
nor U705 (N_705,N_621,N_647);
nor U706 (N_706,N_652,N_658);
and U707 (N_707,N_612,N_601);
and U708 (N_708,N_621,N_640);
nor U709 (N_709,N_622,N_651);
xnor U710 (N_710,N_624,N_607);
xnor U711 (N_711,N_637,N_612);
and U712 (N_712,N_616,N_628);
xor U713 (N_713,N_644,N_652);
and U714 (N_714,N_640,N_627);
or U715 (N_715,N_605,N_643);
xor U716 (N_716,N_619,N_643);
or U717 (N_717,N_625,N_643);
and U718 (N_718,N_635,N_639);
and U719 (N_719,N_639,N_616);
nor U720 (N_720,N_685,N_705);
xor U721 (N_721,N_686,N_690);
or U722 (N_722,N_694,N_672);
xor U723 (N_723,N_661,N_689);
nor U724 (N_724,N_717,N_714);
nor U725 (N_725,N_691,N_680);
or U726 (N_726,N_668,N_676);
nand U727 (N_727,N_679,N_687);
nor U728 (N_728,N_681,N_677);
and U729 (N_729,N_667,N_709);
xnor U730 (N_730,N_684,N_660);
xor U731 (N_731,N_696,N_700);
and U732 (N_732,N_693,N_704);
xnor U733 (N_733,N_719,N_718);
xnor U734 (N_734,N_715,N_669);
xor U735 (N_735,N_670,N_711);
nor U736 (N_736,N_697,N_713);
xnor U737 (N_737,N_708,N_707);
or U738 (N_738,N_688,N_706);
nand U739 (N_739,N_678,N_682);
or U740 (N_740,N_683,N_699);
and U741 (N_741,N_710,N_692);
nand U742 (N_742,N_712,N_665);
and U743 (N_743,N_664,N_695);
or U744 (N_744,N_675,N_663);
or U745 (N_745,N_674,N_662);
or U746 (N_746,N_673,N_671);
nand U747 (N_747,N_702,N_701);
or U748 (N_748,N_698,N_716);
nor U749 (N_749,N_703,N_666);
nor U750 (N_750,N_676,N_693);
nand U751 (N_751,N_684,N_673);
and U752 (N_752,N_670,N_682);
nor U753 (N_753,N_691,N_700);
nand U754 (N_754,N_665,N_692);
nor U755 (N_755,N_718,N_665);
and U756 (N_756,N_710,N_686);
nand U757 (N_757,N_701,N_666);
nand U758 (N_758,N_689,N_702);
and U759 (N_759,N_695,N_700);
and U760 (N_760,N_696,N_682);
and U761 (N_761,N_709,N_692);
or U762 (N_762,N_671,N_663);
and U763 (N_763,N_694,N_678);
and U764 (N_764,N_717,N_708);
or U765 (N_765,N_679,N_715);
xnor U766 (N_766,N_702,N_683);
nor U767 (N_767,N_701,N_692);
xnor U768 (N_768,N_711,N_668);
xnor U769 (N_769,N_718,N_683);
nor U770 (N_770,N_694,N_666);
nor U771 (N_771,N_679,N_713);
and U772 (N_772,N_671,N_698);
and U773 (N_773,N_674,N_717);
and U774 (N_774,N_681,N_714);
or U775 (N_775,N_684,N_717);
nor U776 (N_776,N_661,N_676);
xor U777 (N_777,N_685,N_663);
xor U778 (N_778,N_675,N_699);
nand U779 (N_779,N_708,N_718);
nor U780 (N_780,N_731,N_749);
or U781 (N_781,N_722,N_759);
nor U782 (N_782,N_756,N_767);
nand U783 (N_783,N_771,N_779);
nand U784 (N_784,N_758,N_729);
xor U785 (N_785,N_755,N_770);
nand U786 (N_786,N_740,N_764);
xor U787 (N_787,N_768,N_721);
xor U788 (N_788,N_774,N_744);
and U789 (N_789,N_723,N_736);
nor U790 (N_790,N_761,N_735);
xor U791 (N_791,N_752,N_742);
nor U792 (N_792,N_747,N_753);
or U793 (N_793,N_777,N_750);
nand U794 (N_794,N_724,N_727);
nand U795 (N_795,N_772,N_776);
nand U796 (N_796,N_741,N_760);
nor U797 (N_797,N_726,N_757);
or U798 (N_798,N_769,N_743);
nand U799 (N_799,N_751,N_745);
xor U800 (N_800,N_739,N_754);
or U801 (N_801,N_733,N_738);
nor U802 (N_802,N_734,N_746);
nor U803 (N_803,N_728,N_737);
nor U804 (N_804,N_732,N_748);
xor U805 (N_805,N_766,N_775);
xor U806 (N_806,N_730,N_773);
xor U807 (N_807,N_763,N_778);
nand U808 (N_808,N_725,N_765);
xor U809 (N_809,N_762,N_720);
xnor U810 (N_810,N_744,N_757);
nand U811 (N_811,N_723,N_757);
and U812 (N_812,N_770,N_737);
and U813 (N_813,N_749,N_773);
xor U814 (N_814,N_726,N_735);
nand U815 (N_815,N_720,N_731);
xnor U816 (N_816,N_750,N_728);
and U817 (N_817,N_732,N_733);
xor U818 (N_818,N_748,N_721);
nor U819 (N_819,N_772,N_741);
or U820 (N_820,N_728,N_768);
and U821 (N_821,N_733,N_722);
nand U822 (N_822,N_766,N_724);
xor U823 (N_823,N_735,N_752);
xor U824 (N_824,N_763,N_744);
nand U825 (N_825,N_779,N_762);
and U826 (N_826,N_742,N_747);
nor U827 (N_827,N_740,N_766);
and U828 (N_828,N_775,N_756);
xor U829 (N_829,N_756,N_741);
nor U830 (N_830,N_737,N_721);
and U831 (N_831,N_755,N_729);
nor U832 (N_832,N_738,N_773);
and U833 (N_833,N_763,N_773);
xnor U834 (N_834,N_736,N_778);
or U835 (N_835,N_767,N_727);
xor U836 (N_836,N_721,N_745);
xnor U837 (N_837,N_769,N_767);
or U838 (N_838,N_753,N_736);
xor U839 (N_839,N_724,N_720);
xnor U840 (N_840,N_814,N_819);
nor U841 (N_841,N_830,N_794);
or U842 (N_842,N_829,N_782);
or U843 (N_843,N_820,N_811);
nand U844 (N_844,N_800,N_783);
and U845 (N_845,N_831,N_833);
nor U846 (N_846,N_804,N_788);
and U847 (N_847,N_787,N_836);
nand U848 (N_848,N_780,N_810);
xor U849 (N_849,N_796,N_824);
xnor U850 (N_850,N_827,N_817);
nand U851 (N_851,N_795,N_812);
nand U852 (N_852,N_781,N_818);
nand U853 (N_853,N_813,N_791);
or U854 (N_854,N_805,N_789);
and U855 (N_855,N_799,N_816);
nand U856 (N_856,N_792,N_821);
nor U857 (N_857,N_803,N_784);
or U858 (N_858,N_807,N_823);
xnor U859 (N_859,N_838,N_822);
nand U860 (N_860,N_809,N_798);
nor U861 (N_861,N_828,N_785);
or U862 (N_862,N_815,N_832);
and U863 (N_863,N_802,N_835);
nor U864 (N_864,N_825,N_839);
nand U865 (N_865,N_808,N_834);
nand U866 (N_866,N_806,N_790);
nor U867 (N_867,N_837,N_826);
or U868 (N_868,N_786,N_793);
nand U869 (N_869,N_801,N_797);
and U870 (N_870,N_811,N_793);
xnor U871 (N_871,N_787,N_823);
nor U872 (N_872,N_811,N_795);
nor U873 (N_873,N_833,N_830);
or U874 (N_874,N_784,N_836);
nor U875 (N_875,N_801,N_782);
xnor U876 (N_876,N_787,N_799);
nor U877 (N_877,N_782,N_819);
and U878 (N_878,N_834,N_790);
xor U879 (N_879,N_823,N_831);
nand U880 (N_880,N_786,N_822);
or U881 (N_881,N_806,N_830);
nand U882 (N_882,N_822,N_834);
nor U883 (N_883,N_784,N_801);
or U884 (N_884,N_802,N_797);
xor U885 (N_885,N_800,N_790);
and U886 (N_886,N_821,N_836);
or U887 (N_887,N_813,N_823);
or U888 (N_888,N_834,N_786);
nand U889 (N_889,N_798,N_797);
xnor U890 (N_890,N_780,N_815);
nor U891 (N_891,N_783,N_803);
xor U892 (N_892,N_832,N_787);
xnor U893 (N_893,N_786,N_804);
and U894 (N_894,N_794,N_811);
or U895 (N_895,N_780,N_830);
and U896 (N_896,N_817,N_828);
and U897 (N_897,N_821,N_780);
and U898 (N_898,N_837,N_838);
or U899 (N_899,N_781,N_816);
xor U900 (N_900,N_849,N_852);
nand U901 (N_901,N_865,N_877);
or U902 (N_902,N_872,N_892);
xor U903 (N_903,N_853,N_889);
nand U904 (N_904,N_841,N_869);
and U905 (N_905,N_898,N_842);
or U906 (N_906,N_878,N_850);
nor U907 (N_907,N_864,N_848);
or U908 (N_908,N_887,N_891);
nand U909 (N_909,N_870,N_884);
nor U910 (N_910,N_885,N_890);
nand U911 (N_911,N_847,N_896);
xor U912 (N_912,N_899,N_863);
nand U913 (N_913,N_873,N_893);
nor U914 (N_914,N_851,N_846);
or U915 (N_915,N_845,N_876);
and U916 (N_916,N_857,N_855);
nor U917 (N_917,N_861,N_844);
or U918 (N_918,N_840,N_880);
or U919 (N_919,N_866,N_874);
nand U920 (N_920,N_856,N_886);
nor U921 (N_921,N_860,N_882);
nor U922 (N_922,N_862,N_871);
or U923 (N_923,N_897,N_881);
nor U924 (N_924,N_858,N_867);
or U925 (N_925,N_883,N_879);
xnor U926 (N_926,N_895,N_875);
and U927 (N_927,N_843,N_894);
nor U928 (N_928,N_868,N_888);
or U929 (N_929,N_854,N_859);
and U930 (N_930,N_884,N_840);
nand U931 (N_931,N_891,N_841);
or U932 (N_932,N_846,N_865);
nand U933 (N_933,N_847,N_858);
and U934 (N_934,N_875,N_845);
nor U935 (N_935,N_878,N_868);
and U936 (N_936,N_884,N_856);
nand U937 (N_937,N_863,N_884);
xor U938 (N_938,N_874,N_883);
nand U939 (N_939,N_856,N_883);
and U940 (N_940,N_871,N_896);
nand U941 (N_941,N_865,N_842);
or U942 (N_942,N_853,N_860);
or U943 (N_943,N_866,N_873);
nor U944 (N_944,N_888,N_882);
or U945 (N_945,N_873,N_872);
nand U946 (N_946,N_878,N_889);
or U947 (N_947,N_899,N_867);
or U948 (N_948,N_847,N_845);
nand U949 (N_949,N_854,N_884);
and U950 (N_950,N_853,N_847);
or U951 (N_951,N_874,N_871);
and U952 (N_952,N_883,N_846);
nand U953 (N_953,N_845,N_852);
nor U954 (N_954,N_844,N_862);
and U955 (N_955,N_862,N_896);
and U956 (N_956,N_851,N_840);
xnor U957 (N_957,N_842,N_840);
or U958 (N_958,N_876,N_843);
nor U959 (N_959,N_858,N_844);
nor U960 (N_960,N_931,N_929);
and U961 (N_961,N_915,N_909);
nand U962 (N_962,N_954,N_932);
xnor U963 (N_963,N_925,N_952);
or U964 (N_964,N_911,N_907);
nand U965 (N_965,N_935,N_937);
xnor U966 (N_966,N_945,N_936);
or U967 (N_967,N_928,N_922);
or U968 (N_968,N_951,N_948);
nand U969 (N_969,N_939,N_953);
nand U970 (N_970,N_920,N_905);
and U971 (N_971,N_901,N_956);
or U972 (N_972,N_902,N_950);
xor U973 (N_973,N_918,N_941);
and U974 (N_974,N_927,N_944);
xor U975 (N_975,N_930,N_946);
or U976 (N_976,N_933,N_913);
nand U977 (N_977,N_959,N_934);
nand U978 (N_978,N_908,N_943);
nor U979 (N_979,N_949,N_916);
nor U980 (N_980,N_906,N_924);
and U981 (N_981,N_904,N_940);
xor U982 (N_982,N_921,N_914);
or U983 (N_983,N_942,N_903);
nand U984 (N_984,N_957,N_900);
nand U985 (N_985,N_958,N_910);
nor U986 (N_986,N_917,N_938);
or U987 (N_987,N_955,N_947);
xnor U988 (N_988,N_912,N_919);
or U989 (N_989,N_923,N_926);
xor U990 (N_990,N_925,N_959);
or U991 (N_991,N_947,N_908);
nor U992 (N_992,N_911,N_914);
xnor U993 (N_993,N_947,N_907);
nand U994 (N_994,N_944,N_952);
nand U995 (N_995,N_928,N_904);
nand U996 (N_996,N_942,N_900);
or U997 (N_997,N_957,N_931);
and U998 (N_998,N_932,N_917);
or U999 (N_999,N_905,N_913);
nor U1000 (N_1000,N_902,N_958);
or U1001 (N_1001,N_947,N_917);
or U1002 (N_1002,N_903,N_927);
xor U1003 (N_1003,N_957,N_927);
xor U1004 (N_1004,N_934,N_929);
nand U1005 (N_1005,N_945,N_920);
nor U1006 (N_1006,N_935,N_914);
nor U1007 (N_1007,N_932,N_922);
nand U1008 (N_1008,N_913,N_939);
nand U1009 (N_1009,N_916,N_904);
or U1010 (N_1010,N_927,N_954);
xnor U1011 (N_1011,N_933,N_932);
nor U1012 (N_1012,N_940,N_948);
nand U1013 (N_1013,N_906,N_939);
xor U1014 (N_1014,N_918,N_915);
nand U1015 (N_1015,N_959,N_917);
xnor U1016 (N_1016,N_923,N_929);
nor U1017 (N_1017,N_959,N_922);
nor U1018 (N_1018,N_953,N_942);
xor U1019 (N_1019,N_903,N_934);
nand U1020 (N_1020,N_986,N_969);
xnor U1021 (N_1021,N_1006,N_1008);
xor U1022 (N_1022,N_1001,N_976);
nor U1023 (N_1023,N_987,N_1017);
or U1024 (N_1024,N_979,N_981);
xor U1025 (N_1025,N_998,N_988);
nor U1026 (N_1026,N_968,N_965);
or U1027 (N_1027,N_1018,N_996);
nand U1028 (N_1028,N_962,N_1015);
nor U1029 (N_1029,N_993,N_1009);
xor U1030 (N_1030,N_994,N_1014);
xnor U1031 (N_1031,N_991,N_974);
nor U1032 (N_1032,N_997,N_999);
xor U1033 (N_1033,N_990,N_978);
and U1034 (N_1034,N_972,N_984);
or U1035 (N_1035,N_1002,N_960);
xnor U1036 (N_1036,N_985,N_992);
or U1037 (N_1037,N_973,N_975);
or U1038 (N_1038,N_982,N_1004);
nor U1039 (N_1039,N_970,N_977);
or U1040 (N_1040,N_963,N_1000);
nand U1041 (N_1041,N_971,N_983);
or U1042 (N_1042,N_967,N_1013);
nor U1043 (N_1043,N_1016,N_980);
nand U1044 (N_1044,N_1005,N_1011);
nand U1045 (N_1045,N_1003,N_1007);
or U1046 (N_1046,N_1019,N_961);
or U1047 (N_1047,N_1010,N_989);
nand U1048 (N_1048,N_966,N_1012);
and U1049 (N_1049,N_964,N_995);
nor U1050 (N_1050,N_992,N_999);
or U1051 (N_1051,N_970,N_974);
nor U1052 (N_1052,N_988,N_1009);
nor U1053 (N_1053,N_1004,N_970);
and U1054 (N_1054,N_1006,N_1012);
or U1055 (N_1055,N_981,N_982);
and U1056 (N_1056,N_1015,N_997);
and U1057 (N_1057,N_995,N_962);
nor U1058 (N_1058,N_985,N_1017);
and U1059 (N_1059,N_1004,N_975);
xnor U1060 (N_1060,N_963,N_967);
xnor U1061 (N_1061,N_982,N_991);
nand U1062 (N_1062,N_1011,N_981);
nand U1063 (N_1063,N_1008,N_968);
or U1064 (N_1064,N_1005,N_990);
nor U1065 (N_1065,N_983,N_1009);
nor U1066 (N_1066,N_963,N_1011);
xor U1067 (N_1067,N_982,N_968);
xnor U1068 (N_1068,N_984,N_977);
nand U1069 (N_1069,N_1009,N_973);
nor U1070 (N_1070,N_976,N_1016);
and U1071 (N_1071,N_1006,N_976);
nand U1072 (N_1072,N_1011,N_971);
nor U1073 (N_1073,N_998,N_1003);
and U1074 (N_1074,N_991,N_962);
or U1075 (N_1075,N_999,N_1006);
or U1076 (N_1076,N_981,N_983);
and U1077 (N_1077,N_991,N_1019);
and U1078 (N_1078,N_976,N_1005);
nand U1079 (N_1079,N_985,N_995);
and U1080 (N_1080,N_1040,N_1064);
and U1081 (N_1081,N_1050,N_1069);
nor U1082 (N_1082,N_1072,N_1079);
and U1083 (N_1083,N_1066,N_1051);
nand U1084 (N_1084,N_1061,N_1043);
nand U1085 (N_1085,N_1023,N_1026);
nor U1086 (N_1086,N_1034,N_1029);
and U1087 (N_1087,N_1062,N_1057);
and U1088 (N_1088,N_1045,N_1049);
xnor U1089 (N_1089,N_1065,N_1058);
or U1090 (N_1090,N_1036,N_1059);
and U1091 (N_1091,N_1042,N_1028);
nor U1092 (N_1092,N_1021,N_1077);
nor U1093 (N_1093,N_1022,N_1070);
nand U1094 (N_1094,N_1027,N_1046);
and U1095 (N_1095,N_1033,N_1030);
nor U1096 (N_1096,N_1025,N_1054);
nor U1097 (N_1097,N_1048,N_1044);
nor U1098 (N_1098,N_1055,N_1071);
nor U1099 (N_1099,N_1053,N_1067);
nor U1100 (N_1100,N_1035,N_1024);
nand U1101 (N_1101,N_1031,N_1039);
nand U1102 (N_1102,N_1060,N_1063);
nand U1103 (N_1103,N_1075,N_1041);
or U1104 (N_1104,N_1073,N_1076);
nand U1105 (N_1105,N_1037,N_1078);
and U1106 (N_1106,N_1020,N_1074);
and U1107 (N_1107,N_1038,N_1047);
nand U1108 (N_1108,N_1032,N_1056);
or U1109 (N_1109,N_1068,N_1052);
and U1110 (N_1110,N_1051,N_1045);
and U1111 (N_1111,N_1040,N_1072);
or U1112 (N_1112,N_1029,N_1055);
or U1113 (N_1113,N_1029,N_1050);
and U1114 (N_1114,N_1068,N_1022);
nor U1115 (N_1115,N_1074,N_1030);
and U1116 (N_1116,N_1022,N_1074);
xnor U1117 (N_1117,N_1063,N_1054);
and U1118 (N_1118,N_1047,N_1024);
nor U1119 (N_1119,N_1062,N_1073);
nand U1120 (N_1120,N_1044,N_1062);
nand U1121 (N_1121,N_1022,N_1058);
or U1122 (N_1122,N_1071,N_1046);
nor U1123 (N_1123,N_1046,N_1073);
xnor U1124 (N_1124,N_1020,N_1046);
and U1125 (N_1125,N_1075,N_1020);
and U1126 (N_1126,N_1022,N_1063);
nor U1127 (N_1127,N_1050,N_1020);
xor U1128 (N_1128,N_1052,N_1057);
xnor U1129 (N_1129,N_1074,N_1058);
nor U1130 (N_1130,N_1057,N_1060);
nor U1131 (N_1131,N_1043,N_1068);
nor U1132 (N_1132,N_1058,N_1030);
and U1133 (N_1133,N_1062,N_1072);
and U1134 (N_1134,N_1066,N_1048);
and U1135 (N_1135,N_1072,N_1022);
nand U1136 (N_1136,N_1060,N_1073);
xnor U1137 (N_1137,N_1031,N_1077);
and U1138 (N_1138,N_1059,N_1045);
nand U1139 (N_1139,N_1048,N_1022);
xor U1140 (N_1140,N_1120,N_1119);
xnor U1141 (N_1141,N_1088,N_1096);
or U1142 (N_1142,N_1128,N_1130);
and U1143 (N_1143,N_1103,N_1115);
or U1144 (N_1144,N_1129,N_1097);
or U1145 (N_1145,N_1126,N_1091);
xnor U1146 (N_1146,N_1089,N_1122);
and U1147 (N_1147,N_1139,N_1102);
nand U1148 (N_1148,N_1098,N_1117);
xnor U1149 (N_1149,N_1116,N_1106);
and U1150 (N_1150,N_1092,N_1086);
xnor U1151 (N_1151,N_1111,N_1087);
xor U1152 (N_1152,N_1137,N_1124);
nor U1153 (N_1153,N_1107,N_1095);
and U1154 (N_1154,N_1082,N_1108);
or U1155 (N_1155,N_1125,N_1080);
or U1156 (N_1156,N_1100,N_1118);
nor U1157 (N_1157,N_1099,N_1112);
nor U1158 (N_1158,N_1114,N_1127);
and U1159 (N_1159,N_1136,N_1135);
xor U1160 (N_1160,N_1083,N_1134);
nand U1161 (N_1161,N_1131,N_1093);
nand U1162 (N_1162,N_1081,N_1104);
nor U1163 (N_1163,N_1094,N_1121);
nor U1164 (N_1164,N_1084,N_1085);
xnor U1165 (N_1165,N_1113,N_1133);
or U1166 (N_1166,N_1109,N_1101);
xor U1167 (N_1167,N_1123,N_1138);
nor U1168 (N_1168,N_1110,N_1090);
xnor U1169 (N_1169,N_1132,N_1105);
nor U1170 (N_1170,N_1089,N_1102);
and U1171 (N_1171,N_1098,N_1087);
or U1172 (N_1172,N_1125,N_1133);
nand U1173 (N_1173,N_1138,N_1116);
nand U1174 (N_1174,N_1108,N_1097);
nand U1175 (N_1175,N_1112,N_1089);
nor U1176 (N_1176,N_1121,N_1081);
and U1177 (N_1177,N_1119,N_1091);
nor U1178 (N_1178,N_1089,N_1107);
xnor U1179 (N_1179,N_1116,N_1111);
nand U1180 (N_1180,N_1132,N_1137);
and U1181 (N_1181,N_1089,N_1127);
xor U1182 (N_1182,N_1101,N_1122);
nor U1183 (N_1183,N_1112,N_1085);
nand U1184 (N_1184,N_1086,N_1107);
nand U1185 (N_1185,N_1089,N_1081);
nor U1186 (N_1186,N_1131,N_1105);
nor U1187 (N_1187,N_1094,N_1123);
or U1188 (N_1188,N_1130,N_1108);
nand U1189 (N_1189,N_1084,N_1137);
nand U1190 (N_1190,N_1108,N_1087);
nor U1191 (N_1191,N_1116,N_1133);
nor U1192 (N_1192,N_1133,N_1080);
nor U1193 (N_1193,N_1120,N_1103);
nor U1194 (N_1194,N_1086,N_1130);
nand U1195 (N_1195,N_1116,N_1103);
and U1196 (N_1196,N_1118,N_1138);
or U1197 (N_1197,N_1112,N_1106);
nor U1198 (N_1198,N_1088,N_1105);
and U1199 (N_1199,N_1137,N_1113);
nor U1200 (N_1200,N_1170,N_1175);
and U1201 (N_1201,N_1174,N_1166);
xor U1202 (N_1202,N_1150,N_1161);
nand U1203 (N_1203,N_1171,N_1146);
nor U1204 (N_1204,N_1158,N_1197);
and U1205 (N_1205,N_1156,N_1173);
or U1206 (N_1206,N_1167,N_1178);
nor U1207 (N_1207,N_1148,N_1194);
nor U1208 (N_1208,N_1196,N_1177);
or U1209 (N_1209,N_1169,N_1140);
and U1210 (N_1210,N_1151,N_1183);
and U1211 (N_1211,N_1188,N_1155);
and U1212 (N_1212,N_1162,N_1142);
xor U1213 (N_1213,N_1182,N_1143);
or U1214 (N_1214,N_1149,N_1186);
nand U1215 (N_1215,N_1168,N_1198);
nand U1216 (N_1216,N_1144,N_1154);
and U1217 (N_1217,N_1185,N_1187);
nor U1218 (N_1218,N_1145,N_1181);
and U1219 (N_1219,N_1180,N_1152);
nor U1220 (N_1220,N_1164,N_1184);
or U1221 (N_1221,N_1147,N_1179);
xor U1222 (N_1222,N_1189,N_1193);
xor U1223 (N_1223,N_1163,N_1192);
nor U1224 (N_1224,N_1195,N_1141);
xor U1225 (N_1225,N_1165,N_1157);
or U1226 (N_1226,N_1176,N_1153);
nand U1227 (N_1227,N_1199,N_1172);
nand U1228 (N_1228,N_1160,N_1159);
nor U1229 (N_1229,N_1191,N_1190);
nand U1230 (N_1230,N_1156,N_1192);
nand U1231 (N_1231,N_1144,N_1196);
xor U1232 (N_1232,N_1183,N_1196);
or U1233 (N_1233,N_1149,N_1195);
nor U1234 (N_1234,N_1145,N_1195);
nor U1235 (N_1235,N_1142,N_1192);
or U1236 (N_1236,N_1181,N_1156);
nor U1237 (N_1237,N_1160,N_1148);
nand U1238 (N_1238,N_1184,N_1147);
and U1239 (N_1239,N_1194,N_1152);
and U1240 (N_1240,N_1195,N_1177);
nor U1241 (N_1241,N_1177,N_1155);
nand U1242 (N_1242,N_1161,N_1145);
xor U1243 (N_1243,N_1140,N_1197);
nand U1244 (N_1244,N_1168,N_1179);
or U1245 (N_1245,N_1170,N_1159);
and U1246 (N_1246,N_1184,N_1173);
or U1247 (N_1247,N_1154,N_1165);
and U1248 (N_1248,N_1165,N_1180);
nor U1249 (N_1249,N_1195,N_1163);
or U1250 (N_1250,N_1173,N_1145);
nor U1251 (N_1251,N_1180,N_1174);
nand U1252 (N_1252,N_1199,N_1167);
nor U1253 (N_1253,N_1146,N_1165);
xnor U1254 (N_1254,N_1169,N_1163);
nor U1255 (N_1255,N_1155,N_1183);
nand U1256 (N_1256,N_1146,N_1147);
nor U1257 (N_1257,N_1198,N_1147);
nor U1258 (N_1258,N_1173,N_1141);
or U1259 (N_1259,N_1165,N_1142);
and U1260 (N_1260,N_1253,N_1210);
nor U1261 (N_1261,N_1220,N_1231);
and U1262 (N_1262,N_1205,N_1201);
xor U1263 (N_1263,N_1238,N_1219);
or U1264 (N_1264,N_1208,N_1254);
xnor U1265 (N_1265,N_1256,N_1239);
nand U1266 (N_1266,N_1243,N_1246);
nand U1267 (N_1267,N_1224,N_1222);
nand U1268 (N_1268,N_1211,N_1200);
or U1269 (N_1269,N_1218,N_1226);
nor U1270 (N_1270,N_1229,N_1241);
xnor U1271 (N_1271,N_1251,N_1202);
and U1272 (N_1272,N_1255,N_1209);
nor U1273 (N_1273,N_1221,N_1257);
nand U1274 (N_1274,N_1237,N_1204);
nand U1275 (N_1275,N_1234,N_1242);
nand U1276 (N_1276,N_1216,N_1259);
and U1277 (N_1277,N_1244,N_1225);
nor U1278 (N_1278,N_1258,N_1232);
nand U1279 (N_1279,N_1245,N_1215);
xnor U1280 (N_1280,N_1230,N_1228);
or U1281 (N_1281,N_1240,N_1207);
nand U1282 (N_1282,N_1203,N_1212);
and U1283 (N_1283,N_1249,N_1235);
xnor U1284 (N_1284,N_1248,N_1217);
xor U1285 (N_1285,N_1214,N_1236);
nand U1286 (N_1286,N_1252,N_1233);
xnor U1287 (N_1287,N_1213,N_1250);
or U1288 (N_1288,N_1227,N_1206);
nand U1289 (N_1289,N_1223,N_1247);
or U1290 (N_1290,N_1239,N_1237);
nor U1291 (N_1291,N_1242,N_1246);
nor U1292 (N_1292,N_1207,N_1219);
or U1293 (N_1293,N_1246,N_1254);
nand U1294 (N_1294,N_1221,N_1209);
or U1295 (N_1295,N_1222,N_1203);
xor U1296 (N_1296,N_1225,N_1234);
xor U1297 (N_1297,N_1221,N_1206);
and U1298 (N_1298,N_1214,N_1220);
xor U1299 (N_1299,N_1239,N_1201);
nor U1300 (N_1300,N_1252,N_1218);
nand U1301 (N_1301,N_1255,N_1238);
nand U1302 (N_1302,N_1200,N_1209);
xor U1303 (N_1303,N_1214,N_1246);
nand U1304 (N_1304,N_1229,N_1222);
xnor U1305 (N_1305,N_1211,N_1233);
xor U1306 (N_1306,N_1217,N_1219);
nor U1307 (N_1307,N_1257,N_1230);
and U1308 (N_1308,N_1231,N_1201);
xor U1309 (N_1309,N_1233,N_1238);
xor U1310 (N_1310,N_1235,N_1218);
and U1311 (N_1311,N_1237,N_1232);
nor U1312 (N_1312,N_1219,N_1237);
xor U1313 (N_1313,N_1205,N_1204);
and U1314 (N_1314,N_1218,N_1257);
xnor U1315 (N_1315,N_1234,N_1228);
or U1316 (N_1316,N_1213,N_1208);
xor U1317 (N_1317,N_1218,N_1255);
nand U1318 (N_1318,N_1218,N_1212);
nand U1319 (N_1319,N_1245,N_1233);
xnor U1320 (N_1320,N_1304,N_1270);
xnor U1321 (N_1321,N_1293,N_1268);
nor U1322 (N_1322,N_1271,N_1280);
and U1323 (N_1323,N_1262,N_1283);
nand U1324 (N_1324,N_1299,N_1263);
xnor U1325 (N_1325,N_1290,N_1286);
xnor U1326 (N_1326,N_1285,N_1296);
or U1327 (N_1327,N_1273,N_1277);
xnor U1328 (N_1328,N_1301,N_1303);
nand U1329 (N_1329,N_1316,N_1300);
and U1330 (N_1330,N_1305,N_1289);
and U1331 (N_1331,N_1306,N_1312);
or U1332 (N_1332,N_1274,N_1317);
nor U1333 (N_1333,N_1264,N_1295);
nand U1334 (N_1334,N_1261,N_1294);
and U1335 (N_1335,N_1309,N_1298);
or U1336 (N_1336,N_1287,N_1313);
nor U1337 (N_1337,N_1291,N_1310);
and U1338 (N_1338,N_1292,N_1269);
xnor U1339 (N_1339,N_1276,N_1318);
or U1340 (N_1340,N_1319,N_1260);
and U1341 (N_1341,N_1266,N_1308);
xor U1342 (N_1342,N_1315,N_1275);
nor U1343 (N_1343,N_1288,N_1279);
nand U1344 (N_1344,N_1314,N_1282);
and U1345 (N_1345,N_1297,N_1307);
xor U1346 (N_1346,N_1265,N_1302);
nand U1347 (N_1347,N_1281,N_1284);
nand U1348 (N_1348,N_1272,N_1267);
nand U1349 (N_1349,N_1278,N_1311);
or U1350 (N_1350,N_1298,N_1273);
and U1351 (N_1351,N_1281,N_1274);
xnor U1352 (N_1352,N_1282,N_1280);
xnor U1353 (N_1353,N_1318,N_1290);
nor U1354 (N_1354,N_1296,N_1307);
xnor U1355 (N_1355,N_1281,N_1305);
nor U1356 (N_1356,N_1285,N_1300);
or U1357 (N_1357,N_1276,N_1268);
nor U1358 (N_1358,N_1280,N_1269);
xnor U1359 (N_1359,N_1292,N_1309);
nor U1360 (N_1360,N_1291,N_1301);
or U1361 (N_1361,N_1316,N_1278);
or U1362 (N_1362,N_1303,N_1272);
and U1363 (N_1363,N_1265,N_1285);
nor U1364 (N_1364,N_1317,N_1314);
and U1365 (N_1365,N_1318,N_1296);
nand U1366 (N_1366,N_1303,N_1316);
and U1367 (N_1367,N_1309,N_1262);
xor U1368 (N_1368,N_1302,N_1304);
and U1369 (N_1369,N_1268,N_1287);
xnor U1370 (N_1370,N_1260,N_1300);
xor U1371 (N_1371,N_1276,N_1306);
nand U1372 (N_1372,N_1278,N_1312);
nand U1373 (N_1373,N_1316,N_1293);
xnor U1374 (N_1374,N_1314,N_1268);
xor U1375 (N_1375,N_1319,N_1271);
and U1376 (N_1376,N_1275,N_1287);
nor U1377 (N_1377,N_1289,N_1315);
nor U1378 (N_1378,N_1278,N_1272);
xor U1379 (N_1379,N_1269,N_1312);
and U1380 (N_1380,N_1355,N_1344);
nor U1381 (N_1381,N_1370,N_1360);
and U1382 (N_1382,N_1333,N_1377);
nand U1383 (N_1383,N_1369,N_1363);
nor U1384 (N_1384,N_1329,N_1375);
and U1385 (N_1385,N_1320,N_1335);
nor U1386 (N_1386,N_1366,N_1350);
xor U1387 (N_1387,N_1345,N_1374);
nor U1388 (N_1388,N_1361,N_1372);
or U1389 (N_1389,N_1376,N_1368);
nor U1390 (N_1390,N_1354,N_1327);
xnor U1391 (N_1391,N_1356,N_1353);
nor U1392 (N_1392,N_1379,N_1347);
nor U1393 (N_1393,N_1351,N_1346);
nand U1394 (N_1394,N_1334,N_1362);
and U1395 (N_1395,N_1326,N_1359);
nand U1396 (N_1396,N_1328,N_1340);
or U1397 (N_1397,N_1339,N_1341);
nor U1398 (N_1398,N_1325,N_1371);
and U1399 (N_1399,N_1373,N_1323);
and U1400 (N_1400,N_1324,N_1332);
nor U1401 (N_1401,N_1358,N_1357);
and U1402 (N_1402,N_1352,N_1321);
or U1403 (N_1403,N_1337,N_1336);
or U1404 (N_1404,N_1378,N_1330);
xor U1405 (N_1405,N_1367,N_1365);
xor U1406 (N_1406,N_1322,N_1364);
or U1407 (N_1407,N_1349,N_1342);
nand U1408 (N_1408,N_1331,N_1343);
nor U1409 (N_1409,N_1338,N_1348);
nor U1410 (N_1410,N_1347,N_1341);
xnor U1411 (N_1411,N_1365,N_1362);
xor U1412 (N_1412,N_1324,N_1325);
xnor U1413 (N_1413,N_1323,N_1350);
nand U1414 (N_1414,N_1347,N_1335);
and U1415 (N_1415,N_1372,N_1320);
and U1416 (N_1416,N_1333,N_1360);
xnor U1417 (N_1417,N_1372,N_1332);
or U1418 (N_1418,N_1342,N_1366);
xnor U1419 (N_1419,N_1375,N_1363);
nand U1420 (N_1420,N_1342,N_1345);
nand U1421 (N_1421,N_1369,N_1347);
nand U1422 (N_1422,N_1335,N_1328);
xor U1423 (N_1423,N_1335,N_1365);
nand U1424 (N_1424,N_1322,N_1368);
nand U1425 (N_1425,N_1337,N_1362);
and U1426 (N_1426,N_1361,N_1330);
nor U1427 (N_1427,N_1357,N_1320);
nor U1428 (N_1428,N_1368,N_1366);
and U1429 (N_1429,N_1344,N_1357);
xnor U1430 (N_1430,N_1321,N_1372);
or U1431 (N_1431,N_1335,N_1369);
or U1432 (N_1432,N_1359,N_1344);
nand U1433 (N_1433,N_1373,N_1378);
or U1434 (N_1434,N_1320,N_1374);
and U1435 (N_1435,N_1334,N_1340);
nor U1436 (N_1436,N_1348,N_1351);
xnor U1437 (N_1437,N_1355,N_1373);
nand U1438 (N_1438,N_1368,N_1345);
and U1439 (N_1439,N_1363,N_1326);
nor U1440 (N_1440,N_1423,N_1392);
xnor U1441 (N_1441,N_1386,N_1430);
and U1442 (N_1442,N_1398,N_1432);
nor U1443 (N_1443,N_1435,N_1418);
nand U1444 (N_1444,N_1391,N_1407);
nand U1445 (N_1445,N_1401,N_1381);
and U1446 (N_1446,N_1417,N_1404);
xor U1447 (N_1447,N_1439,N_1406);
or U1448 (N_1448,N_1411,N_1410);
nor U1449 (N_1449,N_1408,N_1403);
xor U1450 (N_1450,N_1389,N_1426);
nor U1451 (N_1451,N_1420,N_1436);
nand U1452 (N_1452,N_1390,N_1425);
or U1453 (N_1453,N_1429,N_1393);
nand U1454 (N_1454,N_1431,N_1382);
nor U1455 (N_1455,N_1412,N_1383);
and U1456 (N_1456,N_1413,N_1400);
nor U1457 (N_1457,N_1409,N_1422);
xor U1458 (N_1458,N_1419,N_1387);
nor U1459 (N_1459,N_1434,N_1384);
or U1460 (N_1460,N_1415,N_1416);
xnor U1461 (N_1461,N_1414,N_1399);
or U1462 (N_1462,N_1428,N_1427);
xnor U1463 (N_1463,N_1397,N_1380);
and U1464 (N_1464,N_1437,N_1385);
xor U1465 (N_1465,N_1438,N_1421);
nor U1466 (N_1466,N_1395,N_1388);
nand U1467 (N_1467,N_1405,N_1424);
and U1468 (N_1468,N_1396,N_1433);
and U1469 (N_1469,N_1402,N_1394);
or U1470 (N_1470,N_1414,N_1432);
and U1471 (N_1471,N_1390,N_1406);
nand U1472 (N_1472,N_1400,N_1414);
xor U1473 (N_1473,N_1428,N_1385);
xnor U1474 (N_1474,N_1402,N_1404);
and U1475 (N_1475,N_1396,N_1407);
and U1476 (N_1476,N_1419,N_1420);
and U1477 (N_1477,N_1434,N_1389);
nor U1478 (N_1478,N_1400,N_1405);
nor U1479 (N_1479,N_1410,N_1421);
or U1480 (N_1480,N_1402,N_1415);
and U1481 (N_1481,N_1426,N_1384);
and U1482 (N_1482,N_1394,N_1435);
xor U1483 (N_1483,N_1396,N_1415);
nor U1484 (N_1484,N_1381,N_1390);
or U1485 (N_1485,N_1433,N_1435);
and U1486 (N_1486,N_1430,N_1383);
nand U1487 (N_1487,N_1395,N_1404);
nor U1488 (N_1488,N_1431,N_1411);
and U1489 (N_1489,N_1439,N_1385);
xnor U1490 (N_1490,N_1412,N_1404);
xor U1491 (N_1491,N_1391,N_1388);
and U1492 (N_1492,N_1401,N_1397);
or U1493 (N_1493,N_1435,N_1430);
xor U1494 (N_1494,N_1429,N_1430);
and U1495 (N_1495,N_1432,N_1435);
nor U1496 (N_1496,N_1430,N_1415);
and U1497 (N_1497,N_1383,N_1410);
nand U1498 (N_1498,N_1401,N_1422);
and U1499 (N_1499,N_1419,N_1382);
xor U1500 (N_1500,N_1497,N_1455);
or U1501 (N_1501,N_1492,N_1460);
and U1502 (N_1502,N_1468,N_1490);
and U1503 (N_1503,N_1463,N_1484);
or U1504 (N_1504,N_1486,N_1465);
xnor U1505 (N_1505,N_1440,N_1444);
nand U1506 (N_1506,N_1472,N_1443);
and U1507 (N_1507,N_1451,N_1489);
and U1508 (N_1508,N_1488,N_1446);
nor U1509 (N_1509,N_1485,N_1473);
and U1510 (N_1510,N_1464,N_1493);
xor U1511 (N_1511,N_1442,N_1498);
xnor U1512 (N_1512,N_1494,N_1441);
nand U1513 (N_1513,N_1457,N_1479);
and U1514 (N_1514,N_1459,N_1454);
or U1515 (N_1515,N_1483,N_1458);
nor U1516 (N_1516,N_1480,N_1456);
xor U1517 (N_1517,N_1448,N_1469);
or U1518 (N_1518,N_1474,N_1453);
or U1519 (N_1519,N_1449,N_1471);
and U1520 (N_1520,N_1475,N_1466);
and U1521 (N_1521,N_1477,N_1495);
xor U1522 (N_1522,N_1467,N_1452);
nand U1523 (N_1523,N_1450,N_1496);
nor U1524 (N_1524,N_1487,N_1461);
and U1525 (N_1525,N_1478,N_1481);
and U1526 (N_1526,N_1470,N_1445);
and U1527 (N_1527,N_1499,N_1476);
and U1528 (N_1528,N_1462,N_1482);
nor U1529 (N_1529,N_1447,N_1491);
or U1530 (N_1530,N_1489,N_1472);
xor U1531 (N_1531,N_1494,N_1479);
nor U1532 (N_1532,N_1468,N_1451);
nor U1533 (N_1533,N_1454,N_1456);
and U1534 (N_1534,N_1498,N_1449);
xor U1535 (N_1535,N_1456,N_1465);
xor U1536 (N_1536,N_1442,N_1472);
and U1537 (N_1537,N_1450,N_1469);
nand U1538 (N_1538,N_1482,N_1490);
or U1539 (N_1539,N_1484,N_1442);
xnor U1540 (N_1540,N_1484,N_1472);
and U1541 (N_1541,N_1448,N_1478);
and U1542 (N_1542,N_1464,N_1498);
and U1543 (N_1543,N_1448,N_1483);
nor U1544 (N_1544,N_1480,N_1469);
or U1545 (N_1545,N_1488,N_1478);
and U1546 (N_1546,N_1461,N_1485);
or U1547 (N_1547,N_1462,N_1447);
and U1548 (N_1548,N_1476,N_1460);
xnor U1549 (N_1549,N_1499,N_1446);
nor U1550 (N_1550,N_1446,N_1477);
xor U1551 (N_1551,N_1455,N_1491);
and U1552 (N_1552,N_1496,N_1455);
and U1553 (N_1553,N_1445,N_1460);
or U1554 (N_1554,N_1483,N_1471);
nor U1555 (N_1555,N_1440,N_1450);
nor U1556 (N_1556,N_1447,N_1464);
xor U1557 (N_1557,N_1470,N_1496);
nor U1558 (N_1558,N_1497,N_1481);
xnor U1559 (N_1559,N_1488,N_1492);
nor U1560 (N_1560,N_1511,N_1509);
xnor U1561 (N_1561,N_1559,N_1522);
nand U1562 (N_1562,N_1533,N_1500);
or U1563 (N_1563,N_1534,N_1526);
nand U1564 (N_1564,N_1540,N_1515);
and U1565 (N_1565,N_1553,N_1524);
and U1566 (N_1566,N_1537,N_1546);
nand U1567 (N_1567,N_1527,N_1512);
nor U1568 (N_1568,N_1556,N_1513);
nor U1569 (N_1569,N_1508,N_1528);
xor U1570 (N_1570,N_1504,N_1501);
or U1571 (N_1571,N_1521,N_1503);
nand U1572 (N_1572,N_1536,N_1514);
and U1573 (N_1573,N_1550,N_1523);
xnor U1574 (N_1574,N_1545,N_1510);
or U1575 (N_1575,N_1518,N_1554);
nor U1576 (N_1576,N_1530,N_1543);
and U1577 (N_1577,N_1519,N_1531);
xor U1578 (N_1578,N_1529,N_1542);
or U1579 (N_1579,N_1548,N_1547);
or U1580 (N_1580,N_1538,N_1551);
nand U1581 (N_1581,N_1557,N_1544);
xor U1582 (N_1582,N_1558,N_1541);
and U1583 (N_1583,N_1506,N_1539);
or U1584 (N_1584,N_1549,N_1505);
and U1585 (N_1585,N_1516,N_1502);
or U1586 (N_1586,N_1555,N_1517);
xor U1587 (N_1587,N_1532,N_1552);
and U1588 (N_1588,N_1507,N_1525);
or U1589 (N_1589,N_1520,N_1535);
xor U1590 (N_1590,N_1520,N_1557);
and U1591 (N_1591,N_1525,N_1528);
xnor U1592 (N_1592,N_1510,N_1539);
or U1593 (N_1593,N_1509,N_1547);
and U1594 (N_1594,N_1509,N_1516);
and U1595 (N_1595,N_1541,N_1509);
or U1596 (N_1596,N_1540,N_1554);
xnor U1597 (N_1597,N_1516,N_1538);
nor U1598 (N_1598,N_1536,N_1551);
and U1599 (N_1599,N_1557,N_1516);
or U1600 (N_1600,N_1509,N_1542);
nand U1601 (N_1601,N_1558,N_1513);
or U1602 (N_1602,N_1533,N_1506);
and U1603 (N_1603,N_1551,N_1506);
or U1604 (N_1604,N_1504,N_1502);
xnor U1605 (N_1605,N_1553,N_1532);
and U1606 (N_1606,N_1520,N_1544);
nor U1607 (N_1607,N_1534,N_1542);
nor U1608 (N_1608,N_1503,N_1549);
xnor U1609 (N_1609,N_1504,N_1548);
xor U1610 (N_1610,N_1520,N_1553);
xnor U1611 (N_1611,N_1546,N_1502);
nor U1612 (N_1612,N_1506,N_1518);
and U1613 (N_1613,N_1534,N_1506);
or U1614 (N_1614,N_1546,N_1549);
nor U1615 (N_1615,N_1520,N_1527);
and U1616 (N_1616,N_1557,N_1508);
nor U1617 (N_1617,N_1527,N_1537);
nor U1618 (N_1618,N_1540,N_1533);
xor U1619 (N_1619,N_1530,N_1549);
nand U1620 (N_1620,N_1588,N_1592);
xor U1621 (N_1621,N_1574,N_1583);
nor U1622 (N_1622,N_1585,N_1614);
and U1623 (N_1623,N_1598,N_1569);
nand U1624 (N_1624,N_1566,N_1613);
nor U1625 (N_1625,N_1595,N_1608);
xor U1626 (N_1626,N_1611,N_1603);
xor U1627 (N_1627,N_1571,N_1573);
nor U1628 (N_1628,N_1577,N_1560);
nand U1629 (N_1629,N_1582,N_1580);
or U1630 (N_1630,N_1581,N_1572);
and U1631 (N_1631,N_1570,N_1586);
nor U1632 (N_1632,N_1562,N_1590);
and U1633 (N_1633,N_1619,N_1578);
xnor U1634 (N_1634,N_1616,N_1596);
nor U1635 (N_1635,N_1593,N_1564);
nor U1636 (N_1636,N_1612,N_1605);
nor U1637 (N_1637,N_1579,N_1615);
nand U1638 (N_1638,N_1587,N_1607);
nor U1639 (N_1639,N_1563,N_1604);
or U1640 (N_1640,N_1601,N_1617);
or U1641 (N_1641,N_1589,N_1567);
xor U1642 (N_1642,N_1602,N_1597);
nand U1643 (N_1643,N_1561,N_1610);
nor U1644 (N_1644,N_1576,N_1568);
xnor U1645 (N_1645,N_1606,N_1575);
nor U1646 (N_1646,N_1591,N_1565);
nor U1647 (N_1647,N_1600,N_1594);
nand U1648 (N_1648,N_1599,N_1584);
or U1649 (N_1649,N_1609,N_1618);
nand U1650 (N_1650,N_1611,N_1610);
and U1651 (N_1651,N_1567,N_1618);
or U1652 (N_1652,N_1565,N_1597);
and U1653 (N_1653,N_1594,N_1565);
nor U1654 (N_1654,N_1606,N_1560);
and U1655 (N_1655,N_1570,N_1567);
or U1656 (N_1656,N_1576,N_1575);
and U1657 (N_1657,N_1601,N_1605);
or U1658 (N_1658,N_1605,N_1615);
xor U1659 (N_1659,N_1588,N_1587);
nand U1660 (N_1660,N_1585,N_1583);
nand U1661 (N_1661,N_1609,N_1579);
nand U1662 (N_1662,N_1588,N_1561);
nand U1663 (N_1663,N_1606,N_1600);
and U1664 (N_1664,N_1608,N_1594);
xnor U1665 (N_1665,N_1570,N_1579);
nand U1666 (N_1666,N_1590,N_1591);
or U1667 (N_1667,N_1589,N_1569);
nand U1668 (N_1668,N_1593,N_1585);
nand U1669 (N_1669,N_1618,N_1579);
and U1670 (N_1670,N_1575,N_1562);
nand U1671 (N_1671,N_1595,N_1578);
xnor U1672 (N_1672,N_1586,N_1563);
xnor U1673 (N_1673,N_1598,N_1615);
xor U1674 (N_1674,N_1578,N_1596);
xor U1675 (N_1675,N_1571,N_1578);
xnor U1676 (N_1676,N_1597,N_1585);
nor U1677 (N_1677,N_1571,N_1569);
or U1678 (N_1678,N_1591,N_1594);
xnor U1679 (N_1679,N_1590,N_1598);
xor U1680 (N_1680,N_1677,N_1664);
xnor U1681 (N_1681,N_1621,N_1662);
nand U1682 (N_1682,N_1669,N_1646);
nand U1683 (N_1683,N_1625,N_1673);
xnor U1684 (N_1684,N_1626,N_1630);
nor U1685 (N_1685,N_1657,N_1635);
nor U1686 (N_1686,N_1656,N_1676);
xnor U1687 (N_1687,N_1661,N_1620);
nand U1688 (N_1688,N_1629,N_1674);
nor U1689 (N_1689,N_1670,N_1652);
nor U1690 (N_1690,N_1639,N_1647);
nor U1691 (N_1691,N_1643,N_1651);
and U1692 (N_1692,N_1667,N_1632);
xor U1693 (N_1693,N_1679,N_1660);
xnor U1694 (N_1694,N_1678,N_1636);
or U1695 (N_1695,N_1644,N_1655);
and U1696 (N_1696,N_1638,N_1653);
or U1697 (N_1697,N_1665,N_1658);
nand U1698 (N_1698,N_1648,N_1623);
xnor U1699 (N_1699,N_1672,N_1671);
nand U1700 (N_1700,N_1633,N_1663);
nor U1701 (N_1701,N_1627,N_1634);
and U1702 (N_1702,N_1640,N_1666);
nand U1703 (N_1703,N_1628,N_1668);
or U1704 (N_1704,N_1641,N_1654);
nor U1705 (N_1705,N_1675,N_1624);
nand U1706 (N_1706,N_1637,N_1659);
or U1707 (N_1707,N_1645,N_1631);
or U1708 (N_1708,N_1622,N_1642);
nand U1709 (N_1709,N_1649,N_1650);
and U1710 (N_1710,N_1670,N_1631);
nand U1711 (N_1711,N_1667,N_1661);
or U1712 (N_1712,N_1635,N_1634);
and U1713 (N_1713,N_1675,N_1679);
and U1714 (N_1714,N_1632,N_1678);
nand U1715 (N_1715,N_1620,N_1675);
xnor U1716 (N_1716,N_1652,N_1633);
or U1717 (N_1717,N_1655,N_1624);
or U1718 (N_1718,N_1643,N_1635);
xnor U1719 (N_1719,N_1646,N_1649);
xnor U1720 (N_1720,N_1627,N_1641);
xnor U1721 (N_1721,N_1633,N_1662);
xor U1722 (N_1722,N_1677,N_1640);
nor U1723 (N_1723,N_1666,N_1662);
nor U1724 (N_1724,N_1662,N_1634);
or U1725 (N_1725,N_1666,N_1643);
nand U1726 (N_1726,N_1660,N_1623);
nor U1727 (N_1727,N_1657,N_1623);
nor U1728 (N_1728,N_1632,N_1644);
and U1729 (N_1729,N_1670,N_1677);
nand U1730 (N_1730,N_1632,N_1641);
nor U1731 (N_1731,N_1632,N_1653);
xor U1732 (N_1732,N_1638,N_1647);
nor U1733 (N_1733,N_1646,N_1637);
and U1734 (N_1734,N_1637,N_1677);
nand U1735 (N_1735,N_1624,N_1679);
xor U1736 (N_1736,N_1658,N_1674);
and U1737 (N_1737,N_1632,N_1626);
xnor U1738 (N_1738,N_1661,N_1672);
or U1739 (N_1739,N_1658,N_1664);
xor U1740 (N_1740,N_1687,N_1705);
nor U1741 (N_1741,N_1697,N_1688);
xor U1742 (N_1742,N_1704,N_1690);
nand U1743 (N_1743,N_1739,N_1732);
nand U1744 (N_1744,N_1699,N_1680);
or U1745 (N_1745,N_1736,N_1713);
or U1746 (N_1746,N_1708,N_1737);
xor U1747 (N_1747,N_1714,N_1683);
xor U1748 (N_1748,N_1720,N_1716);
nand U1749 (N_1749,N_1681,N_1684);
and U1750 (N_1750,N_1682,N_1695);
nand U1751 (N_1751,N_1733,N_1724);
or U1752 (N_1752,N_1731,N_1700);
nand U1753 (N_1753,N_1735,N_1717);
xor U1754 (N_1754,N_1712,N_1718);
and U1755 (N_1755,N_1711,N_1728);
xor U1756 (N_1756,N_1722,N_1685);
or U1757 (N_1757,N_1721,N_1702);
and U1758 (N_1758,N_1715,N_1701);
and U1759 (N_1759,N_1725,N_1706);
nor U1760 (N_1760,N_1696,N_1707);
nor U1761 (N_1761,N_1738,N_1734);
nand U1762 (N_1762,N_1723,N_1689);
or U1763 (N_1763,N_1710,N_1729);
nand U1764 (N_1764,N_1698,N_1726);
xor U1765 (N_1765,N_1692,N_1686);
or U1766 (N_1766,N_1693,N_1730);
nor U1767 (N_1767,N_1709,N_1694);
or U1768 (N_1768,N_1691,N_1727);
and U1769 (N_1769,N_1719,N_1703);
nor U1770 (N_1770,N_1714,N_1680);
or U1771 (N_1771,N_1739,N_1687);
xor U1772 (N_1772,N_1681,N_1701);
xnor U1773 (N_1773,N_1703,N_1732);
xnor U1774 (N_1774,N_1720,N_1693);
xor U1775 (N_1775,N_1696,N_1701);
or U1776 (N_1776,N_1684,N_1711);
xor U1777 (N_1777,N_1688,N_1739);
nor U1778 (N_1778,N_1689,N_1691);
and U1779 (N_1779,N_1714,N_1710);
nor U1780 (N_1780,N_1700,N_1712);
nand U1781 (N_1781,N_1695,N_1696);
xnor U1782 (N_1782,N_1686,N_1680);
nand U1783 (N_1783,N_1727,N_1725);
and U1784 (N_1784,N_1706,N_1718);
nor U1785 (N_1785,N_1724,N_1691);
nor U1786 (N_1786,N_1683,N_1689);
and U1787 (N_1787,N_1687,N_1689);
xor U1788 (N_1788,N_1739,N_1738);
or U1789 (N_1789,N_1684,N_1693);
xnor U1790 (N_1790,N_1684,N_1710);
and U1791 (N_1791,N_1711,N_1696);
xor U1792 (N_1792,N_1689,N_1722);
or U1793 (N_1793,N_1735,N_1696);
nand U1794 (N_1794,N_1716,N_1693);
nor U1795 (N_1795,N_1738,N_1723);
nand U1796 (N_1796,N_1697,N_1691);
xnor U1797 (N_1797,N_1713,N_1691);
nor U1798 (N_1798,N_1712,N_1685);
nor U1799 (N_1799,N_1736,N_1701);
and U1800 (N_1800,N_1794,N_1780);
nand U1801 (N_1801,N_1751,N_1758);
xor U1802 (N_1802,N_1777,N_1752);
nor U1803 (N_1803,N_1768,N_1767);
and U1804 (N_1804,N_1742,N_1798);
and U1805 (N_1805,N_1796,N_1782);
xor U1806 (N_1806,N_1792,N_1781);
and U1807 (N_1807,N_1771,N_1764);
and U1808 (N_1808,N_1799,N_1743);
nor U1809 (N_1809,N_1749,N_1740);
xnor U1810 (N_1810,N_1754,N_1773);
or U1811 (N_1811,N_1783,N_1759);
xor U1812 (N_1812,N_1763,N_1776);
nand U1813 (N_1813,N_1795,N_1772);
nor U1814 (N_1814,N_1774,N_1761);
nand U1815 (N_1815,N_1793,N_1779);
or U1816 (N_1816,N_1787,N_1750);
and U1817 (N_1817,N_1770,N_1762);
nand U1818 (N_1818,N_1756,N_1788);
xor U1819 (N_1819,N_1747,N_1785);
and U1820 (N_1820,N_1766,N_1791);
nor U1821 (N_1821,N_1748,N_1755);
nor U1822 (N_1822,N_1790,N_1789);
xnor U1823 (N_1823,N_1745,N_1784);
nor U1824 (N_1824,N_1741,N_1746);
or U1825 (N_1825,N_1769,N_1797);
or U1826 (N_1826,N_1757,N_1753);
nor U1827 (N_1827,N_1786,N_1744);
nor U1828 (N_1828,N_1760,N_1778);
and U1829 (N_1829,N_1775,N_1765);
xor U1830 (N_1830,N_1796,N_1752);
xor U1831 (N_1831,N_1766,N_1798);
nor U1832 (N_1832,N_1751,N_1781);
xor U1833 (N_1833,N_1755,N_1744);
or U1834 (N_1834,N_1772,N_1789);
nor U1835 (N_1835,N_1799,N_1794);
nand U1836 (N_1836,N_1771,N_1795);
or U1837 (N_1837,N_1785,N_1763);
nor U1838 (N_1838,N_1778,N_1749);
or U1839 (N_1839,N_1758,N_1760);
nor U1840 (N_1840,N_1744,N_1766);
and U1841 (N_1841,N_1775,N_1794);
or U1842 (N_1842,N_1768,N_1784);
and U1843 (N_1843,N_1782,N_1798);
nand U1844 (N_1844,N_1749,N_1746);
and U1845 (N_1845,N_1793,N_1754);
or U1846 (N_1846,N_1743,N_1775);
nand U1847 (N_1847,N_1769,N_1795);
nand U1848 (N_1848,N_1773,N_1794);
and U1849 (N_1849,N_1796,N_1750);
nand U1850 (N_1850,N_1752,N_1761);
nor U1851 (N_1851,N_1761,N_1796);
or U1852 (N_1852,N_1741,N_1795);
nor U1853 (N_1853,N_1750,N_1783);
xor U1854 (N_1854,N_1752,N_1769);
nor U1855 (N_1855,N_1743,N_1770);
nor U1856 (N_1856,N_1751,N_1791);
xnor U1857 (N_1857,N_1761,N_1745);
nor U1858 (N_1858,N_1797,N_1767);
or U1859 (N_1859,N_1756,N_1748);
xnor U1860 (N_1860,N_1846,N_1819);
nand U1861 (N_1861,N_1854,N_1815);
nand U1862 (N_1862,N_1805,N_1829);
nand U1863 (N_1863,N_1824,N_1850);
xnor U1864 (N_1864,N_1844,N_1807);
xor U1865 (N_1865,N_1823,N_1848);
and U1866 (N_1866,N_1813,N_1826);
nor U1867 (N_1867,N_1858,N_1810);
nor U1868 (N_1868,N_1801,N_1821);
nand U1869 (N_1869,N_1840,N_1835);
nand U1870 (N_1870,N_1841,N_1837);
or U1871 (N_1871,N_1806,N_1847);
nor U1872 (N_1872,N_1852,N_1849);
nor U1873 (N_1873,N_1831,N_1842);
or U1874 (N_1874,N_1839,N_1836);
xnor U1875 (N_1875,N_1857,N_1800);
and U1876 (N_1876,N_1851,N_1830);
or U1877 (N_1877,N_1845,N_1820);
and U1878 (N_1878,N_1833,N_1818);
or U1879 (N_1879,N_1812,N_1803);
xnor U1880 (N_1880,N_1804,N_1838);
and U1881 (N_1881,N_1834,N_1808);
or U1882 (N_1882,N_1855,N_1832);
nand U1883 (N_1883,N_1827,N_1828);
xnor U1884 (N_1884,N_1859,N_1802);
or U1885 (N_1885,N_1853,N_1825);
nand U1886 (N_1886,N_1817,N_1811);
nand U1887 (N_1887,N_1814,N_1809);
and U1888 (N_1888,N_1843,N_1822);
nand U1889 (N_1889,N_1816,N_1856);
xor U1890 (N_1890,N_1849,N_1822);
and U1891 (N_1891,N_1832,N_1821);
and U1892 (N_1892,N_1817,N_1818);
nor U1893 (N_1893,N_1856,N_1833);
nor U1894 (N_1894,N_1839,N_1826);
nand U1895 (N_1895,N_1820,N_1804);
and U1896 (N_1896,N_1834,N_1801);
xnor U1897 (N_1897,N_1813,N_1806);
nor U1898 (N_1898,N_1809,N_1832);
or U1899 (N_1899,N_1804,N_1837);
and U1900 (N_1900,N_1827,N_1854);
xnor U1901 (N_1901,N_1853,N_1833);
nor U1902 (N_1902,N_1847,N_1836);
or U1903 (N_1903,N_1821,N_1825);
or U1904 (N_1904,N_1818,N_1852);
or U1905 (N_1905,N_1830,N_1859);
or U1906 (N_1906,N_1850,N_1852);
xor U1907 (N_1907,N_1832,N_1849);
and U1908 (N_1908,N_1850,N_1829);
or U1909 (N_1909,N_1807,N_1838);
xor U1910 (N_1910,N_1850,N_1818);
nor U1911 (N_1911,N_1806,N_1830);
nand U1912 (N_1912,N_1822,N_1820);
nand U1913 (N_1913,N_1805,N_1812);
nor U1914 (N_1914,N_1825,N_1808);
nand U1915 (N_1915,N_1827,N_1811);
nand U1916 (N_1916,N_1819,N_1859);
or U1917 (N_1917,N_1858,N_1838);
nor U1918 (N_1918,N_1806,N_1851);
and U1919 (N_1919,N_1817,N_1806);
nand U1920 (N_1920,N_1893,N_1904);
nor U1921 (N_1921,N_1872,N_1886);
xnor U1922 (N_1922,N_1860,N_1883);
nor U1923 (N_1923,N_1877,N_1888);
xor U1924 (N_1924,N_1891,N_1876);
xor U1925 (N_1925,N_1884,N_1890);
or U1926 (N_1926,N_1913,N_1885);
xnor U1927 (N_1927,N_1879,N_1896);
or U1928 (N_1928,N_1869,N_1894);
or U1929 (N_1929,N_1916,N_1887);
nand U1930 (N_1930,N_1919,N_1902);
or U1931 (N_1931,N_1863,N_1912);
and U1932 (N_1932,N_1905,N_1903);
and U1933 (N_1933,N_1865,N_1909);
nand U1934 (N_1934,N_1908,N_1901);
nand U1935 (N_1935,N_1898,N_1914);
xor U1936 (N_1936,N_1917,N_1862);
xnor U1937 (N_1937,N_1866,N_1892);
nand U1938 (N_1938,N_1889,N_1910);
xor U1939 (N_1939,N_1918,N_1880);
xnor U1940 (N_1940,N_1864,N_1897);
xnor U1941 (N_1941,N_1878,N_1873);
nor U1942 (N_1942,N_1861,N_1881);
and U1943 (N_1943,N_1907,N_1906);
xor U1944 (N_1944,N_1875,N_1895);
nand U1945 (N_1945,N_1868,N_1915);
nand U1946 (N_1946,N_1900,N_1867);
nor U1947 (N_1947,N_1911,N_1871);
nand U1948 (N_1948,N_1882,N_1874);
nor U1949 (N_1949,N_1899,N_1870);
xor U1950 (N_1950,N_1880,N_1904);
xnor U1951 (N_1951,N_1863,N_1884);
xnor U1952 (N_1952,N_1891,N_1900);
nand U1953 (N_1953,N_1878,N_1912);
or U1954 (N_1954,N_1900,N_1912);
nand U1955 (N_1955,N_1887,N_1893);
xnor U1956 (N_1956,N_1900,N_1896);
xor U1957 (N_1957,N_1888,N_1902);
nand U1958 (N_1958,N_1917,N_1899);
nand U1959 (N_1959,N_1869,N_1879);
nor U1960 (N_1960,N_1882,N_1891);
xnor U1961 (N_1961,N_1892,N_1877);
or U1962 (N_1962,N_1913,N_1886);
or U1963 (N_1963,N_1868,N_1862);
xor U1964 (N_1964,N_1910,N_1888);
nand U1965 (N_1965,N_1898,N_1891);
or U1966 (N_1966,N_1883,N_1870);
and U1967 (N_1967,N_1860,N_1864);
xnor U1968 (N_1968,N_1908,N_1871);
nor U1969 (N_1969,N_1919,N_1874);
and U1970 (N_1970,N_1879,N_1881);
nand U1971 (N_1971,N_1877,N_1904);
xor U1972 (N_1972,N_1907,N_1894);
xor U1973 (N_1973,N_1864,N_1895);
and U1974 (N_1974,N_1901,N_1870);
or U1975 (N_1975,N_1918,N_1897);
and U1976 (N_1976,N_1860,N_1910);
xnor U1977 (N_1977,N_1895,N_1907);
or U1978 (N_1978,N_1874,N_1894);
xor U1979 (N_1979,N_1883,N_1919);
or U1980 (N_1980,N_1946,N_1922);
nand U1981 (N_1981,N_1920,N_1947);
nand U1982 (N_1982,N_1940,N_1978);
or U1983 (N_1983,N_1964,N_1973);
and U1984 (N_1984,N_1969,N_1933);
nor U1985 (N_1985,N_1935,N_1953);
nand U1986 (N_1986,N_1932,N_1948);
and U1987 (N_1987,N_1921,N_1923);
xnor U1988 (N_1988,N_1941,N_1967);
xor U1989 (N_1989,N_1950,N_1958);
and U1990 (N_1990,N_1936,N_1979);
or U1991 (N_1991,N_1942,N_1951);
and U1992 (N_1992,N_1970,N_1930);
xor U1993 (N_1993,N_1959,N_1968);
xor U1994 (N_1994,N_1928,N_1957);
and U1995 (N_1995,N_1974,N_1961);
nor U1996 (N_1996,N_1934,N_1943);
nor U1997 (N_1997,N_1963,N_1952);
nor U1998 (N_1998,N_1965,N_1945);
nor U1999 (N_1999,N_1927,N_1962);
and U2000 (N_2000,N_1944,N_1972);
xnor U2001 (N_2001,N_1966,N_1975);
nand U2002 (N_2002,N_1937,N_1939);
or U2003 (N_2003,N_1931,N_1949);
and U2004 (N_2004,N_1971,N_1938);
and U2005 (N_2005,N_1926,N_1977);
and U2006 (N_2006,N_1960,N_1954);
xor U2007 (N_2007,N_1924,N_1925);
xnor U2008 (N_2008,N_1955,N_1976);
or U2009 (N_2009,N_1956,N_1929);
nor U2010 (N_2010,N_1933,N_1963);
and U2011 (N_2011,N_1920,N_1976);
nand U2012 (N_2012,N_1947,N_1928);
or U2013 (N_2013,N_1936,N_1956);
xor U2014 (N_2014,N_1940,N_1962);
and U2015 (N_2015,N_1967,N_1930);
xnor U2016 (N_2016,N_1936,N_1950);
nand U2017 (N_2017,N_1953,N_1929);
xor U2018 (N_2018,N_1922,N_1941);
and U2019 (N_2019,N_1949,N_1928);
or U2020 (N_2020,N_1975,N_1942);
or U2021 (N_2021,N_1952,N_1946);
nand U2022 (N_2022,N_1972,N_1941);
xnor U2023 (N_2023,N_1969,N_1937);
nand U2024 (N_2024,N_1930,N_1950);
and U2025 (N_2025,N_1964,N_1931);
nor U2026 (N_2026,N_1961,N_1933);
nand U2027 (N_2027,N_1971,N_1969);
xnor U2028 (N_2028,N_1945,N_1938);
and U2029 (N_2029,N_1930,N_1954);
or U2030 (N_2030,N_1934,N_1973);
xnor U2031 (N_2031,N_1942,N_1924);
and U2032 (N_2032,N_1926,N_1943);
or U2033 (N_2033,N_1971,N_1948);
nand U2034 (N_2034,N_1964,N_1953);
and U2035 (N_2035,N_1923,N_1941);
nor U2036 (N_2036,N_1959,N_1966);
and U2037 (N_2037,N_1935,N_1941);
xnor U2038 (N_2038,N_1958,N_1923);
xor U2039 (N_2039,N_1979,N_1974);
and U2040 (N_2040,N_1980,N_2013);
or U2041 (N_2041,N_2032,N_1987);
and U2042 (N_2042,N_2038,N_2039);
and U2043 (N_2043,N_2020,N_2036);
nand U2044 (N_2044,N_1985,N_1994);
and U2045 (N_2045,N_1988,N_2012);
nor U2046 (N_2046,N_2027,N_2023);
nor U2047 (N_2047,N_2009,N_1984);
nor U2048 (N_2048,N_1981,N_2014);
or U2049 (N_2049,N_2019,N_2029);
nor U2050 (N_2050,N_1996,N_1993);
nand U2051 (N_2051,N_1986,N_1983);
nor U2052 (N_2052,N_1992,N_2021);
or U2053 (N_2053,N_2031,N_2022);
or U2054 (N_2054,N_2024,N_1997);
xnor U2055 (N_2055,N_2030,N_2008);
xor U2056 (N_2056,N_2003,N_2010);
or U2057 (N_2057,N_1989,N_2025);
and U2058 (N_2058,N_2028,N_2011);
nand U2059 (N_2059,N_2035,N_1982);
nand U2060 (N_2060,N_2034,N_2007);
nor U2061 (N_2061,N_1990,N_2000);
or U2062 (N_2062,N_1995,N_2018);
or U2063 (N_2063,N_2033,N_2015);
nand U2064 (N_2064,N_2006,N_2037);
nor U2065 (N_2065,N_2017,N_1991);
or U2066 (N_2066,N_1999,N_2002);
xor U2067 (N_2067,N_2026,N_2004);
nand U2068 (N_2068,N_2005,N_2016);
nand U2069 (N_2069,N_2001,N_1998);
or U2070 (N_2070,N_2017,N_1989);
nor U2071 (N_2071,N_2028,N_2031);
or U2072 (N_2072,N_1980,N_1988);
and U2073 (N_2073,N_1993,N_2038);
or U2074 (N_2074,N_2030,N_2032);
nor U2075 (N_2075,N_2022,N_1992);
or U2076 (N_2076,N_1991,N_2022);
nor U2077 (N_2077,N_2012,N_2016);
and U2078 (N_2078,N_1988,N_1984);
nand U2079 (N_2079,N_2006,N_2004);
nor U2080 (N_2080,N_1998,N_2007);
or U2081 (N_2081,N_1985,N_1995);
and U2082 (N_2082,N_2007,N_2002);
xnor U2083 (N_2083,N_2033,N_2030);
or U2084 (N_2084,N_1987,N_1988);
or U2085 (N_2085,N_1996,N_2031);
and U2086 (N_2086,N_1983,N_1997);
nor U2087 (N_2087,N_1986,N_2006);
or U2088 (N_2088,N_2018,N_1986);
xnor U2089 (N_2089,N_1991,N_2034);
or U2090 (N_2090,N_2022,N_2018);
nor U2091 (N_2091,N_2006,N_2027);
and U2092 (N_2092,N_2036,N_2022);
xnor U2093 (N_2093,N_2039,N_2001);
nor U2094 (N_2094,N_1990,N_2027);
xor U2095 (N_2095,N_2009,N_1985);
nand U2096 (N_2096,N_1980,N_2001);
nand U2097 (N_2097,N_2000,N_2016);
nor U2098 (N_2098,N_1988,N_2002);
or U2099 (N_2099,N_2002,N_2010);
xnor U2100 (N_2100,N_2079,N_2069);
and U2101 (N_2101,N_2040,N_2046);
nor U2102 (N_2102,N_2089,N_2044);
xnor U2103 (N_2103,N_2058,N_2052);
or U2104 (N_2104,N_2051,N_2073);
xnor U2105 (N_2105,N_2070,N_2041);
or U2106 (N_2106,N_2071,N_2067);
nand U2107 (N_2107,N_2054,N_2099);
nor U2108 (N_2108,N_2057,N_2095);
xor U2109 (N_2109,N_2068,N_2065);
xnor U2110 (N_2110,N_2093,N_2087);
nand U2111 (N_2111,N_2091,N_2060);
xnor U2112 (N_2112,N_2085,N_2047);
nand U2113 (N_2113,N_2078,N_2076);
nand U2114 (N_2114,N_2098,N_2050);
or U2115 (N_2115,N_2092,N_2042);
and U2116 (N_2116,N_2045,N_2086);
xor U2117 (N_2117,N_2049,N_2097);
nor U2118 (N_2118,N_2062,N_2059);
or U2119 (N_2119,N_2096,N_2084);
nor U2120 (N_2120,N_2083,N_2063);
nand U2121 (N_2121,N_2075,N_2090);
and U2122 (N_2122,N_2082,N_2088);
xnor U2123 (N_2123,N_2077,N_2061);
xor U2124 (N_2124,N_2072,N_2043);
nand U2125 (N_2125,N_2056,N_2053);
xor U2126 (N_2126,N_2081,N_2055);
or U2127 (N_2127,N_2094,N_2048);
nand U2128 (N_2128,N_2074,N_2066);
nand U2129 (N_2129,N_2064,N_2080);
nand U2130 (N_2130,N_2049,N_2069);
nor U2131 (N_2131,N_2072,N_2068);
xor U2132 (N_2132,N_2089,N_2083);
nand U2133 (N_2133,N_2068,N_2071);
nand U2134 (N_2134,N_2081,N_2043);
and U2135 (N_2135,N_2058,N_2047);
and U2136 (N_2136,N_2086,N_2069);
xnor U2137 (N_2137,N_2057,N_2052);
nor U2138 (N_2138,N_2049,N_2066);
or U2139 (N_2139,N_2051,N_2046);
and U2140 (N_2140,N_2063,N_2042);
and U2141 (N_2141,N_2050,N_2044);
xor U2142 (N_2142,N_2062,N_2091);
and U2143 (N_2143,N_2093,N_2065);
xnor U2144 (N_2144,N_2046,N_2090);
xnor U2145 (N_2145,N_2050,N_2092);
nor U2146 (N_2146,N_2069,N_2066);
or U2147 (N_2147,N_2068,N_2045);
nor U2148 (N_2148,N_2078,N_2083);
or U2149 (N_2149,N_2059,N_2099);
nor U2150 (N_2150,N_2058,N_2074);
nand U2151 (N_2151,N_2052,N_2070);
and U2152 (N_2152,N_2098,N_2051);
xor U2153 (N_2153,N_2053,N_2096);
or U2154 (N_2154,N_2080,N_2079);
xor U2155 (N_2155,N_2077,N_2042);
or U2156 (N_2156,N_2072,N_2058);
nor U2157 (N_2157,N_2094,N_2075);
nor U2158 (N_2158,N_2093,N_2041);
and U2159 (N_2159,N_2096,N_2078);
nand U2160 (N_2160,N_2143,N_2158);
nor U2161 (N_2161,N_2115,N_2117);
nor U2162 (N_2162,N_2156,N_2153);
or U2163 (N_2163,N_2155,N_2109);
xor U2164 (N_2164,N_2123,N_2141);
nor U2165 (N_2165,N_2140,N_2131);
and U2166 (N_2166,N_2135,N_2151);
nand U2167 (N_2167,N_2100,N_2105);
nor U2168 (N_2168,N_2107,N_2114);
nor U2169 (N_2169,N_2152,N_2129);
or U2170 (N_2170,N_2134,N_2121);
nand U2171 (N_2171,N_2122,N_2118);
and U2172 (N_2172,N_2142,N_2149);
and U2173 (N_2173,N_2120,N_2159);
and U2174 (N_2174,N_2154,N_2116);
or U2175 (N_2175,N_2148,N_2130);
nand U2176 (N_2176,N_2111,N_2106);
nand U2177 (N_2177,N_2127,N_2128);
or U2178 (N_2178,N_2144,N_2132);
and U2179 (N_2179,N_2147,N_2101);
and U2180 (N_2180,N_2119,N_2103);
or U2181 (N_2181,N_2104,N_2102);
or U2182 (N_2182,N_2125,N_2112);
xnor U2183 (N_2183,N_2145,N_2146);
and U2184 (N_2184,N_2136,N_2138);
xnor U2185 (N_2185,N_2139,N_2108);
or U2186 (N_2186,N_2133,N_2110);
nor U2187 (N_2187,N_2124,N_2137);
xor U2188 (N_2188,N_2126,N_2150);
nor U2189 (N_2189,N_2157,N_2113);
xnor U2190 (N_2190,N_2126,N_2132);
and U2191 (N_2191,N_2137,N_2114);
nand U2192 (N_2192,N_2123,N_2129);
nor U2193 (N_2193,N_2128,N_2158);
or U2194 (N_2194,N_2103,N_2112);
xnor U2195 (N_2195,N_2126,N_2136);
or U2196 (N_2196,N_2131,N_2139);
nand U2197 (N_2197,N_2114,N_2119);
nor U2198 (N_2198,N_2107,N_2108);
xor U2199 (N_2199,N_2144,N_2115);
and U2200 (N_2200,N_2132,N_2113);
xnor U2201 (N_2201,N_2134,N_2128);
and U2202 (N_2202,N_2114,N_2134);
or U2203 (N_2203,N_2146,N_2117);
xor U2204 (N_2204,N_2130,N_2131);
nor U2205 (N_2205,N_2144,N_2121);
nor U2206 (N_2206,N_2130,N_2152);
xnor U2207 (N_2207,N_2125,N_2144);
or U2208 (N_2208,N_2128,N_2152);
xor U2209 (N_2209,N_2101,N_2126);
nand U2210 (N_2210,N_2151,N_2110);
or U2211 (N_2211,N_2132,N_2149);
or U2212 (N_2212,N_2150,N_2101);
and U2213 (N_2213,N_2158,N_2125);
and U2214 (N_2214,N_2104,N_2140);
or U2215 (N_2215,N_2130,N_2119);
nor U2216 (N_2216,N_2138,N_2120);
or U2217 (N_2217,N_2117,N_2105);
nand U2218 (N_2218,N_2106,N_2127);
xor U2219 (N_2219,N_2127,N_2146);
nand U2220 (N_2220,N_2215,N_2171);
or U2221 (N_2221,N_2195,N_2197);
nor U2222 (N_2222,N_2167,N_2210);
nor U2223 (N_2223,N_2175,N_2176);
nor U2224 (N_2224,N_2207,N_2165);
or U2225 (N_2225,N_2181,N_2202);
and U2226 (N_2226,N_2194,N_2177);
or U2227 (N_2227,N_2164,N_2173);
nand U2228 (N_2228,N_2160,N_2208);
or U2229 (N_2229,N_2183,N_2166);
xnor U2230 (N_2230,N_2161,N_2188);
xor U2231 (N_2231,N_2172,N_2193);
nand U2232 (N_2232,N_2191,N_2196);
nand U2233 (N_2233,N_2168,N_2217);
and U2234 (N_2234,N_2205,N_2182);
nor U2235 (N_2235,N_2189,N_2211);
and U2236 (N_2236,N_2212,N_2199);
xor U2237 (N_2237,N_2179,N_2200);
nand U2238 (N_2238,N_2184,N_2216);
nor U2239 (N_2239,N_2203,N_2178);
nand U2240 (N_2240,N_2214,N_2170);
nand U2241 (N_2241,N_2190,N_2192);
xnor U2242 (N_2242,N_2209,N_2206);
or U2243 (N_2243,N_2219,N_2174);
or U2244 (N_2244,N_2163,N_2169);
nand U2245 (N_2245,N_2180,N_2201);
nand U2246 (N_2246,N_2162,N_2218);
or U2247 (N_2247,N_2187,N_2198);
or U2248 (N_2248,N_2186,N_2185);
and U2249 (N_2249,N_2213,N_2204);
or U2250 (N_2250,N_2187,N_2164);
xnor U2251 (N_2251,N_2200,N_2170);
nor U2252 (N_2252,N_2168,N_2209);
xor U2253 (N_2253,N_2219,N_2216);
xnor U2254 (N_2254,N_2196,N_2165);
nor U2255 (N_2255,N_2208,N_2185);
or U2256 (N_2256,N_2206,N_2178);
nor U2257 (N_2257,N_2181,N_2211);
and U2258 (N_2258,N_2204,N_2201);
nor U2259 (N_2259,N_2199,N_2216);
or U2260 (N_2260,N_2200,N_2183);
xnor U2261 (N_2261,N_2186,N_2191);
nor U2262 (N_2262,N_2210,N_2208);
nor U2263 (N_2263,N_2197,N_2181);
and U2264 (N_2264,N_2210,N_2170);
nand U2265 (N_2265,N_2180,N_2188);
nand U2266 (N_2266,N_2214,N_2187);
and U2267 (N_2267,N_2168,N_2189);
nand U2268 (N_2268,N_2203,N_2198);
and U2269 (N_2269,N_2184,N_2199);
or U2270 (N_2270,N_2199,N_2213);
and U2271 (N_2271,N_2161,N_2197);
and U2272 (N_2272,N_2214,N_2177);
or U2273 (N_2273,N_2165,N_2182);
nor U2274 (N_2274,N_2166,N_2164);
nand U2275 (N_2275,N_2202,N_2191);
or U2276 (N_2276,N_2216,N_2175);
xor U2277 (N_2277,N_2208,N_2181);
nor U2278 (N_2278,N_2199,N_2167);
xor U2279 (N_2279,N_2163,N_2202);
xor U2280 (N_2280,N_2273,N_2233);
nand U2281 (N_2281,N_2229,N_2263);
nand U2282 (N_2282,N_2268,N_2222);
nor U2283 (N_2283,N_2243,N_2259);
or U2284 (N_2284,N_2251,N_2250);
nor U2285 (N_2285,N_2255,N_2254);
or U2286 (N_2286,N_2221,N_2244);
nand U2287 (N_2287,N_2258,N_2260);
or U2288 (N_2288,N_2266,N_2270);
nor U2289 (N_2289,N_2252,N_2274);
or U2290 (N_2290,N_2248,N_2240);
nand U2291 (N_2291,N_2230,N_2247);
nor U2292 (N_2292,N_2242,N_2239);
or U2293 (N_2293,N_2265,N_2238);
xor U2294 (N_2294,N_2275,N_2225);
or U2295 (N_2295,N_2223,N_2231);
nand U2296 (N_2296,N_2278,N_2235);
nand U2297 (N_2297,N_2236,N_2227);
nand U2298 (N_2298,N_2276,N_2245);
or U2299 (N_2299,N_2256,N_2261);
xor U2300 (N_2300,N_2253,N_2277);
nand U2301 (N_2301,N_2257,N_2279);
nor U2302 (N_2302,N_2228,N_2232);
nor U2303 (N_2303,N_2226,N_2271);
and U2304 (N_2304,N_2220,N_2262);
nor U2305 (N_2305,N_2249,N_2224);
xor U2306 (N_2306,N_2234,N_2267);
nor U2307 (N_2307,N_2269,N_2246);
xor U2308 (N_2308,N_2264,N_2241);
or U2309 (N_2309,N_2237,N_2272);
or U2310 (N_2310,N_2254,N_2220);
or U2311 (N_2311,N_2248,N_2279);
nor U2312 (N_2312,N_2279,N_2251);
nand U2313 (N_2313,N_2236,N_2233);
nand U2314 (N_2314,N_2276,N_2267);
nor U2315 (N_2315,N_2241,N_2250);
xor U2316 (N_2316,N_2223,N_2224);
or U2317 (N_2317,N_2252,N_2250);
xor U2318 (N_2318,N_2246,N_2240);
nand U2319 (N_2319,N_2230,N_2233);
and U2320 (N_2320,N_2237,N_2248);
nand U2321 (N_2321,N_2262,N_2232);
or U2322 (N_2322,N_2259,N_2251);
and U2323 (N_2323,N_2279,N_2250);
or U2324 (N_2324,N_2257,N_2258);
or U2325 (N_2325,N_2265,N_2239);
xnor U2326 (N_2326,N_2245,N_2250);
nor U2327 (N_2327,N_2252,N_2264);
xnor U2328 (N_2328,N_2240,N_2227);
xor U2329 (N_2329,N_2264,N_2232);
or U2330 (N_2330,N_2245,N_2234);
nand U2331 (N_2331,N_2239,N_2253);
nor U2332 (N_2332,N_2266,N_2234);
and U2333 (N_2333,N_2228,N_2241);
xnor U2334 (N_2334,N_2251,N_2252);
and U2335 (N_2335,N_2248,N_2275);
nand U2336 (N_2336,N_2279,N_2240);
or U2337 (N_2337,N_2279,N_2232);
or U2338 (N_2338,N_2277,N_2249);
or U2339 (N_2339,N_2264,N_2268);
xnor U2340 (N_2340,N_2285,N_2309);
or U2341 (N_2341,N_2288,N_2324);
xnor U2342 (N_2342,N_2291,N_2300);
xor U2343 (N_2343,N_2305,N_2330);
nand U2344 (N_2344,N_2289,N_2328);
xor U2345 (N_2345,N_2307,N_2283);
and U2346 (N_2346,N_2331,N_2335);
nand U2347 (N_2347,N_2336,N_2284);
and U2348 (N_2348,N_2281,N_2329);
nand U2349 (N_2349,N_2317,N_2327);
nor U2350 (N_2350,N_2310,N_2293);
nand U2351 (N_2351,N_2294,N_2312);
nand U2352 (N_2352,N_2304,N_2286);
xnor U2353 (N_2353,N_2318,N_2296);
and U2354 (N_2354,N_2326,N_2299);
nor U2355 (N_2355,N_2321,N_2303);
nand U2356 (N_2356,N_2306,N_2316);
and U2357 (N_2357,N_2280,N_2297);
nor U2358 (N_2358,N_2302,N_2298);
nor U2359 (N_2359,N_2313,N_2332);
xor U2360 (N_2360,N_2337,N_2333);
xnor U2361 (N_2361,N_2314,N_2323);
xnor U2362 (N_2362,N_2282,N_2339);
nor U2363 (N_2363,N_2338,N_2322);
and U2364 (N_2364,N_2290,N_2325);
xor U2365 (N_2365,N_2287,N_2292);
or U2366 (N_2366,N_2320,N_2311);
nor U2367 (N_2367,N_2334,N_2315);
and U2368 (N_2368,N_2301,N_2295);
or U2369 (N_2369,N_2308,N_2319);
nand U2370 (N_2370,N_2293,N_2285);
nand U2371 (N_2371,N_2296,N_2308);
xor U2372 (N_2372,N_2327,N_2296);
or U2373 (N_2373,N_2329,N_2286);
xnor U2374 (N_2374,N_2303,N_2286);
nor U2375 (N_2375,N_2314,N_2320);
or U2376 (N_2376,N_2309,N_2293);
xor U2377 (N_2377,N_2283,N_2280);
and U2378 (N_2378,N_2304,N_2290);
or U2379 (N_2379,N_2305,N_2311);
and U2380 (N_2380,N_2313,N_2283);
nand U2381 (N_2381,N_2306,N_2320);
nand U2382 (N_2382,N_2307,N_2298);
and U2383 (N_2383,N_2290,N_2322);
and U2384 (N_2384,N_2299,N_2304);
or U2385 (N_2385,N_2289,N_2299);
or U2386 (N_2386,N_2330,N_2298);
nand U2387 (N_2387,N_2296,N_2295);
and U2388 (N_2388,N_2330,N_2280);
or U2389 (N_2389,N_2313,N_2281);
nand U2390 (N_2390,N_2324,N_2292);
and U2391 (N_2391,N_2318,N_2325);
xor U2392 (N_2392,N_2297,N_2308);
nor U2393 (N_2393,N_2307,N_2282);
nor U2394 (N_2394,N_2293,N_2328);
or U2395 (N_2395,N_2301,N_2310);
or U2396 (N_2396,N_2282,N_2310);
and U2397 (N_2397,N_2313,N_2322);
or U2398 (N_2398,N_2287,N_2329);
nand U2399 (N_2399,N_2328,N_2315);
xor U2400 (N_2400,N_2395,N_2359);
or U2401 (N_2401,N_2362,N_2367);
or U2402 (N_2402,N_2392,N_2341);
nor U2403 (N_2403,N_2391,N_2348);
nor U2404 (N_2404,N_2388,N_2393);
nand U2405 (N_2405,N_2396,N_2352);
or U2406 (N_2406,N_2378,N_2371);
nor U2407 (N_2407,N_2376,N_2343);
or U2408 (N_2408,N_2353,N_2363);
xor U2409 (N_2409,N_2394,N_2345);
nor U2410 (N_2410,N_2383,N_2344);
nand U2411 (N_2411,N_2342,N_2364);
and U2412 (N_2412,N_2356,N_2357);
and U2413 (N_2413,N_2368,N_2372);
nor U2414 (N_2414,N_2350,N_2397);
and U2415 (N_2415,N_2369,N_2349);
xnor U2416 (N_2416,N_2387,N_2389);
nor U2417 (N_2417,N_2358,N_2360);
or U2418 (N_2418,N_2384,N_2361);
nor U2419 (N_2419,N_2399,N_2355);
xnor U2420 (N_2420,N_2381,N_2386);
nand U2421 (N_2421,N_2380,N_2373);
nor U2422 (N_2422,N_2377,N_2385);
and U2423 (N_2423,N_2366,N_2382);
or U2424 (N_2424,N_2374,N_2390);
nor U2425 (N_2425,N_2379,N_2365);
and U2426 (N_2426,N_2340,N_2375);
or U2427 (N_2427,N_2351,N_2398);
and U2428 (N_2428,N_2370,N_2346);
xor U2429 (N_2429,N_2347,N_2354);
nor U2430 (N_2430,N_2351,N_2381);
nand U2431 (N_2431,N_2390,N_2342);
nor U2432 (N_2432,N_2360,N_2344);
or U2433 (N_2433,N_2343,N_2371);
xnor U2434 (N_2434,N_2357,N_2346);
nand U2435 (N_2435,N_2340,N_2358);
nor U2436 (N_2436,N_2386,N_2389);
and U2437 (N_2437,N_2343,N_2356);
and U2438 (N_2438,N_2371,N_2398);
nand U2439 (N_2439,N_2381,N_2348);
nor U2440 (N_2440,N_2364,N_2375);
or U2441 (N_2441,N_2377,N_2388);
nor U2442 (N_2442,N_2351,N_2361);
nand U2443 (N_2443,N_2361,N_2341);
xnor U2444 (N_2444,N_2373,N_2377);
or U2445 (N_2445,N_2362,N_2351);
nand U2446 (N_2446,N_2371,N_2380);
xor U2447 (N_2447,N_2357,N_2393);
or U2448 (N_2448,N_2347,N_2371);
and U2449 (N_2449,N_2352,N_2357);
or U2450 (N_2450,N_2340,N_2371);
or U2451 (N_2451,N_2366,N_2394);
nor U2452 (N_2452,N_2378,N_2355);
and U2453 (N_2453,N_2395,N_2349);
nor U2454 (N_2454,N_2380,N_2391);
or U2455 (N_2455,N_2354,N_2348);
or U2456 (N_2456,N_2398,N_2392);
and U2457 (N_2457,N_2378,N_2350);
nand U2458 (N_2458,N_2364,N_2350);
or U2459 (N_2459,N_2399,N_2374);
or U2460 (N_2460,N_2459,N_2435);
or U2461 (N_2461,N_2422,N_2413);
or U2462 (N_2462,N_2442,N_2444);
or U2463 (N_2463,N_2423,N_2428);
xnor U2464 (N_2464,N_2402,N_2457);
and U2465 (N_2465,N_2434,N_2433);
or U2466 (N_2466,N_2401,N_2409);
nand U2467 (N_2467,N_2418,N_2412);
xor U2468 (N_2468,N_2431,N_2455);
nor U2469 (N_2469,N_2443,N_2452);
nor U2470 (N_2470,N_2449,N_2440);
xnor U2471 (N_2471,N_2439,N_2403);
xor U2472 (N_2472,N_2424,N_2432);
nor U2473 (N_2473,N_2407,N_2414);
or U2474 (N_2474,N_2420,N_2400);
xor U2475 (N_2475,N_2415,N_2430);
and U2476 (N_2476,N_2410,N_2408);
xnor U2477 (N_2477,N_2450,N_2448);
xor U2478 (N_2478,N_2437,N_2436);
or U2479 (N_2479,N_2438,N_2411);
nor U2480 (N_2480,N_2454,N_2404);
nand U2481 (N_2481,N_2456,N_2416);
or U2482 (N_2482,N_2458,N_2426);
or U2483 (N_2483,N_2405,N_2421);
nor U2484 (N_2484,N_2427,N_2445);
xnor U2485 (N_2485,N_2417,N_2429);
nor U2486 (N_2486,N_2453,N_2451);
nor U2487 (N_2487,N_2447,N_2419);
nand U2488 (N_2488,N_2446,N_2425);
nand U2489 (N_2489,N_2406,N_2441);
or U2490 (N_2490,N_2443,N_2434);
xnor U2491 (N_2491,N_2401,N_2431);
xor U2492 (N_2492,N_2457,N_2453);
nand U2493 (N_2493,N_2412,N_2442);
nor U2494 (N_2494,N_2443,N_2403);
nor U2495 (N_2495,N_2450,N_2440);
nand U2496 (N_2496,N_2441,N_2411);
nand U2497 (N_2497,N_2417,N_2406);
or U2498 (N_2498,N_2403,N_2407);
nand U2499 (N_2499,N_2427,N_2440);
xor U2500 (N_2500,N_2454,N_2402);
nand U2501 (N_2501,N_2450,N_2427);
or U2502 (N_2502,N_2435,N_2434);
and U2503 (N_2503,N_2408,N_2430);
nand U2504 (N_2504,N_2420,N_2427);
nand U2505 (N_2505,N_2437,N_2432);
or U2506 (N_2506,N_2419,N_2416);
or U2507 (N_2507,N_2406,N_2434);
nor U2508 (N_2508,N_2436,N_2404);
nand U2509 (N_2509,N_2447,N_2453);
or U2510 (N_2510,N_2421,N_2432);
or U2511 (N_2511,N_2410,N_2417);
nor U2512 (N_2512,N_2427,N_2406);
xor U2513 (N_2513,N_2415,N_2414);
xor U2514 (N_2514,N_2403,N_2412);
xnor U2515 (N_2515,N_2435,N_2443);
nor U2516 (N_2516,N_2457,N_2445);
nor U2517 (N_2517,N_2430,N_2431);
and U2518 (N_2518,N_2407,N_2432);
or U2519 (N_2519,N_2413,N_2411);
or U2520 (N_2520,N_2499,N_2507);
and U2521 (N_2521,N_2490,N_2519);
nor U2522 (N_2522,N_2506,N_2512);
xnor U2523 (N_2523,N_2476,N_2518);
nor U2524 (N_2524,N_2473,N_2464);
nor U2525 (N_2525,N_2466,N_2500);
or U2526 (N_2526,N_2493,N_2460);
nor U2527 (N_2527,N_2517,N_2513);
nand U2528 (N_2528,N_2477,N_2467);
xor U2529 (N_2529,N_2480,N_2487);
nand U2530 (N_2530,N_2488,N_2462);
or U2531 (N_2531,N_2516,N_2468);
nand U2532 (N_2532,N_2510,N_2486);
or U2533 (N_2533,N_2491,N_2463);
xnor U2534 (N_2534,N_2472,N_2502);
xnor U2535 (N_2535,N_2485,N_2503);
xnor U2536 (N_2536,N_2494,N_2479);
or U2537 (N_2537,N_2470,N_2471);
xnor U2538 (N_2538,N_2492,N_2482);
or U2539 (N_2539,N_2505,N_2496);
and U2540 (N_2540,N_2508,N_2501);
or U2541 (N_2541,N_2483,N_2478);
nor U2542 (N_2542,N_2504,N_2495);
nor U2543 (N_2543,N_2511,N_2475);
and U2544 (N_2544,N_2484,N_2481);
and U2545 (N_2545,N_2514,N_2465);
or U2546 (N_2546,N_2509,N_2461);
and U2547 (N_2547,N_2474,N_2489);
and U2548 (N_2548,N_2515,N_2497);
and U2549 (N_2549,N_2498,N_2469);
and U2550 (N_2550,N_2467,N_2510);
nor U2551 (N_2551,N_2490,N_2513);
nand U2552 (N_2552,N_2503,N_2518);
xnor U2553 (N_2553,N_2501,N_2518);
nor U2554 (N_2554,N_2485,N_2478);
nor U2555 (N_2555,N_2469,N_2494);
nand U2556 (N_2556,N_2467,N_2511);
nor U2557 (N_2557,N_2468,N_2509);
xor U2558 (N_2558,N_2477,N_2479);
and U2559 (N_2559,N_2465,N_2473);
and U2560 (N_2560,N_2483,N_2493);
nand U2561 (N_2561,N_2499,N_2475);
nand U2562 (N_2562,N_2491,N_2506);
xnor U2563 (N_2563,N_2465,N_2472);
xor U2564 (N_2564,N_2511,N_2503);
or U2565 (N_2565,N_2503,N_2519);
and U2566 (N_2566,N_2485,N_2468);
or U2567 (N_2567,N_2516,N_2476);
or U2568 (N_2568,N_2462,N_2504);
nand U2569 (N_2569,N_2501,N_2496);
nand U2570 (N_2570,N_2519,N_2496);
or U2571 (N_2571,N_2463,N_2466);
xor U2572 (N_2572,N_2476,N_2477);
and U2573 (N_2573,N_2510,N_2519);
xnor U2574 (N_2574,N_2500,N_2486);
or U2575 (N_2575,N_2514,N_2513);
and U2576 (N_2576,N_2497,N_2512);
nor U2577 (N_2577,N_2489,N_2483);
and U2578 (N_2578,N_2503,N_2472);
and U2579 (N_2579,N_2494,N_2484);
and U2580 (N_2580,N_2545,N_2544);
nor U2581 (N_2581,N_2551,N_2566);
nor U2582 (N_2582,N_2571,N_2560);
xnor U2583 (N_2583,N_2552,N_2557);
nand U2584 (N_2584,N_2577,N_2568);
xor U2585 (N_2585,N_2525,N_2549);
nand U2586 (N_2586,N_2541,N_2530);
nand U2587 (N_2587,N_2567,N_2556);
or U2588 (N_2588,N_2526,N_2535);
xnor U2589 (N_2589,N_2537,N_2520);
or U2590 (N_2590,N_2536,N_2575);
and U2591 (N_2591,N_2579,N_2561);
nor U2592 (N_2592,N_2538,N_2555);
or U2593 (N_2593,N_2563,N_2546);
or U2594 (N_2594,N_2531,N_2564);
or U2595 (N_2595,N_2527,N_2524);
nor U2596 (N_2596,N_2523,N_2570);
nor U2597 (N_2597,N_2578,N_2574);
nand U2598 (N_2598,N_2543,N_2573);
xnor U2599 (N_2599,N_2565,N_2554);
nand U2600 (N_2600,N_2576,N_2528);
and U2601 (N_2601,N_2548,N_2532);
nand U2602 (N_2602,N_2522,N_2562);
and U2603 (N_2603,N_2533,N_2529);
nand U2604 (N_2604,N_2559,N_2539);
nor U2605 (N_2605,N_2540,N_2521);
or U2606 (N_2606,N_2558,N_2547);
and U2607 (N_2607,N_2569,N_2553);
nand U2608 (N_2608,N_2550,N_2534);
and U2609 (N_2609,N_2542,N_2572);
nor U2610 (N_2610,N_2522,N_2533);
nand U2611 (N_2611,N_2554,N_2560);
nor U2612 (N_2612,N_2568,N_2570);
xnor U2613 (N_2613,N_2540,N_2565);
and U2614 (N_2614,N_2570,N_2564);
nor U2615 (N_2615,N_2560,N_2529);
xor U2616 (N_2616,N_2558,N_2539);
and U2617 (N_2617,N_2532,N_2544);
or U2618 (N_2618,N_2523,N_2575);
xor U2619 (N_2619,N_2539,N_2536);
or U2620 (N_2620,N_2578,N_2547);
xor U2621 (N_2621,N_2570,N_2529);
nor U2622 (N_2622,N_2573,N_2574);
nor U2623 (N_2623,N_2562,N_2533);
nor U2624 (N_2624,N_2535,N_2554);
and U2625 (N_2625,N_2554,N_2562);
nand U2626 (N_2626,N_2529,N_2556);
nand U2627 (N_2627,N_2537,N_2556);
nand U2628 (N_2628,N_2551,N_2530);
nand U2629 (N_2629,N_2535,N_2551);
xor U2630 (N_2630,N_2577,N_2540);
xor U2631 (N_2631,N_2536,N_2579);
and U2632 (N_2632,N_2544,N_2534);
nor U2633 (N_2633,N_2548,N_2576);
xor U2634 (N_2634,N_2544,N_2567);
and U2635 (N_2635,N_2579,N_2550);
nand U2636 (N_2636,N_2550,N_2522);
nand U2637 (N_2637,N_2540,N_2529);
nand U2638 (N_2638,N_2525,N_2560);
nand U2639 (N_2639,N_2531,N_2555);
xor U2640 (N_2640,N_2595,N_2586);
nor U2641 (N_2641,N_2626,N_2610);
or U2642 (N_2642,N_2617,N_2600);
or U2643 (N_2643,N_2614,N_2583);
and U2644 (N_2644,N_2594,N_2604);
or U2645 (N_2645,N_2580,N_2591);
and U2646 (N_2646,N_2625,N_2588);
xnor U2647 (N_2647,N_2602,N_2593);
xnor U2648 (N_2648,N_2613,N_2605);
xor U2649 (N_2649,N_2609,N_2599);
nand U2650 (N_2650,N_2606,N_2603);
or U2651 (N_2651,N_2621,N_2611);
or U2652 (N_2652,N_2608,N_2601);
nand U2653 (N_2653,N_2635,N_2582);
nand U2654 (N_2654,N_2636,N_2585);
and U2655 (N_2655,N_2619,N_2607);
or U2656 (N_2656,N_2596,N_2616);
nand U2657 (N_2657,N_2634,N_2587);
or U2658 (N_2658,N_2622,N_2632);
nor U2659 (N_2659,N_2618,N_2629);
or U2660 (N_2660,N_2598,N_2623);
or U2661 (N_2661,N_2637,N_2633);
or U2662 (N_2662,N_2627,N_2630);
nor U2663 (N_2663,N_2615,N_2612);
or U2664 (N_2664,N_2584,N_2624);
nor U2665 (N_2665,N_2628,N_2597);
nor U2666 (N_2666,N_2620,N_2581);
and U2667 (N_2667,N_2631,N_2590);
nor U2668 (N_2668,N_2639,N_2589);
nor U2669 (N_2669,N_2638,N_2592);
nor U2670 (N_2670,N_2591,N_2619);
xor U2671 (N_2671,N_2584,N_2630);
or U2672 (N_2672,N_2597,N_2624);
xnor U2673 (N_2673,N_2622,N_2610);
and U2674 (N_2674,N_2604,N_2588);
nor U2675 (N_2675,N_2625,N_2602);
xor U2676 (N_2676,N_2610,N_2616);
nor U2677 (N_2677,N_2584,N_2611);
nand U2678 (N_2678,N_2587,N_2602);
nand U2679 (N_2679,N_2580,N_2609);
nand U2680 (N_2680,N_2628,N_2637);
nor U2681 (N_2681,N_2602,N_2605);
xnor U2682 (N_2682,N_2622,N_2584);
xor U2683 (N_2683,N_2616,N_2629);
and U2684 (N_2684,N_2588,N_2603);
xnor U2685 (N_2685,N_2619,N_2635);
xor U2686 (N_2686,N_2610,N_2637);
and U2687 (N_2687,N_2600,N_2631);
xor U2688 (N_2688,N_2636,N_2584);
or U2689 (N_2689,N_2619,N_2581);
xor U2690 (N_2690,N_2582,N_2618);
xor U2691 (N_2691,N_2623,N_2622);
nor U2692 (N_2692,N_2602,N_2607);
nand U2693 (N_2693,N_2592,N_2624);
nand U2694 (N_2694,N_2605,N_2589);
nor U2695 (N_2695,N_2606,N_2601);
xnor U2696 (N_2696,N_2621,N_2591);
and U2697 (N_2697,N_2605,N_2581);
or U2698 (N_2698,N_2639,N_2614);
nor U2699 (N_2699,N_2615,N_2616);
nand U2700 (N_2700,N_2668,N_2656);
nand U2701 (N_2701,N_2644,N_2654);
or U2702 (N_2702,N_2642,N_2667);
nand U2703 (N_2703,N_2681,N_2678);
nor U2704 (N_2704,N_2679,N_2673);
nor U2705 (N_2705,N_2658,N_2641);
nor U2706 (N_2706,N_2670,N_2694);
xnor U2707 (N_2707,N_2690,N_2698);
or U2708 (N_2708,N_2671,N_2655);
nand U2709 (N_2709,N_2652,N_2651);
and U2710 (N_2710,N_2640,N_2688);
or U2711 (N_2711,N_2643,N_2669);
xor U2712 (N_2712,N_2657,N_2692);
nor U2713 (N_2713,N_2696,N_2680);
nand U2714 (N_2714,N_2661,N_2693);
nor U2715 (N_2715,N_2672,N_2663);
nor U2716 (N_2716,N_2659,N_2699);
or U2717 (N_2717,N_2660,N_2695);
or U2718 (N_2718,N_2676,N_2687);
nand U2719 (N_2719,N_2686,N_2677);
and U2720 (N_2720,N_2649,N_2666);
and U2721 (N_2721,N_2653,N_2664);
xor U2722 (N_2722,N_2645,N_2662);
nor U2723 (N_2723,N_2647,N_2650);
nor U2724 (N_2724,N_2683,N_2689);
or U2725 (N_2725,N_2691,N_2674);
or U2726 (N_2726,N_2675,N_2665);
nor U2727 (N_2727,N_2646,N_2684);
nand U2728 (N_2728,N_2685,N_2682);
nor U2729 (N_2729,N_2648,N_2697);
and U2730 (N_2730,N_2673,N_2685);
nand U2731 (N_2731,N_2646,N_2664);
xnor U2732 (N_2732,N_2640,N_2644);
nor U2733 (N_2733,N_2686,N_2669);
nand U2734 (N_2734,N_2655,N_2686);
or U2735 (N_2735,N_2676,N_2651);
nand U2736 (N_2736,N_2645,N_2660);
or U2737 (N_2737,N_2680,N_2676);
nand U2738 (N_2738,N_2655,N_2651);
nor U2739 (N_2739,N_2696,N_2685);
and U2740 (N_2740,N_2686,N_2678);
nand U2741 (N_2741,N_2675,N_2660);
nor U2742 (N_2742,N_2676,N_2690);
nor U2743 (N_2743,N_2656,N_2699);
nand U2744 (N_2744,N_2672,N_2698);
nand U2745 (N_2745,N_2645,N_2695);
xnor U2746 (N_2746,N_2686,N_2649);
xor U2747 (N_2747,N_2680,N_2656);
nor U2748 (N_2748,N_2677,N_2695);
or U2749 (N_2749,N_2652,N_2686);
or U2750 (N_2750,N_2677,N_2641);
and U2751 (N_2751,N_2670,N_2688);
or U2752 (N_2752,N_2676,N_2641);
and U2753 (N_2753,N_2685,N_2674);
xnor U2754 (N_2754,N_2654,N_2655);
nor U2755 (N_2755,N_2673,N_2675);
xnor U2756 (N_2756,N_2677,N_2649);
nand U2757 (N_2757,N_2655,N_2680);
and U2758 (N_2758,N_2640,N_2651);
xnor U2759 (N_2759,N_2656,N_2653);
nand U2760 (N_2760,N_2732,N_2731);
and U2761 (N_2761,N_2729,N_2752);
and U2762 (N_2762,N_2747,N_2745);
xnor U2763 (N_2763,N_2759,N_2719);
nand U2764 (N_2764,N_2749,N_2733);
or U2765 (N_2765,N_2751,N_2713);
xnor U2766 (N_2766,N_2707,N_2722);
or U2767 (N_2767,N_2704,N_2705);
xnor U2768 (N_2768,N_2742,N_2754);
or U2769 (N_2769,N_2725,N_2700);
and U2770 (N_2770,N_2723,N_2726);
nor U2771 (N_2771,N_2748,N_2735);
or U2772 (N_2772,N_2756,N_2746);
nor U2773 (N_2773,N_2741,N_2712);
nor U2774 (N_2774,N_2727,N_2743);
or U2775 (N_2775,N_2708,N_2724);
xnor U2776 (N_2776,N_2717,N_2701);
nor U2777 (N_2777,N_2737,N_2753);
nor U2778 (N_2778,N_2715,N_2734);
nand U2779 (N_2779,N_2721,N_2718);
and U2780 (N_2780,N_2716,N_2744);
nand U2781 (N_2781,N_2730,N_2720);
xor U2782 (N_2782,N_2736,N_2702);
and U2783 (N_2783,N_2703,N_2706);
xnor U2784 (N_2784,N_2757,N_2738);
and U2785 (N_2785,N_2755,N_2758);
or U2786 (N_2786,N_2714,N_2709);
and U2787 (N_2787,N_2750,N_2740);
nor U2788 (N_2788,N_2728,N_2711);
nor U2789 (N_2789,N_2739,N_2710);
or U2790 (N_2790,N_2755,N_2706);
and U2791 (N_2791,N_2736,N_2711);
nand U2792 (N_2792,N_2749,N_2737);
xnor U2793 (N_2793,N_2737,N_2701);
or U2794 (N_2794,N_2722,N_2730);
or U2795 (N_2795,N_2748,N_2734);
and U2796 (N_2796,N_2748,N_2722);
and U2797 (N_2797,N_2736,N_2727);
and U2798 (N_2798,N_2744,N_2726);
xor U2799 (N_2799,N_2745,N_2713);
or U2800 (N_2800,N_2742,N_2703);
nand U2801 (N_2801,N_2727,N_2711);
or U2802 (N_2802,N_2710,N_2748);
nand U2803 (N_2803,N_2759,N_2714);
xnor U2804 (N_2804,N_2716,N_2750);
or U2805 (N_2805,N_2743,N_2755);
nor U2806 (N_2806,N_2733,N_2711);
xnor U2807 (N_2807,N_2713,N_2712);
xor U2808 (N_2808,N_2705,N_2742);
or U2809 (N_2809,N_2739,N_2740);
or U2810 (N_2810,N_2757,N_2707);
and U2811 (N_2811,N_2714,N_2737);
nand U2812 (N_2812,N_2729,N_2727);
xor U2813 (N_2813,N_2754,N_2713);
or U2814 (N_2814,N_2729,N_2757);
nor U2815 (N_2815,N_2713,N_2738);
nand U2816 (N_2816,N_2713,N_2737);
or U2817 (N_2817,N_2709,N_2748);
or U2818 (N_2818,N_2701,N_2711);
nand U2819 (N_2819,N_2710,N_2726);
nor U2820 (N_2820,N_2792,N_2797);
xor U2821 (N_2821,N_2802,N_2814);
xnor U2822 (N_2822,N_2807,N_2805);
xor U2823 (N_2823,N_2794,N_2786);
xnor U2824 (N_2824,N_2793,N_2763);
or U2825 (N_2825,N_2795,N_2774);
or U2826 (N_2826,N_2808,N_2790);
nor U2827 (N_2827,N_2776,N_2815);
or U2828 (N_2828,N_2767,N_2768);
nor U2829 (N_2829,N_2804,N_2778);
or U2830 (N_2830,N_2806,N_2765);
nand U2831 (N_2831,N_2784,N_2800);
xnor U2832 (N_2832,N_2809,N_2801);
nor U2833 (N_2833,N_2769,N_2782);
nor U2834 (N_2834,N_2785,N_2798);
and U2835 (N_2835,N_2789,N_2787);
or U2836 (N_2836,N_2779,N_2811);
and U2837 (N_2837,N_2780,N_2818);
and U2838 (N_2838,N_2816,N_2817);
nand U2839 (N_2839,N_2812,N_2766);
and U2840 (N_2840,N_2773,N_2760);
xor U2841 (N_2841,N_2777,N_2781);
nor U2842 (N_2842,N_2761,N_2775);
nor U2843 (N_2843,N_2799,N_2783);
and U2844 (N_2844,N_2772,N_2813);
nor U2845 (N_2845,N_2819,N_2796);
or U2846 (N_2846,N_2791,N_2764);
nand U2847 (N_2847,N_2803,N_2788);
or U2848 (N_2848,N_2770,N_2810);
xor U2849 (N_2849,N_2771,N_2762);
nor U2850 (N_2850,N_2809,N_2785);
nand U2851 (N_2851,N_2786,N_2775);
and U2852 (N_2852,N_2789,N_2815);
nand U2853 (N_2853,N_2805,N_2771);
nor U2854 (N_2854,N_2774,N_2790);
nand U2855 (N_2855,N_2767,N_2793);
nor U2856 (N_2856,N_2767,N_2781);
or U2857 (N_2857,N_2792,N_2769);
nand U2858 (N_2858,N_2790,N_2813);
or U2859 (N_2859,N_2818,N_2795);
or U2860 (N_2860,N_2813,N_2788);
xor U2861 (N_2861,N_2802,N_2815);
and U2862 (N_2862,N_2786,N_2784);
and U2863 (N_2863,N_2762,N_2770);
nand U2864 (N_2864,N_2785,N_2810);
or U2865 (N_2865,N_2799,N_2790);
nand U2866 (N_2866,N_2815,N_2766);
nor U2867 (N_2867,N_2788,N_2775);
xor U2868 (N_2868,N_2812,N_2793);
nor U2869 (N_2869,N_2760,N_2812);
xnor U2870 (N_2870,N_2768,N_2789);
or U2871 (N_2871,N_2779,N_2762);
and U2872 (N_2872,N_2805,N_2794);
nand U2873 (N_2873,N_2801,N_2798);
xnor U2874 (N_2874,N_2782,N_2785);
and U2875 (N_2875,N_2764,N_2783);
or U2876 (N_2876,N_2809,N_2818);
nor U2877 (N_2877,N_2806,N_2778);
or U2878 (N_2878,N_2778,N_2807);
and U2879 (N_2879,N_2816,N_2795);
or U2880 (N_2880,N_2826,N_2823);
or U2881 (N_2881,N_2830,N_2844);
xnor U2882 (N_2882,N_2836,N_2854);
nor U2883 (N_2883,N_2852,N_2842);
xor U2884 (N_2884,N_2860,N_2874);
or U2885 (N_2885,N_2845,N_2853);
and U2886 (N_2886,N_2829,N_2879);
or U2887 (N_2887,N_2850,N_2847);
or U2888 (N_2888,N_2871,N_2820);
xor U2889 (N_2889,N_2877,N_2869);
nand U2890 (N_2890,N_2848,N_2878);
xor U2891 (N_2891,N_2855,N_2846);
nand U2892 (N_2892,N_2849,N_2873);
nor U2893 (N_2893,N_2828,N_2835);
xor U2894 (N_2894,N_2864,N_2862);
xnor U2895 (N_2895,N_2876,N_2839);
xnor U2896 (N_2896,N_2838,N_2851);
xnor U2897 (N_2897,N_2834,N_2863);
nand U2898 (N_2898,N_2821,N_2861);
or U2899 (N_2899,N_2857,N_2872);
and U2900 (N_2900,N_2840,N_2837);
and U2901 (N_2901,N_2822,N_2868);
or U2902 (N_2902,N_2824,N_2875);
and U2903 (N_2903,N_2865,N_2825);
nand U2904 (N_2904,N_2827,N_2870);
nor U2905 (N_2905,N_2843,N_2832);
xor U2906 (N_2906,N_2866,N_2831);
and U2907 (N_2907,N_2867,N_2841);
and U2908 (N_2908,N_2856,N_2833);
and U2909 (N_2909,N_2859,N_2858);
xnor U2910 (N_2910,N_2822,N_2846);
xnor U2911 (N_2911,N_2848,N_2854);
nor U2912 (N_2912,N_2859,N_2823);
and U2913 (N_2913,N_2838,N_2834);
or U2914 (N_2914,N_2820,N_2867);
or U2915 (N_2915,N_2828,N_2857);
and U2916 (N_2916,N_2842,N_2829);
and U2917 (N_2917,N_2857,N_2848);
and U2918 (N_2918,N_2876,N_2860);
nor U2919 (N_2919,N_2878,N_2862);
or U2920 (N_2920,N_2870,N_2876);
nor U2921 (N_2921,N_2855,N_2840);
and U2922 (N_2922,N_2839,N_2863);
nor U2923 (N_2923,N_2832,N_2855);
nor U2924 (N_2924,N_2842,N_2840);
xnor U2925 (N_2925,N_2872,N_2840);
nor U2926 (N_2926,N_2828,N_2862);
nand U2927 (N_2927,N_2866,N_2876);
and U2928 (N_2928,N_2879,N_2852);
or U2929 (N_2929,N_2866,N_2843);
and U2930 (N_2930,N_2858,N_2860);
nor U2931 (N_2931,N_2827,N_2879);
xor U2932 (N_2932,N_2879,N_2866);
nor U2933 (N_2933,N_2863,N_2854);
and U2934 (N_2934,N_2867,N_2823);
and U2935 (N_2935,N_2855,N_2871);
or U2936 (N_2936,N_2832,N_2853);
xnor U2937 (N_2937,N_2870,N_2820);
or U2938 (N_2938,N_2862,N_2824);
nor U2939 (N_2939,N_2842,N_2869);
nor U2940 (N_2940,N_2884,N_2939);
xor U2941 (N_2941,N_2931,N_2932);
nand U2942 (N_2942,N_2934,N_2896);
nor U2943 (N_2943,N_2887,N_2905);
nor U2944 (N_2944,N_2936,N_2911);
nor U2945 (N_2945,N_2891,N_2889);
and U2946 (N_2946,N_2910,N_2917);
nand U2947 (N_2947,N_2903,N_2918);
and U2948 (N_2948,N_2895,N_2914);
nor U2949 (N_2949,N_2922,N_2937);
or U2950 (N_2950,N_2893,N_2880);
or U2951 (N_2951,N_2938,N_2927);
nor U2952 (N_2952,N_2898,N_2902);
nor U2953 (N_2953,N_2923,N_2909);
nand U2954 (N_2954,N_2883,N_2920);
or U2955 (N_2955,N_2916,N_2899);
nor U2956 (N_2956,N_2908,N_2892);
or U2957 (N_2957,N_2912,N_2907);
and U2958 (N_2958,N_2886,N_2935);
nor U2959 (N_2959,N_2906,N_2904);
nand U2960 (N_2960,N_2929,N_2890);
and U2961 (N_2961,N_2882,N_2926);
xor U2962 (N_2962,N_2901,N_2933);
xnor U2963 (N_2963,N_2919,N_2897);
and U2964 (N_2964,N_2881,N_2913);
xnor U2965 (N_2965,N_2894,N_2928);
or U2966 (N_2966,N_2925,N_2900);
nand U2967 (N_2967,N_2888,N_2924);
nand U2968 (N_2968,N_2921,N_2930);
or U2969 (N_2969,N_2885,N_2915);
or U2970 (N_2970,N_2886,N_2933);
nor U2971 (N_2971,N_2939,N_2938);
and U2972 (N_2972,N_2933,N_2894);
nor U2973 (N_2973,N_2899,N_2926);
or U2974 (N_2974,N_2921,N_2934);
nand U2975 (N_2975,N_2936,N_2887);
or U2976 (N_2976,N_2882,N_2910);
nor U2977 (N_2977,N_2886,N_2902);
xor U2978 (N_2978,N_2881,N_2894);
nor U2979 (N_2979,N_2881,N_2916);
xnor U2980 (N_2980,N_2912,N_2894);
xnor U2981 (N_2981,N_2923,N_2908);
nor U2982 (N_2982,N_2915,N_2923);
nor U2983 (N_2983,N_2939,N_2905);
nand U2984 (N_2984,N_2895,N_2905);
xor U2985 (N_2985,N_2913,N_2922);
and U2986 (N_2986,N_2881,N_2928);
nand U2987 (N_2987,N_2887,N_2891);
xnor U2988 (N_2988,N_2915,N_2892);
nor U2989 (N_2989,N_2900,N_2939);
nand U2990 (N_2990,N_2890,N_2905);
nor U2991 (N_2991,N_2897,N_2938);
or U2992 (N_2992,N_2920,N_2882);
or U2993 (N_2993,N_2931,N_2881);
xor U2994 (N_2994,N_2909,N_2938);
nand U2995 (N_2995,N_2885,N_2907);
and U2996 (N_2996,N_2919,N_2880);
nor U2997 (N_2997,N_2928,N_2889);
nand U2998 (N_2998,N_2931,N_2896);
or U2999 (N_2999,N_2929,N_2885);
and UO_0 (O_0,N_2940,N_2980);
xnor UO_1 (O_1,N_2971,N_2982);
or UO_2 (O_2,N_2988,N_2972);
xnor UO_3 (O_3,N_2950,N_2973);
nand UO_4 (O_4,N_2998,N_2997);
and UO_5 (O_5,N_2955,N_2953);
xnor UO_6 (O_6,N_2941,N_2974);
xnor UO_7 (O_7,N_2967,N_2978);
or UO_8 (O_8,N_2951,N_2993);
or UO_9 (O_9,N_2994,N_2984);
nor UO_10 (O_10,N_2962,N_2944);
or UO_11 (O_11,N_2987,N_2959);
or UO_12 (O_12,N_2977,N_2956);
or UO_13 (O_13,N_2989,N_2999);
nor UO_14 (O_14,N_2969,N_2983);
xnor UO_15 (O_15,N_2958,N_2986);
or UO_16 (O_16,N_2942,N_2961);
or UO_17 (O_17,N_2992,N_2964);
or UO_18 (O_18,N_2949,N_2991);
and UO_19 (O_19,N_2943,N_2968);
nand UO_20 (O_20,N_2957,N_2975);
nand UO_21 (O_21,N_2995,N_2945);
or UO_22 (O_22,N_2952,N_2946);
or UO_23 (O_23,N_2948,N_2963);
and UO_24 (O_24,N_2965,N_2966);
nor UO_25 (O_25,N_2970,N_2954);
and UO_26 (O_26,N_2985,N_2981);
and UO_27 (O_27,N_2960,N_2990);
nor UO_28 (O_28,N_2976,N_2979);
and UO_29 (O_29,N_2947,N_2996);
nand UO_30 (O_30,N_2943,N_2992);
and UO_31 (O_31,N_2961,N_2996);
and UO_32 (O_32,N_2978,N_2962);
and UO_33 (O_33,N_2980,N_2972);
nor UO_34 (O_34,N_2976,N_2983);
nand UO_35 (O_35,N_2991,N_2947);
and UO_36 (O_36,N_2998,N_2967);
nor UO_37 (O_37,N_2967,N_2985);
xnor UO_38 (O_38,N_2961,N_2981);
nand UO_39 (O_39,N_2962,N_2948);
xnor UO_40 (O_40,N_2979,N_2993);
and UO_41 (O_41,N_2985,N_2999);
nand UO_42 (O_42,N_2947,N_2992);
xor UO_43 (O_43,N_2948,N_2974);
nor UO_44 (O_44,N_2953,N_2942);
and UO_45 (O_45,N_2952,N_2941);
xor UO_46 (O_46,N_2964,N_2941);
xnor UO_47 (O_47,N_2982,N_2962);
nand UO_48 (O_48,N_2979,N_2987);
and UO_49 (O_49,N_2998,N_2979);
xor UO_50 (O_50,N_2969,N_2980);
or UO_51 (O_51,N_2955,N_2951);
nand UO_52 (O_52,N_2997,N_2978);
nand UO_53 (O_53,N_2956,N_2995);
and UO_54 (O_54,N_2951,N_2944);
and UO_55 (O_55,N_2984,N_2989);
nand UO_56 (O_56,N_2980,N_2973);
and UO_57 (O_57,N_2986,N_2996);
or UO_58 (O_58,N_2988,N_2941);
and UO_59 (O_59,N_2976,N_2998);
nor UO_60 (O_60,N_2956,N_2953);
and UO_61 (O_61,N_2951,N_2942);
or UO_62 (O_62,N_2993,N_2982);
or UO_63 (O_63,N_2994,N_2961);
nand UO_64 (O_64,N_2985,N_2974);
nand UO_65 (O_65,N_2978,N_2947);
nand UO_66 (O_66,N_2961,N_2943);
nor UO_67 (O_67,N_2955,N_2982);
xor UO_68 (O_68,N_2949,N_2953);
or UO_69 (O_69,N_2995,N_2946);
and UO_70 (O_70,N_2946,N_2941);
and UO_71 (O_71,N_2978,N_2995);
and UO_72 (O_72,N_2950,N_2992);
xnor UO_73 (O_73,N_2955,N_2949);
nor UO_74 (O_74,N_2946,N_2954);
xnor UO_75 (O_75,N_2946,N_2963);
xor UO_76 (O_76,N_2990,N_2988);
xnor UO_77 (O_77,N_2980,N_2977);
nand UO_78 (O_78,N_2964,N_2977);
and UO_79 (O_79,N_2968,N_2945);
and UO_80 (O_80,N_2966,N_2981);
and UO_81 (O_81,N_2950,N_2944);
and UO_82 (O_82,N_2947,N_2956);
nand UO_83 (O_83,N_2972,N_2976);
nor UO_84 (O_84,N_2970,N_2948);
nor UO_85 (O_85,N_2998,N_2999);
or UO_86 (O_86,N_2985,N_2942);
nor UO_87 (O_87,N_2987,N_2978);
nor UO_88 (O_88,N_2979,N_2950);
and UO_89 (O_89,N_2963,N_2982);
nor UO_90 (O_90,N_2941,N_2970);
or UO_91 (O_91,N_2976,N_2965);
xor UO_92 (O_92,N_2964,N_2945);
nor UO_93 (O_93,N_2958,N_2977);
or UO_94 (O_94,N_2968,N_2948);
nor UO_95 (O_95,N_2956,N_2971);
and UO_96 (O_96,N_2994,N_2944);
nor UO_97 (O_97,N_2977,N_2981);
nand UO_98 (O_98,N_2987,N_2972);
xnor UO_99 (O_99,N_2943,N_2946);
xor UO_100 (O_100,N_2951,N_2969);
nor UO_101 (O_101,N_2998,N_2965);
or UO_102 (O_102,N_2985,N_2969);
xor UO_103 (O_103,N_2972,N_2992);
and UO_104 (O_104,N_2943,N_2950);
nand UO_105 (O_105,N_2985,N_2971);
or UO_106 (O_106,N_2953,N_2984);
nor UO_107 (O_107,N_2954,N_2957);
nor UO_108 (O_108,N_2994,N_2962);
nor UO_109 (O_109,N_2995,N_2958);
nor UO_110 (O_110,N_2981,N_2993);
and UO_111 (O_111,N_2959,N_2971);
xnor UO_112 (O_112,N_2952,N_2955);
nand UO_113 (O_113,N_2972,N_2955);
and UO_114 (O_114,N_2950,N_2951);
or UO_115 (O_115,N_2964,N_2979);
xor UO_116 (O_116,N_2996,N_2988);
or UO_117 (O_117,N_2984,N_2995);
and UO_118 (O_118,N_2971,N_2940);
xnor UO_119 (O_119,N_2949,N_2948);
nand UO_120 (O_120,N_2983,N_2986);
nor UO_121 (O_121,N_2970,N_2949);
and UO_122 (O_122,N_2979,N_2948);
xnor UO_123 (O_123,N_2961,N_2953);
or UO_124 (O_124,N_2984,N_2998);
nor UO_125 (O_125,N_2986,N_2982);
and UO_126 (O_126,N_2992,N_2970);
or UO_127 (O_127,N_2952,N_2969);
nor UO_128 (O_128,N_2984,N_2943);
nand UO_129 (O_129,N_2957,N_2974);
nand UO_130 (O_130,N_2994,N_2951);
nor UO_131 (O_131,N_2982,N_2958);
nor UO_132 (O_132,N_2999,N_2944);
nor UO_133 (O_133,N_2980,N_2963);
xor UO_134 (O_134,N_2966,N_2984);
xor UO_135 (O_135,N_2989,N_2955);
or UO_136 (O_136,N_2963,N_2966);
nand UO_137 (O_137,N_2948,N_2984);
xor UO_138 (O_138,N_2953,N_2983);
or UO_139 (O_139,N_2959,N_2956);
xor UO_140 (O_140,N_2969,N_2971);
xnor UO_141 (O_141,N_2941,N_2978);
nor UO_142 (O_142,N_2949,N_2962);
and UO_143 (O_143,N_2963,N_2945);
nor UO_144 (O_144,N_2961,N_2974);
or UO_145 (O_145,N_2967,N_2945);
nor UO_146 (O_146,N_2971,N_2961);
xnor UO_147 (O_147,N_2987,N_2998);
nor UO_148 (O_148,N_2947,N_2945);
or UO_149 (O_149,N_2945,N_2956);
nor UO_150 (O_150,N_2971,N_2974);
nand UO_151 (O_151,N_2979,N_2986);
nor UO_152 (O_152,N_2962,N_2984);
xnor UO_153 (O_153,N_2949,N_2963);
or UO_154 (O_154,N_2984,N_2979);
nor UO_155 (O_155,N_2977,N_2997);
xnor UO_156 (O_156,N_2963,N_2958);
nand UO_157 (O_157,N_2944,N_2949);
xnor UO_158 (O_158,N_2965,N_2979);
or UO_159 (O_159,N_2974,N_2953);
nand UO_160 (O_160,N_2955,N_2990);
xor UO_161 (O_161,N_2986,N_2948);
or UO_162 (O_162,N_2996,N_2966);
or UO_163 (O_163,N_2970,N_2991);
and UO_164 (O_164,N_2962,N_2940);
and UO_165 (O_165,N_2983,N_2959);
nor UO_166 (O_166,N_2981,N_2957);
xnor UO_167 (O_167,N_2959,N_2978);
nor UO_168 (O_168,N_2973,N_2942);
or UO_169 (O_169,N_2978,N_2958);
nand UO_170 (O_170,N_2992,N_2957);
and UO_171 (O_171,N_2979,N_2981);
and UO_172 (O_172,N_2973,N_2966);
or UO_173 (O_173,N_2948,N_2981);
or UO_174 (O_174,N_2977,N_2982);
xnor UO_175 (O_175,N_2946,N_2988);
nor UO_176 (O_176,N_2965,N_2994);
or UO_177 (O_177,N_2943,N_2967);
and UO_178 (O_178,N_2993,N_2963);
or UO_179 (O_179,N_2992,N_2968);
xnor UO_180 (O_180,N_2962,N_2988);
nand UO_181 (O_181,N_2959,N_2977);
xor UO_182 (O_182,N_2960,N_2969);
or UO_183 (O_183,N_2959,N_2957);
and UO_184 (O_184,N_2969,N_2988);
xor UO_185 (O_185,N_2989,N_2963);
nand UO_186 (O_186,N_2968,N_2961);
nor UO_187 (O_187,N_2958,N_2944);
xor UO_188 (O_188,N_2941,N_2971);
and UO_189 (O_189,N_2974,N_2954);
and UO_190 (O_190,N_2999,N_2966);
nor UO_191 (O_191,N_2971,N_2983);
and UO_192 (O_192,N_2964,N_2983);
or UO_193 (O_193,N_2960,N_2984);
or UO_194 (O_194,N_2983,N_2942);
and UO_195 (O_195,N_2970,N_2956);
and UO_196 (O_196,N_2961,N_2954);
nor UO_197 (O_197,N_2989,N_2956);
and UO_198 (O_198,N_2985,N_2947);
nand UO_199 (O_199,N_2976,N_2969);
nand UO_200 (O_200,N_2975,N_2958);
nand UO_201 (O_201,N_2968,N_2980);
nand UO_202 (O_202,N_2970,N_2976);
nor UO_203 (O_203,N_2998,N_2951);
xor UO_204 (O_204,N_2979,N_2961);
and UO_205 (O_205,N_2947,N_2997);
nor UO_206 (O_206,N_2991,N_2973);
nand UO_207 (O_207,N_2963,N_2960);
or UO_208 (O_208,N_2951,N_2995);
or UO_209 (O_209,N_2984,N_2944);
and UO_210 (O_210,N_2946,N_2986);
or UO_211 (O_211,N_2941,N_2957);
nor UO_212 (O_212,N_2948,N_2998);
nor UO_213 (O_213,N_2959,N_2940);
and UO_214 (O_214,N_2991,N_2980);
and UO_215 (O_215,N_2944,N_2947);
and UO_216 (O_216,N_2960,N_2995);
nand UO_217 (O_217,N_2944,N_2977);
or UO_218 (O_218,N_2979,N_2952);
nor UO_219 (O_219,N_2956,N_2994);
nand UO_220 (O_220,N_2958,N_2956);
and UO_221 (O_221,N_2963,N_2978);
and UO_222 (O_222,N_2996,N_2942);
xor UO_223 (O_223,N_2951,N_2959);
nand UO_224 (O_224,N_2995,N_2974);
nand UO_225 (O_225,N_2947,N_2987);
nand UO_226 (O_226,N_2991,N_2977);
nand UO_227 (O_227,N_2982,N_2984);
and UO_228 (O_228,N_2985,N_2966);
nand UO_229 (O_229,N_2965,N_2956);
or UO_230 (O_230,N_2942,N_2968);
nor UO_231 (O_231,N_2993,N_2998);
nand UO_232 (O_232,N_2950,N_2970);
nand UO_233 (O_233,N_2962,N_2991);
or UO_234 (O_234,N_2948,N_2952);
and UO_235 (O_235,N_2989,N_2966);
xor UO_236 (O_236,N_2998,N_2940);
or UO_237 (O_237,N_2996,N_2952);
and UO_238 (O_238,N_2992,N_2953);
or UO_239 (O_239,N_2950,N_2981);
nor UO_240 (O_240,N_2982,N_2975);
nand UO_241 (O_241,N_2976,N_2995);
xor UO_242 (O_242,N_2954,N_2984);
or UO_243 (O_243,N_2986,N_2998);
or UO_244 (O_244,N_2988,N_2984);
or UO_245 (O_245,N_2990,N_2997);
nand UO_246 (O_246,N_2967,N_2948);
xor UO_247 (O_247,N_2964,N_2968);
xnor UO_248 (O_248,N_2945,N_2944);
nand UO_249 (O_249,N_2964,N_2942);
xor UO_250 (O_250,N_2980,N_2959);
or UO_251 (O_251,N_2987,N_2953);
nand UO_252 (O_252,N_2940,N_2990);
or UO_253 (O_253,N_2993,N_2977);
and UO_254 (O_254,N_2948,N_2997);
xor UO_255 (O_255,N_2947,N_2976);
and UO_256 (O_256,N_2982,N_2989);
xnor UO_257 (O_257,N_2964,N_2958);
nand UO_258 (O_258,N_2971,N_2957);
xor UO_259 (O_259,N_2995,N_2968);
and UO_260 (O_260,N_2979,N_2942);
xnor UO_261 (O_261,N_2963,N_2965);
xor UO_262 (O_262,N_2945,N_2976);
nand UO_263 (O_263,N_2997,N_2975);
or UO_264 (O_264,N_2997,N_2964);
xnor UO_265 (O_265,N_2954,N_2967);
and UO_266 (O_266,N_2974,N_2982);
nand UO_267 (O_267,N_2952,N_2990);
and UO_268 (O_268,N_2975,N_2966);
nor UO_269 (O_269,N_2951,N_2984);
xor UO_270 (O_270,N_2998,N_2981);
nand UO_271 (O_271,N_2970,N_2998);
xor UO_272 (O_272,N_2949,N_2975);
xnor UO_273 (O_273,N_2966,N_2994);
nor UO_274 (O_274,N_2987,N_2961);
xor UO_275 (O_275,N_2980,N_2944);
and UO_276 (O_276,N_2965,N_2952);
and UO_277 (O_277,N_2967,N_2946);
nand UO_278 (O_278,N_2971,N_2942);
nor UO_279 (O_279,N_2998,N_2975);
xor UO_280 (O_280,N_2981,N_2972);
or UO_281 (O_281,N_2941,N_2981);
or UO_282 (O_282,N_2981,N_2986);
nand UO_283 (O_283,N_2983,N_2987);
or UO_284 (O_284,N_2975,N_2992);
and UO_285 (O_285,N_2963,N_2962);
nand UO_286 (O_286,N_2979,N_2958);
nand UO_287 (O_287,N_2995,N_2982);
nand UO_288 (O_288,N_2944,N_2991);
or UO_289 (O_289,N_2968,N_2978);
or UO_290 (O_290,N_2950,N_2958);
nand UO_291 (O_291,N_2974,N_2983);
nor UO_292 (O_292,N_2982,N_2949);
nand UO_293 (O_293,N_2942,N_2988);
or UO_294 (O_294,N_2991,N_2955);
nor UO_295 (O_295,N_2941,N_2994);
or UO_296 (O_296,N_2956,N_2987);
nor UO_297 (O_297,N_2946,N_2972);
or UO_298 (O_298,N_2980,N_2946);
nand UO_299 (O_299,N_2989,N_2997);
nand UO_300 (O_300,N_2945,N_2978);
nand UO_301 (O_301,N_2987,N_2980);
xnor UO_302 (O_302,N_2991,N_2964);
nand UO_303 (O_303,N_2998,N_2943);
nor UO_304 (O_304,N_2946,N_2964);
or UO_305 (O_305,N_2944,N_2971);
and UO_306 (O_306,N_2978,N_2979);
and UO_307 (O_307,N_2945,N_2970);
nand UO_308 (O_308,N_2991,N_2941);
nand UO_309 (O_309,N_2984,N_2958);
and UO_310 (O_310,N_2984,N_2964);
and UO_311 (O_311,N_2971,N_2973);
nand UO_312 (O_312,N_2954,N_2944);
nor UO_313 (O_313,N_2995,N_2994);
or UO_314 (O_314,N_2949,N_2987);
or UO_315 (O_315,N_2977,N_2992);
xor UO_316 (O_316,N_2995,N_2947);
nand UO_317 (O_317,N_2999,N_2951);
and UO_318 (O_318,N_2975,N_2991);
nor UO_319 (O_319,N_2989,N_2995);
nand UO_320 (O_320,N_2944,N_2966);
nor UO_321 (O_321,N_2994,N_2948);
or UO_322 (O_322,N_2990,N_2991);
xnor UO_323 (O_323,N_2968,N_2990);
or UO_324 (O_324,N_2988,N_2952);
nand UO_325 (O_325,N_2943,N_2947);
and UO_326 (O_326,N_2968,N_2952);
nand UO_327 (O_327,N_2962,N_2956);
xnor UO_328 (O_328,N_2986,N_2944);
nand UO_329 (O_329,N_2965,N_2950);
or UO_330 (O_330,N_2953,N_2980);
xnor UO_331 (O_331,N_2980,N_2975);
and UO_332 (O_332,N_2997,N_2976);
and UO_333 (O_333,N_2979,N_2992);
and UO_334 (O_334,N_2991,N_2981);
nand UO_335 (O_335,N_2950,N_2954);
xnor UO_336 (O_336,N_2965,N_2943);
and UO_337 (O_337,N_2971,N_2951);
or UO_338 (O_338,N_2975,N_2965);
or UO_339 (O_339,N_2971,N_2992);
nand UO_340 (O_340,N_2958,N_2943);
nand UO_341 (O_341,N_2974,N_2967);
nand UO_342 (O_342,N_2974,N_2959);
nor UO_343 (O_343,N_2983,N_2965);
nand UO_344 (O_344,N_2962,N_2980);
nand UO_345 (O_345,N_2944,N_2965);
and UO_346 (O_346,N_2996,N_2979);
or UO_347 (O_347,N_2962,N_2964);
nand UO_348 (O_348,N_2955,N_2995);
or UO_349 (O_349,N_2956,N_2990);
nor UO_350 (O_350,N_2993,N_2978);
and UO_351 (O_351,N_2967,N_2963);
xnor UO_352 (O_352,N_2964,N_2987);
or UO_353 (O_353,N_2951,N_2981);
xnor UO_354 (O_354,N_2994,N_2969);
xnor UO_355 (O_355,N_2983,N_2989);
nor UO_356 (O_356,N_2953,N_2990);
nor UO_357 (O_357,N_2988,N_2953);
nor UO_358 (O_358,N_2958,N_2949);
nor UO_359 (O_359,N_2978,N_2972);
and UO_360 (O_360,N_2999,N_2979);
nand UO_361 (O_361,N_2977,N_2978);
xnor UO_362 (O_362,N_2946,N_2999);
xnor UO_363 (O_363,N_2984,N_2972);
or UO_364 (O_364,N_2948,N_2972);
nor UO_365 (O_365,N_2978,N_2940);
nand UO_366 (O_366,N_2996,N_2976);
and UO_367 (O_367,N_2972,N_2968);
nor UO_368 (O_368,N_2944,N_2973);
or UO_369 (O_369,N_2991,N_2948);
and UO_370 (O_370,N_2954,N_2991);
or UO_371 (O_371,N_2977,N_2941);
xor UO_372 (O_372,N_2994,N_2946);
nor UO_373 (O_373,N_2969,N_2944);
nand UO_374 (O_374,N_2994,N_2971);
nand UO_375 (O_375,N_2967,N_2980);
and UO_376 (O_376,N_2986,N_2967);
and UO_377 (O_377,N_2995,N_2990);
xor UO_378 (O_378,N_2968,N_2941);
nand UO_379 (O_379,N_2977,N_2983);
nor UO_380 (O_380,N_2947,N_2949);
or UO_381 (O_381,N_2958,N_2952);
nor UO_382 (O_382,N_2993,N_2965);
or UO_383 (O_383,N_2956,N_2955);
nand UO_384 (O_384,N_2943,N_2949);
nor UO_385 (O_385,N_2960,N_2950);
or UO_386 (O_386,N_2988,N_2977);
nor UO_387 (O_387,N_2991,N_2995);
xor UO_388 (O_388,N_2973,N_2985);
and UO_389 (O_389,N_2968,N_2979);
nor UO_390 (O_390,N_2942,N_2943);
xnor UO_391 (O_391,N_2988,N_2998);
xor UO_392 (O_392,N_2984,N_2980);
xor UO_393 (O_393,N_2994,N_2974);
xor UO_394 (O_394,N_2949,N_2945);
or UO_395 (O_395,N_2956,N_2997);
and UO_396 (O_396,N_2973,N_2945);
xor UO_397 (O_397,N_2965,N_2957);
nor UO_398 (O_398,N_2956,N_2985);
nand UO_399 (O_399,N_2953,N_2951);
xnor UO_400 (O_400,N_2964,N_2980);
nor UO_401 (O_401,N_2966,N_2990);
or UO_402 (O_402,N_2959,N_2942);
or UO_403 (O_403,N_2987,N_2993);
or UO_404 (O_404,N_2941,N_2961);
and UO_405 (O_405,N_2971,N_2958);
xnor UO_406 (O_406,N_2989,N_2980);
nor UO_407 (O_407,N_2946,N_2978);
or UO_408 (O_408,N_2954,N_2973);
nand UO_409 (O_409,N_2980,N_2986);
nand UO_410 (O_410,N_2995,N_2998);
xor UO_411 (O_411,N_2948,N_2942);
or UO_412 (O_412,N_2961,N_2966);
nor UO_413 (O_413,N_2970,N_2940);
nor UO_414 (O_414,N_2949,N_2981);
and UO_415 (O_415,N_2951,N_2978);
xnor UO_416 (O_416,N_2974,N_2960);
or UO_417 (O_417,N_2978,N_2991);
nor UO_418 (O_418,N_2948,N_2990);
xor UO_419 (O_419,N_2958,N_2993);
xnor UO_420 (O_420,N_2950,N_2959);
nor UO_421 (O_421,N_2991,N_2976);
or UO_422 (O_422,N_2946,N_2983);
xor UO_423 (O_423,N_2995,N_2979);
and UO_424 (O_424,N_2941,N_2998);
nand UO_425 (O_425,N_2947,N_2984);
nand UO_426 (O_426,N_2978,N_2943);
nor UO_427 (O_427,N_2942,N_2981);
and UO_428 (O_428,N_2959,N_2988);
xnor UO_429 (O_429,N_2989,N_2944);
xnor UO_430 (O_430,N_2975,N_2978);
nand UO_431 (O_431,N_2991,N_2993);
nand UO_432 (O_432,N_2997,N_2967);
nor UO_433 (O_433,N_2969,N_2987);
xnor UO_434 (O_434,N_2970,N_2977);
xnor UO_435 (O_435,N_2968,N_2984);
or UO_436 (O_436,N_2961,N_2970);
nand UO_437 (O_437,N_2948,N_2958);
xnor UO_438 (O_438,N_2949,N_2941);
and UO_439 (O_439,N_2961,N_2948);
nor UO_440 (O_440,N_2990,N_2975);
and UO_441 (O_441,N_2995,N_2948);
and UO_442 (O_442,N_2949,N_2976);
xor UO_443 (O_443,N_2994,N_2945);
xnor UO_444 (O_444,N_2956,N_2960);
and UO_445 (O_445,N_2948,N_2988);
and UO_446 (O_446,N_2958,N_2945);
and UO_447 (O_447,N_2956,N_2951);
xor UO_448 (O_448,N_2958,N_2957);
and UO_449 (O_449,N_2962,N_2954);
or UO_450 (O_450,N_2954,N_2951);
nand UO_451 (O_451,N_2973,N_2993);
or UO_452 (O_452,N_2966,N_2958);
and UO_453 (O_453,N_2957,N_2964);
or UO_454 (O_454,N_2941,N_2955);
nand UO_455 (O_455,N_2970,N_2985);
xnor UO_456 (O_456,N_2974,N_2979);
xor UO_457 (O_457,N_2943,N_2988);
nand UO_458 (O_458,N_2971,N_2964);
and UO_459 (O_459,N_2961,N_2962);
nor UO_460 (O_460,N_2975,N_2995);
nand UO_461 (O_461,N_2954,N_2964);
nand UO_462 (O_462,N_2998,N_2964);
xnor UO_463 (O_463,N_2947,N_2971);
nor UO_464 (O_464,N_2990,N_2950);
nor UO_465 (O_465,N_2956,N_2996);
and UO_466 (O_466,N_2963,N_2999);
nand UO_467 (O_467,N_2970,N_2968);
or UO_468 (O_468,N_2957,N_2955);
xnor UO_469 (O_469,N_2970,N_2944);
and UO_470 (O_470,N_2973,N_2984);
nand UO_471 (O_471,N_2957,N_2982);
and UO_472 (O_472,N_2986,N_2977);
nand UO_473 (O_473,N_2983,N_2985);
xor UO_474 (O_474,N_2975,N_2996);
or UO_475 (O_475,N_2992,N_2982);
xnor UO_476 (O_476,N_2977,N_2998);
nand UO_477 (O_477,N_2963,N_2968);
or UO_478 (O_478,N_2986,N_2974);
nor UO_479 (O_479,N_2980,N_2997);
or UO_480 (O_480,N_2970,N_2969);
or UO_481 (O_481,N_2982,N_2947);
xnor UO_482 (O_482,N_2966,N_2988);
nor UO_483 (O_483,N_2988,N_2992);
xnor UO_484 (O_484,N_2968,N_2951);
and UO_485 (O_485,N_2975,N_2956);
and UO_486 (O_486,N_2943,N_2975);
or UO_487 (O_487,N_2981,N_2952);
xnor UO_488 (O_488,N_2971,N_2993);
or UO_489 (O_489,N_2965,N_2977);
xnor UO_490 (O_490,N_2979,N_2990);
nand UO_491 (O_491,N_2950,N_2975);
or UO_492 (O_492,N_2962,N_2998);
nor UO_493 (O_493,N_2980,N_2992);
and UO_494 (O_494,N_2950,N_2998);
or UO_495 (O_495,N_2974,N_2964);
nor UO_496 (O_496,N_2948,N_2944);
and UO_497 (O_497,N_2973,N_2975);
or UO_498 (O_498,N_2977,N_2952);
nand UO_499 (O_499,N_2973,N_2982);
endmodule