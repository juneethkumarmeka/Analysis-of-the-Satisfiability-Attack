module basic_500_3000_500_60_levels_5xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_27,In_123);
or U1 (N_1,In_448,In_319);
nand U2 (N_2,In_165,In_79);
or U3 (N_3,In_28,In_9);
and U4 (N_4,In_218,In_174);
or U5 (N_5,In_492,In_45);
xnor U6 (N_6,In_231,In_168);
nand U7 (N_7,In_56,In_294);
nand U8 (N_8,In_110,In_138);
nor U9 (N_9,In_316,In_359);
nand U10 (N_10,In_30,In_118);
or U11 (N_11,In_115,In_190);
nor U12 (N_12,In_83,In_340);
and U13 (N_13,In_212,In_345);
nand U14 (N_14,In_36,In_247);
nand U15 (N_15,In_409,In_251);
xor U16 (N_16,In_362,In_235);
nand U17 (N_17,In_203,In_423);
xor U18 (N_18,In_351,In_390);
xor U19 (N_19,In_446,In_274);
nand U20 (N_20,In_223,In_222);
xor U21 (N_21,In_177,In_140);
or U22 (N_22,In_131,In_93);
and U23 (N_23,In_114,In_263);
xor U24 (N_24,In_332,In_148);
xor U25 (N_25,In_474,In_358);
or U26 (N_26,In_323,In_216);
and U27 (N_27,In_293,In_239);
nand U28 (N_28,In_167,In_98);
and U29 (N_29,In_401,In_169);
and U30 (N_30,In_188,In_387);
nor U31 (N_31,In_443,In_17);
xnor U32 (N_32,In_262,In_346);
nor U33 (N_33,In_145,In_490);
or U34 (N_34,In_287,In_107);
xnor U35 (N_35,In_71,In_483);
or U36 (N_36,In_24,In_399);
and U37 (N_37,In_105,In_26);
nor U38 (N_38,In_19,In_350);
xor U39 (N_39,In_108,In_261);
or U40 (N_40,In_289,In_52);
or U41 (N_41,In_146,In_42);
or U42 (N_42,In_199,In_322);
and U43 (N_43,In_183,In_229);
nor U44 (N_44,In_18,In_248);
and U45 (N_45,In_318,In_429);
or U46 (N_46,In_259,In_102);
and U47 (N_47,In_193,In_435);
xnor U48 (N_48,In_296,In_163);
or U49 (N_49,In_187,In_415);
or U50 (N_50,N_29,In_134);
or U51 (N_51,N_26,In_72);
xnor U52 (N_52,In_40,In_121);
nor U53 (N_53,In_74,In_484);
or U54 (N_54,In_445,In_152);
or U55 (N_55,In_220,In_473);
nor U56 (N_56,In_477,In_325);
nor U57 (N_57,In_170,In_449);
and U58 (N_58,In_1,In_428);
nand U59 (N_59,In_126,In_376);
nor U60 (N_60,In_299,In_256);
nor U61 (N_61,N_2,In_444);
and U62 (N_62,In_315,In_420);
nand U63 (N_63,In_57,In_433);
nor U64 (N_64,In_86,In_275);
nand U65 (N_65,In_156,In_427);
nand U66 (N_66,In_291,In_411);
nand U67 (N_67,In_103,In_354);
nand U68 (N_68,In_61,In_476);
or U69 (N_69,In_150,In_158);
nor U70 (N_70,In_268,In_8);
and U71 (N_71,In_122,In_185);
and U72 (N_72,In_4,In_422);
nand U73 (N_73,In_64,In_491);
nand U74 (N_74,In_392,In_436);
or U75 (N_75,In_374,In_77);
nand U76 (N_76,In_280,In_100);
xor U77 (N_77,In_207,N_45);
or U78 (N_78,N_0,N_27);
and U79 (N_79,In_456,In_246);
nor U80 (N_80,In_394,N_39);
nand U81 (N_81,In_113,In_485);
nor U82 (N_82,In_137,N_41);
nor U83 (N_83,In_157,In_405);
nor U84 (N_84,In_241,In_80);
nor U85 (N_85,In_398,In_92);
or U86 (N_86,N_32,In_69);
and U87 (N_87,In_457,In_230);
xnor U88 (N_88,In_281,In_437);
or U89 (N_89,In_391,In_111);
nor U90 (N_90,In_438,In_499);
xor U91 (N_91,In_78,In_11);
and U92 (N_92,In_303,In_39);
xnor U93 (N_93,In_160,In_87);
nor U94 (N_94,In_141,N_43);
xnor U95 (N_95,In_408,In_482);
or U96 (N_96,In_326,N_46);
nand U97 (N_97,In_224,In_338);
nor U98 (N_98,In_339,In_147);
and U99 (N_99,In_439,In_67);
nor U100 (N_100,N_44,In_35);
or U101 (N_101,N_50,In_356);
nor U102 (N_102,In_16,In_81);
nand U103 (N_103,In_455,In_397);
nand U104 (N_104,In_2,In_305);
nor U105 (N_105,In_43,In_198);
nand U106 (N_106,In_329,In_493);
nor U107 (N_107,In_292,In_426);
xor U108 (N_108,In_347,In_378);
nor U109 (N_109,N_71,In_442);
nand U110 (N_110,In_424,In_191);
and U111 (N_111,In_215,In_37);
and U112 (N_112,N_54,N_90);
or U113 (N_113,In_307,In_125);
xnor U114 (N_114,In_3,In_182);
nand U115 (N_115,In_59,N_67);
nor U116 (N_116,In_380,In_213);
or U117 (N_117,N_56,In_425);
or U118 (N_118,In_400,N_69);
or U119 (N_119,N_13,In_116);
and U120 (N_120,In_388,In_284);
nor U121 (N_121,In_278,In_496);
xor U122 (N_122,In_447,In_10);
nand U123 (N_123,In_166,In_334);
nand U124 (N_124,In_197,In_469);
and U125 (N_125,In_497,In_430);
or U126 (N_126,In_244,N_17);
nor U127 (N_127,In_478,In_498);
nor U128 (N_128,In_300,In_90);
nor U129 (N_129,In_29,In_161);
nand U130 (N_130,N_98,In_369);
xor U131 (N_131,In_432,In_258);
or U132 (N_132,In_253,In_227);
nor U133 (N_133,In_34,In_416);
or U134 (N_134,N_70,In_273);
or U135 (N_135,In_48,In_49);
nand U136 (N_136,In_277,In_310);
nor U137 (N_137,N_61,In_327);
nor U138 (N_138,In_129,In_381);
nand U139 (N_139,In_46,N_95);
or U140 (N_140,In_341,N_87);
nand U141 (N_141,N_58,N_52);
and U142 (N_142,N_30,In_196);
xnor U143 (N_143,In_272,In_384);
nor U144 (N_144,In_88,In_269);
xnor U145 (N_145,N_18,In_421);
nor U146 (N_146,In_266,In_373);
and U147 (N_147,In_379,N_92);
or U148 (N_148,In_342,In_464);
nor U149 (N_149,In_245,In_309);
nor U150 (N_150,N_1,N_109);
nor U151 (N_151,In_142,N_91);
nor U152 (N_152,In_209,N_77);
nor U153 (N_153,In_466,N_53);
or U154 (N_154,N_120,N_135);
and U155 (N_155,In_65,In_252);
nor U156 (N_156,In_402,In_104);
nor U157 (N_157,In_51,N_51);
and U158 (N_158,In_331,In_414);
nor U159 (N_159,N_112,In_431);
and U160 (N_160,In_404,N_94);
and U161 (N_161,In_225,In_73);
nand U162 (N_162,In_479,In_171);
and U163 (N_163,In_130,N_4);
or U164 (N_164,In_386,N_97);
nand U165 (N_165,In_312,N_12);
xnor U166 (N_166,N_142,In_189);
xnor U167 (N_167,N_101,In_58);
and U168 (N_168,In_234,N_100);
nand U169 (N_169,N_78,N_116);
nor U170 (N_170,N_20,In_120);
and U171 (N_171,N_49,In_321);
nand U172 (N_172,In_194,In_205);
nand U173 (N_173,In_418,N_14);
xor U174 (N_174,N_104,In_12);
and U175 (N_175,In_179,In_279);
or U176 (N_176,N_88,In_249);
nand U177 (N_177,N_60,In_270);
or U178 (N_178,In_357,In_144);
or U179 (N_179,In_14,N_7);
or U180 (N_180,In_395,In_460);
nor U181 (N_181,In_192,In_396);
nand U182 (N_182,In_117,N_34);
xnor U183 (N_183,N_106,In_47);
nor U184 (N_184,In_172,In_330);
nand U185 (N_185,In_393,In_463);
nor U186 (N_186,In_176,In_434);
and U187 (N_187,N_121,N_146);
nor U188 (N_188,In_320,In_233);
xnor U189 (N_189,N_108,In_406);
and U190 (N_190,In_481,N_81);
and U191 (N_191,In_462,In_132);
or U192 (N_192,In_385,In_53);
and U193 (N_193,In_154,In_301);
xor U194 (N_194,N_138,N_21);
xnor U195 (N_195,In_295,N_127);
nor U196 (N_196,In_128,In_290);
nor U197 (N_197,In_135,In_186);
nor U198 (N_198,In_89,In_136);
or U199 (N_199,In_201,In_0);
and U200 (N_200,In_271,In_441);
or U201 (N_201,In_200,In_243);
nor U202 (N_202,N_118,In_317);
xnor U203 (N_203,N_10,In_349);
and U204 (N_204,N_181,In_265);
nor U205 (N_205,N_150,In_124);
nand U206 (N_206,In_282,N_131);
nand U207 (N_207,In_459,N_157);
nor U208 (N_208,In_286,In_242);
nand U209 (N_209,In_153,In_23);
nor U210 (N_210,N_66,In_5);
or U211 (N_211,In_276,In_151);
or U212 (N_212,In_335,N_74);
nor U213 (N_213,N_147,N_160);
and U214 (N_214,In_297,In_21);
and U215 (N_215,N_197,N_175);
xnor U216 (N_216,N_130,In_472);
nand U217 (N_217,In_6,In_94);
nor U218 (N_218,N_141,N_174);
xnor U219 (N_219,N_193,In_68);
and U220 (N_220,N_25,N_195);
xnor U221 (N_221,In_375,In_238);
and U222 (N_222,In_368,In_288);
xnor U223 (N_223,In_377,In_97);
and U224 (N_224,In_383,N_96);
and U225 (N_225,N_165,N_166);
or U226 (N_226,In_15,N_75);
and U227 (N_227,In_363,In_236);
and U228 (N_228,N_158,In_344);
nand U229 (N_229,In_311,N_83);
or U230 (N_230,In_336,N_151);
nor U231 (N_231,In_410,N_24);
and U232 (N_232,N_172,In_407);
nor U233 (N_233,In_221,In_210);
nand U234 (N_234,N_185,N_188);
nor U235 (N_235,N_16,In_44);
nand U236 (N_236,In_453,In_264);
or U237 (N_237,N_8,In_181);
nor U238 (N_238,In_159,In_328);
and U239 (N_239,N_136,In_475);
nor U240 (N_240,In_257,N_37);
nor U241 (N_241,In_133,N_125);
nand U242 (N_242,N_62,In_454);
or U243 (N_243,N_113,N_22);
nand U244 (N_244,N_82,N_59);
and U245 (N_245,In_155,In_333);
nand U246 (N_246,In_254,In_458);
nor U247 (N_247,In_31,In_95);
nor U248 (N_248,N_153,In_360);
nor U249 (N_249,N_145,N_171);
or U250 (N_250,N_248,N_202);
or U251 (N_251,N_207,In_467);
nand U252 (N_252,N_216,In_495);
or U253 (N_253,In_109,N_155);
and U254 (N_254,N_240,In_419);
or U255 (N_255,In_149,In_480);
and U256 (N_256,In_285,In_370);
nand U257 (N_257,N_222,N_111);
xor U258 (N_258,N_68,In_139);
xnor U259 (N_259,N_161,N_236);
and U260 (N_260,N_233,N_182);
nor U261 (N_261,In_440,N_184);
or U262 (N_262,N_198,In_451);
nor U263 (N_263,N_93,N_132);
nand U264 (N_264,In_364,In_66);
nor U265 (N_265,In_494,In_240);
nor U266 (N_266,N_215,N_114);
nand U267 (N_267,N_231,In_372);
nor U268 (N_268,N_179,In_412);
and U269 (N_269,In_76,N_128);
or U270 (N_270,In_226,In_33);
and U271 (N_271,In_232,N_177);
nor U272 (N_272,N_249,N_156);
nand U273 (N_273,N_204,In_206);
and U274 (N_274,N_134,N_219);
nand U275 (N_275,N_224,N_201);
and U276 (N_276,In_162,N_119);
nor U277 (N_277,In_417,N_221);
or U278 (N_278,N_103,In_204);
or U279 (N_279,N_140,N_76);
or U280 (N_280,In_403,N_220);
or U281 (N_281,In_313,N_167);
nand U282 (N_282,N_163,N_57);
xnor U283 (N_283,N_169,In_217);
and U284 (N_284,In_308,N_187);
and U285 (N_285,N_123,N_159);
nor U286 (N_286,N_65,N_189);
xor U287 (N_287,N_238,N_143);
and U288 (N_288,In_450,In_348);
and U289 (N_289,In_255,N_206);
or U290 (N_290,In_465,In_20);
or U291 (N_291,In_119,In_382);
nor U292 (N_292,N_168,N_214);
or U293 (N_293,N_162,N_40);
and U294 (N_294,In_70,In_62);
nand U295 (N_295,N_79,In_84);
nor U296 (N_296,N_64,N_102);
nand U297 (N_297,In_260,In_366);
nor U298 (N_298,N_237,In_237);
or U299 (N_299,N_227,N_5);
and U300 (N_300,N_186,In_112);
or U301 (N_301,In_343,In_355);
and U302 (N_302,In_75,N_235);
and U303 (N_303,In_60,N_275);
and U304 (N_304,In_211,N_218);
xor U305 (N_305,In_208,N_242);
nor U306 (N_306,N_38,N_253);
or U307 (N_307,N_288,In_488);
or U308 (N_308,N_85,In_314);
and U309 (N_309,In_32,N_295);
nor U310 (N_310,In_468,N_276);
nor U311 (N_311,N_99,In_54);
and U312 (N_312,N_280,N_164);
nor U313 (N_313,In_195,N_247);
nor U314 (N_314,In_487,In_178);
nor U315 (N_315,N_126,N_234);
and U316 (N_316,N_208,N_265);
and U317 (N_317,In_22,In_470);
nand U318 (N_318,N_272,N_180);
xnor U319 (N_319,In_202,In_214);
and U320 (N_320,In_461,N_255);
nor U321 (N_321,N_11,N_107);
nand U322 (N_322,N_42,N_298);
xnor U323 (N_323,N_285,N_48);
and U324 (N_324,N_84,N_200);
and U325 (N_325,In_25,In_283);
or U326 (N_326,N_190,N_115);
and U327 (N_327,N_261,N_294);
nand U328 (N_328,N_279,N_241);
nor U329 (N_329,N_73,In_471);
or U330 (N_330,N_256,N_258);
and U331 (N_331,N_278,N_252);
nand U332 (N_332,N_270,N_284);
nand U333 (N_333,N_196,In_365);
or U334 (N_334,N_277,N_228);
nor U335 (N_335,N_144,N_243);
xnor U336 (N_336,N_6,In_367);
or U337 (N_337,N_225,N_72);
nor U338 (N_338,In_304,In_452);
nand U339 (N_339,N_229,N_9);
or U340 (N_340,N_210,N_251);
nand U341 (N_341,N_269,N_80);
and U342 (N_342,In_219,N_226);
or U343 (N_343,In_63,N_205);
nor U344 (N_344,In_302,N_290);
and U345 (N_345,N_287,N_263);
nor U346 (N_346,In_352,N_211);
or U347 (N_347,N_35,N_239);
nand U348 (N_348,N_124,N_259);
nand U349 (N_349,In_101,N_289);
or U350 (N_350,In_267,N_105);
and U351 (N_351,N_309,N_331);
nor U352 (N_352,In_85,N_254);
xor U353 (N_353,In_298,In_184);
nor U354 (N_354,N_274,N_203);
nor U355 (N_355,In_353,N_267);
and U356 (N_356,N_329,N_271);
or U357 (N_357,N_273,N_336);
and U358 (N_358,N_301,N_323);
nor U359 (N_359,N_311,N_335);
nand U360 (N_360,N_152,N_347);
nand U361 (N_361,N_86,N_324);
nand U362 (N_362,N_117,N_192);
and U363 (N_363,N_133,N_304);
or U364 (N_364,In_337,In_38);
xor U365 (N_365,N_232,In_164);
nor U366 (N_366,In_106,N_317);
nand U367 (N_367,In_180,N_149);
or U368 (N_368,N_268,N_31);
xor U369 (N_369,In_55,N_310);
and U370 (N_370,N_302,N_313);
nand U371 (N_371,N_318,N_129);
and U372 (N_372,N_303,N_282);
xor U373 (N_373,N_306,N_199);
and U374 (N_374,N_305,N_343);
nor U375 (N_375,In_389,In_96);
nor U376 (N_376,N_346,N_325);
and U377 (N_377,N_348,In_13);
nand U378 (N_378,N_33,N_209);
nand U379 (N_379,N_334,N_3);
or U380 (N_380,N_173,N_63);
or U381 (N_381,N_291,In_306);
and U382 (N_382,In_143,N_191);
nand U383 (N_383,In_175,In_413);
or U384 (N_384,N_296,N_178);
nor U385 (N_385,In_99,N_15);
and U386 (N_386,N_308,N_328);
and U387 (N_387,N_217,N_344);
nor U388 (N_388,N_110,N_300);
nor U389 (N_389,N_330,N_194);
nor U390 (N_390,In_173,In_228);
xnor U391 (N_391,N_257,N_170);
and U392 (N_392,In_7,N_286);
and U393 (N_393,N_339,N_176);
and U394 (N_394,In_361,N_246);
or U395 (N_395,N_212,N_319);
nand U396 (N_396,N_154,N_315);
nand U397 (N_397,N_312,N_321);
xor U398 (N_398,N_139,N_341);
nor U399 (N_399,N_137,N_283);
or U400 (N_400,N_122,In_82);
or U401 (N_401,N_337,N_394);
nand U402 (N_402,N_230,In_50);
nor U403 (N_403,N_342,N_385);
nand U404 (N_404,N_390,N_345);
nor U405 (N_405,In_371,In_250);
nand U406 (N_406,N_362,N_89);
or U407 (N_407,N_371,N_355);
xnor U408 (N_408,In_41,N_387);
nor U409 (N_409,N_250,N_367);
and U410 (N_410,N_380,N_292);
nand U411 (N_411,N_244,N_372);
nor U412 (N_412,N_326,N_322);
and U413 (N_413,N_293,N_327);
xor U414 (N_414,N_213,N_23);
nand U415 (N_415,N_359,N_389);
xnor U416 (N_416,N_375,N_340);
xor U417 (N_417,N_351,N_368);
nor U418 (N_418,In_486,N_382);
and U419 (N_419,N_378,N_245);
and U420 (N_420,N_266,N_379);
nand U421 (N_421,N_47,N_352);
xnor U422 (N_422,N_314,N_338);
nand U423 (N_423,N_395,N_366);
xor U424 (N_424,N_281,N_358);
xnor U425 (N_425,N_384,N_376);
xnor U426 (N_426,N_396,N_307);
or U427 (N_427,N_361,N_360);
xor U428 (N_428,N_388,N_354);
nor U429 (N_429,N_353,In_324);
and U430 (N_430,N_148,N_297);
and U431 (N_431,N_262,In_91);
or U432 (N_432,N_320,N_386);
or U433 (N_433,N_350,N_391);
nand U434 (N_434,N_383,N_28);
and U435 (N_435,N_392,N_260);
and U436 (N_436,N_264,N_223);
or U437 (N_437,In_127,N_393);
and U438 (N_438,In_489,N_349);
xnor U439 (N_439,N_333,N_316);
or U440 (N_440,N_397,N_398);
and U441 (N_441,N_183,N_399);
or U442 (N_442,N_381,N_364);
xor U443 (N_443,N_374,N_369);
or U444 (N_444,N_332,N_299);
and U445 (N_445,N_363,N_370);
nor U446 (N_446,N_356,N_365);
or U447 (N_447,N_377,N_36);
or U448 (N_448,N_55,N_19);
nand U449 (N_449,N_373,N_357);
nand U450 (N_450,N_421,N_402);
or U451 (N_451,N_415,N_418);
or U452 (N_452,N_446,N_419);
and U453 (N_453,N_407,N_440);
or U454 (N_454,N_428,N_430);
and U455 (N_455,N_448,N_444);
nand U456 (N_456,N_412,N_404);
or U457 (N_457,N_423,N_424);
nor U458 (N_458,N_443,N_429);
nand U459 (N_459,N_437,N_401);
and U460 (N_460,N_422,N_433);
xnor U461 (N_461,N_406,N_410);
nor U462 (N_462,N_445,N_434);
xnor U463 (N_463,N_405,N_400);
xor U464 (N_464,N_411,N_439);
or U465 (N_465,N_414,N_432);
or U466 (N_466,N_426,N_425);
or U467 (N_467,N_416,N_413);
or U468 (N_468,N_403,N_420);
or U469 (N_469,N_447,N_417);
nand U470 (N_470,N_438,N_441);
xnor U471 (N_471,N_409,N_449);
nor U472 (N_472,N_435,N_408);
or U473 (N_473,N_427,N_442);
or U474 (N_474,N_436,N_431);
xnor U475 (N_475,N_438,N_418);
nand U476 (N_476,N_449,N_427);
and U477 (N_477,N_434,N_411);
xnor U478 (N_478,N_412,N_445);
nand U479 (N_479,N_441,N_433);
nand U480 (N_480,N_436,N_401);
or U481 (N_481,N_429,N_402);
nand U482 (N_482,N_419,N_428);
nand U483 (N_483,N_423,N_444);
and U484 (N_484,N_406,N_437);
nor U485 (N_485,N_441,N_446);
nor U486 (N_486,N_405,N_428);
nand U487 (N_487,N_400,N_426);
or U488 (N_488,N_438,N_414);
and U489 (N_489,N_403,N_425);
nor U490 (N_490,N_436,N_447);
and U491 (N_491,N_403,N_429);
or U492 (N_492,N_424,N_447);
and U493 (N_493,N_402,N_423);
and U494 (N_494,N_434,N_435);
nor U495 (N_495,N_442,N_426);
or U496 (N_496,N_432,N_411);
and U497 (N_497,N_448,N_423);
and U498 (N_498,N_406,N_418);
nor U499 (N_499,N_403,N_447);
nor U500 (N_500,N_458,N_479);
or U501 (N_501,N_464,N_468);
nor U502 (N_502,N_471,N_470);
nand U503 (N_503,N_491,N_486);
xor U504 (N_504,N_480,N_466);
xor U505 (N_505,N_460,N_498);
or U506 (N_506,N_481,N_459);
nand U507 (N_507,N_482,N_495);
nand U508 (N_508,N_472,N_451);
nor U509 (N_509,N_496,N_478);
or U510 (N_510,N_483,N_477);
nand U511 (N_511,N_493,N_499);
and U512 (N_512,N_474,N_497);
nor U513 (N_513,N_475,N_490);
nand U514 (N_514,N_456,N_467);
nor U515 (N_515,N_488,N_453);
nor U516 (N_516,N_454,N_457);
or U517 (N_517,N_487,N_476);
nor U518 (N_518,N_462,N_485);
nand U519 (N_519,N_461,N_450);
nand U520 (N_520,N_452,N_465);
nand U521 (N_521,N_455,N_494);
nand U522 (N_522,N_473,N_463);
nand U523 (N_523,N_492,N_469);
xnor U524 (N_524,N_484,N_489);
or U525 (N_525,N_476,N_470);
and U526 (N_526,N_477,N_467);
and U527 (N_527,N_493,N_483);
nor U528 (N_528,N_454,N_494);
nand U529 (N_529,N_461,N_465);
and U530 (N_530,N_452,N_478);
or U531 (N_531,N_478,N_477);
or U532 (N_532,N_494,N_468);
xnor U533 (N_533,N_473,N_494);
and U534 (N_534,N_485,N_452);
or U535 (N_535,N_456,N_485);
nand U536 (N_536,N_482,N_475);
or U537 (N_537,N_481,N_498);
or U538 (N_538,N_471,N_484);
and U539 (N_539,N_473,N_452);
or U540 (N_540,N_455,N_499);
nand U541 (N_541,N_496,N_488);
or U542 (N_542,N_454,N_462);
and U543 (N_543,N_454,N_483);
and U544 (N_544,N_458,N_494);
xor U545 (N_545,N_452,N_486);
xnor U546 (N_546,N_460,N_486);
nand U547 (N_547,N_467,N_468);
nor U548 (N_548,N_463,N_484);
and U549 (N_549,N_466,N_494);
nor U550 (N_550,N_538,N_539);
nand U551 (N_551,N_519,N_537);
nor U552 (N_552,N_507,N_506);
nor U553 (N_553,N_517,N_533);
nand U554 (N_554,N_512,N_530);
or U555 (N_555,N_544,N_548);
nand U556 (N_556,N_503,N_514);
nand U557 (N_557,N_535,N_543);
and U558 (N_558,N_545,N_520);
nor U559 (N_559,N_540,N_504);
nand U560 (N_560,N_529,N_528);
nor U561 (N_561,N_527,N_534);
or U562 (N_562,N_511,N_523);
or U563 (N_563,N_521,N_508);
or U564 (N_564,N_541,N_549);
nand U565 (N_565,N_501,N_546);
and U566 (N_566,N_518,N_515);
nand U567 (N_567,N_525,N_524);
nor U568 (N_568,N_505,N_547);
xor U569 (N_569,N_531,N_500);
nor U570 (N_570,N_542,N_502);
and U571 (N_571,N_509,N_522);
nor U572 (N_572,N_536,N_510);
nand U573 (N_573,N_513,N_532);
nor U574 (N_574,N_516,N_526);
and U575 (N_575,N_510,N_526);
nand U576 (N_576,N_505,N_543);
or U577 (N_577,N_532,N_517);
nor U578 (N_578,N_524,N_541);
or U579 (N_579,N_547,N_533);
and U580 (N_580,N_529,N_549);
nor U581 (N_581,N_538,N_531);
nor U582 (N_582,N_544,N_542);
or U583 (N_583,N_501,N_529);
and U584 (N_584,N_538,N_514);
and U585 (N_585,N_505,N_528);
nor U586 (N_586,N_543,N_531);
and U587 (N_587,N_545,N_519);
or U588 (N_588,N_502,N_543);
and U589 (N_589,N_526,N_532);
or U590 (N_590,N_516,N_510);
and U591 (N_591,N_508,N_548);
nand U592 (N_592,N_501,N_549);
and U593 (N_593,N_524,N_519);
nand U594 (N_594,N_522,N_523);
or U595 (N_595,N_511,N_525);
xnor U596 (N_596,N_517,N_541);
and U597 (N_597,N_508,N_532);
or U598 (N_598,N_521,N_545);
nor U599 (N_599,N_514,N_525);
and U600 (N_600,N_559,N_593);
and U601 (N_601,N_592,N_577);
nand U602 (N_602,N_586,N_572);
nand U603 (N_603,N_558,N_589);
or U604 (N_604,N_575,N_571);
or U605 (N_605,N_560,N_595);
nor U606 (N_606,N_569,N_590);
nor U607 (N_607,N_583,N_563);
nor U608 (N_608,N_556,N_562);
and U609 (N_609,N_578,N_599);
and U610 (N_610,N_585,N_566);
and U611 (N_611,N_553,N_552);
or U612 (N_612,N_580,N_551);
nor U613 (N_613,N_565,N_588);
or U614 (N_614,N_557,N_597);
xnor U615 (N_615,N_594,N_576);
or U616 (N_616,N_582,N_554);
nor U617 (N_617,N_567,N_570);
nand U618 (N_618,N_555,N_596);
nand U619 (N_619,N_573,N_598);
and U620 (N_620,N_561,N_581);
nand U621 (N_621,N_591,N_564);
xnor U622 (N_622,N_550,N_568);
or U623 (N_623,N_579,N_584);
nor U624 (N_624,N_587,N_574);
or U625 (N_625,N_588,N_579);
and U626 (N_626,N_594,N_554);
nor U627 (N_627,N_588,N_555);
or U628 (N_628,N_558,N_560);
nor U629 (N_629,N_575,N_583);
and U630 (N_630,N_567,N_588);
nand U631 (N_631,N_576,N_570);
xor U632 (N_632,N_586,N_574);
and U633 (N_633,N_561,N_593);
or U634 (N_634,N_599,N_584);
or U635 (N_635,N_562,N_596);
xnor U636 (N_636,N_594,N_553);
and U637 (N_637,N_594,N_552);
or U638 (N_638,N_591,N_550);
or U639 (N_639,N_578,N_577);
nor U640 (N_640,N_571,N_556);
nand U641 (N_641,N_551,N_572);
nor U642 (N_642,N_587,N_585);
or U643 (N_643,N_564,N_595);
and U644 (N_644,N_556,N_552);
nor U645 (N_645,N_554,N_584);
or U646 (N_646,N_550,N_554);
nor U647 (N_647,N_578,N_560);
nor U648 (N_648,N_590,N_574);
and U649 (N_649,N_564,N_590);
nor U650 (N_650,N_606,N_631);
nand U651 (N_651,N_620,N_637);
and U652 (N_652,N_626,N_628);
or U653 (N_653,N_649,N_627);
nand U654 (N_654,N_608,N_630);
and U655 (N_655,N_621,N_618);
or U656 (N_656,N_646,N_616);
nor U657 (N_657,N_601,N_633);
xor U658 (N_658,N_613,N_619);
nor U659 (N_659,N_625,N_648);
or U660 (N_660,N_639,N_614);
and U661 (N_661,N_605,N_617);
and U662 (N_662,N_632,N_634);
and U663 (N_663,N_623,N_629);
or U664 (N_664,N_647,N_641);
nand U665 (N_665,N_640,N_622);
nand U666 (N_666,N_600,N_642);
nor U667 (N_667,N_611,N_644);
or U668 (N_668,N_615,N_602);
and U669 (N_669,N_607,N_645);
or U670 (N_670,N_604,N_638);
nor U671 (N_671,N_610,N_624);
nand U672 (N_672,N_635,N_643);
and U673 (N_673,N_609,N_603);
or U674 (N_674,N_612,N_636);
nor U675 (N_675,N_610,N_611);
nor U676 (N_676,N_607,N_646);
nand U677 (N_677,N_626,N_621);
or U678 (N_678,N_640,N_633);
nor U679 (N_679,N_639,N_627);
and U680 (N_680,N_620,N_607);
nand U681 (N_681,N_610,N_612);
nor U682 (N_682,N_606,N_644);
and U683 (N_683,N_646,N_640);
nor U684 (N_684,N_606,N_605);
and U685 (N_685,N_622,N_635);
or U686 (N_686,N_615,N_647);
or U687 (N_687,N_611,N_605);
nand U688 (N_688,N_609,N_607);
nand U689 (N_689,N_637,N_608);
nand U690 (N_690,N_608,N_627);
and U691 (N_691,N_632,N_644);
or U692 (N_692,N_619,N_640);
xnor U693 (N_693,N_611,N_600);
or U694 (N_694,N_628,N_644);
nor U695 (N_695,N_623,N_611);
or U696 (N_696,N_608,N_648);
nor U697 (N_697,N_644,N_605);
and U698 (N_698,N_628,N_636);
and U699 (N_699,N_607,N_611);
and U700 (N_700,N_669,N_661);
or U701 (N_701,N_681,N_699);
or U702 (N_702,N_693,N_655);
nor U703 (N_703,N_676,N_663);
nor U704 (N_704,N_660,N_684);
nor U705 (N_705,N_657,N_694);
and U706 (N_706,N_685,N_674);
or U707 (N_707,N_651,N_679);
nor U708 (N_708,N_698,N_672);
nor U709 (N_709,N_652,N_659);
nor U710 (N_710,N_687,N_690);
nand U711 (N_711,N_691,N_678);
xor U712 (N_712,N_664,N_665);
or U713 (N_713,N_667,N_697);
and U714 (N_714,N_668,N_666);
xnor U715 (N_715,N_654,N_695);
nand U716 (N_716,N_673,N_682);
nor U717 (N_717,N_677,N_653);
and U718 (N_718,N_656,N_686);
nor U719 (N_719,N_671,N_688);
xor U720 (N_720,N_658,N_680);
and U721 (N_721,N_675,N_683);
and U722 (N_722,N_696,N_670);
and U723 (N_723,N_662,N_650);
nand U724 (N_724,N_689,N_692);
or U725 (N_725,N_699,N_696);
and U726 (N_726,N_671,N_677);
nand U727 (N_727,N_678,N_658);
or U728 (N_728,N_693,N_654);
nor U729 (N_729,N_660,N_680);
nand U730 (N_730,N_657,N_651);
nor U731 (N_731,N_664,N_660);
and U732 (N_732,N_689,N_686);
and U733 (N_733,N_686,N_672);
or U734 (N_734,N_672,N_688);
nor U735 (N_735,N_689,N_676);
nor U736 (N_736,N_677,N_686);
nor U737 (N_737,N_689,N_661);
nand U738 (N_738,N_653,N_671);
nand U739 (N_739,N_651,N_696);
or U740 (N_740,N_684,N_661);
xor U741 (N_741,N_670,N_656);
nand U742 (N_742,N_670,N_685);
and U743 (N_743,N_675,N_668);
nand U744 (N_744,N_691,N_669);
and U745 (N_745,N_663,N_680);
and U746 (N_746,N_698,N_691);
nor U747 (N_747,N_682,N_652);
or U748 (N_748,N_661,N_691);
xnor U749 (N_749,N_677,N_689);
and U750 (N_750,N_711,N_707);
and U751 (N_751,N_736,N_720);
nor U752 (N_752,N_738,N_705);
nor U753 (N_753,N_748,N_722);
nand U754 (N_754,N_746,N_749);
or U755 (N_755,N_721,N_702);
xnor U756 (N_756,N_709,N_713);
and U757 (N_757,N_739,N_718);
nand U758 (N_758,N_723,N_747);
xnor U759 (N_759,N_715,N_714);
and U760 (N_760,N_712,N_732);
or U761 (N_761,N_725,N_704);
nand U762 (N_762,N_734,N_700);
nor U763 (N_763,N_728,N_741);
and U764 (N_764,N_735,N_719);
nor U765 (N_765,N_710,N_701);
nand U766 (N_766,N_730,N_745);
xor U767 (N_767,N_729,N_717);
nor U768 (N_768,N_708,N_740);
nand U769 (N_769,N_716,N_706);
or U770 (N_770,N_724,N_743);
nor U771 (N_771,N_742,N_731);
xnor U772 (N_772,N_733,N_726);
and U773 (N_773,N_744,N_703);
and U774 (N_774,N_727,N_737);
nand U775 (N_775,N_731,N_741);
xor U776 (N_776,N_707,N_739);
or U777 (N_777,N_729,N_705);
and U778 (N_778,N_732,N_739);
and U779 (N_779,N_745,N_733);
nor U780 (N_780,N_735,N_710);
and U781 (N_781,N_740,N_736);
xnor U782 (N_782,N_724,N_706);
and U783 (N_783,N_730,N_709);
xor U784 (N_784,N_703,N_714);
or U785 (N_785,N_743,N_715);
xor U786 (N_786,N_720,N_704);
nor U787 (N_787,N_709,N_735);
nand U788 (N_788,N_729,N_745);
nand U789 (N_789,N_714,N_749);
and U790 (N_790,N_736,N_725);
or U791 (N_791,N_715,N_748);
nand U792 (N_792,N_723,N_719);
nor U793 (N_793,N_738,N_743);
or U794 (N_794,N_737,N_725);
or U795 (N_795,N_741,N_729);
nor U796 (N_796,N_719,N_727);
nand U797 (N_797,N_742,N_734);
or U798 (N_798,N_739,N_709);
or U799 (N_799,N_738,N_747);
and U800 (N_800,N_791,N_797);
and U801 (N_801,N_760,N_789);
and U802 (N_802,N_781,N_763);
and U803 (N_803,N_771,N_778);
nor U804 (N_804,N_774,N_792);
and U805 (N_805,N_756,N_768);
and U806 (N_806,N_793,N_762);
and U807 (N_807,N_782,N_780);
and U808 (N_808,N_798,N_767);
nor U809 (N_809,N_758,N_775);
or U810 (N_810,N_772,N_752);
nand U811 (N_811,N_794,N_786);
nand U812 (N_812,N_785,N_764);
or U813 (N_813,N_754,N_769);
nor U814 (N_814,N_759,N_787);
nand U815 (N_815,N_765,N_799);
and U816 (N_816,N_796,N_776);
xnor U817 (N_817,N_753,N_766);
nor U818 (N_818,N_757,N_783);
nor U819 (N_819,N_761,N_750);
or U820 (N_820,N_755,N_784);
or U821 (N_821,N_777,N_788);
nand U822 (N_822,N_795,N_779);
and U823 (N_823,N_773,N_770);
nand U824 (N_824,N_751,N_790);
nor U825 (N_825,N_760,N_777);
nor U826 (N_826,N_773,N_762);
nand U827 (N_827,N_774,N_757);
nand U828 (N_828,N_771,N_775);
nand U829 (N_829,N_777,N_783);
and U830 (N_830,N_787,N_760);
and U831 (N_831,N_766,N_797);
and U832 (N_832,N_771,N_790);
or U833 (N_833,N_776,N_767);
nand U834 (N_834,N_771,N_780);
or U835 (N_835,N_786,N_760);
or U836 (N_836,N_778,N_767);
nand U837 (N_837,N_788,N_750);
nand U838 (N_838,N_779,N_753);
nor U839 (N_839,N_771,N_756);
or U840 (N_840,N_770,N_754);
or U841 (N_841,N_793,N_785);
nand U842 (N_842,N_771,N_769);
nor U843 (N_843,N_770,N_783);
nor U844 (N_844,N_788,N_799);
and U845 (N_845,N_751,N_771);
nand U846 (N_846,N_754,N_773);
or U847 (N_847,N_784,N_752);
nor U848 (N_848,N_788,N_794);
and U849 (N_849,N_797,N_798);
or U850 (N_850,N_801,N_826);
and U851 (N_851,N_838,N_837);
xor U852 (N_852,N_827,N_824);
and U853 (N_853,N_807,N_828);
nor U854 (N_854,N_823,N_829);
nand U855 (N_855,N_817,N_839);
or U856 (N_856,N_813,N_805);
or U857 (N_857,N_814,N_822);
or U858 (N_858,N_804,N_845);
nand U859 (N_859,N_815,N_806);
and U860 (N_860,N_848,N_809);
or U861 (N_861,N_846,N_843);
and U862 (N_862,N_832,N_803);
nand U863 (N_863,N_842,N_844);
nor U864 (N_864,N_800,N_825);
or U865 (N_865,N_831,N_811);
nor U866 (N_866,N_816,N_810);
nand U867 (N_867,N_802,N_835);
nand U868 (N_868,N_836,N_820);
and U869 (N_869,N_841,N_833);
nor U870 (N_870,N_834,N_840);
nor U871 (N_871,N_812,N_830);
nand U872 (N_872,N_821,N_808);
nand U873 (N_873,N_847,N_819);
xor U874 (N_874,N_818,N_849);
nor U875 (N_875,N_823,N_819);
nor U876 (N_876,N_808,N_818);
xor U877 (N_877,N_808,N_840);
or U878 (N_878,N_818,N_830);
and U879 (N_879,N_838,N_826);
and U880 (N_880,N_814,N_842);
xor U881 (N_881,N_814,N_801);
nand U882 (N_882,N_828,N_801);
nor U883 (N_883,N_821,N_812);
nor U884 (N_884,N_811,N_835);
nand U885 (N_885,N_832,N_848);
nor U886 (N_886,N_832,N_833);
nor U887 (N_887,N_802,N_816);
nand U888 (N_888,N_816,N_835);
and U889 (N_889,N_834,N_819);
and U890 (N_890,N_810,N_842);
nand U891 (N_891,N_820,N_814);
and U892 (N_892,N_829,N_831);
nor U893 (N_893,N_820,N_804);
nor U894 (N_894,N_841,N_815);
nand U895 (N_895,N_839,N_849);
nor U896 (N_896,N_827,N_804);
and U897 (N_897,N_821,N_841);
and U898 (N_898,N_827,N_819);
nor U899 (N_899,N_833,N_806);
nand U900 (N_900,N_894,N_850);
nor U901 (N_901,N_886,N_860);
or U902 (N_902,N_898,N_881);
or U903 (N_903,N_895,N_896);
and U904 (N_904,N_883,N_852);
xnor U905 (N_905,N_851,N_877);
xor U906 (N_906,N_884,N_855);
xor U907 (N_907,N_859,N_878);
and U908 (N_908,N_888,N_861);
or U909 (N_909,N_863,N_876);
nor U910 (N_910,N_899,N_870);
and U911 (N_911,N_866,N_897);
nand U912 (N_912,N_873,N_875);
and U913 (N_913,N_893,N_889);
or U914 (N_914,N_856,N_853);
and U915 (N_915,N_868,N_857);
and U916 (N_916,N_872,N_880);
or U917 (N_917,N_882,N_862);
nand U918 (N_918,N_879,N_874);
or U919 (N_919,N_891,N_865);
and U920 (N_920,N_867,N_864);
nand U921 (N_921,N_892,N_869);
or U922 (N_922,N_890,N_887);
xnor U923 (N_923,N_858,N_871);
nor U924 (N_924,N_885,N_854);
nor U925 (N_925,N_862,N_854);
and U926 (N_926,N_895,N_857);
xor U927 (N_927,N_886,N_883);
nand U928 (N_928,N_875,N_877);
xor U929 (N_929,N_876,N_869);
and U930 (N_930,N_874,N_851);
or U931 (N_931,N_863,N_895);
nand U932 (N_932,N_885,N_890);
or U933 (N_933,N_874,N_875);
and U934 (N_934,N_858,N_885);
nand U935 (N_935,N_862,N_850);
and U936 (N_936,N_873,N_895);
or U937 (N_937,N_868,N_862);
and U938 (N_938,N_890,N_881);
or U939 (N_939,N_877,N_873);
or U940 (N_940,N_852,N_892);
or U941 (N_941,N_884,N_886);
nand U942 (N_942,N_871,N_888);
or U943 (N_943,N_878,N_857);
nand U944 (N_944,N_860,N_892);
or U945 (N_945,N_850,N_879);
or U946 (N_946,N_883,N_870);
nor U947 (N_947,N_850,N_868);
or U948 (N_948,N_896,N_874);
and U949 (N_949,N_867,N_862);
xnor U950 (N_950,N_918,N_933);
and U951 (N_951,N_907,N_920);
and U952 (N_952,N_927,N_931);
or U953 (N_953,N_929,N_905);
xor U954 (N_954,N_928,N_934);
nand U955 (N_955,N_921,N_943);
and U956 (N_956,N_935,N_902);
xnor U957 (N_957,N_930,N_914);
and U958 (N_958,N_946,N_919);
and U959 (N_959,N_942,N_911);
nand U960 (N_960,N_910,N_913);
or U961 (N_961,N_909,N_925);
or U962 (N_962,N_947,N_903);
nor U963 (N_963,N_923,N_949);
nand U964 (N_964,N_924,N_936);
and U965 (N_965,N_900,N_906);
nand U966 (N_966,N_932,N_915);
nor U967 (N_967,N_940,N_948);
xnor U968 (N_968,N_939,N_926);
nand U969 (N_969,N_916,N_912);
nand U970 (N_970,N_938,N_937);
nand U971 (N_971,N_904,N_944);
and U972 (N_972,N_922,N_917);
nand U973 (N_973,N_941,N_901);
and U974 (N_974,N_908,N_945);
or U975 (N_975,N_941,N_907);
nor U976 (N_976,N_920,N_904);
and U977 (N_977,N_910,N_908);
nor U978 (N_978,N_940,N_906);
and U979 (N_979,N_912,N_918);
nor U980 (N_980,N_935,N_930);
or U981 (N_981,N_943,N_947);
nand U982 (N_982,N_937,N_905);
or U983 (N_983,N_922,N_930);
and U984 (N_984,N_941,N_942);
and U985 (N_985,N_921,N_936);
or U986 (N_986,N_931,N_917);
nand U987 (N_987,N_939,N_913);
xor U988 (N_988,N_949,N_934);
or U989 (N_989,N_937,N_948);
or U990 (N_990,N_936,N_925);
nand U991 (N_991,N_938,N_900);
nand U992 (N_992,N_902,N_900);
nor U993 (N_993,N_905,N_926);
and U994 (N_994,N_928,N_916);
and U995 (N_995,N_913,N_908);
nor U996 (N_996,N_922,N_910);
or U997 (N_997,N_918,N_900);
xnor U998 (N_998,N_947,N_937);
or U999 (N_999,N_940,N_926);
and U1000 (N_1000,N_992,N_952);
nand U1001 (N_1001,N_950,N_975);
xor U1002 (N_1002,N_967,N_964);
nor U1003 (N_1003,N_974,N_960);
and U1004 (N_1004,N_983,N_971);
and U1005 (N_1005,N_986,N_985);
and U1006 (N_1006,N_953,N_987);
xor U1007 (N_1007,N_981,N_991);
and U1008 (N_1008,N_968,N_962);
or U1009 (N_1009,N_990,N_956);
or U1010 (N_1010,N_978,N_969);
nand U1011 (N_1011,N_998,N_977);
nand U1012 (N_1012,N_959,N_995);
or U1013 (N_1013,N_993,N_951);
and U1014 (N_1014,N_973,N_989);
nor U1015 (N_1015,N_970,N_994);
nand U1016 (N_1016,N_996,N_988);
and U1017 (N_1017,N_972,N_955);
nor U1018 (N_1018,N_957,N_979);
and U1019 (N_1019,N_958,N_997);
nand U1020 (N_1020,N_965,N_999);
nor U1021 (N_1021,N_954,N_961);
nor U1022 (N_1022,N_982,N_984);
nor U1023 (N_1023,N_980,N_963);
xor U1024 (N_1024,N_976,N_966);
or U1025 (N_1025,N_951,N_988);
or U1026 (N_1026,N_998,N_956);
nor U1027 (N_1027,N_970,N_953);
nand U1028 (N_1028,N_982,N_957);
and U1029 (N_1029,N_985,N_973);
nor U1030 (N_1030,N_952,N_979);
nor U1031 (N_1031,N_972,N_966);
and U1032 (N_1032,N_964,N_984);
and U1033 (N_1033,N_951,N_961);
or U1034 (N_1034,N_990,N_953);
or U1035 (N_1035,N_980,N_957);
nand U1036 (N_1036,N_975,N_978);
and U1037 (N_1037,N_969,N_994);
nand U1038 (N_1038,N_985,N_965);
or U1039 (N_1039,N_984,N_995);
xnor U1040 (N_1040,N_996,N_955);
and U1041 (N_1041,N_955,N_987);
or U1042 (N_1042,N_952,N_999);
or U1043 (N_1043,N_974,N_992);
or U1044 (N_1044,N_980,N_989);
nand U1045 (N_1045,N_952,N_981);
and U1046 (N_1046,N_956,N_977);
or U1047 (N_1047,N_991,N_963);
and U1048 (N_1048,N_979,N_983);
or U1049 (N_1049,N_998,N_972);
and U1050 (N_1050,N_1000,N_1044);
nand U1051 (N_1051,N_1036,N_1012);
or U1052 (N_1052,N_1040,N_1004);
or U1053 (N_1053,N_1023,N_1041);
nor U1054 (N_1054,N_1031,N_1049);
and U1055 (N_1055,N_1028,N_1003);
nor U1056 (N_1056,N_1019,N_1045);
nand U1057 (N_1057,N_1038,N_1037);
xnor U1058 (N_1058,N_1009,N_1013);
or U1059 (N_1059,N_1001,N_1008);
and U1060 (N_1060,N_1007,N_1042);
nor U1061 (N_1061,N_1005,N_1018);
nand U1062 (N_1062,N_1043,N_1046);
or U1063 (N_1063,N_1039,N_1035);
nand U1064 (N_1064,N_1006,N_1021);
and U1065 (N_1065,N_1016,N_1027);
nor U1066 (N_1066,N_1017,N_1011);
xnor U1067 (N_1067,N_1047,N_1002);
nand U1068 (N_1068,N_1026,N_1032);
nor U1069 (N_1069,N_1029,N_1015);
nor U1070 (N_1070,N_1030,N_1010);
and U1071 (N_1071,N_1025,N_1020);
nand U1072 (N_1072,N_1014,N_1048);
and U1073 (N_1073,N_1022,N_1034);
or U1074 (N_1074,N_1024,N_1033);
nor U1075 (N_1075,N_1017,N_1046);
or U1076 (N_1076,N_1002,N_1012);
and U1077 (N_1077,N_1027,N_1046);
nor U1078 (N_1078,N_1009,N_1005);
or U1079 (N_1079,N_1038,N_1012);
xnor U1080 (N_1080,N_1021,N_1036);
or U1081 (N_1081,N_1011,N_1039);
xnor U1082 (N_1082,N_1010,N_1024);
nor U1083 (N_1083,N_1042,N_1022);
or U1084 (N_1084,N_1013,N_1001);
nand U1085 (N_1085,N_1025,N_1007);
nand U1086 (N_1086,N_1005,N_1004);
or U1087 (N_1087,N_1013,N_1039);
or U1088 (N_1088,N_1038,N_1047);
nor U1089 (N_1089,N_1040,N_1049);
xor U1090 (N_1090,N_1028,N_1031);
xor U1091 (N_1091,N_1013,N_1003);
nand U1092 (N_1092,N_1046,N_1040);
or U1093 (N_1093,N_1013,N_1035);
nor U1094 (N_1094,N_1015,N_1002);
nand U1095 (N_1095,N_1007,N_1048);
and U1096 (N_1096,N_1035,N_1029);
and U1097 (N_1097,N_1001,N_1023);
or U1098 (N_1098,N_1034,N_1019);
or U1099 (N_1099,N_1036,N_1010);
or U1100 (N_1100,N_1059,N_1073);
xnor U1101 (N_1101,N_1061,N_1052);
nor U1102 (N_1102,N_1093,N_1055);
and U1103 (N_1103,N_1057,N_1051);
and U1104 (N_1104,N_1097,N_1077);
nand U1105 (N_1105,N_1079,N_1054);
or U1106 (N_1106,N_1083,N_1070);
or U1107 (N_1107,N_1060,N_1056);
nor U1108 (N_1108,N_1076,N_1089);
nor U1109 (N_1109,N_1072,N_1088);
nand U1110 (N_1110,N_1094,N_1071);
xnor U1111 (N_1111,N_1080,N_1087);
nand U1112 (N_1112,N_1062,N_1074);
nor U1113 (N_1113,N_1082,N_1075);
and U1114 (N_1114,N_1078,N_1066);
xor U1115 (N_1115,N_1069,N_1096);
xnor U1116 (N_1116,N_1084,N_1063);
and U1117 (N_1117,N_1090,N_1098);
nand U1118 (N_1118,N_1091,N_1065);
nand U1119 (N_1119,N_1058,N_1068);
nor U1120 (N_1120,N_1085,N_1067);
nor U1121 (N_1121,N_1050,N_1095);
or U1122 (N_1122,N_1092,N_1081);
nor U1123 (N_1123,N_1064,N_1086);
nand U1124 (N_1124,N_1053,N_1099);
or U1125 (N_1125,N_1063,N_1099);
and U1126 (N_1126,N_1095,N_1058);
or U1127 (N_1127,N_1093,N_1089);
or U1128 (N_1128,N_1058,N_1051);
or U1129 (N_1129,N_1088,N_1087);
or U1130 (N_1130,N_1090,N_1061);
nand U1131 (N_1131,N_1096,N_1055);
nand U1132 (N_1132,N_1074,N_1087);
or U1133 (N_1133,N_1055,N_1078);
or U1134 (N_1134,N_1052,N_1094);
or U1135 (N_1135,N_1093,N_1094);
and U1136 (N_1136,N_1096,N_1087);
nand U1137 (N_1137,N_1058,N_1085);
xor U1138 (N_1138,N_1085,N_1066);
and U1139 (N_1139,N_1059,N_1064);
nand U1140 (N_1140,N_1076,N_1068);
nand U1141 (N_1141,N_1079,N_1056);
nand U1142 (N_1142,N_1089,N_1060);
or U1143 (N_1143,N_1089,N_1068);
nand U1144 (N_1144,N_1057,N_1063);
nor U1145 (N_1145,N_1095,N_1083);
nor U1146 (N_1146,N_1086,N_1070);
nor U1147 (N_1147,N_1060,N_1082);
nor U1148 (N_1148,N_1056,N_1064);
nor U1149 (N_1149,N_1064,N_1097);
or U1150 (N_1150,N_1101,N_1108);
and U1151 (N_1151,N_1146,N_1134);
or U1152 (N_1152,N_1148,N_1114);
nor U1153 (N_1153,N_1144,N_1135);
or U1154 (N_1154,N_1126,N_1131);
nand U1155 (N_1155,N_1102,N_1145);
or U1156 (N_1156,N_1133,N_1137);
and U1157 (N_1157,N_1119,N_1136);
and U1158 (N_1158,N_1129,N_1141);
or U1159 (N_1159,N_1112,N_1113);
nor U1160 (N_1160,N_1123,N_1128);
nor U1161 (N_1161,N_1149,N_1140);
or U1162 (N_1162,N_1103,N_1116);
nor U1163 (N_1163,N_1117,N_1143);
nand U1164 (N_1164,N_1132,N_1121);
or U1165 (N_1165,N_1138,N_1122);
and U1166 (N_1166,N_1124,N_1104);
and U1167 (N_1167,N_1105,N_1139);
nand U1168 (N_1168,N_1106,N_1142);
nand U1169 (N_1169,N_1109,N_1111);
nor U1170 (N_1170,N_1110,N_1127);
nand U1171 (N_1171,N_1147,N_1100);
or U1172 (N_1172,N_1125,N_1107);
nand U1173 (N_1173,N_1118,N_1120);
or U1174 (N_1174,N_1115,N_1130);
and U1175 (N_1175,N_1112,N_1117);
nand U1176 (N_1176,N_1130,N_1125);
or U1177 (N_1177,N_1122,N_1119);
and U1178 (N_1178,N_1116,N_1140);
nor U1179 (N_1179,N_1116,N_1121);
nand U1180 (N_1180,N_1108,N_1100);
nor U1181 (N_1181,N_1144,N_1116);
nor U1182 (N_1182,N_1112,N_1125);
nor U1183 (N_1183,N_1122,N_1133);
nand U1184 (N_1184,N_1120,N_1127);
nand U1185 (N_1185,N_1119,N_1127);
nand U1186 (N_1186,N_1143,N_1129);
and U1187 (N_1187,N_1127,N_1124);
or U1188 (N_1188,N_1107,N_1100);
xnor U1189 (N_1189,N_1110,N_1141);
nand U1190 (N_1190,N_1103,N_1140);
and U1191 (N_1191,N_1114,N_1102);
nor U1192 (N_1192,N_1123,N_1140);
and U1193 (N_1193,N_1113,N_1110);
nor U1194 (N_1194,N_1123,N_1110);
or U1195 (N_1195,N_1124,N_1130);
nand U1196 (N_1196,N_1123,N_1101);
nor U1197 (N_1197,N_1147,N_1116);
nor U1198 (N_1198,N_1123,N_1117);
nand U1199 (N_1199,N_1139,N_1100);
and U1200 (N_1200,N_1158,N_1170);
and U1201 (N_1201,N_1167,N_1197);
xnor U1202 (N_1202,N_1166,N_1150);
and U1203 (N_1203,N_1172,N_1193);
nand U1204 (N_1204,N_1176,N_1174);
or U1205 (N_1205,N_1179,N_1175);
and U1206 (N_1206,N_1195,N_1192);
nor U1207 (N_1207,N_1168,N_1151);
nor U1208 (N_1208,N_1190,N_1191);
nor U1209 (N_1209,N_1162,N_1194);
nor U1210 (N_1210,N_1159,N_1154);
and U1211 (N_1211,N_1164,N_1182);
or U1212 (N_1212,N_1185,N_1178);
nor U1213 (N_1213,N_1163,N_1152);
or U1214 (N_1214,N_1161,N_1180);
nand U1215 (N_1215,N_1169,N_1153);
or U1216 (N_1216,N_1181,N_1177);
nand U1217 (N_1217,N_1157,N_1199);
nor U1218 (N_1218,N_1160,N_1183);
nand U1219 (N_1219,N_1184,N_1187);
nor U1220 (N_1220,N_1171,N_1165);
nor U1221 (N_1221,N_1155,N_1188);
nand U1222 (N_1222,N_1156,N_1198);
nand U1223 (N_1223,N_1196,N_1189);
nor U1224 (N_1224,N_1186,N_1173);
nand U1225 (N_1225,N_1162,N_1180);
xor U1226 (N_1226,N_1170,N_1180);
nor U1227 (N_1227,N_1153,N_1174);
nand U1228 (N_1228,N_1167,N_1174);
nor U1229 (N_1229,N_1171,N_1186);
nor U1230 (N_1230,N_1160,N_1177);
nor U1231 (N_1231,N_1184,N_1173);
xnor U1232 (N_1232,N_1155,N_1193);
xor U1233 (N_1233,N_1181,N_1196);
or U1234 (N_1234,N_1166,N_1188);
nand U1235 (N_1235,N_1162,N_1182);
and U1236 (N_1236,N_1174,N_1194);
and U1237 (N_1237,N_1152,N_1187);
nand U1238 (N_1238,N_1181,N_1186);
nand U1239 (N_1239,N_1188,N_1169);
or U1240 (N_1240,N_1165,N_1198);
nor U1241 (N_1241,N_1158,N_1166);
nand U1242 (N_1242,N_1174,N_1164);
xor U1243 (N_1243,N_1196,N_1182);
or U1244 (N_1244,N_1192,N_1170);
or U1245 (N_1245,N_1199,N_1189);
nand U1246 (N_1246,N_1150,N_1176);
or U1247 (N_1247,N_1194,N_1175);
and U1248 (N_1248,N_1192,N_1185);
nor U1249 (N_1249,N_1169,N_1162);
nor U1250 (N_1250,N_1231,N_1210);
or U1251 (N_1251,N_1200,N_1213);
nand U1252 (N_1252,N_1237,N_1220);
nor U1253 (N_1253,N_1214,N_1216);
nor U1254 (N_1254,N_1206,N_1208);
nor U1255 (N_1255,N_1228,N_1221);
nor U1256 (N_1256,N_1204,N_1247);
or U1257 (N_1257,N_1203,N_1242);
nor U1258 (N_1258,N_1209,N_1211);
or U1259 (N_1259,N_1219,N_1223);
nor U1260 (N_1260,N_1245,N_1218);
nand U1261 (N_1261,N_1226,N_1246);
nor U1262 (N_1262,N_1236,N_1234);
nor U1263 (N_1263,N_1233,N_1225);
nand U1264 (N_1264,N_1224,N_1230);
xor U1265 (N_1265,N_1202,N_1235);
nor U1266 (N_1266,N_1207,N_1238);
or U1267 (N_1267,N_1222,N_1229);
xnor U1268 (N_1268,N_1239,N_1232);
and U1269 (N_1269,N_1212,N_1227);
and U1270 (N_1270,N_1201,N_1241);
and U1271 (N_1271,N_1217,N_1244);
nor U1272 (N_1272,N_1215,N_1243);
or U1273 (N_1273,N_1240,N_1249);
xnor U1274 (N_1274,N_1248,N_1205);
nand U1275 (N_1275,N_1240,N_1202);
nand U1276 (N_1276,N_1233,N_1226);
or U1277 (N_1277,N_1214,N_1248);
nand U1278 (N_1278,N_1238,N_1248);
and U1279 (N_1279,N_1244,N_1230);
nor U1280 (N_1280,N_1219,N_1221);
and U1281 (N_1281,N_1241,N_1211);
or U1282 (N_1282,N_1228,N_1213);
or U1283 (N_1283,N_1215,N_1221);
or U1284 (N_1284,N_1203,N_1238);
xor U1285 (N_1285,N_1228,N_1202);
and U1286 (N_1286,N_1219,N_1227);
and U1287 (N_1287,N_1226,N_1229);
nand U1288 (N_1288,N_1201,N_1230);
or U1289 (N_1289,N_1204,N_1233);
nand U1290 (N_1290,N_1223,N_1211);
nor U1291 (N_1291,N_1235,N_1205);
nor U1292 (N_1292,N_1222,N_1201);
and U1293 (N_1293,N_1240,N_1211);
and U1294 (N_1294,N_1224,N_1212);
nor U1295 (N_1295,N_1243,N_1233);
or U1296 (N_1296,N_1227,N_1244);
nor U1297 (N_1297,N_1227,N_1239);
nand U1298 (N_1298,N_1220,N_1200);
or U1299 (N_1299,N_1224,N_1227);
nor U1300 (N_1300,N_1259,N_1289);
nand U1301 (N_1301,N_1260,N_1280);
and U1302 (N_1302,N_1263,N_1276);
nor U1303 (N_1303,N_1283,N_1251);
or U1304 (N_1304,N_1292,N_1281);
and U1305 (N_1305,N_1253,N_1273);
nor U1306 (N_1306,N_1271,N_1293);
nand U1307 (N_1307,N_1287,N_1255);
xor U1308 (N_1308,N_1256,N_1270);
nand U1309 (N_1309,N_1286,N_1275);
nand U1310 (N_1310,N_1285,N_1272);
or U1311 (N_1311,N_1278,N_1291);
nor U1312 (N_1312,N_1268,N_1269);
and U1313 (N_1313,N_1288,N_1274);
and U1314 (N_1314,N_1284,N_1279);
nand U1315 (N_1315,N_1264,N_1252);
nor U1316 (N_1316,N_1267,N_1250);
xnor U1317 (N_1317,N_1257,N_1277);
and U1318 (N_1318,N_1299,N_1297);
xor U1319 (N_1319,N_1290,N_1262);
or U1320 (N_1320,N_1261,N_1258);
nor U1321 (N_1321,N_1294,N_1295);
nor U1322 (N_1322,N_1298,N_1254);
or U1323 (N_1323,N_1282,N_1296);
and U1324 (N_1324,N_1265,N_1266);
nor U1325 (N_1325,N_1274,N_1287);
and U1326 (N_1326,N_1271,N_1257);
or U1327 (N_1327,N_1282,N_1292);
or U1328 (N_1328,N_1261,N_1287);
nand U1329 (N_1329,N_1253,N_1280);
xnor U1330 (N_1330,N_1270,N_1293);
and U1331 (N_1331,N_1262,N_1276);
nand U1332 (N_1332,N_1267,N_1295);
and U1333 (N_1333,N_1269,N_1292);
nor U1334 (N_1334,N_1275,N_1268);
nor U1335 (N_1335,N_1286,N_1289);
nor U1336 (N_1336,N_1250,N_1253);
nor U1337 (N_1337,N_1282,N_1290);
nand U1338 (N_1338,N_1262,N_1259);
and U1339 (N_1339,N_1278,N_1271);
nor U1340 (N_1340,N_1254,N_1292);
nor U1341 (N_1341,N_1292,N_1276);
nor U1342 (N_1342,N_1252,N_1257);
nor U1343 (N_1343,N_1291,N_1252);
nor U1344 (N_1344,N_1274,N_1265);
or U1345 (N_1345,N_1295,N_1297);
nor U1346 (N_1346,N_1269,N_1263);
nor U1347 (N_1347,N_1263,N_1285);
or U1348 (N_1348,N_1286,N_1298);
and U1349 (N_1349,N_1283,N_1286);
nand U1350 (N_1350,N_1346,N_1324);
nor U1351 (N_1351,N_1322,N_1335);
nand U1352 (N_1352,N_1311,N_1314);
nand U1353 (N_1353,N_1337,N_1349);
and U1354 (N_1354,N_1339,N_1325);
nor U1355 (N_1355,N_1342,N_1301);
nor U1356 (N_1356,N_1345,N_1315);
nor U1357 (N_1357,N_1309,N_1319);
and U1358 (N_1358,N_1327,N_1340);
nor U1359 (N_1359,N_1333,N_1308);
and U1360 (N_1360,N_1347,N_1348);
nand U1361 (N_1361,N_1338,N_1321);
and U1362 (N_1362,N_1331,N_1336);
or U1363 (N_1363,N_1332,N_1329);
nand U1364 (N_1364,N_1302,N_1330);
or U1365 (N_1365,N_1320,N_1343);
nand U1366 (N_1366,N_1317,N_1307);
and U1367 (N_1367,N_1316,N_1300);
nand U1368 (N_1368,N_1334,N_1323);
and U1369 (N_1369,N_1318,N_1304);
nor U1370 (N_1370,N_1328,N_1306);
xor U1371 (N_1371,N_1326,N_1305);
and U1372 (N_1372,N_1303,N_1313);
and U1373 (N_1373,N_1312,N_1344);
and U1374 (N_1374,N_1310,N_1341);
xor U1375 (N_1375,N_1310,N_1312);
xnor U1376 (N_1376,N_1343,N_1331);
nand U1377 (N_1377,N_1316,N_1330);
nor U1378 (N_1378,N_1318,N_1320);
nor U1379 (N_1379,N_1336,N_1335);
nor U1380 (N_1380,N_1309,N_1320);
nand U1381 (N_1381,N_1315,N_1314);
nand U1382 (N_1382,N_1315,N_1301);
xor U1383 (N_1383,N_1302,N_1320);
nand U1384 (N_1384,N_1346,N_1314);
nand U1385 (N_1385,N_1308,N_1339);
nand U1386 (N_1386,N_1323,N_1313);
nor U1387 (N_1387,N_1335,N_1345);
and U1388 (N_1388,N_1309,N_1321);
or U1389 (N_1389,N_1339,N_1344);
or U1390 (N_1390,N_1346,N_1341);
nor U1391 (N_1391,N_1317,N_1308);
and U1392 (N_1392,N_1347,N_1323);
or U1393 (N_1393,N_1305,N_1328);
or U1394 (N_1394,N_1343,N_1313);
xnor U1395 (N_1395,N_1336,N_1312);
and U1396 (N_1396,N_1306,N_1329);
nor U1397 (N_1397,N_1312,N_1315);
nor U1398 (N_1398,N_1323,N_1318);
or U1399 (N_1399,N_1330,N_1339);
or U1400 (N_1400,N_1359,N_1365);
or U1401 (N_1401,N_1391,N_1350);
or U1402 (N_1402,N_1361,N_1363);
nor U1403 (N_1403,N_1370,N_1383);
nand U1404 (N_1404,N_1373,N_1382);
nor U1405 (N_1405,N_1351,N_1394);
nand U1406 (N_1406,N_1385,N_1355);
or U1407 (N_1407,N_1377,N_1367);
or U1408 (N_1408,N_1390,N_1386);
or U1409 (N_1409,N_1371,N_1399);
nor U1410 (N_1410,N_1398,N_1360);
xnor U1411 (N_1411,N_1378,N_1396);
nand U1412 (N_1412,N_1380,N_1364);
or U1413 (N_1413,N_1381,N_1379);
nand U1414 (N_1414,N_1356,N_1354);
nand U1415 (N_1415,N_1352,N_1353);
nor U1416 (N_1416,N_1395,N_1393);
nor U1417 (N_1417,N_1375,N_1376);
or U1418 (N_1418,N_1358,N_1374);
nor U1419 (N_1419,N_1389,N_1366);
xnor U1420 (N_1420,N_1387,N_1372);
and U1421 (N_1421,N_1388,N_1357);
nand U1422 (N_1422,N_1362,N_1369);
nand U1423 (N_1423,N_1368,N_1384);
or U1424 (N_1424,N_1397,N_1392);
and U1425 (N_1425,N_1352,N_1364);
or U1426 (N_1426,N_1380,N_1391);
or U1427 (N_1427,N_1388,N_1363);
nand U1428 (N_1428,N_1380,N_1360);
nor U1429 (N_1429,N_1375,N_1383);
or U1430 (N_1430,N_1395,N_1373);
nor U1431 (N_1431,N_1368,N_1396);
nor U1432 (N_1432,N_1365,N_1357);
or U1433 (N_1433,N_1364,N_1358);
nor U1434 (N_1434,N_1369,N_1398);
or U1435 (N_1435,N_1362,N_1352);
xor U1436 (N_1436,N_1388,N_1390);
or U1437 (N_1437,N_1381,N_1352);
and U1438 (N_1438,N_1392,N_1389);
nand U1439 (N_1439,N_1362,N_1394);
or U1440 (N_1440,N_1389,N_1379);
or U1441 (N_1441,N_1376,N_1356);
or U1442 (N_1442,N_1370,N_1354);
xnor U1443 (N_1443,N_1389,N_1359);
nor U1444 (N_1444,N_1363,N_1379);
or U1445 (N_1445,N_1397,N_1360);
nor U1446 (N_1446,N_1360,N_1370);
and U1447 (N_1447,N_1385,N_1373);
nor U1448 (N_1448,N_1354,N_1394);
nor U1449 (N_1449,N_1384,N_1398);
nor U1450 (N_1450,N_1408,N_1449);
xor U1451 (N_1451,N_1402,N_1421);
xor U1452 (N_1452,N_1424,N_1413);
or U1453 (N_1453,N_1405,N_1414);
nor U1454 (N_1454,N_1422,N_1420);
nor U1455 (N_1455,N_1443,N_1415);
or U1456 (N_1456,N_1432,N_1423);
nand U1457 (N_1457,N_1403,N_1430);
nand U1458 (N_1458,N_1437,N_1431);
or U1459 (N_1459,N_1436,N_1406);
and U1460 (N_1460,N_1448,N_1411);
nor U1461 (N_1461,N_1433,N_1438);
nand U1462 (N_1462,N_1447,N_1410);
nand U1463 (N_1463,N_1435,N_1446);
nor U1464 (N_1464,N_1441,N_1425);
or U1465 (N_1465,N_1434,N_1428);
nand U1466 (N_1466,N_1439,N_1440);
nand U1467 (N_1467,N_1444,N_1427);
nor U1468 (N_1468,N_1426,N_1417);
and U1469 (N_1469,N_1419,N_1442);
xor U1470 (N_1470,N_1418,N_1404);
nand U1471 (N_1471,N_1407,N_1416);
xor U1472 (N_1472,N_1429,N_1412);
or U1473 (N_1473,N_1409,N_1445);
nand U1474 (N_1474,N_1400,N_1401);
nand U1475 (N_1475,N_1425,N_1413);
and U1476 (N_1476,N_1445,N_1438);
xnor U1477 (N_1477,N_1421,N_1436);
and U1478 (N_1478,N_1446,N_1424);
and U1479 (N_1479,N_1438,N_1403);
or U1480 (N_1480,N_1434,N_1449);
nor U1481 (N_1481,N_1426,N_1428);
xnor U1482 (N_1482,N_1400,N_1434);
nand U1483 (N_1483,N_1435,N_1428);
nor U1484 (N_1484,N_1441,N_1413);
nand U1485 (N_1485,N_1447,N_1406);
and U1486 (N_1486,N_1423,N_1427);
nand U1487 (N_1487,N_1415,N_1448);
nand U1488 (N_1488,N_1405,N_1435);
nand U1489 (N_1489,N_1448,N_1445);
and U1490 (N_1490,N_1443,N_1442);
nand U1491 (N_1491,N_1412,N_1404);
and U1492 (N_1492,N_1416,N_1438);
nor U1493 (N_1493,N_1420,N_1406);
or U1494 (N_1494,N_1448,N_1431);
nor U1495 (N_1495,N_1422,N_1417);
nor U1496 (N_1496,N_1414,N_1440);
nand U1497 (N_1497,N_1403,N_1426);
and U1498 (N_1498,N_1400,N_1420);
nor U1499 (N_1499,N_1448,N_1425);
and U1500 (N_1500,N_1477,N_1470);
or U1501 (N_1501,N_1494,N_1491);
nor U1502 (N_1502,N_1453,N_1481);
nand U1503 (N_1503,N_1460,N_1451);
or U1504 (N_1504,N_1457,N_1468);
and U1505 (N_1505,N_1450,N_1472);
nor U1506 (N_1506,N_1492,N_1493);
or U1507 (N_1507,N_1496,N_1464);
nor U1508 (N_1508,N_1465,N_1498);
nand U1509 (N_1509,N_1476,N_1467);
nand U1510 (N_1510,N_1483,N_1466);
and U1511 (N_1511,N_1462,N_1454);
and U1512 (N_1512,N_1490,N_1480);
nand U1513 (N_1513,N_1473,N_1452);
xnor U1514 (N_1514,N_1456,N_1463);
and U1515 (N_1515,N_1459,N_1461);
and U1516 (N_1516,N_1479,N_1486);
or U1517 (N_1517,N_1474,N_1499);
nor U1518 (N_1518,N_1469,N_1485);
or U1519 (N_1519,N_1471,N_1487);
and U1520 (N_1520,N_1495,N_1455);
xor U1521 (N_1521,N_1475,N_1458);
and U1522 (N_1522,N_1489,N_1488);
nor U1523 (N_1523,N_1478,N_1497);
nor U1524 (N_1524,N_1482,N_1484);
or U1525 (N_1525,N_1463,N_1476);
or U1526 (N_1526,N_1453,N_1491);
nand U1527 (N_1527,N_1496,N_1473);
nor U1528 (N_1528,N_1482,N_1475);
and U1529 (N_1529,N_1483,N_1456);
nor U1530 (N_1530,N_1460,N_1489);
or U1531 (N_1531,N_1452,N_1477);
nor U1532 (N_1532,N_1465,N_1452);
nand U1533 (N_1533,N_1471,N_1472);
nor U1534 (N_1534,N_1470,N_1475);
nand U1535 (N_1535,N_1464,N_1495);
xor U1536 (N_1536,N_1470,N_1493);
xor U1537 (N_1537,N_1462,N_1468);
or U1538 (N_1538,N_1487,N_1473);
nor U1539 (N_1539,N_1454,N_1483);
nand U1540 (N_1540,N_1484,N_1469);
and U1541 (N_1541,N_1485,N_1487);
nand U1542 (N_1542,N_1475,N_1465);
nand U1543 (N_1543,N_1450,N_1470);
and U1544 (N_1544,N_1497,N_1452);
nand U1545 (N_1545,N_1499,N_1460);
nor U1546 (N_1546,N_1479,N_1497);
or U1547 (N_1547,N_1450,N_1499);
nor U1548 (N_1548,N_1499,N_1472);
nor U1549 (N_1549,N_1476,N_1453);
and U1550 (N_1550,N_1542,N_1513);
nand U1551 (N_1551,N_1532,N_1521);
or U1552 (N_1552,N_1509,N_1501);
xor U1553 (N_1553,N_1538,N_1549);
xnor U1554 (N_1554,N_1508,N_1541);
or U1555 (N_1555,N_1547,N_1526);
nand U1556 (N_1556,N_1545,N_1540);
or U1557 (N_1557,N_1528,N_1503);
nand U1558 (N_1558,N_1548,N_1524);
xnor U1559 (N_1559,N_1525,N_1536);
nand U1560 (N_1560,N_1520,N_1515);
nand U1561 (N_1561,N_1533,N_1527);
nor U1562 (N_1562,N_1534,N_1516);
nand U1563 (N_1563,N_1510,N_1504);
nor U1564 (N_1564,N_1530,N_1505);
nor U1565 (N_1565,N_1543,N_1502);
or U1566 (N_1566,N_1519,N_1514);
nor U1567 (N_1567,N_1523,N_1522);
xor U1568 (N_1568,N_1535,N_1544);
and U1569 (N_1569,N_1539,N_1511);
and U1570 (N_1570,N_1529,N_1500);
or U1571 (N_1571,N_1507,N_1517);
and U1572 (N_1572,N_1546,N_1512);
nor U1573 (N_1573,N_1506,N_1531);
xor U1574 (N_1574,N_1518,N_1537);
or U1575 (N_1575,N_1538,N_1525);
xnor U1576 (N_1576,N_1513,N_1503);
nand U1577 (N_1577,N_1522,N_1515);
nand U1578 (N_1578,N_1538,N_1523);
nand U1579 (N_1579,N_1516,N_1502);
nor U1580 (N_1580,N_1502,N_1501);
or U1581 (N_1581,N_1549,N_1547);
xor U1582 (N_1582,N_1523,N_1529);
nor U1583 (N_1583,N_1501,N_1527);
or U1584 (N_1584,N_1517,N_1523);
nand U1585 (N_1585,N_1529,N_1539);
or U1586 (N_1586,N_1543,N_1517);
nand U1587 (N_1587,N_1539,N_1519);
or U1588 (N_1588,N_1534,N_1503);
nand U1589 (N_1589,N_1522,N_1518);
nand U1590 (N_1590,N_1504,N_1503);
nor U1591 (N_1591,N_1523,N_1531);
nand U1592 (N_1592,N_1531,N_1537);
nand U1593 (N_1593,N_1528,N_1516);
nand U1594 (N_1594,N_1517,N_1502);
nor U1595 (N_1595,N_1531,N_1539);
nand U1596 (N_1596,N_1543,N_1526);
and U1597 (N_1597,N_1504,N_1537);
nor U1598 (N_1598,N_1545,N_1510);
nand U1599 (N_1599,N_1517,N_1540);
nor U1600 (N_1600,N_1566,N_1554);
and U1601 (N_1601,N_1560,N_1580);
and U1602 (N_1602,N_1591,N_1590);
nor U1603 (N_1603,N_1567,N_1573);
nand U1604 (N_1604,N_1579,N_1581);
xnor U1605 (N_1605,N_1572,N_1588);
or U1606 (N_1606,N_1582,N_1561);
and U1607 (N_1607,N_1575,N_1576);
nand U1608 (N_1608,N_1583,N_1563);
and U1609 (N_1609,N_1569,N_1562);
and U1610 (N_1610,N_1558,N_1599);
or U1611 (N_1611,N_1586,N_1550);
nor U1612 (N_1612,N_1593,N_1557);
xnor U1613 (N_1613,N_1578,N_1565);
or U1614 (N_1614,N_1559,N_1598);
nor U1615 (N_1615,N_1585,N_1552);
nor U1616 (N_1616,N_1592,N_1596);
nor U1617 (N_1617,N_1589,N_1551);
or U1618 (N_1618,N_1597,N_1577);
and U1619 (N_1619,N_1570,N_1571);
nor U1620 (N_1620,N_1555,N_1574);
or U1621 (N_1621,N_1553,N_1556);
and U1622 (N_1622,N_1595,N_1587);
and U1623 (N_1623,N_1564,N_1594);
or U1624 (N_1624,N_1568,N_1584);
nor U1625 (N_1625,N_1594,N_1598);
and U1626 (N_1626,N_1592,N_1570);
xor U1627 (N_1627,N_1551,N_1558);
and U1628 (N_1628,N_1580,N_1561);
nor U1629 (N_1629,N_1574,N_1567);
and U1630 (N_1630,N_1598,N_1563);
or U1631 (N_1631,N_1571,N_1554);
xor U1632 (N_1632,N_1566,N_1553);
or U1633 (N_1633,N_1568,N_1591);
nand U1634 (N_1634,N_1570,N_1574);
and U1635 (N_1635,N_1572,N_1591);
or U1636 (N_1636,N_1580,N_1595);
nor U1637 (N_1637,N_1596,N_1586);
and U1638 (N_1638,N_1599,N_1568);
nor U1639 (N_1639,N_1589,N_1586);
xnor U1640 (N_1640,N_1573,N_1581);
nand U1641 (N_1641,N_1576,N_1560);
nor U1642 (N_1642,N_1562,N_1588);
or U1643 (N_1643,N_1597,N_1596);
nor U1644 (N_1644,N_1592,N_1580);
nor U1645 (N_1645,N_1577,N_1573);
or U1646 (N_1646,N_1576,N_1591);
nor U1647 (N_1647,N_1593,N_1564);
and U1648 (N_1648,N_1598,N_1573);
xor U1649 (N_1649,N_1557,N_1597);
nand U1650 (N_1650,N_1627,N_1646);
nor U1651 (N_1651,N_1636,N_1610);
and U1652 (N_1652,N_1619,N_1647);
and U1653 (N_1653,N_1640,N_1609);
or U1654 (N_1654,N_1631,N_1614);
or U1655 (N_1655,N_1633,N_1606);
nor U1656 (N_1656,N_1613,N_1634);
or U1657 (N_1657,N_1616,N_1630);
and U1658 (N_1658,N_1611,N_1620);
and U1659 (N_1659,N_1604,N_1608);
or U1660 (N_1660,N_1629,N_1635);
nand U1661 (N_1661,N_1643,N_1645);
nand U1662 (N_1662,N_1621,N_1628);
nand U1663 (N_1663,N_1607,N_1623);
nand U1664 (N_1664,N_1626,N_1632);
or U1665 (N_1665,N_1641,N_1639);
or U1666 (N_1666,N_1644,N_1601);
xnor U1667 (N_1667,N_1602,N_1617);
nor U1668 (N_1668,N_1612,N_1622);
and U1669 (N_1669,N_1618,N_1637);
or U1670 (N_1670,N_1624,N_1625);
xnor U1671 (N_1671,N_1649,N_1648);
and U1672 (N_1672,N_1603,N_1605);
and U1673 (N_1673,N_1638,N_1615);
and U1674 (N_1674,N_1642,N_1600);
and U1675 (N_1675,N_1607,N_1611);
xor U1676 (N_1676,N_1628,N_1607);
or U1677 (N_1677,N_1628,N_1636);
nand U1678 (N_1678,N_1604,N_1606);
nand U1679 (N_1679,N_1632,N_1649);
or U1680 (N_1680,N_1646,N_1621);
and U1681 (N_1681,N_1622,N_1626);
and U1682 (N_1682,N_1645,N_1631);
and U1683 (N_1683,N_1637,N_1620);
nand U1684 (N_1684,N_1628,N_1639);
nand U1685 (N_1685,N_1604,N_1642);
nand U1686 (N_1686,N_1617,N_1634);
nand U1687 (N_1687,N_1602,N_1609);
nand U1688 (N_1688,N_1600,N_1621);
or U1689 (N_1689,N_1617,N_1641);
nand U1690 (N_1690,N_1639,N_1629);
nand U1691 (N_1691,N_1627,N_1603);
or U1692 (N_1692,N_1611,N_1635);
nand U1693 (N_1693,N_1619,N_1608);
nand U1694 (N_1694,N_1621,N_1627);
nor U1695 (N_1695,N_1639,N_1647);
or U1696 (N_1696,N_1600,N_1634);
nor U1697 (N_1697,N_1619,N_1602);
nand U1698 (N_1698,N_1625,N_1616);
nand U1699 (N_1699,N_1617,N_1649);
nand U1700 (N_1700,N_1657,N_1673);
nand U1701 (N_1701,N_1699,N_1693);
and U1702 (N_1702,N_1653,N_1690);
and U1703 (N_1703,N_1664,N_1669);
xnor U1704 (N_1704,N_1679,N_1680);
or U1705 (N_1705,N_1691,N_1674);
and U1706 (N_1706,N_1697,N_1666);
nor U1707 (N_1707,N_1668,N_1652);
or U1708 (N_1708,N_1687,N_1692);
nand U1709 (N_1709,N_1658,N_1689);
and U1710 (N_1710,N_1681,N_1671);
xor U1711 (N_1711,N_1660,N_1663);
nor U1712 (N_1712,N_1698,N_1650);
nor U1713 (N_1713,N_1676,N_1686);
nand U1714 (N_1714,N_1675,N_1684);
xnor U1715 (N_1715,N_1670,N_1688);
and U1716 (N_1716,N_1685,N_1694);
or U1717 (N_1717,N_1654,N_1678);
or U1718 (N_1718,N_1682,N_1667);
or U1719 (N_1719,N_1656,N_1683);
nor U1720 (N_1720,N_1659,N_1672);
nand U1721 (N_1721,N_1655,N_1665);
nor U1722 (N_1722,N_1695,N_1661);
or U1723 (N_1723,N_1696,N_1651);
nand U1724 (N_1724,N_1662,N_1677);
and U1725 (N_1725,N_1694,N_1690);
or U1726 (N_1726,N_1689,N_1656);
and U1727 (N_1727,N_1696,N_1683);
and U1728 (N_1728,N_1695,N_1699);
nand U1729 (N_1729,N_1678,N_1692);
nand U1730 (N_1730,N_1677,N_1665);
nor U1731 (N_1731,N_1686,N_1655);
and U1732 (N_1732,N_1697,N_1680);
nand U1733 (N_1733,N_1674,N_1653);
xor U1734 (N_1734,N_1679,N_1663);
or U1735 (N_1735,N_1663,N_1682);
xnor U1736 (N_1736,N_1674,N_1654);
nor U1737 (N_1737,N_1675,N_1654);
nand U1738 (N_1738,N_1665,N_1667);
xor U1739 (N_1739,N_1697,N_1691);
and U1740 (N_1740,N_1651,N_1695);
and U1741 (N_1741,N_1662,N_1696);
xor U1742 (N_1742,N_1661,N_1669);
or U1743 (N_1743,N_1677,N_1690);
or U1744 (N_1744,N_1697,N_1674);
nor U1745 (N_1745,N_1652,N_1669);
and U1746 (N_1746,N_1690,N_1669);
and U1747 (N_1747,N_1658,N_1681);
or U1748 (N_1748,N_1678,N_1682);
nor U1749 (N_1749,N_1693,N_1688);
xor U1750 (N_1750,N_1705,N_1745);
and U1751 (N_1751,N_1719,N_1744);
or U1752 (N_1752,N_1747,N_1704);
xor U1753 (N_1753,N_1712,N_1721);
and U1754 (N_1754,N_1739,N_1713);
nor U1755 (N_1755,N_1735,N_1722);
or U1756 (N_1756,N_1715,N_1740);
nand U1757 (N_1757,N_1720,N_1724);
and U1758 (N_1758,N_1732,N_1706);
or U1759 (N_1759,N_1727,N_1726);
and U1760 (N_1760,N_1738,N_1718);
nand U1761 (N_1761,N_1702,N_1734);
nor U1762 (N_1762,N_1742,N_1749);
and U1763 (N_1763,N_1736,N_1717);
and U1764 (N_1764,N_1730,N_1743);
and U1765 (N_1765,N_1707,N_1737);
and U1766 (N_1766,N_1714,N_1700);
and U1767 (N_1767,N_1733,N_1748);
or U1768 (N_1768,N_1741,N_1708);
and U1769 (N_1769,N_1728,N_1701);
nor U1770 (N_1770,N_1731,N_1716);
and U1771 (N_1771,N_1725,N_1711);
or U1772 (N_1772,N_1710,N_1729);
xor U1773 (N_1773,N_1709,N_1703);
or U1774 (N_1774,N_1746,N_1723);
nor U1775 (N_1775,N_1740,N_1741);
and U1776 (N_1776,N_1738,N_1709);
and U1777 (N_1777,N_1741,N_1710);
xnor U1778 (N_1778,N_1710,N_1723);
or U1779 (N_1779,N_1718,N_1740);
nor U1780 (N_1780,N_1717,N_1738);
or U1781 (N_1781,N_1735,N_1704);
nand U1782 (N_1782,N_1729,N_1706);
nand U1783 (N_1783,N_1711,N_1747);
and U1784 (N_1784,N_1713,N_1746);
xor U1785 (N_1785,N_1708,N_1701);
nor U1786 (N_1786,N_1731,N_1744);
nor U1787 (N_1787,N_1719,N_1741);
and U1788 (N_1788,N_1738,N_1740);
or U1789 (N_1789,N_1717,N_1703);
nor U1790 (N_1790,N_1710,N_1717);
nor U1791 (N_1791,N_1742,N_1714);
and U1792 (N_1792,N_1720,N_1725);
and U1793 (N_1793,N_1711,N_1744);
xor U1794 (N_1794,N_1746,N_1743);
nand U1795 (N_1795,N_1700,N_1724);
or U1796 (N_1796,N_1747,N_1717);
or U1797 (N_1797,N_1728,N_1743);
nor U1798 (N_1798,N_1739,N_1735);
nand U1799 (N_1799,N_1723,N_1729);
and U1800 (N_1800,N_1759,N_1765);
nor U1801 (N_1801,N_1751,N_1761);
xnor U1802 (N_1802,N_1769,N_1758);
and U1803 (N_1803,N_1754,N_1787);
nand U1804 (N_1804,N_1762,N_1779);
and U1805 (N_1805,N_1768,N_1777);
nor U1806 (N_1806,N_1753,N_1797);
or U1807 (N_1807,N_1792,N_1752);
or U1808 (N_1808,N_1794,N_1788);
nor U1809 (N_1809,N_1774,N_1763);
or U1810 (N_1810,N_1795,N_1781);
and U1811 (N_1811,N_1785,N_1796);
nand U1812 (N_1812,N_1783,N_1772);
and U1813 (N_1813,N_1789,N_1764);
xor U1814 (N_1814,N_1793,N_1750);
nand U1815 (N_1815,N_1798,N_1757);
nor U1816 (N_1816,N_1767,N_1775);
and U1817 (N_1817,N_1799,N_1755);
and U1818 (N_1818,N_1766,N_1778);
or U1819 (N_1819,N_1780,N_1784);
nand U1820 (N_1820,N_1760,N_1773);
nand U1821 (N_1821,N_1771,N_1791);
nor U1822 (N_1822,N_1770,N_1756);
nand U1823 (N_1823,N_1776,N_1790);
nand U1824 (N_1824,N_1786,N_1782);
nor U1825 (N_1825,N_1763,N_1766);
or U1826 (N_1826,N_1754,N_1795);
or U1827 (N_1827,N_1796,N_1778);
xnor U1828 (N_1828,N_1783,N_1796);
and U1829 (N_1829,N_1760,N_1798);
nor U1830 (N_1830,N_1761,N_1769);
or U1831 (N_1831,N_1761,N_1770);
and U1832 (N_1832,N_1759,N_1774);
and U1833 (N_1833,N_1783,N_1795);
and U1834 (N_1834,N_1753,N_1776);
nand U1835 (N_1835,N_1794,N_1795);
nand U1836 (N_1836,N_1780,N_1770);
nand U1837 (N_1837,N_1785,N_1754);
nor U1838 (N_1838,N_1787,N_1790);
or U1839 (N_1839,N_1790,N_1767);
or U1840 (N_1840,N_1775,N_1784);
or U1841 (N_1841,N_1755,N_1786);
or U1842 (N_1842,N_1787,N_1782);
nand U1843 (N_1843,N_1799,N_1788);
or U1844 (N_1844,N_1769,N_1797);
nor U1845 (N_1845,N_1759,N_1794);
xor U1846 (N_1846,N_1784,N_1755);
nor U1847 (N_1847,N_1759,N_1755);
xnor U1848 (N_1848,N_1771,N_1763);
or U1849 (N_1849,N_1788,N_1766);
and U1850 (N_1850,N_1809,N_1844);
nand U1851 (N_1851,N_1814,N_1837);
and U1852 (N_1852,N_1813,N_1817);
xor U1853 (N_1853,N_1802,N_1832);
nor U1854 (N_1854,N_1831,N_1821);
and U1855 (N_1855,N_1845,N_1807);
and U1856 (N_1856,N_1824,N_1825);
nor U1857 (N_1857,N_1808,N_1841);
and U1858 (N_1858,N_1826,N_1833);
or U1859 (N_1859,N_1812,N_1849);
nand U1860 (N_1860,N_1847,N_1838);
xnor U1861 (N_1861,N_1835,N_1818);
nand U1862 (N_1862,N_1840,N_1804);
or U1863 (N_1863,N_1806,N_1842);
and U1864 (N_1864,N_1811,N_1800);
or U1865 (N_1865,N_1822,N_1815);
nor U1866 (N_1866,N_1819,N_1830);
xor U1867 (N_1867,N_1846,N_1848);
or U1868 (N_1868,N_1836,N_1843);
or U1869 (N_1869,N_1839,N_1823);
xnor U1870 (N_1870,N_1805,N_1827);
and U1871 (N_1871,N_1816,N_1829);
nand U1872 (N_1872,N_1803,N_1828);
xor U1873 (N_1873,N_1834,N_1801);
nand U1874 (N_1874,N_1810,N_1820);
nor U1875 (N_1875,N_1813,N_1843);
nor U1876 (N_1876,N_1808,N_1807);
and U1877 (N_1877,N_1808,N_1843);
or U1878 (N_1878,N_1810,N_1812);
nor U1879 (N_1879,N_1823,N_1849);
or U1880 (N_1880,N_1807,N_1818);
nand U1881 (N_1881,N_1803,N_1809);
nor U1882 (N_1882,N_1815,N_1824);
nor U1883 (N_1883,N_1802,N_1834);
and U1884 (N_1884,N_1838,N_1830);
nand U1885 (N_1885,N_1822,N_1826);
or U1886 (N_1886,N_1836,N_1818);
or U1887 (N_1887,N_1826,N_1800);
xor U1888 (N_1888,N_1835,N_1844);
or U1889 (N_1889,N_1843,N_1816);
xor U1890 (N_1890,N_1835,N_1829);
nand U1891 (N_1891,N_1836,N_1819);
nor U1892 (N_1892,N_1837,N_1817);
or U1893 (N_1893,N_1836,N_1814);
or U1894 (N_1894,N_1828,N_1811);
xor U1895 (N_1895,N_1814,N_1845);
and U1896 (N_1896,N_1834,N_1848);
nor U1897 (N_1897,N_1827,N_1821);
nand U1898 (N_1898,N_1821,N_1834);
nor U1899 (N_1899,N_1813,N_1812);
nor U1900 (N_1900,N_1891,N_1854);
or U1901 (N_1901,N_1894,N_1874);
nor U1902 (N_1902,N_1888,N_1859);
nand U1903 (N_1903,N_1872,N_1850);
and U1904 (N_1904,N_1879,N_1892);
or U1905 (N_1905,N_1885,N_1878);
and U1906 (N_1906,N_1883,N_1898);
and U1907 (N_1907,N_1896,N_1856);
nand U1908 (N_1908,N_1866,N_1857);
nor U1909 (N_1909,N_1870,N_1876);
nand U1910 (N_1910,N_1877,N_1873);
and U1911 (N_1911,N_1890,N_1893);
nor U1912 (N_1912,N_1886,N_1862);
nor U1913 (N_1913,N_1882,N_1875);
and U1914 (N_1914,N_1895,N_1861);
or U1915 (N_1915,N_1851,N_1865);
nor U1916 (N_1916,N_1852,N_1863);
xnor U1917 (N_1917,N_1881,N_1887);
or U1918 (N_1918,N_1867,N_1860);
nor U1919 (N_1919,N_1864,N_1899);
or U1920 (N_1920,N_1897,N_1884);
nand U1921 (N_1921,N_1858,N_1853);
and U1922 (N_1922,N_1869,N_1880);
nor U1923 (N_1923,N_1868,N_1855);
xor U1924 (N_1924,N_1889,N_1871);
xor U1925 (N_1925,N_1866,N_1859);
nand U1926 (N_1926,N_1860,N_1896);
nand U1927 (N_1927,N_1873,N_1854);
xor U1928 (N_1928,N_1881,N_1884);
and U1929 (N_1929,N_1867,N_1895);
or U1930 (N_1930,N_1866,N_1871);
or U1931 (N_1931,N_1876,N_1869);
nor U1932 (N_1932,N_1851,N_1858);
or U1933 (N_1933,N_1867,N_1881);
or U1934 (N_1934,N_1888,N_1854);
nand U1935 (N_1935,N_1856,N_1887);
and U1936 (N_1936,N_1859,N_1872);
nand U1937 (N_1937,N_1854,N_1876);
nand U1938 (N_1938,N_1894,N_1886);
nor U1939 (N_1939,N_1870,N_1873);
and U1940 (N_1940,N_1853,N_1893);
nand U1941 (N_1941,N_1882,N_1857);
or U1942 (N_1942,N_1898,N_1884);
nor U1943 (N_1943,N_1875,N_1860);
nand U1944 (N_1944,N_1875,N_1872);
nor U1945 (N_1945,N_1899,N_1878);
and U1946 (N_1946,N_1856,N_1874);
nor U1947 (N_1947,N_1881,N_1888);
and U1948 (N_1948,N_1869,N_1867);
nand U1949 (N_1949,N_1885,N_1899);
and U1950 (N_1950,N_1939,N_1928);
nor U1951 (N_1951,N_1937,N_1948);
or U1952 (N_1952,N_1903,N_1940);
nor U1953 (N_1953,N_1925,N_1936);
and U1954 (N_1954,N_1929,N_1949);
or U1955 (N_1955,N_1917,N_1941);
and U1956 (N_1956,N_1918,N_1911);
nor U1957 (N_1957,N_1942,N_1902);
nor U1958 (N_1958,N_1913,N_1904);
and U1959 (N_1959,N_1923,N_1931);
xor U1960 (N_1960,N_1915,N_1921);
nor U1961 (N_1961,N_1910,N_1926);
or U1962 (N_1962,N_1900,N_1907);
nand U1963 (N_1963,N_1909,N_1934);
xor U1964 (N_1964,N_1922,N_1944);
nor U1965 (N_1965,N_1927,N_1908);
nand U1966 (N_1966,N_1920,N_1938);
and U1967 (N_1967,N_1905,N_1933);
nand U1968 (N_1968,N_1924,N_1912);
or U1969 (N_1969,N_1914,N_1947);
nand U1970 (N_1970,N_1901,N_1946);
nand U1971 (N_1971,N_1916,N_1919);
nor U1972 (N_1972,N_1906,N_1935);
and U1973 (N_1973,N_1932,N_1930);
or U1974 (N_1974,N_1943,N_1945);
nand U1975 (N_1975,N_1934,N_1921);
xnor U1976 (N_1976,N_1928,N_1906);
xor U1977 (N_1977,N_1932,N_1915);
and U1978 (N_1978,N_1908,N_1913);
nand U1979 (N_1979,N_1920,N_1944);
nor U1980 (N_1980,N_1901,N_1935);
nor U1981 (N_1981,N_1928,N_1934);
nand U1982 (N_1982,N_1932,N_1947);
nand U1983 (N_1983,N_1908,N_1924);
xnor U1984 (N_1984,N_1924,N_1929);
nand U1985 (N_1985,N_1944,N_1913);
nor U1986 (N_1986,N_1917,N_1915);
and U1987 (N_1987,N_1940,N_1915);
and U1988 (N_1988,N_1943,N_1924);
xor U1989 (N_1989,N_1908,N_1925);
or U1990 (N_1990,N_1917,N_1948);
or U1991 (N_1991,N_1941,N_1945);
or U1992 (N_1992,N_1902,N_1900);
nor U1993 (N_1993,N_1911,N_1939);
nor U1994 (N_1994,N_1927,N_1912);
nand U1995 (N_1995,N_1943,N_1935);
nand U1996 (N_1996,N_1923,N_1917);
nand U1997 (N_1997,N_1939,N_1902);
xor U1998 (N_1998,N_1915,N_1926);
and U1999 (N_1999,N_1919,N_1905);
nand U2000 (N_2000,N_1957,N_1978);
nand U2001 (N_2001,N_1966,N_1996);
nor U2002 (N_2002,N_1988,N_1963);
and U2003 (N_2003,N_1953,N_1961);
nor U2004 (N_2004,N_1955,N_1975);
and U2005 (N_2005,N_1981,N_1999);
nor U2006 (N_2006,N_1979,N_1984);
or U2007 (N_2007,N_1980,N_1990);
nand U2008 (N_2008,N_1985,N_1967);
nand U2009 (N_2009,N_1962,N_1974);
nor U2010 (N_2010,N_1993,N_1994);
or U2011 (N_2011,N_1965,N_1951);
nor U2012 (N_2012,N_1973,N_1956);
nand U2013 (N_2013,N_1998,N_1960);
nor U2014 (N_2014,N_1986,N_1952);
nand U2015 (N_2015,N_1982,N_1995);
nor U2016 (N_2016,N_1977,N_1954);
nor U2017 (N_2017,N_1950,N_1991);
nor U2018 (N_2018,N_1970,N_1969);
or U2019 (N_2019,N_1987,N_1976);
or U2020 (N_2020,N_1983,N_1972);
or U2021 (N_2021,N_1958,N_1997);
and U2022 (N_2022,N_1992,N_1989);
or U2023 (N_2023,N_1971,N_1959);
nor U2024 (N_2024,N_1964,N_1968);
nor U2025 (N_2025,N_1977,N_1980);
xor U2026 (N_2026,N_1952,N_1970);
and U2027 (N_2027,N_1966,N_1953);
nor U2028 (N_2028,N_1996,N_1964);
and U2029 (N_2029,N_1968,N_1996);
or U2030 (N_2030,N_1981,N_1976);
or U2031 (N_2031,N_1993,N_1972);
or U2032 (N_2032,N_1957,N_1994);
or U2033 (N_2033,N_1978,N_1998);
and U2034 (N_2034,N_1979,N_1972);
and U2035 (N_2035,N_1978,N_1996);
nand U2036 (N_2036,N_1985,N_1990);
nand U2037 (N_2037,N_1977,N_1994);
or U2038 (N_2038,N_1972,N_1987);
or U2039 (N_2039,N_1961,N_1968);
nor U2040 (N_2040,N_1964,N_1973);
or U2041 (N_2041,N_1986,N_1987);
nand U2042 (N_2042,N_1960,N_1967);
xnor U2043 (N_2043,N_1959,N_1974);
or U2044 (N_2044,N_1961,N_1954);
nor U2045 (N_2045,N_1958,N_1961);
and U2046 (N_2046,N_1982,N_1955);
nand U2047 (N_2047,N_1984,N_1962);
and U2048 (N_2048,N_1961,N_1988);
nor U2049 (N_2049,N_1995,N_1974);
nor U2050 (N_2050,N_2026,N_2035);
xnor U2051 (N_2051,N_2009,N_2016);
nor U2052 (N_2052,N_2012,N_2030);
nor U2053 (N_2053,N_2046,N_2023);
xor U2054 (N_2054,N_2040,N_2025);
nor U2055 (N_2055,N_2029,N_2011);
or U2056 (N_2056,N_2001,N_2047);
nand U2057 (N_2057,N_2015,N_2013);
or U2058 (N_2058,N_2049,N_2042);
or U2059 (N_2059,N_2036,N_2045);
and U2060 (N_2060,N_2028,N_2043);
and U2061 (N_2061,N_2006,N_2004);
or U2062 (N_2062,N_2031,N_2021);
nand U2063 (N_2063,N_2003,N_2022);
nand U2064 (N_2064,N_2048,N_2000);
and U2065 (N_2065,N_2017,N_2010);
nand U2066 (N_2066,N_2037,N_2018);
nand U2067 (N_2067,N_2038,N_2020);
or U2068 (N_2068,N_2019,N_2032);
xnor U2069 (N_2069,N_2014,N_2033);
or U2070 (N_2070,N_2005,N_2007);
and U2071 (N_2071,N_2002,N_2044);
or U2072 (N_2072,N_2008,N_2041);
and U2073 (N_2073,N_2024,N_2034);
and U2074 (N_2074,N_2027,N_2039);
xor U2075 (N_2075,N_2028,N_2026);
nor U2076 (N_2076,N_2022,N_2043);
nand U2077 (N_2077,N_2026,N_2011);
nor U2078 (N_2078,N_2029,N_2049);
nor U2079 (N_2079,N_2010,N_2012);
nor U2080 (N_2080,N_2002,N_2034);
and U2081 (N_2081,N_2009,N_2040);
nor U2082 (N_2082,N_2017,N_2003);
or U2083 (N_2083,N_2030,N_2048);
nand U2084 (N_2084,N_2049,N_2046);
nor U2085 (N_2085,N_2044,N_2021);
nand U2086 (N_2086,N_2049,N_2013);
nor U2087 (N_2087,N_2041,N_2037);
nand U2088 (N_2088,N_2028,N_2044);
nand U2089 (N_2089,N_2040,N_2010);
xnor U2090 (N_2090,N_2005,N_2011);
and U2091 (N_2091,N_2043,N_2000);
xor U2092 (N_2092,N_2049,N_2005);
and U2093 (N_2093,N_2038,N_2049);
and U2094 (N_2094,N_2023,N_2047);
nand U2095 (N_2095,N_2003,N_2023);
or U2096 (N_2096,N_2014,N_2032);
or U2097 (N_2097,N_2004,N_2020);
nand U2098 (N_2098,N_2039,N_2046);
and U2099 (N_2099,N_2047,N_2041);
and U2100 (N_2100,N_2094,N_2092);
nand U2101 (N_2101,N_2051,N_2093);
or U2102 (N_2102,N_2074,N_2052);
or U2103 (N_2103,N_2055,N_2063);
and U2104 (N_2104,N_2061,N_2058);
nand U2105 (N_2105,N_2067,N_2065);
and U2106 (N_2106,N_2082,N_2070);
or U2107 (N_2107,N_2097,N_2075);
nor U2108 (N_2108,N_2066,N_2096);
and U2109 (N_2109,N_2083,N_2077);
or U2110 (N_2110,N_2091,N_2099);
xor U2111 (N_2111,N_2086,N_2059);
and U2112 (N_2112,N_2087,N_2088);
xnor U2113 (N_2113,N_2085,N_2098);
and U2114 (N_2114,N_2069,N_2050);
and U2115 (N_2115,N_2054,N_2089);
or U2116 (N_2116,N_2084,N_2081);
or U2117 (N_2117,N_2080,N_2073);
xnor U2118 (N_2118,N_2056,N_2060);
and U2119 (N_2119,N_2072,N_2057);
or U2120 (N_2120,N_2076,N_2071);
nand U2121 (N_2121,N_2090,N_2064);
nor U2122 (N_2122,N_2068,N_2062);
xor U2123 (N_2123,N_2079,N_2095);
or U2124 (N_2124,N_2053,N_2078);
nor U2125 (N_2125,N_2060,N_2090);
and U2126 (N_2126,N_2050,N_2067);
or U2127 (N_2127,N_2066,N_2073);
nand U2128 (N_2128,N_2076,N_2059);
or U2129 (N_2129,N_2090,N_2089);
nand U2130 (N_2130,N_2092,N_2085);
nor U2131 (N_2131,N_2063,N_2059);
nand U2132 (N_2132,N_2096,N_2068);
nand U2133 (N_2133,N_2058,N_2066);
and U2134 (N_2134,N_2070,N_2068);
or U2135 (N_2135,N_2098,N_2061);
and U2136 (N_2136,N_2077,N_2074);
or U2137 (N_2137,N_2060,N_2078);
nand U2138 (N_2138,N_2087,N_2074);
nand U2139 (N_2139,N_2055,N_2094);
or U2140 (N_2140,N_2062,N_2064);
nor U2141 (N_2141,N_2089,N_2098);
or U2142 (N_2142,N_2094,N_2089);
nand U2143 (N_2143,N_2082,N_2076);
and U2144 (N_2144,N_2054,N_2063);
nand U2145 (N_2145,N_2065,N_2079);
nor U2146 (N_2146,N_2089,N_2066);
and U2147 (N_2147,N_2072,N_2090);
and U2148 (N_2148,N_2079,N_2091);
and U2149 (N_2149,N_2078,N_2052);
nor U2150 (N_2150,N_2122,N_2116);
or U2151 (N_2151,N_2140,N_2109);
nand U2152 (N_2152,N_2126,N_2139);
and U2153 (N_2153,N_2117,N_2100);
nor U2154 (N_2154,N_2136,N_2135);
or U2155 (N_2155,N_2111,N_2113);
nor U2156 (N_2156,N_2147,N_2106);
nor U2157 (N_2157,N_2123,N_2132);
nor U2158 (N_2158,N_2115,N_2102);
and U2159 (N_2159,N_2138,N_2114);
nor U2160 (N_2160,N_2149,N_2118);
nand U2161 (N_2161,N_2137,N_2131);
nor U2162 (N_2162,N_2112,N_2124);
nor U2163 (N_2163,N_2143,N_2134);
nor U2164 (N_2164,N_2105,N_2141);
nor U2165 (N_2165,N_2129,N_2144);
and U2166 (N_2166,N_2130,N_2148);
or U2167 (N_2167,N_2107,N_2103);
nand U2168 (N_2168,N_2120,N_2128);
and U2169 (N_2169,N_2108,N_2142);
xnor U2170 (N_2170,N_2146,N_2133);
nand U2171 (N_2171,N_2121,N_2127);
xnor U2172 (N_2172,N_2145,N_2119);
or U2173 (N_2173,N_2110,N_2125);
xnor U2174 (N_2174,N_2101,N_2104);
nand U2175 (N_2175,N_2114,N_2143);
nand U2176 (N_2176,N_2149,N_2140);
or U2177 (N_2177,N_2139,N_2142);
and U2178 (N_2178,N_2136,N_2138);
xnor U2179 (N_2179,N_2108,N_2136);
or U2180 (N_2180,N_2100,N_2127);
xnor U2181 (N_2181,N_2130,N_2121);
nor U2182 (N_2182,N_2147,N_2127);
and U2183 (N_2183,N_2139,N_2148);
and U2184 (N_2184,N_2144,N_2113);
nand U2185 (N_2185,N_2131,N_2141);
nor U2186 (N_2186,N_2146,N_2103);
nor U2187 (N_2187,N_2101,N_2116);
nor U2188 (N_2188,N_2129,N_2113);
nand U2189 (N_2189,N_2105,N_2117);
nand U2190 (N_2190,N_2127,N_2148);
nor U2191 (N_2191,N_2109,N_2102);
xnor U2192 (N_2192,N_2116,N_2147);
nand U2193 (N_2193,N_2121,N_2120);
nor U2194 (N_2194,N_2112,N_2118);
nor U2195 (N_2195,N_2105,N_2146);
nor U2196 (N_2196,N_2140,N_2142);
or U2197 (N_2197,N_2141,N_2135);
nand U2198 (N_2198,N_2131,N_2140);
nand U2199 (N_2199,N_2107,N_2118);
nor U2200 (N_2200,N_2182,N_2163);
or U2201 (N_2201,N_2162,N_2160);
nand U2202 (N_2202,N_2188,N_2150);
and U2203 (N_2203,N_2152,N_2154);
nor U2204 (N_2204,N_2186,N_2166);
nor U2205 (N_2205,N_2151,N_2155);
and U2206 (N_2206,N_2176,N_2180);
or U2207 (N_2207,N_2170,N_2183);
nor U2208 (N_2208,N_2194,N_2175);
nand U2209 (N_2209,N_2187,N_2164);
or U2210 (N_2210,N_2173,N_2185);
or U2211 (N_2211,N_2196,N_2177);
or U2212 (N_2212,N_2197,N_2178);
nor U2213 (N_2213,N_2159,N_2165);
nor U2214 (N_2214,N_2192,N_2168);
nor U2215 (N_2215,N_2184,N_2156);
nand U2216 (N_2216,N_2199,N_2157);
nor U2217 (N_2217,N_2195,N_2161);
or U2218 (N_2218,N_2172,N_2158);
or U2219 (N_2219,N_2167,N_2179);
nand U2220 (N_2220,N_2171,N_2190);
nor U2221 (N_2221,N_2181,N_2198);
xnor U2222 (N_2222,N_2193,N_2169);
nand U2223 (N_2223,N_2153,N_2189);
nand U2224 (N_2224,N_2174,N_2191);
xor U2225 (N_2225,N_2184,N_2192);
nand U2226 (N_2226,N_2186,N_2159);
nor U2227 (N_2227,N_2188,N_2193);
and U2228 (N_2228,N_2163,N_2184);
and U2229 (N_2229,N_2159,N_2197);
or U2230 (N_2230,N_2184,N_2160);
or U2231 (N_2231,N_2166,N_2171);
nand U2232 (N_2232,N_2152,N_2175);
nor U2233 (N_2233,N_2164,N_2157);
or U2234 (N_2234,N_2166,N_2172);
nor U2235 (N_2235,N_2157,N_2172);
nor U2236 (N_2236,N_2197,N_2155);
or U2237 (N_2237,N_2165,N_2186);
or U2238 (N_2238,N_2158,N_2151);
and U2239 (N_2239,N_2186,N_2194);
nor U2240 (N_2240,N_2167,N_2162);
xor U2241 (N_2241,N_2185,N_2150);
nand U2242 (N_2242,N_2188,N_2187);
or U2243 (N_2243,N_2159,N_2177);
nor U2244 (N_2244,N_2158,N_2155);
nor U2245 (N_2245,N_2150,N_2187);
nand U2246 (N_2246,N_2182,N_2194);
nor U2247 (N_2247,N_2189,N_2163);
or U2248 (N_2248,N_2157,N_2196);
and U2249 (N_2249,N_2156,N_2197);
nor U2250 (N_2250,N_2240,N_2218);
nor U2251 (N_2251,N_2245,N_2223);
nor U2252 (N_2252,N_2239,N_2230);
nor U2253 (N_2253,N_2248,N_2211);
or U2254 (N_2254,N_2222,N_2204);
or U2255 (N_2255,N_2241,N_2238);
nor U2256 (N_2256,N_2208,N_2203);
and U2257 (N_2257,N_2214,N_2215);
and U2258 (N_2258,N_2234,N_2201);
and U2259 (N_2259,N_2237,N_2207);
nor U2260 (N_2260,N_2231,N_2206);
xor U2261 (N_2261,N_2226,N_2220);
and U2262 (N_2262,N_2247,N_2243);
or U2263 (N_2263,N_2209,N_2228);
or U2264 (N_2264,N_2219,N_2229);
nor U2265 (N_2265,N_2249,N_2210);
and U2266 (N_2266,N_2205,N_2221);
or U2267 (N_2267,N_2217,N_2236);
nor U2268 (N_2268,N_2246,N_2202);
nor U2269 (N_2269,N_2227,N_2244);
nor U2270 (N_2270,N_2213,N_2225);
or U2271 (N_2271,N_2235,N_2232);
nand U2272 (N_2272,N_2224,N_2212);
and U2273 (N_2273,N_2216,N_2242);
or U2274 (N_2274,N_2233,N_2200);
and U2275 (N_2275,N_2239,N_2240);
or U2276 (N_2276,N_2233,N_2228);
and U2277 (N_2277,N_2233,N_2221);
and U2278 (N_2278,N_2249,N_2215);
or U2279 (N_2279,N_2210,N_2234);
or U2280 (N_2280,N_2231,N_2223);
or U2281 (N_2281,N_2224,N_2240);
xor U2282 (N_2282,N_2214,N_2231);
xor U2283 (N_2283,N_2217,N_2246);
or U2284 (N_2284,N_2226,N_2222);
xor U2285 (N_2285,N_2203,N_2210);
nor U2286 (N_2286,N_2205,N_2218);
or U2287 (N_2287,N_2205,N_2241);
and U2288 (N_2288,N_2203,N_2234);
nand U2289 (N_2289,N_2206,N_2220);
nor U2290 (N_2290,N_2210,N_2213);
or U2291 (N_2291,N_2238,N_2230);
nor U2292 (N_2292,N_2247,N_2249);
nor U2293 (N_2293,N_2230,N_2223);
and U2294 (N_2294,N_2248,N_2237);
or U2295 (N_2295,N_2220,N_2224);
xnor U2296 (N_2296,N_2230,N_2205);
xnor U2297 (N_2297,N_2225,N_2239);
nand U2298 (N_2298,N_2236,N_2212);
or U2299 (N_2299,N_2206,N_2228);
or U2300 (N_2300,N_2260,N_2261);
or U2301 (N_2301,N_2282,N_2268);
and U2302 (N_2302,N_2286,N_2293);
nand U2303 (N_2303,N_2287,N_2256);
or U2304 (N_2304,N_2252,N_2298);
nand U2305 (N_2305,N_2295,N_2264);
nand U2306 (N_2306,N_2284,N_2299);
xnor U2307 (N_2307,N_2270,N_2262);
and U2308 (N_2308,N_2276,N_2250);
nand U2309 (N_2309,N_2257,N_2280);
nand U2310 (N_2310,N_2253,N_2275);
nand U2311 (N_2311,N_2297,N_2283);
nand U2312 (N_2312,N_2266,N_2289);
and U2313 (N_2313,N_2259,N_2294);
or U2314 (N_2314,N_2278,N_2269);
and U2315 (N_2315,N_2271,N_2274);
or U2316 (N_2316,N_2273,N_2255);
nor U2317 (N_2317,N_2263,N_2292);
nor U2318 (N_2318,N_2285,N_2281);
nor U2319 (N_2319,N_2296,N_2267);
nor U2320 (N_2320,N_2265,N_2272);
or U2321 (N_2321,N_2258,N_2290);
nand U2322 (N_2322,N_2291,N_2288);
nor U2323 (N_2323,N_2254,N_2251);
nor U2324 (N_2324,N_2279,N_2277);
nand U2325 (N_2325,N_2258,N_2264);
nor U2326 (N_2326,N_2293,N_2268);
nand U2327 (N_2327,N_2266,N_2250);
or U2328 (N_2328,N_2251,N_2294);
nor U2329 (N_2329,N_2268,N_2279);
nand U2330 (N_2330,N_2282,N_2259);
nor U2331 (N_2331,N_2273,N_2266);
nor U2332 (N_2332,N_2270,N_2287);
nor U2333 (N_2333,N_2251,N_2278);
xor U2334 (N_2334,N_2274,N_2293);
nand U2335 (N_2335,N_2287,N_2299);
or U2336 (N_2336,N_2289,N_2285);
or U2337 (N_2337,N_2252,N_2273);
nand U2338 (N_2338,N_2275,N_2281);
nor U2339 (N_2339,N_2280,N_2250);
and U2340 (N_2340,N_2261,N_2254);
or U2341 (N_2341,N_2295,N_2287);
nor U2342 (N_2342,N_2283,N_2282);
and U2343 (N_2343,N_2281,N_2273);
and U2344 (N_2344,N_2250,N_2265);
nand U2345 (N_2345,N_2279,N_2253);
nand U2346 (N_2346,N_2285,N_2254);
nor U2347 (N_2347,N_2265,N_2252);
xor U2348 (N_2348,N_2251,N_2269);
and U2349 (N_2349,N_2264,N_2257);
nand U2350 (N_2350,N_2313,N_2335);
nor U2351 (N_2351,N_2346,N_2312);
nand U2352 (N_2352,N_2323,N_2334);
nor U2353 (N_2353,N_2318,N_2310);
nand U2354 (N_2354,N_2314,N_2304);
or U2355 (N_2355,N_2326,N_2329);
nor U2356 (N_2356,N_2344,N_2302);
nand U2357 (N_2357,N_2316,N_2336);
and U2358 (N_2358,N_2320,N_2337);
nor U2359 (N_2359,N_2309,N_2348);
nand U2360 (N_2360,N_2324,N_2325);
nand U2361 (N_2361,N_2315,N_2328);
xnor U2362 (N_2362,N_2343,N_2340);
nor U2363 (N_2363,N_2300,N_2341);
xor U2364 (N_2364,N_2322,N_2317);
nand U2365 (N_2365,N_2347,N_2333);
and U2366 (N_2366,N_2306,N_2319);
nand U2367 (N_2367,N_2327,N_2308);
nand U2368 (N_2368,N_2338,N_2307);
nand U2369 (N_2369,N_2321,N_2345);
or U2370 (N_2370,N_2342,N_2301);
nand U2371 (N_2371,N_2332,N_2303);
or U2372 (N_2372,N_2331,N_2311);
nor U2373 (N_2373,N_2330,N_2349);
nor U2374 (N_2374,N_2305,N_2339);
and U2375 (N_2375,N_2323,N_2312);
nand U2376 (N_2376,N_2322,N_2305);
nor U2377 (N_2377,N_2349,N_2329);
nor U2378 (N_2378,N_2316,N_2349);
nor U2379 (N_2379,N_2346,N_2328);
and U2380 (N_2380,N_2340,N_2344);
or U2381 (N_2381,N_2303,N_2335);
nor U2382 (N_2382,N_2319,N_2324);
nor U2383 (N_2383,N_2343,N_2306);
nor U2384 (N_2384,N_2324,N_2333);
xor U2385 (N_2385,N_2319,N_2302);
nor U2386 (N_2386,N_2339,N_2321);
and U2387 (N_2387,N_2337,N_2309);
and U2388 (N_2388,N_2344,N_2333);
nor U2389 (N_2389,N_2301,N_2330);
or U2390 (N_2390,N_2333,N_2310);
nand U2391 (N_2391,N_2308,N_2315);
or U2392 (N_2392,N_2341,N_2302);
or U2393 (N_2393,N_2327,N_2318);
nor U2394 (N_2394,N_2313,N_2315);
nand U2395 (N_2395,N_2329,N_2301);
nor U2396 (N_2396,N_2334,N_2346);
nor U2397 (N_2397,N_2311,N_2307);
nand U2398 (N_2398,N_2316,N_2320);
nand U2399 (N_2399,N_2309,N_2305);
xor U2400 (N_2400,N_2354,N_2364);
and U2401 (N_2401,N_2373,N_2377);
or U2402 (N_2402,N_2357,N_2362);
and U2403 (N_2403,N_2397,N_2351);
or U2404 (N_2404,N_2398,N_2381);
nor U2405 (N_2405,N_2389,N_2352);
and U2406 (N_2406,N_2359,N_2395);
or U2407 (N_2407,N_2366,N_2392);
nand U2408 (N_2408,N_2369,N_2382);
nor U2409 (N_2409,N_2386,N_2380);
nor U2410 (N_2410,N_2383,N_2376);
nor U2411 (N_2411,N_2368,N_2391);
nor U2412 (N_2412,N_2378,N_2393);
xor U2413 (N_2413,N_2387,N_2356);
nor U2414 (N_2414,N_2363,N_2358);
nand U2415 (N_2415,N_2367,N_2360);
and U2416 (N_2416,N_2353,N_2396);
and U2417 (N_2417,N_2394,N_2361);
nor U2418 (N_2418,N_2388,N_2385);
and U2419 (N_2419,N_2371,N_2355);
or U2420 (N_2420,N_2374,N_2350);
or U2421 (N_2421,N_2375,N_2390);
nor U2422 (N_2422,N_2399,N_2379);
nand U2423 (N_2423,N_2370,N_2365);
or U2424 (N_2424,N_2384,N_2372);
nor U2425 (N_2425,N_2355,N_2376);
xor U2426 (N_2426,N_2354,N_2375);
nand U2427 (N_2427,N_2357,N_2358);
and U2428 (N_2428,N_2398,N_2360);
nand U2429 (N_2429,N_2351,N_2390);
nand U2430 (N_2430,N_2375,N_2386);
or U2431 (N_2431,N_2365,N_2357);
nor U2432 (N_2432,N_2353,N_2369);
nor U2433 (N_2433,N_2373,N_2390);
nand U2434 (N_2434,N_2352,N_2364);
nand U2435 (N_2435,N_2374,N_2390);
nor U2436 (N_2436,N_2367,N_2395);
nand U2437 (N_2437,N_2374,N_2382);
or U2438 (N_2438,N_2398,N_2366);
or U2439 (N_2439,N_2361,N_2358);
nand U2440 (N_2440,N_2367,N_2380);
nand U2441 (N_2441,N_2386,N_2378);
nor U2442 (N_2442,N_2379,N_2357);
nand U2443 (N_2443,N_2383,N_2398);
nor U2444 (N_2444,N_2371,N_2374);
or U2445 (N_2445,N_2385,N_2363);
or U2446 (N_2446,N_2358,N_2371);
or U2447 (N_2447,N_2378,N_2376);
and U2448 (N_2448,N_2379,N_2355);
nand U2449 (N_2449,N_2378,N_2355);
nand U2450 (N_2450,N_2417,N_2413);
xor U2451 (N_2451,N_2423,N_2422);
nand U2452 (N_2452,N_2434,N_2438);
nor U2453 (N_2453,N_2446,N_2430);
and U2454 (N_2454,N_2401,N_2443);
or U2455 (N_2455,N_2400,N_2442);
xnor U2456 (N_2456,N_2420,N_2445);
nor U2457 (N_2457,N_2416,N_2402);
and U2458 (N_2458,N_2439,N_2435);
nand U2459 (N_2459,N_2426,N_2441);
xnor U2460 (N_2460,N_2415,N_2428);
nor U2461 (N_2461,N_2421,N_2447);
and U2462 (N_2462,N_2440,N_2444);
xor U2463 (N_2463,N_2425,N_2404);
and U2464 (N_2464,N_2427,N_2414);
nor U2465 (N_2465,N_2405,N_2411);
nor U2466 (N_2466,N_2419,N_2429);
or U2467 (N_2467,N_2410,N_2407);
and U2468 (N_2468,N_2403,N_2432);
and U2469 (N_2469,N_2418,N_2449);
or U2470 (N_2470,N_2412,N_2437);
nor U2471 (N_2471,N_2424,N_2406);
nor U2472 (N_2472,N_2408,N_2436);
nand U2473 (N_2473,N_2431,N_2409);
nor U2474 (N_2474,N_2448,N_2433);
xor U2475 (N_2475,N_2414,N_2403);
xor U2476 (N_2476,N_2427,N_2419);
and U2477 (N_2477,N_2421,N_2429);
or U2478 (N_2478,N_2416,N_2433);
nor U2479 (N_2479,N_2410,N_2414);
or U2480 (N_2480,N_2423,N_2438);
xor U2481 (N_2481,N_2434,N_2422);
and U2482 (N_2482,N_2444,N_2417);
nand U2483 (N_2483,N_2414,N_2436);
nand U2484 (N_2484,N_2402,N_2400);
nand U2485 (N_2485,N_2430,N_2424);
and U2486 (N_2486,N_2425,N_2436);
or U2487 (N_2487,N_2415,N_2432);
nor U2488 (N_2488,N_2410,N_2429);
xor U2489 (N_2489,N_2443,N_2422);
or U2490 (N_2490,N_2407,N_2445);
and U2491 (N_2491,N_2406,N_2416);
or U2492 (N_2492,N_2440,N_2403);
nand U2493 (N_2493,N_2402,N_2441);
and U2494 (N_2494,N_2413,N_2436);
nor U2495 (N_2495,N_2430,N_2426);
nand U2496 (N_2496,N_2429,N_2416);
nand U2497 (N_2497,N_2437,N_2400);
and U2498 (N_2498,N_2444,N_2407);
xor U2499 (N_2499,N_2406,N_2400);
nor U2500 (N_2500,N_2461,N_2481);
nor U2501 (N_2501,N_2484,N_2454);
nor U2502 (N_2502,N_2494,N_2491);
xnor U2503 (N_2503,N_2470,N_2462);
nor U2504 (N_2504,N_2460,N_2450);
and U2505 (N_2505,N_2485,N_2453);
nor U2506 (N_2506,N_2469,N_2490);
or U2507 (N_2507,N_2487,N_2475);
nand U2508 (N_2508,N_2467,N_2473);
nor U2509 (N_2509,N_2489,N_2472);
nand U2510 (N_2510,N_2495,N_2464);
or U2511 (N_2511,N_2480,N_2497);
or U2512 (N_2512,N_2455,N_2478);
nand U2513 (N_2513,N_2477,N_2457);
nand U2514 (N_2514,N_2463,N_2482);
or U2515 (N_2515,N_2488,N_2498);
and U2516 (N_2516,N_2465,N_2466);
nand U2517 (N_2517,N_2474,N_2458);
nand U2518 (N_2518,N_2496,N_2476);
or U2519 (N_2519,N_2483,N_2499);
and U2520 (N_2520,N_2452,N_2451);
and U2521 (N_2521,N_2459,N_2479);
or U2522 (N_2522,N_2468,N_2493);
nand U2523 (N_2523,N_2486,N_2492);
and U2524 (N_2524,N_2471,N_2456);
or U2525 (N_2525,N_2477,N_2468);
nand U2526 (N_2526,N_2485,N_2486);
nor U2527 (N_2527,N_2454,N_2477);
or U2528 (N_2528,N_2487,N_2479);
xor U2529 (N_2529,N_2481,N_2457);
or U2530 (N_2530,N_2472,N_2473);
and U2531 (N_2531,N_2489,N_2488);
or U2532 (N_2532,N_2466,N_2454);
nor U2533 (N_2533,N_2455,N_2490);
nand U2534 (N_2534,N_2456,N_2495);
xnor U2535 (N_2535,N_2497,N_2481);
nor U2536 (N_2536,N_2492,N_2479);
nand U2537 (N_2537,N_2479,N_2455);
and U2538 (N_2538,N_2494,N_2485);
or U2539 (N_2539,N_2457,N_2465);
or U2540 (N_2540,N_2482,N_2452);
nand U2541 (N_2541,N_2454,N_2481);
nand U2542 (N_2542,N_2486,N_2471);
xor U2543 (N_2543,N_2466,N_2470);
nand U2544 (N_2544,N_2466,N_2452);
nand U2545 (N_2545,N_2453,N_2463);
or U2546 (N_2546,N_2470,N_2489);
nor U2547 (N_2547,N_2451,N_2455);
nor U2548 (N_2548,N_2451,N_2478);
xor U2549 (N_2549,N_2468,N_2486);
or U2550 (N_2550,N_2508,N_2542);
nor U2551 (N_2551,N_2543,N_2513);
nand U2552 (N_2552,N_2537,N_2519);
or U2553 (N_2553,N_2527,N_2532);
nor U2554 (N_2554,N_2547,N_2533);
nand U2555 (N_2555,N_2548,N_2515);
or U2556 (N_2556,N_2523,N_2514);
or U2557 (N_2557,N_2506,N_2539);
or U2558 (N_2558,N_2518,N_2510);
xor U2559 (N_2559,N_2531,N_2522);
nand U2560 (N_2560,N_2528,N_2505);
nor U2561 (N_2561,N_2530,N_2520);
or U2562 (N_2562,N_2546,N_2509);
nand U2563 (N_2563,N_2535,N_2524);
xor U2564 (N_2564,N_2500,N_2525);
xor U2565 (N_2565,N_2541,N_2544);
nand U2566 (N_2566,N_2545,N_2512);
xor U2567 (N_2567,N_2503,N_2529);
nor U2568 (N_2568,N_2536,N_2502);
nand U2569 (N_2569,N_2526,N_2516);
and U2570 (N_2570,N_2511,N_2538);
and U2571 (N_2571,N_2507,N_2501);
nor U2572 (N_2572,N_2517,N_2549);
xnor U2573 (N_2573,N_2540,N_2504);
nand U2574 (N_2574,N_2521,N_2534);
and U2575 (N_2575,N_2522,N_2532);
nor U2576 (N_2576,N_2543,N_2504);
and U2577 (N_2577,N_2525,N_2529);
nor U2578 (N_2578,N_2531,N_2541);
or U2579 (N_2579,N_2500,N_2530);
nand U2580 (N_2580,N_2502,N_2503);
nor U2581 (N_2581,N_2535,N_2533);
nor U2582 (N_2582,N_2535,N_2511);
and U2583 (N_2583,N_2538,N_2520);
and U2584 (N_2584,N_2510,N_2512);
nor U2585 (N_2585,N_2536,N_2512);
nor U2586 (N_2586,N_2512,N_2505);
nor U2587 (N_2587,N_2544,N_2503);
nor U2588 (N_2588,N_2511,N_2536);
and U2589 (N_2589,N_2518,N_2521);
xor U2590 (N_2590,N_2526,N_2511);
and U2591 (N_2591,N_2546,N_2527);
nand U2592 (N_2592,N_2503,N_2548);
xnor U2593 (N_2593,N_2522,N_2538);
and U2594 (N_2594,N_2509,N_2504);
nor U2595 (N_2595,N_2511,N_2510);
and U2596 (N_2596,N_2534,N_2532);
and U2597 (N_2597,N_2509,N_2544);
xor U2598 (N_2598,N_2547,N_2542);
or U2599 (N_2599,N_2501,N_2534);
xnor U2600 (N_2600,N_2573,N_2575);
nand U2601 (N_2601,N_2566,N_2559);
xnor U2602 (N_2602,N_2587,N_2585);
nor U2603 (N_2603,N_2577,N_2599);
nand U2604 (N_2604,N_2574,N_2561);
nor U2605 (N_2605,N_2591,N_2563);
nand U2606 (N_2606,N_2576,N_2564);
or U2607 (N_2607,N_2594,N_2592);
and U2608 (N_2608,N_2593,N_2554);
xnor U2609 (N_2609,N_2578,N_2583);
xnor U2610 (N_2610,N_2551,N_2560);
xnor U2611 (N_2611,N_2582,N_2590);
nand U2612 (N_2612,N_2568,N_2584);
nand U2613 (N_2613,N_2555,N_2562);
nand U2614 (N_2614,N_2581,N_2571);
and U2615 (N_2615,N_2589,N_2580);
nand U2616 (N_2616,N_2588,N_2567);
nand U2617 (N_2617,N_2579,N_2570);
or U2618 (N_2618,N_2598,N_2552);
or U2619 (N_2619,N_2572,N_2595);
nor U2620 (N_2620,N_2569,N_2553);
nand U2621 (N_2621,N_2597,N_2556);
nand U2622 (N_2622,N_2586,N_2565);
xor U2623 (N_2623,N_2550,N_2558);
and U2624 (N_2624,N_2557,N_2596);
and U2625 (N_2625,N_2577,N_2579);
nor U2626 (N_2626,N_2571,N_2586);
or U2627 (N_2627,N_2554,N_2551);
or U2628 (N_2628,N_2582,N_2574);
and U2629 (N_2629,N_2553,N_2565);
nor U2630 (N_2630,N_2573,N_2565);
xor U2631 (N_2631,N_2574,N_2585);
and U2632 (N_2632,N_2561,N_2590);
xor U2633 (N_2633,N_2570,N_2580);
and U2634 (N_2634,N_2561,N_2579);
and U2635 (N_2635,N_2579,N_2560);
or U2636 (N_2636,N_2575,N_2567);
and U2637 (N_2637,N_2566,N_2550);
and U2638 (N_2638,N_2552,N_2566);
xor U2639 (N_2639,N_2587,N_2573);
xnor U2640 (N_2640,N_2563,N_2597);
nor U2641 (N_2641,N_2581,N_2597);
and U2642 (N_2642,N_2565,N_2593);
and U2643 (N_2643,N_2580,N_2599);
and U2644 (N_2644,N_2572,N_2565);
or U2645 (N_2645,N_2557,N_2572);
or U2646 (N_2646,N_2550,N_2597);
nand U2647 (N_2647,N_2556,N_2593);
and U2648 (N_2648,N_2595,N_2596);
nor U2649 (N_2649,N_2552,N_2595);
and U2650 (N_2650,N_2605,N_2647);
nor U2651 (N_2651,N_2620,N_2631);
or U2652 (N_2652,N_2626,N_2628);
and U2653 (N_2653,N_2643,N_2609);
nand U2654 (N_2654,N_2627,N_2601);
nand U2655 (N_2655,N_2607,N_2610);
and U2656 (N_2656,N_2639,N_2611);
nand U2657 (N_2657,N_2640,N_2648);
nand U2658 (N_2658,N_2617,N_2613);
and U2659 (N_2659,N_2632,N_2641);
nor U2660 (N_2660,N_2604,N_2634);
and U2661 (N_2661,N_2649,N_2629);
and U2662 (N_2662,N_2614,N_2630);
nor U2663 (N_2663,N_2618,N_2635);
and U2664 (N_2664,N_2642,N_2622);
nand U2665 (N_2665,N_2645,N_2625);
or U2666 (N_2666,N_2637,N_2621);
nand U2667 (N_2667,N_2619,N_2606);
and U2668 (N_2668,N_2636,N_2646);
and U2669 (N_2669,N_2600,N_2602);
nand U2670 (N_2670,N_2612,N_2624);
nand U2671 (N_2671,N_2615,N_2633);
or U2672 (N_2672,N_2608,N_2623);
xor U2673 (N_2673,N_2644,N_2638);
nand U2674 (N_2674,N_2603,N_2616);
nor U2675 (N_2675,N_2636,N_2620);
nand U2676 (N_2676,N_2635,N_2620);
nor U2677 (N_2677,N_2622,N_2608);
nor U2678 (N_2678,N_2629,N_2647);
or U2679 (N_2679,N_2642,N_2624);
nand U2680 (N_2680,N_2620,N_2641);
nor U2681 (N_2681,N_2642,N_2626);
and U2682 (N_2682,N_2607,N_2619);
nand U2683 (N_2683,N_2642,N_2610);
nor U2684 (N_2684,N_2631,N_2649);
xor U2685 (N_2685,N_2622,N_2618);
nor U2686 (N_2686,N_2616,N_2604);
nand U2687 (N_2687,N_2603,N_2621);
nor U2688 (N_2688,N_2606,N_2640);
nor U2689 (N_2689,N_2643,N_2634);
nand U2690 (N_2690,N_2637,N_2606);
and U2691 (N_2691,N_2623,N_2630);
nor U2692 (N_2692,N_2601,N_2649);
or U2693 (N_2693,N_2622,N_2648);
or U2694 (N_2694,N_2648,N_2630);
nor U2695 (N_2695,N_2635,N_2616);
or U2696 (N_2696,N_2619,N_2616);
nor U2697 (N_2697,N_2641,N_2630);
or U2698 (N_2698,N_2621,N_2644);
nor U2699 (N_2699,N_2649,N_2642);
nor U2700 (N_2700,N_2674,N_2673);
nand U2701 (N_2701,N_2651,N_2683);
or U2702 (N_2702,N_2677,N_2672);
nand U2703 (N_2703,N_2685,N_2653);
or U2704 (N_2704,N_2692,N_2675);
nor U2705 (N_2705,N_2662,N_2689);
xnor U2706 (N_2706,N_2658,N_2688);
and U2707 (N_2707,N_2657,N_2699);
nor U2708 (N_2708,N_2678,N_2666);
nand U2709 (N_2709,N_2690,N_2696);
and U2710 (N_2710,N_2667,N_2686);
or U2711 (N_2711,N_2679,N_2695);
nand U2712 (N_2712,N_2684,N_2693);
or U2713 (N_2713,N_2655,N_2691);
or U2714 (N_2714,N_2652,N_2668);
nor U2715 (N_2715,N_2697,N_2664);
or U2716 (N_2716,N_2671,N_2698);
or U2717 (N_2717,N_2682,N_2694);
and U2718 (N_2718,N_2665,N_2681);
and U2719 (N_2719,N_2654,N_2656);
or U2720 (N_2720,N_2659,N_2687);
or U2721 (N_2721,N_2663,N_2660);
or U2722 (N_2722,N_2661,N_2676);
nand U2723 (N_2723,N_2670,N_2669);
nor U2724 (N_2724,N_2680,N_2650);
and U2725 (N_2725,N_2677,N_2695);
and U2726 (N_2726,N_2688,N_2664);
xor U2727 (N_2727,N_2673,N_2664);
and U2728 (N_2728,N_2692,N_2670);
or U2729 (N_2729,N_2673,N_2681);
nand U2730 (N_2730,N_2664,N_2652);
xor U2731 (N_2731,N_2674,N_2672);
or U2732 (N_2732,N_2685,N_2663);
nand U2733 (N_2733,N_2653,N_2670);
nor U2734 (N_2734,N_2684,N_2668);
nor U2735 (N_2735,N_2655,N_2696);
and U2736 (N_2736,N_2657,N_2679);
and U2737 (N_2737,N_2688,N_2695);
and U2738 (N_2738,N_2679,N_2672);
or U2739 (N_2739,N_2688,N_2674);
nor U2740 (N_2740,N_2670,N_2681);
nor U2741 (N_2741,N_2675,N_2697);
and U2742 (N_2742,N_2654,N_2663);
and U2743 (N_2743,N_2673,N_2669);
and U2744 (N_2744,N_2695,N_2675);
or U2745 (N_2745,N_2664,N_2675);
and U2746 (N_2746,N_2675,N_2688);
nor U2747 (N_2747,N_2655,N_2652);
nand U2748 (N_2748,N_2657,N_2691);
and U2749 (N_2749,N_2674,N_2659);
nand U2750 (N_2750,N_2716,N_2715);
and U2751 (N_2751,N_2724,N_2700);
nand U2752 (N_2752,N_2729,N_2705);
nand U2753 (N_2753,N_2725,N_2722);
xnor U2754 (N_2754,N_2708,N_2745);
and U2755 (N_2755,N_2718,N_2742);
xnor U2756 (N_2756,N_2703,N_2720);
or U2757 (N_2757,N_2736,N_2732);
xnor U2758 (N_2758,N_2749,N_2748);
and U2759 (N_2759,N_2728,N_2740);
and U2760 (N_2760,N_2701,N_2731);
or U2761 (N_2761,N_2738,N_2741);
or U2762 (N_2762,N_2704,N_2712);
or U2763 (N_2763,N_2730,N_2723);
nor U2764 (N_2764,N_2717,N_2719);
or U2765 (N_2765,N_2727,N_2714);
nor U2766 (N_2766,N_2746,N_2743);
and U2767 (N_2767,N_2711,N_2747);
xnor U2768 (N_2768,N_2709,N_2737);
nand U2769 (N_2769,N_2733,N_2710);
and U2770 (N_2770,N_2702,N_2734);
nand U2771 (N_2771,N_2721,N_2707);
xnor U2772 (N_2772,N_2735,N_2744);
nor U2773 (N_2773,N_2726,N_2706);
xor U2774 (N_2774,N_2739,N_2713);
and U2775 (N_2775,N_2706,N_2703);
and U2776 (N_2776,N_2749,N_2725);
nor U2777 (N_2777,N_2745,N_2740);
and U2778 (N_2778,N_2747,N_2703);
and U2779 (N_2779,N_2706,N_2744);
xor U2780 (N_2780,N_2727,N_2702);
and U2781 (N_2781,N_2720,N_2729);
or U2782 (N_2782,N_2713,N_2717);
and U2783 (N_2783,N_2713,N_2743);
or U2784 (N_2784,N_2749,N_2734);
xor U2785 (N_2785,N_2703,N_2744);
nor U2786 (N_2786,N_2707,N_2702);
and U2787 (N_2787,N_2726,N_2721);
and U2788 (N_2788,N_2702,N_2740);
or U2789 (N_2789,N_2727,N_2717);
and U2790 (N_2790,N_2723,N_2705);
nor U2791 (N_2791,N_2727,N_2740);
and U2792 (N_2792,N_2714,N_2743);
nor U2793 (N_2793,N_2745,N_2743);
and U2794 (N_2794,N_2702,N_2737);
and U2795 (N_2795,N_2738,N_2713);
and U2796 (N_2796,N_2700,N_2726);
nor U2797 (N_2797,N_2707,N_2743);
nand U2798 (N_2798,N_2737,N_2723);
nor U2799 (N_2799,N_2717,N_2714);
nand U2800 (N_2800,N_2786,N_2753);
nor U2801 (N_2801,N_2783,N_2751);
xnor U2802 (N_2802,N_2770,N_2794);
xnor U2803 (N_2803,N_2764,N_2789);
nor U2804 (N_2804,N_2769,N_2774);
and U2805 (N_2805,N_2780,N_2756);
or U2806 (N_2806,N_2779,N_2787);
or U2807 (N_2807,N_2799,N_2798);
or U2808 (N_2808,N_2791,N_2781);
and U2809 (N_2809,N_2792,N_2758);
nand U2810 (N_2810,N_2752,N_2775);
nand U2811 (N_2811,N_2777,N_2790);
nor U2812 (N_2812,N_2795,N_2761);
or U2813 (N_2813,N_2785,N_2755);
and U2814 (N_2814,N_2762,N_2760);
and U2815 (N_2815,N_2793,N_2788);
or U2816 (N_2816,N_2797,N_2771);
and U2817 (N_2817,N_2750,N_2757);
nand U2818 (N_2818,N_2763,N_2776);
nor U2819 (N_2819,N_2772,N_2765);
nand U2820 (N_2820,N_2782,N_2796);
and U2821 (N_2821,N_2766,N_2754);
nor U2822 (N_2822,N_2778,N_2773);
xor U2823 (N_2823,N_2767,N_2759);
nand U2824 (N_2824,N_2784,N_2768);
nor U2825 (N_2825,N_2755,N_2799);
xnor U2826 (N_2826,N_2784,N_2790);
xnor U2827 (N_2827,N_2798,N_2763);
nand U2828 (N_2828,N_2756,N_2795);
and U2829 (N_2829,N_2797,N_2793);
nor U2830 (N_2830,N_2787,N_2786);
and U2831 (N_2831,N_2774,N_2763);
xnor U2832 (N_2832,N_2768,N_2797);
xor U2833 (N_2833,N_2773,N_2764);
nor U2834 (N_2834,N_2761,N_2765);
or U2835 (N_2835,N_2780,N_2796);
nor U2836 (N_2836,N_2753,N_2765);
nor U2837 (N_2837,N_2779,N_2776);
nor U2838 (N_2838,N_2783,N_2797);
nand U2839 (N_2839,N_2771,N_2763);
nor U2840 (N_2840,N_2770,N_2773);
nor U2841 (N_2841,N_2796,N_2797);
and U2842 (N_2842,N_2761,N_2787);
nand U2843 (N_2843,N_2778,N_2751);
nand U2844 (N_2844,N_2760,N_2750);
and U2845 (N_2845,N_2781,N_2795);
nor U2846 (N_2846,N_2790,N_2769);
or U2847 (N_2847,N_2761,N_2797);
xor U2848 (N_2848,N_2788,N_2778);
nand U2849 (N_2849,N_2753,N_2754);
or U2850 (N_2850,N_2812,N_2832);
or U2851 (N_2851,N_2819,N_2806);
nand U2852 (N_2852,N_2826,N_2838);
or U2853 (N_2853,N_2827,N_2801);
or U2854 (N_2854,N_2811,N_2816);
and U2855 (N_2855,N_2808,N_2814);
xor U2856 (N_2856,N_2820,N_2818);
and U2857 (N_2857,N_2817,N_2829);
or U2858 (N_2858,N_2846,N_2805);
xor U2859 (N_2859,N_2833,N_2830);
nand U2860 (N_2860,N_2839,N_2803);
or U2861 (N_2861,N_2822,N_2800);
nand U2862 (N_2862,N_2810,N_2845);
and U2863 (N_2863,N_2824,N_2807);
xnor U2864 (N_2864,N_2847,N_2802);
nand U2865 (N_2865,N_2831,N_2842);
nand U2866 (N_2866,N_2804,N_2813);
nand U2867 (N_2867,N_2844,N_2821);
nor U2868 (N_2868,N_2848,N_2837);
nor U2869 (N_2869,N_2849,N_2834);
nand U2870 (N_2870,N_2809,N_2836);
and U2871 (N_2871,N_2825,N_2823);
nand U2872 (N_2872,N_2828,N_2840);
and U2873 (N_2873,N_2843,N_2841);
nand U2874 (N_2874,N_2815,N_2835);
and U2875 (N_2875,N_2813,N_2837);
xnor U2876 (N_2876,N_2844,N_2806);
nand U2877 (N_2877,N_2825,N_2803);
nand U2878 (N_2878,N_2829,N_2802);
nand U2879 (N_2879,N_2804,N_2839);
nand U2880 (N_2880,N_2839,N_2829);
and U2881 (N_2881,N_2802,N_2826);
and U2882 (N_2882,N_2829,N_2844);
and U2883 (N_2883,N_2806,N_2817);
xor U2884 (N_2884,N_2821,N_2807);
and U2885 (N_2885,N_2819,N_2836);
nor U2886 (N_2886,N_2819,N_2818);
nor U2887 (N_2887,N_2849,N_2847);
and U2888 (N_2888,N_2807,N_2810);
and U2889 (N_2889,N_2841,N_2837);
nor U2890 (N_2890,N_2839,N_2847);
nor U2891 (N_2891,N_2800,N_2807);
and U2892 (N_2892,N_2800,N_2804);
or U2893 (N_2893,N_2803,N_2844);
nand U2894 (N_2894,N_2833,N_2837);
or U2895 (N_2895,N_2824,N_2819);
or U2896 (N_2896,N_2834,N_2807);
nor U2897 (N_2897,N_2822,N_2829);
nand U2898 (N_2898,N_2839,N_2832);
or U2899 (N_2899,N_2827,N_2830);
xnor U2900 (N_2900,N_2894,N_2852);
and U2901 (N_2901,N_2868,N_2885);
or U2902 (N_2902,N_2865,N_2891);
nor U2903 (N_2903,N_2864,N_2850);
nand U2904 (N_2904,N_2887,N_2869);
nand U2905 (N_2905,N_2862,N_2866);
nor U2906 (N_2906,N_2898,N_2878);
nor U2907 (N_2907,N_2892,N_2870);
xor U2908 (N_2908,N_2879,N_2875);
nor U2909 (N_2909,N_2880,N_2882);
nand U2910 (N_2910,N_2859,N_2874);
and U2911 (N_2911,N_2883,N_2863);
nand U2912 (N_2912,N_2881,N_2896);
nor U2913 (N_2913,N_2855,N_2872);
or U2914 (N_2914,N_2873,N_2876);
nor U2915 (N_2915,N_2888,N_2871);
nor U2916 (N_2916,N_2886,N_2861);
nor U2917 (N_2917,N_2858,N_2897);
nor U2918 (N_2918,N_2877,N_2851);
xor U2919 (N_2919,N_2893,N_2853);
or U2920 (N_2920,N_2860,N_2854);
nand U2921 (N_2921,N_2867,N_2889);
and U2922 (N_2922,N_2884,N_2899);
or U2923 (N_2923,N_2857,N_2856);
xnor U2924 (N_2924,N_2890,N_2895);
or U2925 (N_2925,N_2887,N_2894);
nor U2926 (N_2926,N_2875,N_2865);
nand U2927 (N_2927,N_2887,N_2874);
or U2928 (N_2928,N_2893,N_2852);
nor U2929 (N_2929,N_2894,N_2888);
nand U2930 (N_2930,N_2877,N_2856);
nor U2931 (N_2931,N_2896,N_2880);
nand U2932 (N_2932,N_2863,N_2850);
and U2933 (N_2933,N_2876,N_2858);
nand U2934 (N_2934,N_2851,N_2874);
nand U2935 (N_2935,N_2871,N_2884);
xnor U2936 (N_2936,N_2898,N_2852);
nand U2937 (N_2937,N_2877,N_2889);
nor U2938 (N_2938,N_2896,N_2860);
nor U2939 (N_2939,N_2853,N_2874);
and U2940 (N_2940,N_2884,N_2896);
or U2941 (N_2941,N_2891,N_2854);
nand U2942 (N_2942,N_2893,N_2891);
nor U2943 (N_2943,N_2866,N_2874);
and U2944 (N_2944,N_2886,N_2894);
nor U2945 (N_2945,N_2898,N_2862);
nor U2946 (N_2946,N_2852,N_2883);
or U2947 (N_2947,N_2865,N_2864);
and U2948 (N_2948,N_2869,N_2881);
nand U2949 (N_2949,N_2882,N_2852);
or U2950 (N_2950,N_2915,N_2939);
nor U2951 (N_2951,N_2938,N_2925);
and U2952 (N_2952,N_2913,N_2947);
xor U2953 (N_2953,N_2910,N_2936);
and U2954 (N_2954,N_2904,N_2905);
xor U2955 (N_2955,N_2914,N_2909);
xor U2956 (N_2956,N_2900,N_2912);
and U2957 (N_2957,N_2930,N_2942);
and U2958 (N_2958,N_2921,N_2906);
and U2959 (N_2959,N_2908,N_2924);
or U2960 (N_2960,N_2923,N_2911);
nor U2961 (N_2961,N_2944,N_2902);
nor U2962 (N_2962,N_2920,N_2918);
nand U2963 (N_2963,N_2934,N_2946);
and U2964 (N_2964,N_2941,N_2937);
nand U2965 (N_2965,N_2928,N_2901);
or U2966 (N_2966,N_2919,N_2943);
xnor U2967 (N_2967,N_2916,N_2931);
or U2968 (N_2968,N_2940,N_2933);
or U2969 (N_2969,N_2949,N_2935);
nor U2970 (N_2970,N_2926,N_2903);
and U2971 (N_2971,N_2929,N_2945);
and U2972 (N_2972,N_2948,N_2917);
nand U2973 (N_2973,N_2922,N_2907);
and U2974 (N_2974,N_2927,N_2932);
or U2975 (N_2975,N_2925,N_2916);
and U2976 (N_2976,N_2933,N_2936);
or U2977 (N_2977,N_2936,N_2914);
nor U2978 (N_2978,N_2911,N_2914);
or U2979 (N_2979,N_2935,N_2932);
and U2980 (N_2980,N_2937,N_2935);
or U2981 (N_2981,N_2928,N_2945);
nor U2982 (N_2982,N_2900,N_2946);
or U2983 (N_2983,N_2902,N_2935);
and U2984 (N_2984,N_2929,N_2904);
nand U2985 (N_2985,N_2948,N_2901);
nor U2986 (N_2986,N_2933,N_2916);
and U2987 (N_2987,N_2904,N_2949);
or U2988 (N_2988,N_2928,N_2926);
nor U2989 (N_2989,N_2929,N_2911);
nand U2990 (N_2990,N_2909,N_2922);
or U2991 (N_2991,N_2925,N_2927);
nor U2992 (N_2992,N_2903,N_2915);
and U2993 (N_2993,N_2949,N_2911);
and U2994 (N_2994,N_2904,N_2908);
nand U2995 (N_2995,N_2906,N_2939);
nand U2996 (N_2996,N_2929,N_2909);
or U2997 (N_2997,N_2915,N_2914);
and U2998 (N_2998,N_2900,N_2923);
and U2999 (N_2999,N_2933,N_2921);
and UO_0 (O_0,N_2969,N_2963);
nand UO_1 (O_1,N_2962,N_2966);
xor UO_2 (O_2,N_2961,N_2957);
xnor UO_3 (O_3,N_2965,N_2998);
nor UO_4 (O_4,N_2972,N_2968);
xor UO_5 (O_5,N_2979,N_2992);
xor UO_6 (O_6,N_2984,N_2970);
or UO_7 (O_7,N_2991,N_2959);
or UO_8 (O_8,N_2950,N_2952);
or UO_9 (O_9,N_2956,N_2983);
nand UO_10 (O_10,N_2988,N_2996);
nor UO_11 (O_11,N_2980,N_2995);
nand UO_12 (O_12,N_2977,N_2960);
xnor UO_13 (O_13,N_2982,N_2974);
nor UO_14 (O_14,N_2981,N_2997);
nand UO_15 (O_15,N_2989,N_2967);
nand UO_16 (O_16,N_2953,N_2987);
nand UO_17 (O_17,N_2964,N_2958);
or UO_18 (O_18,N_2999,N_2955);
xnor UO_19 (O_19,N_2973,N_2990);
nand UO_20 (O_20,N_2985,N_2976);
nand UO_21 (O_21,N_2986,N_2993);
nor UO_22 (O_22,N_2971,N_2994);
nor UO_23 (O_23,N_2978,N_2975);
nand UO_24 (O_24,N_2951,N_2954);
nor UO_25 (O_25,N_2998,N_2969);
xnor UO_26 (O_26,N_2990,N_2992);
nand UO_27 (O_27,N_2951,N_2974);
nor UO_28 (O_28,N_2956,N_2985);
and UO_29 (O_29,N_2967,N_2984);
and UO_30 (O_30,N_2999,N_2952);
nand UO_31 (O_31,N_2992,N_2965);
and UO_32 (O_32,N_2987,N_2984);
nor UO_33 (O_33,N_2985,N_2992);
xnor UO_34 (O_34,N_2950,N_2999);
or UO_35 (O_35,N_2966,N_2981);
and UO_36 (O_36,N_2982,N_2993);
or UO_37 (O_37,N_2985,N_2954);
and UO_38 (O_38,N_2983,N_2951);
nor UO_39 (O_39,N_2956,N_2988);
and UO_40 (O_40,N_2997,N_2954);
and UO_41 (O_41,N_2969,N_2995);
nor UO_42 (O_42,N_2960,N_2995);
and UO_43 (O_43,N_2955,N_2992);
xnor UO_44 (O_44,N_2969,N_2954);
and UO_45 (O_45,N_2974,N_2984);
or UO_46 (O_46,N_2964,N_2959);
nand UO_47 (O_47,N_2973,N_2951);
and UO_48 (O_48,N_2958,N_2967);
or UO_49 (O_49,N_2992,N_2956);
nor UO_50 (O_50,N_2964,N_2986);
or UO_51 (O_51,N_2978,N_2959);
nor UO_52 (O_52,N_2996,N_2980);
and UO_53 (O_53,N_2994,N_2979);
or UO_54 (O_54,N_2972,N_2979);
nor UO_55 (O_55,N_2990,N_2960);
or UO_56 (O_56,N_2990,N_2968);
nand UO_57 (O_57,N_2968,N_2997);
and UO_58 (O_58,N_2988,N_2961);
nand UO_59 (O_59,N_2987,N_2995);
nor UO_60 (O_60,N_2958,N_2969);
and UO_61 (O_61,N_2970,N_2971);
nand UO_62 (O_62,N_2991,N_2978);
nor UO_63 (O_63,N_2969,N_2951);
and UO_64 (O_64,N_2950,N_2955);
nor UO_65 (O_65,N_2964,N_2982);
nor UO_66 (O_66,N_2956,N_2973);
or UO_67 (O_67,N_2996,N_2982);
nand UO_68 (O_68,N_2973,N_2957);
nand UO_69 (O_69,N_2977,N_2989);
nor UO_70 (O_70,N_2961,N_2994);
xnor UO_71 (O_71,N_2950,N_2980);
nand UO_72 (O_72,N_2952,N_2951);
nand UO_73 (O_73,N_2994,N_2967);
nand UO_74 (O_74,N_2992,N_2996);
and UO_75 (O_75,N_2955,N_2967);
nand UO_76 (O_76,N_2961,N_2984);
or UO_77 (O_77,N_2991,N_2961);
or UO_78 (O_78,N_2989,N_2990);
or UO_79 (O_79,N_2990,N_2952);
or UO_80 (O_80,N_2954,N_2959);
and UO_81 (O_81,N_2997,N_2999);
nor UO_82 (O_82,N_2959,N_2996);
nor UO_83 (O_83,N_2962,N_2990);
xor UO_84 (O_84,N_2952,N_2953);
nand UO_85 (O_85,N_2993,N_2983);
nor UO_86 (O_86,N_2963,N_2967);
and UO_87 (O_87,N_2989,N_2965);
nor UO_88 (O_88,N_2972,N_2999);
nand UO_89 (O_89,N_2995,N_2966);
nor UO_90 (O_90,N_2997,N_2974);
and UO_91 (O_91,N_2999,N_2982);
and UO_92 (O_92,N_2976,N_2956);
and UO_93 (O_93,N_2962,N_2986);
nand UO_94 (O_94,N_2994,N_2982);
or UO_95 (O_95,N_2954,N_2965);
or UO_96 (O_96,N_2994,N_2958);
or UO_97 (O_97,N_2957,N_2978);
or UO_98 (O_98,N_2954,N_2998);
xor UO_99 (O_99,N_2996,N_2978);
and UO_100 (O_100,N_2967,N_2971);
nor UO_101 (O_101,N_2988,N_2965);
and UO_102 (O_102,N_2981,N_2951);
or UO_103 (O_103,N_2968,N_2963);
and UO_104 (O_104,N_2973,N_2969);
nand UO_105 (O_105,N_2994,N_2959);
or UO_106 (O_106,N_2951,N_2998);
and UO_107 (O_107,N_2969,N_2950);
nand UO_108 (O_108,N_2984,N_2972);
nand UO_109 (O_109,N_2972,N_2986);
or UO_110 (O_110,N_2978,N_2983);
or UO_111 (O_111,N_2959,N_2997);
nand UO_112 (O_112,N_2974,N_2968);
and UO_113 (O_113,N_2978,N_2968);
nor UO_114 (O_114,N_2996,N_2952);
or UO_115 (O_115,N_2957,N_2969);
xor UO_116 (O_116,N_2968,N_2973);
nor UO_117 (O_117,N_2977,N_2991);
or UO_118 (O_118,N_2972,N_2973);
nor UO_119 (O_119,N_2968,N_2967);
nor UO_120 (O_120,N_2988,N_2968);
and UO_121 (O_121,N_2966,N_2961);
nand UO_122 (O_122,N_2974,N_2971);
or UO_123 (O_123,N_2970,N_2988);
and UO_124 (O_124,N_2954,N_2981);
or UO_125 (O_125,N_2950,N_2987);
nor UO_126 (O_126,N_2990,N_2994);
and UO_127 (O_127,N_2997,N_2988);
nand UO_128 (O_128,N_2973,N_2953);
and UO_129 (O_129,N_2991,N_2962);
xor UO_130 (O_130,N_2990,N_2954);
or UO_131 (O_131,N_2997,N_2970);
or UO_132 (O_132,N_2952,N_2966);
nor UO_133 (O_133,N_2969,N_2976);
nor UO_134 (O_134,N_2951,N_2985);
or UO_135 (O_135,N_2981,N_2960);
or UO_136 (O_136,N_2989,N_2974);
or UO_137 (O_137,N_2998,N_2950);
nand UO_138 (O_138,N_2971,N_2977);
nand UO_139 (O_139,N_2962,N_2952);
or UO_140 (O_140,N_2998,N_2957);
or UO_141 (O_141,N_2960,N_2996);
xor UO_142 (O_142,N_2995,N_2999);
nand UO_143 (O_143,N_2984,N_2999);
or UO_144 (O_144,N_2979,N_2982);
xnor UO_145 (O_145,N_2962,N_2975);
and UO_146 (O_146,N_2971,N_2969);
xnor UO_147 (O_147,N_2956,N_2984);
or UO_148 (O_148,N_2976,N_2962);
nand UO_149 (O_149,N_2987,N_2999);
and UO_150 (O_150,N_2988,N_2953);
and UO_151 (O_151,N_2963,N_2971);
nand UO_152 (O_152,N_2972,N_2953);
or UO_153 (O_153,N_2993,N_2954);
or UO_154 (O_154,N_2953,N_2968);
xnor UO_155 (O_155,N_2980,N_2992);
nand UO_156 (O_156,N_2993,N_2958);
nor UO_157 (O_157,N_2970,N_2979);
and UO_158 (O_158,N_2954,N_2964);
nor UO_159 (O_159,N_2956,N_2958);
xor UO_160 (O_160,N_2960,N_2961);
nand UO_161 (O_161,N_2950,N_2968);
nand UO_162 (O_162,N_2975,N_2952);
nand UO_163 (O_163,N_2961,N_2963);
nand UO_164 (O_164,N_2986,N_2990);
nand UO_165 (O_165,N_2952,N_2954);
and UO_166 (O_166,N_2985,N_2959);
or UO_167 (O_167,N_2961,N_2952);
and UO_168 (O_168,N_2991,N_2966);
nor UO_169 (O_169,N_2990,N_2976);
and UO_170 (O_170,N_2999,N_2983);
nand UO_171 (O_171,N_2988,N_2969);
nor UO_172 (O_172,N_2964,N_2962);
and UO_173 (O_173,N_2960,N_2957);
nand UO_174 (O_174,N_2970,N_2960);
nand UO_175 (O_175,N_2961,N_2992);
nor UO_176 (O_176,N_2979,N_2997);
or UO_177 (O_177,N_2994,N_2980);
nand UO_178 (O_178,N_2958,N_2988);
or UO_179 (O_179,N_2959,N_2998);
or UO_180 (O_180,N_2987,N_2954);
nand UO_181 (O_181,N_2986,N_2987);
or UO_182 (O_182,N_2958,N_2978);
and UO_183 (O_183,N_2955,N_2973);
or UO_184 (O_184,N_2980,N_2966);
nor UO_185 (O_185,N_2991,N_2976);
or UO_186 (O_186,N_2964,N_2998);
or UO_187 (O_187,N_2991,N_2953);
nand UO_188 (O_188,N_2962,N_2993);
nand UO_189 (O_189,N_2974,N_2978);
nor UO_190 (O_190,N_2983,N_2987);
nand UO_191 (O_191,N_2960,N_2971);
xnor UO_192 (O_192,N_2950,N_2982);
nand UO_193 (O_193,N_2967,N_2965);
or UO_194 (O_194,N_2958,N_2950);
and UO_195 (O_195,N_2999,N_2991);
and UO_196 (O_196,N_2993,N_2978);
nand UO_197 (O_197,N_2955,N_2978);
or UO_198 (O_198,N_2964,N_2960);
and UO_199 (O_199,N_2962,N_2977);
and UO_200 (O_200,N_2991,N_2989);
nand UO_201 (O_201,N_2983,N_2990);
or UO_202 (O_202,N_2990,N_2995);
nand UO_203 (O_203,N_2980,N_2964);
nor UO_204 (O_204,N_2981,N_2990);
nor UO_205 (O_205,N_2995,N_2953);
nand UO_206 (O_206,N_2996,N_2986);
xnor UO_207 (O_207,N_2976,N_2970);
and UO_208 (O_208,N_2955,N_2953);
nor UO_209 (O_209,N_2981,N_2973);
or UO_210 (O_210,N_2988,N_2989);
nor UO_211 (O_211,N_2966,N_2956);
xnor UO_212 (O_212,N_2973,N_2985);
or UO_213 (O_213,N_2951,N_2968);
and UO_214 (O_214,N_2962,N_2988);
and UO_215 (O_215,N_2996,N_2990);
or UO_216 (O_216,N_2950,N_2970);
nor UO_217 (O_217,N_2998,N_2973);
or UO_218 (O_218,N_2960,N_2954);
nand UO_219 (O_219,N_2972,N_2974);
and UO_220 (O_220,N_2966,N_2987);
and UO_221 (O_221,N_2983,N_2957);
xnor UO_222 (O_222,N_2972,N_2956);
or UO_223 (O_223,N_2958,N_2983);
and UO_224 (O_224,N_2977,N_2975);
nand UO_225 (O_225,N_2970,N_2957);
and UO_226 (O_226,N_2967,N_2995);
nor UO_227 (O_227,N_2961,N_2989);
nor UO_228 (O_228,N_2963,N_2989);
nor UO_229 (O_229,N_2960,N_2980);
nor UO_230 (O_230,N_2996,N_2967);
nor UO_231 (O_231,N_2988,N_2974);
or UO_232 (O_232,N_2988,N_2963);
nand UO_233 (O_233,N_2981,N_2980);
or UO_234 (O_234,N_2966,N_2968);
and UO_235 (O_235,N_2990,N_2998);
or UO_236 (O_236,N_2976,N_2981);
nor UO_237 (O_237,N_2956,N_2994);
or UO_238 (O_238,N_2991,N_2973);
xor UO_239 (O_239,N_2992,N_2976);
and UO_240 (O_240,N_2964,N_2995);
xor UO_241 (O_241,N_2961,N_2974);
and UO_242 (O_242,N_2969,N_2986);
nand UO_243 (O_243,N_2955,N_2972);
and UO_244 (O_244,N_2972,N_2971);
nor UO_245 (O_245,N_2989,N_2952);
or UO_246 (O_246,N_2967,N_2974);
and UO_247 (O_247,N_2965,N_2968);
or UO_248 (O_248,N_2991,N_2986);
xor UO_249 (O_249,N_2952,N_2995);
or UO_250 (O_250,N_2994,N_2972);
nand UO_251 (O_251,N_2995,N_2998);
and UO_252 (O_252,N_2958,N_2972);
xnor UO_253 (O_253,N_2962,N_2997);
nor UO_254 (O_254,N_2962,N_2999);
nand UO_255 (O_255,N_2971,N_2988);
nand UO_256 (O_256,N_2954,N_2957);
nand UO_257 (O_257,N_2979,N_2960);
or UO_258 (O_258,N_2993,N_2991);
nand UO_259 (O_259,N_2967,N_2998);
and UO_260 (O_260,N_2961,N_2954);
xor UO_261 (O_261,N_2955,N_2990);
or UO_262 (O_262,N_2965,N_2994);
and UO_263 (O_263,N_2974,N_2957);
xor UO_264 (O_264,N_2990,N_2980);
and UO_265 (O_265,N_2993,N_2988);
nand UO_266 (O_266,N_2975,N_2953);
and UO_267 (O_267,N_2955,N_2991);
and UO_268 (O_268,N_2989,N_2984);
or UO_269 (O_269,N_2984,N_2965);
and UO_270 (O_270,N_2974,N_2964);
nor UO_271 (O_271,N_2961,N_2979);
nor UO_272 (O_272,N_2968,N_2962);
nand UO_273 (O_273,N_2999,N_2957);
nand UO_274 (O_274,N_2970,N_2990);
xnor UO_275 (O_275,N_2979,N_2988);
xor UO_276 (O_276,N_2978,N_2956);
or UO_277 (O_277,N_2994,N_2970);
nand UO_278 (O_278,N_2994,N_2986);
nor UO_279 (O_279,N_2967,N_2973);
and UO_280 (O_280,N_2962,N_2972);
and UO_281 (O_281,N_2964,N_2981);
nand UO_282 (O_282,N_2950,N_2976);
and UO_283 (O_283,N_2982,N_2956);
and UO_284 (O_284,N_2952,N_2955);
nor UO_285 (O_285,N_2966,N_2963);
xor UO_286 (O_286,N_2982,N_2965);
nand UO_287 (O_287,N_2999,N_2966);
nor UO_288 (O_288,N_2966,N_2978);
xnor UO_289 (O_289,N_2955,N_2996);
nand UO_290 (O_290,N_2964,N_2965);
nand UO_291 (O_291,N_2958,N_2980);
and UO_292 (O_292,N_2983,N_2989);
nor UO_293 (O_293,N_2976,N_2967);
nor UO_294 (O_294,N_2968,N_2989);
or UO_295 (O_295,N_2998,N_2955);
nor UO_296 (O_296,N_2971,N_2965);
or UO_297 (O_297,N_2996,N_2974);
and UO_298 (O_298,N_2952,N_2997);
xor UO_299 (O_299,N_2988,N_2959);
xnor UO_300 (O_300,N_2983,N_2959);
or UO_301 (O_301,N_2992,N_2958);
or UO_302 (O_302,N_2977,N_2987);
nand UO_303 (O_303,N_2997,N_2985);
and UO_304 (O_304,N_2972,N_2995);
and UO_305 (O_305,N_2965,N_2976);
or UO_306 (O_306,N_2977,N_2964);
nor UO_307 (O_307,N_2967,N_2979);
nand UO_308 (O_308,N_2992,N_2998);
and UO_309 (O_309,N_2995,N_2961);
nand UO_310 (O_310,N_2983,N_2963);
xor UO_311 (O_311,N_2998,N_2993);
or UO_312 (O_312,N_2968,N_2969);
nand UO_313 (O_313,N_2960,N_2983);
or UO_314 (O_314,N_2965,N_2980);
and UO_315 (O_315,N_2991,N_2965);
nor UO_316 (O_316,N_2951,N_2988);
nor UO_317 (O_317,N_2996,N_2969);
nor UO_318 (O_318,N_2984,N_2988);
nor UO_319 (O_319,N_2969,N_2977);
and UO_320 (O_320,N_2979,N_2963);
or UO_321 (O_321,N_2995,N_2979);
or UO_322 (O_322,N_2981,N_2979);
and UO_323 (O_323,N_2965,N_2956);
and UO_324 (O_324,N_2950,N_2975);
or UO_325 (O_325,N_2955,N_2976);
nor UO_326 (O_326,N_2977,N_2980);
nor UO_327 (O_327,N_2959,N_2992);
or UO_328 (O_328,N_2960,N_2987);
or UO_329 (O_329,N_2998,N_2956);
or UO_330 (O_330,N_2997,N_2990);
or UO_331 (O_331,N_2994,N_2960);
or UO_332 (O_332,N_2980,N_2961);
nand UO_333 (O_333,N_2987,N_2982);
nor UO_334 (O_334,N_2996,N_2993);
nor UO_335 (O_335,N_2955,N_2993);
or UO_336 (O_336,N_2978,N_2999);
and UO_337 (O_337,N_2951,N_2980);
and UO_338 (O_338,N_2977,N_2963);
nor UO_339 (O_339,N_2954,N_2986);
nand UO_340 (O_340,N_2998,N_2974);
or UO_341 (O_341,N_2973,N_2989);
nor UO_342 (O_342,N_2962,N_2958);
and UO_343 (O_343,N_2987,N_2972);
nor UO_344 (O_344,N_2953,N_2998);
and UO_345 (O_345,N_2998,N_2986);
xor UO_346 (O_346,N_2980,N_2959);
nor UO_347 (O_347,N_2956,N_2987);
nand UO_348 (O_348,N_2956,N_2991);
nor UO_349 (O_349,N_2963,N_2994);
and UO_350 (O_350,N_2952,N_2971);
and UO_351 (O_351,N_2994,N_2992);
nand UO_352 (O_352,N_2955,N_2984);
or UO_353 (O_353,N_2952,N_2959);
or UO_354 (O_354,N_2980,N_2963);
nand UO_355 (O_355,N_2970,N_2995);
or UO_356 (O_356,N_2992,N_2970);
xor UO_357 (O_357,N_2954,N_2991);
nor UO_358 (O_358,N_2970,N_2980);
xnor UO_359 (O_359,N_2981,N_2965);
xnor UO_360 (O_360,N_2985,N_2953);
nand UO_361 (O_361,N_2984,N_2986);
and UO_362 (O_362,N_2960,N_2993);
nor UO_363 (O_363,N_2970,N_2986);
and UO_364 (O_364,N_2956,N_2979);
nand UO_365 (O_365,N_2952,N_2978);
and UO_366 (O_366,N_2986,N_2963);
nor UO_367 (O_367,N_2984,N_2975);
xor UO_368 (O_368,N_2954,N_2994);
and UO_369 (O_369,N_2986,N_2958);
or UO_370 (O_370,N_2990,N_2964);
or UO_371 (O_371,N_2956,N_2959);
nor UO_372 (O_372,N_2955,N_2997);
or UO_373 (O_373,N_2954,N_2989);
nor UO_374 (O_374,N_2994,N_2996);
nand UO_375 (O_375,N_2985,N_2967);
nor UO_376 (O_376,N_2964,N_2993);
and UO_377 (O_377,N_2974,N_2981);
nand UO_378 (O_378,N_2980,N_2953);
or UO_379 (O_379,N_2984,N_2997);
nand UO_380 (O_380,N_2962,N_2982);
and UO_381 (O_381,N_2950,N_2974);
nor UO_382 (O_382,N_2954,N_2953);
nor UO_383 (O_383,N_2953,N_2994);
xnor UO_384 (O_384,N_2973,N_2979);
nor UO_385 (O_385,N_2959,N_2958);
and UO_386 (O_386,N_2983,N_2971);
nand UO_387 (O_387,N_2967,N_2981);
nand UO_388 (O_388,N_2998,N_2976);
nor UO_389 (O_389,N_2997,N_2966);
xnor UO_390 (O_390,N_2952,N_2969);
nand UO_391 (O_391,N_2984,N_2950);
or UO_392 (O_392,N_2987,N_2964);
nand UO_393 (O_393,N_2951,N_2972);
nand UO_394 (O_394,N_2996,N_2984);
and UO_395 (O_395,N_2971,N_2981);
nor UO_396 (O_396,N_2966,N_2976);
and UO_397 (O_397,N_2984,N_2981);
nor UO_398 (O_398,N_2958,N_2960);
xor UO_399 (O_399,N_2951,N_2989);
nand UO_400 (O_400,N_2975,N_2957);
nor UO_401 (O_401,N_2975,N_2955);
nand UO_402 (O_402,N_2995,N_2996);
or UO_403 (O_403,N_2999,N_2967);
or UO_404 (O_404,N_2975,N_2990);
or UO_405 (O_405,N_2973,N_2997);
or UO_406 (O_406,N_2955,N_2956);
nor UO_407 (O_407,N_2989,N_2993);
nand UO_408 (O_408,N_2958,N_2973);
nor UO_409 (O_409,N_2973,N_2996);
nor UO_410 (O_410,N_2968,N_2977);
xor UO_411 (O_411,N_2999,N_2998);
or UO_412 (O_412,N_2987,N_2976);
or UO_413 (O_413,N_2951,N_2987);
and UO_414 (O_414,N_2964,N_2996);
xor UO_415 (O_415,N_2967,N_2960);
nand UO_416 (O_416,N_2977,N_2955);
nor UO_417 (O_417,N_2963,N_2982);
and UO_418 (O_418,N_2972,N_2976);
or UO_419 (O_419,N_2959,N_2987);
or UO_420 (O_420,N_2961,N_2983);
or UO_421 (O_421,N_2993,N_2979);
or UO_422 (O_422,N_2996,N_2977);
and UO_423 (O_423,N_2968,N_2976);
or UO_424 (O_424,N_2959,N_2957);
nor UO_425 (O_425,N_2950,N_2966);
nor UO_426 (O_426,N_2981,N_2968);
or UO_427 (O_427,N_2953,N_2956);
nand UO_428 (O_428,N_2983,N_2968);
and UO_429 (O_429,N_2972,N_2964);
nor UO_430 (O_430,N_2991,N_2987);
and UO_431 (O_431,N_2974,N_2962);
and UO_432 (O_432,N_2971,N_2978);
and UO_433 (O_433,N_2978,N_2982);
nor UO_434 (O_434,N_2951,N_2956);
nor UO_435 (O_435,N_2993,N_2992);
nor UO_436 (O_436,N_2984,N_2977);
nand UO_437 (O_437,N_2969,N_2962);
nand UO_438 (O_438,N_2969,N_2965);
and UO_439 (O_439,N_2973,N_2974);
nand UO_440 (O_440,N_2972,N_2991);
nand UO_441 (O_441,N_2950,N_2971);
nor UO_442 (O_442,N_2967,N_2954);
nand UO_443 (O_443,N_2989,N_2987);
nand UO_444 (O_444,N_2975,N_2965);
nor UO_445 (O_445,N_2987,N_2981);
and UO_446 (O_446,N_2988,N_2987);
xnor UO_447 (O_447,N_2991,N_2950);
or UO_448 (O_448,N_2957,N_2964);
or UO_449 (O_449,N_2960,N_2973);
and UO_450 (O_450,N_2993,N_2961);
or UO_451 (O_451,N_2958,N_2952);
or UO_452 (O_452,N_2957,N_2955);
nor UO_453 (O_453,N_2972,N_2993);
or UO_454 (O_454,N_2963,N_2972);
xor UO_455 (O_455,N_2976,N_2960);
or UO_456 (O_456,N_2985,N_2966);
nand UO_457 (O_457,N_2986,N_2953);
nor UO_458 (O_458,N_2959,N_2953);
or UO_459 (O_459,N_2965,N_2985);
xnor UO_460 (O_460,N_2952,N_2956);
xor UO_461 (O_461,N_2959,N_2979);
or UO_462 (O_462,N_2988,N_2995);
and UO_463 (O_463,N_2953,N_2982);
nor UO_464 (O_464,N_2955,N_2982);
nor UO_465 (O_465,N_2955,N_2963);
and UO_466 (O_466,N_2957,N_2986);
or UO_467 (O_467,N_2983,N_2980);
nand UO_468 (O_468,N_2970,N_2968);
and UO_469 (O_469,N_2991,N_2990);
or UO_470 (O_470,N_2985,N_2950);
nand UO_471 (O_471,N_2989,N_2953);
xnor UO_472 (O_472,N_2988,N_2967);
and UO_473 (O_473,N_2977,N_2954);
xnor UO_474 (O_474,N_2978,N_2981);
nor UO_475 (O_475,N_2985,N_2977);
nand UO_476 (O_476,N_2986,N_2983);
nand UO_477 (O_477,N_2976,N_2975);
nand UO_478 (O_478,N_2963,N_2991);
xor UO_479 (O_479,N_2956,N_2954);
or UO_480 (O_480,N_2962,N_2973);
nand UO_481 (O_481,N_2975,N_2994);
and UO_482 (O_482,N_2975,N_2956);
nor UO_483 (O_483,N_2952,N_2982);
nand UO_484 (O_484,N_2985,N_2979);
nor UO_485 (O_485,N_2993,N_2995);
nand UO_486 (O_486,N_2996,N_2951);
nand UO_487 (O_487,N_2961,N_2997);
or UO_488 (O_488,N_2992,N_2991);
or UO_489 (O_489,N_2964,N_2961);
and UO_490 (O_490,N_2967,N_2951);
and UO_491 (O_491,N_2997,N_2996);
xor UO_492 (O_492,N_2965,N_2995);
and UO_493 (O_493,N_2989,N_2956);
nor UO_494 (O_494,N_2980,N_2975);
or UO_495 (O_495,N_2990,N_2978);
nor UO_496 (O_496,N_2969,N_2975);
or UO_497 (O_497,N_2981,N_2982);
or UO_498 (O_498,N_2959,N_2982);
and UO_499 (O_499,N_2996,N_2970);
endmodule