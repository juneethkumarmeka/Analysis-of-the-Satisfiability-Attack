module basic_500_3000_500_5_levels_2xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_383,In_46);
and U1 (N_1,In_370,In_374);
and U2 (N_2,In_495,In_283);
or U3 (N_3,In_470,In_291);
nor U4 (N_4,In_323,In_103);
nor U5 (N_5,In_250,In_366);
or U6 (N_6,In_429,In_392);
or U7 (N_7,In_7,In_113);
or U8 (N_8,In_20,In_116);
nand U9 (N_9,In_346,In_410);
xnor U10 (N_10,In_231,In_152);
nand U11 (N_11,In_436,In_271);
nor U12 (N_12,In_57,In_237);
nor U13 (N_13,In_300,In_398);
and U14 (N_14,In_428,In_0);
nand U15 (N_15,In_453,In_320);
or U16 (N_16,In_361,In_365);
and U17 (N_17,In_308,In_13);
or U18 (N_18,In_432,In_350);
or U19 (N_19,In_490,In_50);
nand U20 (N_20,In_336,In_142);
nand U21 (N_21,In_433,In_232);
nand U22 (N_22,In_315,In_148);
nor U23 (N_23,In_264,In_90);
nor U24 (N_24,In_397,In_497);
nand U25 (N_25,In_440,In_401);
or U26 (N_26,In_62,In_419);
nor U27 (N_27,In_130,In_168);
nor U28 (N_28,In_171,In_89);
nand U29 (N_29,In_377,In_9);
or U30 (N_30,In_468,In_267);
nand U31 (N_31,In_489,In_40);
or U32 (N_32,In_212,In_159);
nand U33 (N_33,In_27,In_73);
nand U34 (N_34,In_394,In_345);
xnor U35 (N_35,In_165,In_303);
nand U36 (N_36,In_480,In_25);
or U37 (N_37,In_127,In_106);
and U38 (N_38,In_329,In_150);
or U39 (N_39,In_281,In_71);
or U40 (N_40,In_227,In_176);
and U41 (N_41,In_200,In_177);
and U42 (N_42,In_287,In_339);
nand U43 (N_43,In_249,In_282);
or U44 (N_44,In_342,In_349);
or U45 (N_45,In_298,In_33);
xor U46 (N_46,In_252,In_412);
and U47 (N_47,In_322,In_403);
nor U48 (N_48,In_402,In_121);
nor U49 (N_49,In_373,In_238);
nor U50 (N_50,In_385,In_460);
or U51 (N_51,In_133,In_347);
and U52 (N_52,In_371,In_301);
nand U53 (N_53,In_156,In_333);
or U54 (N_54,In_78,In_484);
nor U55 (N_55,In_293,In_262);
or U56 (N_56,In_414,In_265);
and U57 (N_57,In_444,In_155);
nand U58 (N_58,In_486,In_457);
nand U59 (N_59,In_306,In_359);
nand U60 (N_60,In_325,In_270);
nand U61 (N_61,In_216,In_154);
and U62 (N_62,In_491,In_230);
nor U63 (N_63,In_188,In_307);
nand U64 (N_64,In_132,In_96);
or U65 (N_65,In_151,In_74);
or U66 (N_66,In_215,In_77);
and U67 (N_67,In_245,In_338);
nand U68 (N_68,In_37,In_26);
nor U69 (N_69,In_290,In_161);
xor U70 (N_70,In_426,In_275);
or U71 (N_71,In_467,In_239);
nand U72 (N_72,In_81,In_311);
nor U73 (N_73,In_4,In_29);
and U74 (N_74,In_337,In_424);
or U75 (N_75,In_368,In_167);
and U76 (N_76,In_102,In_362);
nand U77 (N_77,In_475,In_418);
and U78 (N_78,In_114,In_134);
nand U79 (N_79,In_382,In_60);
nor U80 (N_80,In_242,In_97);
nor U81 (N_81,In_446,In_68);
or U82 (N_82,In_465,In_421);
nor U83 (N_83,In_15,In_408);
and U84 (N_84,In_56,In_69);
nand U85 (N_85,In_273,In_482);
nand U86 (N_86,In_105,In_492);
nor U87 (N_87,In_254,In_318);
or U88 (N_88,In_478,In_272);
or U89 (N_89,In_386,In_246);
nand U90 (N_90,In_358,In_51);
nand U91 (N_91,In_198,In_376);
nor U92 (N_92,In_352,In_396);
nor U93 (N_93,In_181,In_115);
or U94 (N_94,In_431,In_34);
and U95 (N_95,In_76,In_416);
xnor U96 (N_96,In_261,In_296);
nand U97 (N_97,In_191,In_192);
nor U98 (N_98,In_448,In_80);
nor U99 (N_99,In_472,In_248);
nand U100 (N_100,In_205,In_217);
xor U101 (N_101,In_479,In_119);
nand U102 (N_102,In_354,In_356);
or U103 (N_103,In_257,In_277);
xor U104 (N_104,In_206,In_314);
nand U105 (N_105,In_1,In_48);
nor U106 (N_106,In_251,In_118);
nand U107 (N_107,In_294,In_331);
or U108 (N_108,In_125,In_201);
nor U109 (N_109,In_445,In_407);
nor U110 (N_110,In_185,In_340);
nand U111 (N_111,In_169,In_391);
nand U112 (N_112,In_44,In_88);
or U113 (N_113,In_499,In_312);
nor U114 (N_114,In_461,In_143);
xor U115 (N_115,In_24,In_422);
nor U116 (N_116,In_138,In_321);
or U117 (N_117,In_12,In_65);
nand U118 (N_118,In_140,In_413);
nand U119 (N_119,In_14,In_86);
nor U120 (N_120,In_43,In_434);
nor U121 (N_121,In_63,In_190);
and U122 (N_122,In_128,In_47);
nand U123 (N_123,In_483,In_111);
nand U124 (N_124,In_91,In_149);
and U125 (N_125,In_10,In_243);
nor U126 (N_126,In_268,In_124);
or U127 (N_127,In_450,In_225);
nand U128 (N_128,In_488,In_469);
nand U129 (N_129,In_59,In_112);
nand U130 (N_130,In_35,In_335);
nand U131 (N_131,In_5,In_305);
and U132 (N_132,In_313,In_195);
and U133 (N_133,In_420,In_375);
nor U134 (N_134,In_255,In_18);
nor U135 (N_135,In_45,In_395);
nor U136 (N_136,In_438,In_187);
and U137 (N_137,In_92,In_477);
xor U138 (N_138,In_297,In_266);
or U139 (N_139,In_213,In_344);
or U140 (N_140,In_388,In_202);
nand U141 (N_141,In_302,In_456);
nor U142 (N_142,In_330,In_380);
or U143 (N_143,In_61,In_295);
or U144 (N_144,In_332,In_226);
nand U145 (N_145,In_8,In_348);
and U146 (N_146,In_109,In_53);
nor U147 (N_147,In_170,In_28);
or U148 (N_148,In_363,In_279);
nor U149 (N_149,In_274,In_319);
and U150 (N_150,In_441,In_487);
and U151 (N_151,In_99,In_235);
nor U152 (N_152,In_471,In_343);
or U153 (N_153,In_415,In_430);
nor U154 (N_154,In_459,In_87);
or U155 (N_155,In_107,In_316);
nor U156 (N_156,In_276,In_442);
or U157 (N_157,In_400,In_357);
nor U158 (N_158,In_207,In_135);
nand U159 (N_159,In_208,In_104);
or U160 (N_160,In_199,In_222);
nor U161 (N_161,In_427,In_58);
nor U162 (N_162,In_189,In_153);
nor U163 (N_163,In_146,In_6);
nand U164 (N_164,In_258,In_79);
and U165 (N_165,In_304,In_32);
xnor U166 (N_166,In_317,In_67);
or U167 (N_167,In_66,In_209);
nor U168 (N_168,In_259,In_141);
nor U169 (N_169,In_117,In_131);
nor U170 (N_170,In_42,In_224);
and U171 (N_171,In_341,In_164);
or U172 (N_172,In_405,In_372);
nand U173 (N_173,In_95,In_203);
nand U174 (N_174,In_379,In_41);
and U175 (N_175,In_204,In_473);
and U176 (N_176,In_485,In_23);
nand U177 (N_177,In_183,In_389);
nor U178 (N_178,In_98,In_417);
and U179 (N_179,In_21,In_334);
or U180 (N_180,In_455,In_129);
or U181 (N_181,In_292,In_476);
or U182 (N_182,In_145,In_197);
nand U183 (N_183,In_233,In_411);
and U184 (N_184,In_423,In_22);
nand U185 (N_185,In_299,In_184);
and U186 (N_186,In_240,In_289);
or U187 (N_187,In_174,In_481);
or U188 (N_188,In_173,In_30);
nand U189 (N_189,In_218,In_166);
nand U190 (N_190,In_280,In_452);
or U191 (N_191,In_136,In_496);
nand U192 (N_192,In_193,In_82);
nor U193 (N_193,In_384,In_228);
xor U194 (N_194,In_369,In_162);
or U195 (N_195,In_406,In_180);
and U196 (N_196,In_223,In_494);
and U197 (N_197,In_75,In_234);
and U198 (N_198,In_221,In_85);
nor U199 (N_199,In_309,In_55);
and U200 (N_200,In_443,In_84);
or U201 (N_201,In_2,In_70);
nor U202 (N_202,In_381,In_404);
nand U203 (N_203,In_360,In_178);
nand U204 (N_204,In_94,In_54);
xnor U205 (N_205,In_182,In_186);
or U206 (N_206,In_244,In_463);
nand U207 (N_207,In_462,In_458);
nor U208 (N_208,In_286,In_474);
nand U209 (N_209,In_367,In_11);
or U210 (N_210,In_172,In_253);
or U211 (N_211,In_324,In_210);
nor U212 (N_212,In_437,In_236);
and U213 (N_213,In_123,In_49);
and U214 (N_214,In_52,In_100);
or U215 (N_215,In_241,In_327);
or U216 (N_216,In_285,In_256);
nand U217 (N_217,In_93,In_110);
nand U218 (N_218,In_158,In_409);
and U219 (N_219,In_390,In_364);
nor U220 (N_220,In_399,In_16);
or U221 (N_221,In_72,In_260);
nand U222 (N_222,In_31,In_144);
and U223 (N_223,In_38,In_326);
or U224 (N_224,In_263,In_464);
nor U225 (N_225,In_83,In_449);
or U226 (N_226,In_175,In_220);
and U227 (N_227,In_157,In_310);
nor U228 (N_228,In_126,In_196);
nor U229 (N_229,In_179,In_328);
or U230 (N_230,In_351,In_387);
nand U231 (N_231,In_425,In_439);
or U232 (N_232,In_39,In_108);
and U233 (N_233,In_120,In_493);
and U234 (N_234,In_211,In_355);
nand U235 (N_235,In_447,In_19);
and U236 (N_236,In_214,In_101);
or U237 (N_237,In_160,In_284);
nor U238 (N_238,In_17,In_353);
nand U239 (N_239,In_451,In_219);
nand U240 (N_240,In_194,In_269);
or U241 (N_241,In_137,In_139);
and U242 (N_242,In_454,In_36);
and U243 (N_243,In_147,In_229);
nor U244 (N_244,In_3,In_278);
nand U245 (N_245,In_466,In_378);
or U246 (N_246,In_122,In_435);
nand U247 (N_247,In_163,In_393);
and U248 (N_248,In_247,In_64);
and U249 (N_249,In_288,In_498);
nor U250 (N_250,In_113,In_339);
nor U251 (N_251,In_56,In_362);
nand U252 (N_252,In_19,In_68);
nor U253 (N_253,In_406,In_142);
nand U254 (N_254,In_480,In_483);
nand U255 (N_255,In_351,In_135);
nand U256 (N_256,In_358,In_497);
and U257 (N_257,In_468,In_40);
or U258 (N_258,In_403,In_288);
nand U259 (N_259,In_122,In_296);
and U260 (N_260,In_71,In_70);
and U261 (N_261,In_433,In_159);
and U262 (N_262,In_180,In_288);
nand U263 (N_263,In_254,In_32);
nor U264 (N_264,In_90,In_266);
nor U265 (N_265,In_446,In_196);
nor U266 (N_266,In_143,In_13);
and U267 (N_267,In_358,In_355);
nand U268 (N_268,In_216,In_466);
nand U269 (N_269,In_234,In_63);
nor U270 (N_270,In_404,In_155);
or U271 (N_271,In_329,In_17);
and U272 (N_272,In_378,In_260);
nand U273 (N_273,In_307,In_453);
nand U274 (N_274,In_242,In_212);
xor U275 (N_275,In_191,In_19);
or U276 (N_276,In_471,In_487);
xnor U277 (N_277,In_472,In_45);
or U278 (N_278,In_318,In_327);
and U279 (N_279,In_246,In_131);
nor U280 (N_280,In_310,In_134);
or U281 (N_281,In_387,In_136);
nor U282 (N_282,In_51,In_472);
nand U283 (N_283,In_138,In_342);
nand U284 (N_284,In_200,In_413);
and U285 (N_285,In_203,In_468);
and U286 (N_286,In_80,In_481);
or U287 (N_287,In_474,In_182);
nor U288 (N_288,In_417,In_175);
nor U289 (N_289,In_119,In_323);
and U290 (N_290,In_235,In_109);
xor U291 (N_291,In_289,In_414);
nand U292 (N_292,In_342,In_403);
nor U293 (N_293,In_296,In_72);
or U294 (N_294,In_301,In_320);
or U295 (N_295,In_11,In_495);
nand U296 (N_296,In_385,In_495);
nor U297 (N_297,In_252,In_379);
and U298 (N_298,In_9,In_177);
nand U299 (N_299,In_299,In_257);
nor U300 (N_300,In_297,In_26);
nand U301 (N_301,In_379,In_6);
and U302 (N_302,In_115,In_497);
nand U303 (N_303,In_389,In_261);
and U304 (N_304,In_66,In_116);
nand U305 (N_305,In_196,In_339);
or U306 (N_306,In_10,In_452);
and U307 (N_307,In_235,In_438);
and U308 (N_308,In_418,In_41);
and U309 (N_309,In_203,In_352);
or U310 (N_310,In_415,In_165);
or U311 (N_311,In_12,In_290);
nand U312 (N_312,In_469,In_246);
nor U313 (N_313,In_439,In_192);
and U314 (N_314,In_176,In_300);
nand U315 (N_315,In_26,In_62);
or U316 (N_316,In_157,In_188);
or U317 (N_317,In_77,In_19);
nand U318 (N_318,In_487,In_220);
nand U319 (N_319,In_231,In_393);
nor U320 (N_320,In_418,In_431);
nor U321 (N_321,In_411,In_68);
or U322 (N_322,In_61,In_57);
nand U323 (N_323,In_470,In_160);
nand U324 (N_324,In_263,In_329);
nor U325 (N_325,In_164,In_2);
and U326 (N_326,In_22,In_392);
and U327 (N_327,In_351,In_226);
nand U328 (N_328,In_349,In_237);
nor U329 (N_329,In_403,In_413);
nor U330 (N_330,In_71,In_258);
and U331 (N_331,In_320,In_394);
nor U332 (N_332,In_438,In_24);
nand U333 (N_333,In_4,In_115);
nand U334 (N_334,In_395,In_105);
and U335 (N_335,In_56,In_230);
nand U336 (N_336,In_245,In_471);
and U337 (N_337,In_411,In_105);
and U338 (N_338,In_439,In_355);
or U339 (N_339,In_122,In_481);
nand U340 (N_340,In_297,In_369);
or U341 (N_341,In_344,In_305);
or U342 (N_342,In_129,In_352);
nor U343 (N_343,In_475,In_221);
and U344 (N_344,In_272,In_353);
and U345 (N_345,In_120,In_477);
nand U346 (N_346,In_383,In_391);
nand U347 (N_347,In_59,In_54);
and U348 (N_348,In_79,In_67);
nor U349 (N_349,In_487,In_69);
or U350 (N_350,In_196,In_329);
nor U351 (N_351,In_237,In_193);
or U352 (N_352,In_457,In_36);
nor U353 (N_353,In_13,In_293);
or U354 (N_354,In_53,In_247);
nand U355 (N_355,In_318,In_213);
xor U356 (N_356,In_130,In_347);
or U357 (N_357,In_176,In_448);
or U358 (N_358,In_160,In_24);
nor U359 (N_359,In_269,In_87);
nor U360 (N_360,In_265,In_85);
nand U361 (N_361,In_401,In_458);
nor U362 (N_362,In_187,In_434);
nand U363 (N_363,In_241,In_334);
nor U364 (N_364,In_107,In_407);
nand U365 (N_365,In_160,In_229);
nand U366 (N_366,In_317,In_205);
nor U367 (N_367,In_322,In_247);
or U368 (N_368,In_292,In_156);
and U369 (N_369,In_395,In_316);
nand U370 (N_370,In_432,In_28);
nand U371 (N_371,In_496,In_464);
nor U372 (N_372,In_17,In_342);
nand U373 (N_373,In_247,In_424);
nor U374 (N_374,In_133,In_432);
nor U375 (N_375,In_125,In_442);
or U376 (N_376,In_6,In_277);
nor U377 (N_377,In_70,In_225);
and U378 (N_378,In_248,In_368);
nor U379 (N_379,In_412,In_426);
nor U380 (N_380,In_231,In_409);
nand U381 (N_381,In_13,In_80);
and U382 (N_382,In_88,In_55);
nand U383 (N_383,In_255,In_10);
nor U384 (N_384,In_58,In_99);
nor U385 (N_385,In_227,In_90);
xnor U386 (N_386,In_462,In_175);
nor U387 (N_387,In_40,In_205);
nand U388 (N_388,In_468,In_430);
nor U389 (N_389,In_380,In_185);
or U390 (N_390,In_4,In_114);
or U391 (N_391,In_166,In_221);
nor U392 (N_392,In_146,In_468);
and U393 (N_393,In_380,In_102);
nand U394 (N_394,In_279,In_492);
or U395 (N_395,In_242,In_292);
nor U396 (N_396,In_340,In_130);
nand U397 (N_397,In_458,In_259);
nor U398 (N_398,In_173,In_446);
or U399 (N_399,In_43,In_386);
or U400 (N_400,In_399,In_49);
and U401 (N_401,In_90,In_330);
and U402 (N_402,In_341,In_159);
and U403 (N_403,In_369,In_486);
or U404 (N_404,In_371,In_133);
and U405 (N_405,In_422,In_232);
nand U406 (N_406,In_363,In_158);
and U407 (N_407,In_311,In_115);
nand U408 (N_408,In_49,In_47);
nor U409 (N_409,In_17,In_190);
and U410 (N_410,In_186,In_151);
nand U411 (N_411,In_311,In_210);
nor U412 (N_412,In_480,In_335);
nor U413 (N_413,In_36,In_181);
nor U414 (N_414,In_435,In_79);
or U415 (N_415,In_417,In_387);
or U416 (N_416,In_177,In_385);
nand U417 (N_417,In_364,In_21);
nand U418 (N_418,In_140,In_208);
and U419 (N_419,In_179,In_475);
and U420 (N_420,In_0,In_427);
or U421 (N_421,In_211,In_143);
nand U422 (N_422,In_446,In_58);
or U423 (N_423,In_147,In_218);
nand U424 (N_424,In_165,In_36);
and U425 (N_425,In_426,In_318);
nor U426 (N_426,In_212,In_137);
or U427 (N_427,In_289,In_99);
or U428 (N_428,In_262,In_426);
nor U429 (N_429,In_385,In_473);
and U430 (N_430,In_405,In_44);
or U431 (N_431,In_320,In_90);
and U432 (N_432,In_448,In_38);
and U433 (N_433,In_208,In_362);
and U434 (N_434,In_49,In_320);
nor U435 (N_435,In_401,In_236);
or U436 (N_436,In_478,In_49);
nand U437 (N_437,In_82,In_116);
nor U438 (N_438,In_432,In_490);
nand U439 (N_439,In_474,In_265);
or U440 (N_440,In_397,In_17);
nor U441 (N_441,In_450,In_336);
and U442 (N_442,In_436,In_397);
xor U443 (N_443,In_432,In_69);
and U444 (N_444,In_168,In_4);
nand U445 (N_445,In_241,In_53);
or U446 (N_446,In_310,In_475);
and U447 (N_447,In_98,In_452);
nor U448 (N_448,In_430,In_363);
nor U449 (N_449,In_134,In_463);
or U450 (N_450,In_57,In_258);
xor U451 (N_451,In_19,In_83);
nand U452 (N_452,In_277,In_136);
nor U453 (N_453,In_16,In_25);
or U454 (N_454,In_452,In_116);
nor U455 (N_455,In_499,In_187);
and U456 (N_456,In_18,In_321);
or U457 (N_457,In_0,In_193);
and U458 (N_458,In_359,In_339);
nand U459 (N_459,In_295,In_50);
nor U460 (N_460,In_300,In_334);
and U461 (N_461,In_477,In_435);
nor U462 (N_462,In_335,In_366);
nor U463 (N_463,In_78,In_294);
or U464 (N_464,In_159,In_302);
nand U465 (N_465,In_156,In_152);
or U466 (N_466,In_173,In_309);
nand U467 (N_467,In_225,In_390);
nand U468 (N_468,In_174,In_55);
nand U469 (N_469,In_66,In_23);
or U470 (N_470,In_275,In_245);
or U471 (N_471,In_332,In_54);
nand U472 (N_472,In_429,In_485);
and U473 (N_473,In_134,In_394);
or U474 (N_474,In_335,In_189);
nand U475 (N_475,In_404,In_410);
nor U476 (N_476,In_393,In_48);
nor U477 (N_477,In_489,In_93);
and U478 (N_478,In_181,In_195);
nor U479 (N_479,In_239,In_266);
nor U480 (N_480,In_59,In_57);
or U481 (N_481,In_168,In_42);
nor U482 (N_482,In_243,In_224);
xnor U483 (N_483,In_296,In_394);
nor U484 (N_484,In_211,In_127);
and U485 (N_485,In_107,In_53);
nand U486 (N_486,In_283,In_233);
nor U487 (N_487,In_174,In_94);
nor U488 (N_488,In_64,In_294);
nor U489 (N_489,In_397,In_420);
nand U490 (N_490,In_442,In_244);
xnor U491 (N_491,In_314,In_238);
or U492 (N_492,In_282,In_341);
nand U493 (N_493,In_422,In_260);
nor U494 (N_494,In_259,In_203);
or U495 (N_495,In_122,In_107);
and U496 (N_496,In_447,In_13);
nor U497 (N_497,In_231,In_404);
or U498 (N_498,In_281,In_98);
or U499 (N_499,In_249,In_56);
and U500 (N_500,In_284,In_177);
nand U501 (N_501,In_439,In_148);
nand U502 (N_502,In_308,In_260);
nand U503 (N_503,In_203,In_47);
or U504 (N_504,In_420,In_244);
or U505 (N_505,In_387,In_241);
and U506 (N_506,In_425,In_429);
nand U507 (N_507,In_338,In_399);
nor U508 (N_508,In_461,In_241);
or U509 (N_509,In_47,In_391);
nand U510 (N_510,In_49,In_135);
or U511 (N_511,In_137,In_28);
nand U512 (N_512,In_274,In_266);
or U513 (N_513,In_307,In_128);
nor U514 (N_514,In_310,In_311);
nor U515 (N_515,In_80,In_39);
nor U516 (N_516,In_128,In_424);
and U517 (N_517,In_326,In_451);
or U518 (N_518,In_479,In_157);
nand U519 (N_519,In_249,In_231);
nand U520 (N_520,In_321,In_464);
nand U521 (N_521,In_491,In_395);
or U522 (N_522,In_324,In_299);
nor U523 (N_523,In_454,In_0);
or U524 (N_524,In_322,In_113);
nor U525 (N_525,In_64,In_346);
and U526 (N_526,In_224,In_262);
xnor U527 (N_527,In_141,In_70);
and U528 (N_528,In_435,In_123);
nor U529 (N_529,In_130,In_149);
and U530 (N_530,In_141,In_473);
or U531 (N_531,In_365,In_299);
and U532 (N_532,In_7,In_289);
nand U533 (N_533,In_265,In_250);
and U534 (N_534,In_38,In_338);
nor U535 (N_535,In_130,In_283);
nand U536 (N_536,In_286,In_157);
and U537 (N_537,In_11,In_414);
and U538 (N_538,In_201,In_250);
and U539 (N_539,In_101,In_171);
nand U540 (N_540,In_219,In_203);
and U541 (N_541,In_39,In_136);
and U542 (N_542,In_394,In_369);
nor U543 (N_543,In_297,In_258);
or U544 (N_544,In_218,In_213);
nand U545 (N_545,In_451,In_421);
or U546 (N_546,In_315,In_443);
or U547 (N_547,In_22,In_102);
or U548 (N_548,In_251,In_339);
and U549 (N_549,In_360,In_100);
and U550 (N_550,In_46,In_497);
or U551 (N_551,In_316,In_172);
nor U552 (N_552,In_110,In_412);
nand U553 (N_553,In_67,In_338);
nor U554 (N_554,In_304,In_137);
or U555 (N_555,In_353,In_118);
or U556 (N_556,In_176,In_96);
nor U557 (N_557,In_337,In_313);
or U558 (N_558,In_154,In_384);
nor U559 (N_559,In_264,In_295);
nand U560 (N_560,In_281,In_295);
nor U561 (N_561,In_256,In_225);
and U562 (N_562,In_165,In_146);
nor U563 (N_563,In_453,In_425);
or U564 (N_564,In_85,In_424);
nand U565 (N_565,In_146,In_443);
and U566 (N_566,In_279,In_165);
nor U567 (N_567,In_332,In_18);
nor U568 (N_568,In_422,In_156);
and U569 (N_569,In_476,In_361);
nand U570 (N_570,In_420,In_176);
and U571 (N_571,In_59,In_192);
or U572 (N_572,In_343,In_342);
nor U573 (N_573,In_339,In_121);
nor U574 (N_574,In_193,In_153);
nand U575 (N_575,In_94,In_411);
and U576 (N_576,In_33,In_452);
nor U577 (N_577,In_285,In_478);
or U578 (N_578,In_230,In_60);
nand U579 (N_579,In_456,In_401);
nand U580 (N_580,In_41,In_125);
or U581 (N_581,In_67,In_18);
nor U582 (N_582,In_488,In_72);
or U583 (N_583,In_248,In_184);
and U584 (N_584,In_152,In_335);
nor U585 (N_585,In_11,In_399);
or U586 (N_586,In_75,In_210);
nand U587 (N_587,In_453,In_12);
and U588 (N_588,In_279,In_151);
nor U589 (N_589,In_167,In_39);
or U590 (N_590,In_161,In_201);
nand U591 (N_591,In_430,In_94);
or U592 (N_592,In_347,In_213);
or U593 (N_593,In_177,In_213);
and U594 (N_594,In_256,In_240);
nand U595 (N_595,In_192,In_49);
nor U596 (N_596,In_338,In_256);
and U597 (N_597,In_441,In_447);
and U598 (N_598,In_434,In_293);
nand U599 (N_599,In_136,In_99);
and U600 (N_600,N_391,N_88);
nand U601 (N_601,N_148,N_465);
or U602 (N_602,N_228,N_274);
nand U603 (N_603,N_389,N_255);
and U604 (N_604,N_76,N_422);
nor U605 (N_605,N_382,N_435);
and U606 (N_606,N_183,N_512);
or U607 (N_607,N_226,N_533);
nand U608 (N_608,N_262,N_544);
nor U609 (N_609,N_19,N_338);
nor U610 (N_610,N_361,N_251);
nor U611 (N_611,N_116,N_588);
or U612 (N_612,N_252,N_46);
and U613 (N_613,N_464,N_28);
nand U614 (N_614,N_488,N_161);
nor U615 (N_615,N_453,N_528);
xor U616 (N_616,N_295,N_296);
or U617 (N_617,N_253,N_147);
xnor U618 (N_618,N_135,N_16);
and U619 (N_619,N_366,N_142);
nor U620 (N_620,N_564,N_312);
nor U621 (N_621,N_530,N_188);
and U622 (N_622,N_98,N_423);
nand U623 (N_623,N_534,N_95);
and U624 (N_624,N_106,N_208);
nor U625 (N_625,N_586,N_129);
and U626 (N_626,N_200,N_470);
and U627 (N_627,N_47,N_196);
nand U628 (N_628,N_75,N_340);
or U629 (N_629,N_539,N_450);
or U630 (N_630,N_568,N_314);
nor U631 (N_631,N_258,N_431);
and U632 (N_632,N_25,N_275);
or U633 (N_633,N_288,N_5);
nor U634 (N_634,N_364,N_91);
or U635 (N_635,N_572,N_466);
nor U636 (N_636,N_21,N_43);
nor U637 (N_637,N_59,N_281);
and U638 (N_638,N_357,N_204);
and U639 (N_639,N_407,N_497);
nand U640 (N_640,N_526,N_119);
nand U641 (N_641,N_158,N_137);
or U642 (N_642,N_176,N_42);
or U643 (N_643,N_362,N_334);
and U644 (N_644,N_273,N_136);
and U645 (N_645,N_233,N_493);
nand U646 (N_646,N_324,N_489);
nor U647 (N_647,N_220,N_92);
or U648 (N_648,N_579,N_311);
or U649 (N_649,N_294,N_202);
nand U650 (N_650,N_229,N_261);
and U651 (N_651,N_557,N_399);
nand U652 (N_652,N_452,N_286);
or U653 (N_653,N_303,N_521);
and U654 (N_654,N_553,N_484);
and U655 (N_655,N_440,N_141);
nand U656 (N_656,N_309,N_12);
and U657 (N_657,N_214,N_112);
nand U658 (N_658,N_83,N_426);
and U659 (N_659,N_160,N_90);
and U660 (N_660,N_495,N_175);
or U661 (N_661,N_498,N_271);
nand U662 (N_662,N_0,N_87);
and U663 (N_663,N_344,N_9);
and U664 (N_664,N_561,N_577);
and U665 (N_665,N_367,N_241);
nand U666 (N_666,N_406,N_347);
and U667 (N_667,N_243,N_118);
or U668 (N_668,N_545,N_245);
xnor U669 (N_669,N_173,N_123);
and U670 (N_670,N_581,N_172);
and U671 (N_671,N_380,N_52);
or U672 (N_672,N_86,N_502);
xor U673 (N_673,N_235,N_201);
and U674 (N_674,N_384,N_72);
nor U675 (N_675,N_506,N_523);
and U676 (N_676,N_349,N_33);
nand U677 (N_677,N_479,N_491);
and U678 (N_678,N_571,N_218);
or U679 (N_679,N_4,N_240);
nor U680 (N_680,N_400,N_205);
or U681 (N_681,N_266,N_532);
nor U682 (N_682,N_313,N_556);
or U683 (N_683,N_103,N_215);
and U684 (N_684,N_331,N_584);
nor U685 (N_685,N_414,N_327);
and U686 (N_686,N_394,N_50);
nor U687 (N_687,N_385,N_336);
nand U688 (N_688,N_69,N_429);
or U689 (N_689,N_569,N_78);
nor U690 (N_690,N_140,N_131);
or U691 (N_691,N_476,N_443);
nor U692 (N_692,N_139,N_93);
nor U693 (N_693,N_471,N_174);
or U694 (N_694,N_287,N_146);
or U695 (N_695,N_437,N_89);
xor U696 (N_696,N_594,N_449);
nand U697 (N_697,N_24,N_531);
nand U698 (N_698,N_345,N_84);
nor U699 (N_699,N_456,N_388);
nor U700 (N_700,N_31,N_254);
nand U701 (N_701,N_291,N_583);
nor U702 (N_702,N_282,N_335);
or U703 (N_703,N_97,N_510);
or U704 (N_704,N_66,N_224);
nand U705 (N_705,N_150,N_515);
nor U706 (N_706,N_15,N_328);
nand U707 (N_707,N_513,N_580);
nor U708 (N_708,N_591,N_138);
and U709 (N_709,N_166,N_297);
or U710 (N_710,N_58,N_427);
or U711 (N_711,N_494,N_540);
and U712 (N_712,N_430,N_8);
nor U713 (N_713,N_80,N_153);
nand U714 (N_714,N_375,N_82);
and U715 (N_715,N_249,N_403);
and U716 (N_716,N_96,N_321);
nand U717 (N_717,N_216,N_487);
or U718 (N_718,N_325,N_246);
and U719 (N_719,N_3,N_565);
nor U720 (N_720,N_458,N_469);
nor U721 (N_721,N_221,N_451);
or U722 (N_722,N_223,N_276);
or U723 (N_723,N_289,N_317);
nor U724 (N_724,N_468,N_193);
nand U725 (N_725,N_219,N_270);
and U726 (N_726,N_596,N_593);
or U727 (N_727,N_298,N_222);
or U728 (N_728,N_597,N_197);
nand U729 (N_729,N_555,N_390);
nand U730 (N_730,N_34,N_501);
and U731 (N_731,N_121,N_272);
and U732 (N_732,N_169,N_381);
nand U733 (N_733,N_283,N_17);
nor U734 (N_734,N_575,N_191);
nor U735 (N_735,N_529,N_104);
and U736 (N_736,N_401,N_444);
or U737 (N_737,N_448,N_304);
nor U738 (N_738,N_524,N_373);
nor U739 (N_739,N_459,N_419);
nor U740 (N_740,N_306,N_307);
nor U741 (N_741,N_333,N_549);
and U742 (N_742,N_117,N_370);
nand U743 (N_743,N_144,N_473);
xor U744 (N_744,N_590,N_463);
nand U745 (N_745,N_111,N_411);
or U746 (N_746,N_360,N_554);
nand U747 (N_747,N_499,N_32);
or U748 (N_748,N_29,N_64);
or U749 (N_749,N_238,N_165);
or U750 (N_750,N_192,N_18);
or U751 (N_751,N_374,N_280);
and U752 (N_752,N_301,N_461);
nor U753 (N_753,N_27,N_23);
xor U754 (N_754,N_424,N_14);
nor U755 (N_755,N_536,N_70);
nor U756 (N_756,N_396,N_212);
nand U757 (N_757,N_578,N_170);
and U758 (N_758,N_481,N_413);
and U759 (N_759,N_355,N_30);
and U760 (N_760,N_35,N_81);
nand U761 (N_761,N_329,N_439);
nand U762 (N_762,N_386,N_154);
or U763 (N_763,N_559,N_483);
and U764 (N_764,N_363,N_163);
and U765 (N_765,N_299,N_482);
nand U766 (N_766,N_421,N_376);
xnor U767 (N_767,N_207,N_548);
and U768 (N_768,N_518,N_38);
or U769 (N_769,N_124,N_108);
nor U770 (N_770,N_412,N_113);
nor U771 (N_771,N_567,N_293);
nand U772 (N_772,N_351,N_284);
or U773 (N_773,N_36,N_213);
nor U774 (N_774,N_560,N_558);
or U775 (N_775,N_457,N_178);
and U776 (N_776,N_500,N_589);
nor U777 (N_777,N_26,N_592);
or U778 (N_778,N_41,N_542);
nand U779 (N_779,N_190,N_65);
nor U780 (N_780,N_210,N_408);
nor U781 (N_781,N_441,N_496);
nand U782 (N_782,N_315,N_405);
nand U783 (N_783,N_45,N_455);
or U784 (N_784,N_551,N_356);
nor U785 (N_785,N_79,N_341);
xnor U786 (N_786,N_425,N_199);
nand U787 (N_787,N_134,N_447);
nor U788 (N_788,N_547,N_475);
nand U789 (N_789,N_109,N_257);
or U790 (N_790,N_263,N_132);
and U791 (N_791,N_420,N_326);
and U792 (N_792,N_445,N_102);
nor U793 (N_793,N_48,N_478);
and U794 (N_794,N_209,N_53);
nand U795 (N_795,N_320,N_377);
or U796 (N_796,N_392,N_181);
xnor U797 (N_797,N_11,N_342);
and U798 (N_798,N_267,N_179);
and U799 (N_799,N_231,N_265);
nor U800 (N_800,N_62,N_516);
and U801 (N_801,N_279,N_250);
nand U802 (N_802,N_120,N_285);
nor U803 (N_803,N_462,N_107);
and U804 (N_804,N_114,N_162);
or U805 (N_805,N_509,N_187);
and U806 (N_806,N_387,N_379);
and U807 (N_807,N_352,N_348);
and U808 (N_808,N_77,N_305);
nor U809 (N_809,N_101,N_39);
nor U810 (N_810,N_74,N_230);
and U811 (N_811,N_346,N_247);
nand U812 (N_812,N_490,N_63);
nand U813 (N_813,N_159,N_13);
nor U814 (N_814,N_55,N_156);
nor U815 (N_815,N_599,N_308);
nor U816 (N_816,N_508,N_51);
and U817 (N_817,N_177,N_402);
nor U818 (N_818,N_598,N_264);
or U819 (N_819,N_268,N_409);
nor U820 (N_820,N_474,N_480);
or U821 (N_821,N_353,N_7);
nor U822 (N_822,N_507,N_185);
or U823 (N_823,N_168,N_527);
nand U824 (N_824,N_383,N_573);
or U825 (N_825,N_505,N_511);
and U826 (N_826,N_432,N_189);
nor U827 (N_827,N_60,N_57);
nand U828 (N_828,N_73,N_37);
nand U829 (N_829,N_541,N_472);
or U830 (N_830,N_446,N_186);
and U831 (N_831,N_368,N_359);
or U832 (N_832,N_492,N_167);
nand U833 (N_833,N_467,N_416);
and U834 (N_834,N_203,N_85);
nor U835 (N_835,N_486,N_155);
nand U836 (N_836,N_126,N_316);
nor U837 (N_837,N_587,N_369);
or U838 (N_838,N_40,N_180);
or U839 (N_839,N_239,N_550);
and U840 (N_840,N_438,N_256);
nand U841 (N_841,N_485,N_418);
or U842 (N_842,N_145,N_514);
or U843 (N_843,N_595,N_71);
or U844 (N_844,N_22,N_519);
nor U845 (N_845,N_225,N_94);
xnor U846 (N_846,N_54,N_503);
nor U847 (N_847,N_290,N_152);
and U848 (N_848,N_227,N_99);
and U849 (N_849,N_417,N_198);
and U850 (N_850,N_397,N_127);
nand U851 (N_851,N_322,N_566);
and U852 (N_852,N_151,N_194);
nor U853 (N_853,N_522,N_436);
or U854 (N_854,N_277,N_350);
nand U855 (N_855,N_323,N_582);
nand U856 (N_856,N_410,N_105);
nand U857 (N_857,N_20,N_393);
nand U858 (N_858,N_454,N_130);
and U859 (N_859,N_211,N_570);
and U860 (N_860,N_337,N_100);
and U861 (N_861,N_68,N_576);
nand U862 (N_862,N_477,N_260);
or U863 (N_863,N_182,N_259);
nand U864 (N_864,N_56,N_110);
or U865 (N_865,N_244,N_504);
or U866 (N_866,N_61,N_563);
nand U867 (N_867,N_115,N_10);
nand U868 (N_868,N_44,N_434);
or U869 (N_869,N_237,N_310);
nand U870 (N_870,N_433,N_195);
and U871 (N_871,N_537,N_242);
and U872 (N_872,N_122,N_354);
and U873 (N_873,N_538,N_269);
nand U874 (N_874,N_535,N_171);
and U875 (N_875,N_206,N_143);
nand U876 (N_876,N_460,N_1);
or U877 (N_877,N_428,N_552);
nor U878 (N_878,N_292,N_343);
or U879 (N_879,N_232,N_184);
nand U880 (N_880,N_330,N_157);
nand U881 (N_881,N_149,N_164);
and U882 (N_882,N_395,N_372);
and U883 (N_883,N_248,N_415);
nor U884 (N_884,N_442,N_234);
nand U885 (N_885,N_358,N_546);
or U886 (N_886,N_2,N_525);
nor U887 (N_887,N_128,N_133);
or U888 (N_888,N_404,N_236);
xnor U889 (N_889,N_543,N_398);
nor U890 (N_890,N_339,N_300);
nand U891 (N_891,N_562,N_6);
or U892 (N_892,N_302,N_371);
or U893 (N_893,N_217,N_278);
nor U894 (N_894,N_378,N_574);
nor U895 (N_895,N_585,N_319);
or U896 (N_896,N_318,N_517);
nand U897 (N_897,N_125,N_332);
xor U898 (N_898,N_365,N_67);
nor U899 (N_899,N_520,N_49);
and U900 (N_900,N_254,N_93);
nand U901 (N_901,N_255,N_282);
or U902 (N_902,N_147,N_262);
nor U903 (N_903,N_366,N_90);
nand U904 (N_904,N_346,N_165);
nand U905 (N_905,N_292,N_13);
nor U906 (N_906,N_115,N_348);
nor U907 (N_907,N_553,N_44);
nor U908 (N_908,N_69,N_383);
and U909 (N_909,N_241,N_86);
nand U910 (N_910,N_221,N_438);
nor U911 (N_911,N_538,N_285);
nand U912 (N_912,N_525,N_240);
nand U913 (N_913,N_297,N_574);
nand U914 (N_914,N_529,N_303);
and U915 (N_915,N_244,N_306);
or U916 (N_916,N_383,N_338);
nand U917 (N_917,N_356,N_591);
nand U918 (N_918,N_332,N_109);
nor U919 (N_919,N_166,N_321);
nor U920 (N_920,N_64,N_140);
nand U921 (N_921,N_59,N_62);
or U922 (N_922,N_408,N_205);
nand U923 (N_923,N_471,N_271);
or U924 (N_924,N_356,N_289);
or U925 (N_925,N_112,N_358);
or U926 (N_926,N_154,N_39);
and U927 (N_927,N_432,N_503);
nand U928 (N_928,N_402,N_162);
nand U929 (N_929,N_323,N_307);
nor U930 (N_930,N_20,N_486);
or U931 (N_931,N_33,N_485);
nor U932 (N_932,N_503,N_546);
and U933 (N_933,N_536,N_157);
and U934 (N_934,N_337,N_549);
nor U935 (N_935,N_152,N_574);
and U936 (N_936,N_208,N_327);
nor U937 (N_937,N_561,N_31);
or U938 (N_938,N_202,N_577);
nand U939 (N_939,N_157,N_306);
nand U940 (N_940,N_279,N_258);
or U941 (N_941,N_208,N_337);
nand U942 (N_942,N_391,N_144);
or U943 (N_943,N_351,N_73);
nand U944 (N_944,N_392,N_434);
and U945 (N_945,N_378,N_209);
or U946 (N_946,N_213,N_166);
nor U947 (N_947,N_442,N_444);
or U948 (N_948,N_573,N_369);
nand U949 (N_949,N_165,N_567);
and U950 (N_950,N_406,N_576);
and U951 (N_951,N_355,N_135);
nor U952 (N_952,N_174,N_240);
nand U953 (N_953,N_478,N_417);
or U954 (N_954,N_531,N_499);
or U955 (N_955,N_230,N_176);
and U956 (N_956,N_233,N_258);
nor U957 (N_957,N_523,N_473);
nor U958 (N_958,N_478,N_570);
or U959 (N_959,N_194,N_206);
and U960 (N_960,N_276,N_465);
or U961 (N_961,N_277,N_206);
and U962 (N_962,N_138,N_379);
nor U963 (N_963,N_485,N_19);
and U964 (N_964,N_539,N_83);
nand U965 (N_965,N_381,N_489);
nand U966 (N_966,N_595,N_557);
nand U967 (N_967,N_389,N_535);
nand U968 (N_968,N_149,N_81);
and U969 (N_969,N_294,N_240);
and U970 (N_970,N_514,N_482);
nor U971 (N_971,N_18,N_340);
or U972 (N_972,N_128,N_555);
or U973 (N_973,N_290,N_82);
or U974 (N_974,N_491,N_486);
nor U975 (N_975,N_414,N_502);
nor U976 (N_976,N_141,N_68);
or U977 (N_977,N_6,N_571);
nor U978 (N_978,N_41,N_2);
and U979 (N_979,N_521,N_240);
nor U980 (N_980,N_586,N_521);
or U981 (N_981,N_597,N_68);
and U982 (N_982,N_393,N_583);
or U983 (N_983,N_23,N_216);
nor U984 (N_984,N_130,N_358);
nor U985 (N_985,N_235,N_316);
and U986 (N_986,N_297,N_200);
nor U987 (N_987,N_449,N_439);
nand U988 (N_988,N_516,N_523);
nand U989 (N_989,N_502,N_369);
nor U990 (N_990,N_89,N_263);
nand U991 (N_991,N_84,N_132);
and U992 (N_992,N_1,N_263);
nor U993 (N_993,N_45,N_269);
and U994 (N_994,N_125,N_145);
and U995 (N_995,N_256,N_177);
and U996 (N_996,N_452,N_132);
nand U997 (N_997,N_23,N_439);
nor U998 (N_998,N_96,N_472);
nand U999 (N_999,N_106,N_68);
nor U1000 (N_1000,N_525,N_250);
nor U1001 (N_1001,N_433,N_521);
nand U1002 (N_1002,N_494,N_372);
nor U1003 (N_1003,N_4,N_17);
or U1004 (N_1004,N_274,N_336);
nor U1005 (N_1005,N_58,N_252);
and U1006 (N_1006,N_467,N_536);
nor U1007 (N_1007,N_7,N_479);
and U1008 (N_1008,N_248,N_530);
nor U1009 (N_1009,N_258,N_123);
and U1010 (N_1010,N_443,N_307);
or U1011 (N_1011,N_325,N_156);
or U1012 (N_1012,N_334,N_124);
and U1013 (N_1013,N_348,N_511);
or U1014 (N_1014,N_535,N_258);
or U1015 (N_1015,N_440,N_469);
and U1016 (N_1016,N_470,N_359);
and U1017 (N_1017,N_173,N_434);
and U1018 (N_1018,N_523,N_340);
or U1019 (N_1019,N_259,N_513);
nor U1020 (N_1020,N_166,N_232);
nor U1021 (N_1021,N_480,N_519);
nand U1022 (N_1022,N_242,N_573);
or U1023 (N_1023,N_359,N_7);
nand U1024 (N_1024,N_73,N_278);
nor U1025 (N_1025,N_173,N_393);
and U1026 (N_1026,N_486,N_268);
and U1027 (N_1027,N_77,N_248);
or U1028 (N_1028,N_248,N_403);
nand U1029 (N_1029,N_311,N_146);
nand U1030 (N_1030,N_225,N_136);
or U1031 (N_1031,N_487,N_592);
nand U1032 (N_1032,N_122,N_504);
or U1033 (N_1033,N_167,N_422);
and U1034 (N_1034,N_510,N_426);
nand U1035 (N_1035,N_542,N_402);
and U1036 (N_1036,N_448,N_297);
xnor U1037 (N_1037,N_243,N_417);
xor U1038 (N_1038,N_578,N_139);
or U1039 (N_1039,N_284,N_593);
nor U1040 (N_1040,N_77,N_117);
nand U1041 (N_1041,N_401,N_318);
nor U1042 (N_1042,N_517,N_497);
or U1043 (N_1043,N_178,N_115);
and U1044 (N_1044,N_536,N_537);
nor U1045 (N_1045,N_115,N_492);
nand U1046 (N_1046,N_555,N_376);
or U1047 (N_1047,N_249,N_44);
nor U1048 (N_1048,N_407,N_189);
nand U1049 (N_1049,N_68,N_545);
and U1050 (N_1050,N_200,N_400);
nand U1051 (N_1051,N_35,N_128);
nand U1052 (N_1052,N_472,N_64);
and U1053 (N_1053,N_336,N_511);
nand U1054 (N_1054,N_69,N_474);
or U1055 (N_1055,N_169,N_366);
or U1056 (N_1056,N_517,N_84);
and U1057 (N_1057,N_462,N_464);
nor U1058 (N_1058,N_379,N_221);
nor U1059 (N_1059,N_437,N_189);
or U1060 (N_1060,N_290,N_50);
and U1061 (N_1061,N_521,N_428);
and U1062 (N_1062,N_381,N_101);
nor U1063 (N_1063,N_476,N_342);
nor U1064 (N_1064,N_148,N_213);
or U1065 (N_1065,N_533,N_276);
or U1066 (N_1066,N_418,N_202);
nand U1067 (N_1067,N_400,N_357);
nor U1068 (N_1068,N_229,N_128);
nor U1069 (N_1069,N_65,N_512);
nor U1070 (N_1070,N_277,N_177);
nand U1071 (N_1071,N_428,N_562);
or U1072 (N_1072,N_179,N_145);
nor U1073 (N_1073,N_554,N_371);
nor U1074 (N_1074,N_458,N_238);
nor U1075 (N_1075,N_19,N_501);
or U1076 (N_1076,N_487,N_252);
or U1077 (N_1077,N_441,N_545);
nand U1078 (N_1078,N_242,N_570);
and U1079 (N_1079,N_499,N_3);
nor U1080 (N_1080,N_19,N_5);
nand U1081 (N_1081,N_23,N_344);
nand U1082 (N_1082,N_34,N_420);
and U1083 (N_1083,N_189,N_255);
or U1084 (N_1084,N_516,N_478);
or U1085 (N_1085,N_41,N_288);
nor U1086 (N_1086,N_412,N_523);
and U1087 (N_1087,N_2,N_560);
nor U1088 (N_1088,N_385,N_229);
xnor U1089 (N_1089,N_563,N_456);
nand U1090 (N_1090,N_598,N_195);
nand U1091 (N_1091,N_403,N_444);
and U1092 (N_1092,N_425,N_45);
and U1093 (N_1093,N_192,N_153);
and U1094 (N_1094,N_130,N_463);
xnor U1095 (N_1095,N_419,N_24);
nor U1096 (N_1096,N_292,N_515);
or U1097 (N_1097,N_558,N_374);
and U1098 (N_1098,N_6,N_108);
or U1099 (N_1099,N_268,N_215);
and U1100 (N_1100,N_439,N_324);
and U1101 (N_1101,N_30,N_104);
and U1102 (N_1102,N_182,N_459);
or U1103 (N_1103,N_127,N_129);
nand U1104 (N_1104,N_0,N_27);
and U1105 (N_1105,N_360,N_220);
nand U1106 (N_1106,N_535,N_521);
nor U1107 (N_1107,N_88,N_119);
nand U1108 (N_1108,N_492,N_76);
xnor U1109 (N_1109,N_33,N_36);
and U1110 (N_1110,N_538,N_137);
or U1111 (N_1111,N_598,N_367);
xor U1112 (N_1112,N_490,N_575);
nand U1113 (N_1113,N_316,N_582);
nand U1114 (N_1114,N_341,N_590);
and U1115 (N_1115,N_292,N_481);
nor U1116 (N_1116,N_494,N_453);
and U1117 (N_1117,N_156,N_353);
nand U1118 (N_1118,N_404,N_31);
or U1119 (N_1119,N_357,N_207);
nor U1120 (N_1120,N_414,N_528);
nor U1121 (N_1121,N_88,N_170);
nor U1122 (N_1122,N_521,N_402);
or U1123 (N_1123,N_229,N_498);
or U1124 (N_1124,N_411,N_267);
or U1125 (N_1125,N_586,N_277);
or U1126 (N_1126,N_224,N_457);
nand U1127 (N_1127,N_458,N_439);
nand U1128 (N_1128,N_106,N_217);
nand U1129 (N_1129,N_265,N_309);
nand U1130 (N_1130,N_191,N_66);
nor U1131 (N_1131,N_289,N_117);
nor U1132 (N_1132,N_143,N_98);
and U1133 (N_1133,N_445,N_414);
or U1134 (N_1134,N_233,N_554);
nor U1135 (N_1135,N_386,N_42);
or U1136 (N_1136,N_571,N_365);
or U1137 (N_1137,N_209,N_273);
or U1138 (N_1138,N_395,N_354);
nand U1139 (N_1139,N_160,N_536);
or U1140 (N_1140,N_451,N_454);
and U1141 (N_1141,N_437,N_481);
and U1142 (N_1142,N_526,N_491);
or U1143 (N_1143,N_480,N_555);
and U1144 (N_1144,N_245,N_241);
nor U1145 (N_1145,N_404,N_12);
nand U1146 (N_1146,N_359,N_399);
nand U1147 (N_1147,N_67,N_125);
or U1148 (N_1148,N_524,N_212);
or U1149 (N_1149,N_173,N_314);
or U1150 (N_1150,N_424,N_400);
nor U1151 (N_1151,N_40,N_412);
nor U1152 (N_1152,N_459,N_70);
xor U1153 (N_1153,N_340,N_192);
and U1154 (N_1154,N_420,N_283);
or U1155 (N_1155,N_569,N_240);
nor U1156 (N_1156,N_214,N_453);
or U1157 (N_1157,N_421,N_574);
xnor U1158 (N_1158,N_246,N_394);
or U1159 (N_1159,N_407,N_452);
or U1160 (N_1160,N_134,N_301);
or U1161 (N_1161,N_275,N_385);
nand U1162 (N_1162,N_499,N_349);
xnor U1163 (N_1163,N_530,N_136);
nor U1164 (N_1164,N_427,N_337);
and U1165 (N_1165,N_137,N_344);
or U1166 (N_1166,N_423,N_569);
nor U1167 (N_1167,N_382,N_113);
and U1168 (N_1168,N_129,N_471);
and U1169 (N_1169,N_112,N_49);
or U1170 (N_1170,N_336,N_376);
nand U1171 (N_1171,N_72,N_187);
nor U1172 (N_1172,N_580,N_571);
and U1173 (N_1173,N_320,N_2);
nand U1174 (N_1174,N_161,N_578);
nand U1175 (N_1175,N_397,N_357);
nand U1176 (N_1176,N_5,N_176);
nand U1177 (N_1177,N_5,N_230);
or U1178 (N_1178,N_12,N_202);
xnor U1179 (N_1179,N_489,N_105);
and U1180 (N_1180,N_464,N_26);
and U1181 (N_1181,N_229,N_505);
and U1182 (N_1182,N_172,N_551);
nor U1183 (N_1183,N_22,N_455);
nand U1184 (N_1184,N_188,N_173);
or U1185 (N_1185,N_10,N_448);
nor U1186 (N_1186,N_21,N_576);
nand U1187 (N_1187,N_593,N_142);
and U1188 (N_1188,N_71,N_242);
nand U1189 (N_1189,N_356,N_147);
and U1190 (N_1190,N_223,N_107);
or U1191 (N_1191,N_449,N_327);
or U1192 (N_1192,N_589,N_478);
nand U1193 (N_1193,N_551,N_28);
nor U1194 (N_1194,N_404,N_390);
or U1195 (N_1195,N_65,N_270);
and U1196 (N_1196,N_220,N_484);
or U1197 (N_1197,N_486,N_433);
nor U1198 (N_1198,N_99,N_48);
and U1199 (N_1199,N_294,N_360);
or U1200 (N_1200,N_965,N_815);
nor U1201 (N_1201,N_671,N_963);
nand U1202 (N_1202,N_690,N_983);
nor U1203 (N_1203,N_634,N_972);
nor U1204 (N_1204,N_1078,N_1030);
or U1205 (N_1205,N_1086,N_862);
or U1206 (N_1206,N_982,N_1008);
or U1207 (N_1207,N_603,N_1193);
or U1208 (N_1208,N_947,N_922);
nor U1209 (N_1209,N_1142,N_713);
and U1210 (N_1210,N_1091,N_707);
or U1211 (N_1211,N_863,N_886);
and U1212 (N_1212,N_1129,N_1100);
nor U1213 (N_1213,N_724,N_996);
nor U1214 (N_1214,N_741,N_1034);
and U1215 (N_1215,N_788,N_1109);
and U1216 (N_1216,N_643,N_1052);
nand U1217 (N_1217,N_1164,N_638);
or U1218 (N_1218,N_926,N_934);
nor U1219 (N_1219,N_608,N_1069);
or U1220 (N_1220,N_743,N_892);
nor U1221 (N_1221,N_925,N_1158);
nor U1222 (N_1222,N_870,N_842);
and U1223 (N_1223,N_785,N_930);
nand U1224 (N_1224,N_1122,N_903);
or U1225 (N_1225,N_916,N_826);
nor U1226 (N_1226,N_1197,N_878);
nand U1227 (N_1227,N_1110,N_1098);
xor U1228 (N_1228,N_637,N_1104);
and U1229 (N_1229,N_631,N_894);
nor U1230 (N_1230,N_795,N_1181);
or U1231 (N_1231,N_890,N_1134);
nor U1232 (N_1232,N_844,N_812);
and U1233 (N_1233,N_951,N_921);
nor U1234 (N_1234,N_917,N_1066);
nand U1235 (N_1235,N_619,N_821);
xnor U1236 (N_1236,N_1171,N_754);
nand U1237 (N_1237,N_617,N_1195);
and U1238 (N_1238,N_1155,N_918);
nand U1239 (N_1239,N_685,N_1165);
nor U1240 (N_1240,N_764,N_755);
or U1241 (N_1241,N_1126,N_672);
and U1242 (N_1242,N_860,N_745);
or U1243 (N_1243,N_796,N_611);
nor U1244 (N_1244,N_704,N_871);
or U1245 (N_1245,N_1114,N_865);
and U1246 (N_1246,N_737,N_1071);
nand U1247 (N_1247,N_661,N_718);
nand U1248 (N_1248,N_630,N_1037);
nor U1249 (N_1249,N_760,N_1138);
and U1250 (N_1250,N_825,N_1137);
nor U1251 (N_1251,N_786,N_993);
or U1252 (N_1252,N_1026,N_907);
nor U1253 (N_1253,N_877,N_893);
nand U1254 (N_1254,N_1160,N_1179);
nor U1255 (N_1255,N_872,N_1081);
nand U1256 (N_1256,N_814,N_1196);
and U1257 (N_1257,N_984,N_942);
nand U1258 (N_1258,N_652,N_1152);
nand U1259 (N_1259,N_901,N_905);
and U1260 (N_1260,N_615,N_771);
nor U1261 (N_1261,N_882,N_1186);
nand U1262 (N_1262,N_935,N_1185);
and U1263 (N_1263,N_977,N_888);
nor U1264 (N_1264,N_1143,N_1075);
or U1265 (N_1265,N_950,N_750);
nand U1266 (N_1266,N_807,N_884);
or U1267 (N_1267,N_1106,N_902);
nor U1268 (N_1268,N_1020,N_656);
nor U1269 (N_1269,N_1059,N_1116);
and U1270 (N_1270,N_727,N_775);
and U1271 (N_1271,N_1121,N_753);
nand U1272 (N_1272,N_885,N_797);
nand U1273 (N_1273,N_1191,N_846);
or U1274 (N_1274,N_911,N_610);
and U1275 (N_1275,N_845,N_1079);
or U1276 (N_1276,N_1035,N_747);
or U1277 (N_1277,N_999,N_667);
nor U1278 (N_1278,N_1127,N_662);
nand U1279 (N_1279,N_1042,N_809);
or U1280 (N_1280,N_1159,N_959);
nor U1281 (N_1281,N_974,N_1057);
or U1282 (N_1282,N_1172,N_910);
nor U1283 (N_1283,N_783,N_698);
nor U1284 (N_1284,N_699,N_990);
nand U1285 (N_1285,N_723,N_820);
nand U1286 (N_1286,N_876,N_997);
or U1287 (N_1287,N_1007,N_1088);
and U1288 (N_1288,N_1157,N_988);
nand U1289 (N_1289,N_980,N_614);
nor U1290 (N_1290,N_1173,N_879);
nand U1291 (N_1291,N_1107,N_1199);
nor U1292 (N_1292,N_883,N_691);
or U1293 (N_1293,N_1182,N_1189);
nor U1294 (N_1294,N_602,N_897);
nand U1295 (N_1295,N_726,N_835);
nand U1296 (N_1296,N_714,N_734);
and U1297 (N_1297,N_696,N_1183);
nand U1298 (N_1298,N_1187,N_819);
nor U1299 (N_1299,N_843,N_1025);
or U1300 (N_1300,N_712,N_855);
nand U1301 (N_1301,N_1174,N_735);
and U1302 (N_1302,N_1154,N_861);
nand U1303 (N_1303,N_952,N_640);
or U1304 (N_1304,N_1064,N_1198);
or U1305 (N_1305,N_981,N_841);
nor U1306 (N_1306,N_1130,N_649);
and U1307 (N_1307,N_1004,N_628);
and U1308 (N_1308,N_937,N_818);
and U1309 (N_1309,N_1175,N_1153);
nand U1310 (N_1310,N_1060,N_765);
or U1311 (N_1311,N_1169,N_677);
nand U1312 (N_1312,N_1067,N_1039);
nand U1313 (N_1313,N_1013,N_898);
nand U1314 (N_1314,N_927,N_957);
nor U1315 (N_1315,N_1128,N_979);
and U1316 (N_1316,N_995,N_1150);
or U1317 (N_1317,N_768,N_659);
or U1318 (N_1318,N_1046,N_684);
and U1319 (N_1319,N_683,N_978);
nor U1320 (N_1320,N_940,N_1047);
nand U1321 (N_1321,N_848,N_1053);
nand U1322 (N_1322,N_728,N_1135);
or U1323 (N_1323,N_742,N_609);
and U1324 (N_1324,N_645,N_773);
and U1325 (N_1325,N_960,N_715);
nand U1326 (N_1326,N_1001,N_618);
nor U1327 (N_1327,N_675,N_1036);
nand U1328 (N_1328,N_1003,N_1024);
or U1329 (N_1329,N_964,N_782);
nor U1330 (N_1330,N_1119,N_1076);
or U1331 (N_1331,N_1056,N_808);
nor U1332 (N_1332,N_829,N_868);
or U1333 (N_1333,N_1123,N_1167);
and U1334 (N_1334,N_1054,N_1084);
nor U1335 (N_1335,N_772,N_881);
nand U1336 (N_1336,N_804,N_654);
and U1337 (N_1337,N_1015,N_1031);
and U1338 (N_1338,N_607,N_866);
or U1339 (N_1339,N_900,N_823);
or U1340 (N_1340,N_650,N_1090);
nor U1341 (N_1341,N_899,N_803);
or U1342 (N_1342,N_949,N_1111);
nor U1343 (N_1343,N_904,N_1012);
nor U1344 (N_1344,N_732,N_1062);
or U1345 (N_1345,N_817,N_802);
nor U1346 (N_1346,N_780,N_604);
or U1347 (N_1347,N_1161,N_998);
nor U1348 (N_1348,N_941,N_717);
nand U1349 (N_1349,N_931,N_1168);
and U1350 (N_1350,N_669,N_668);
nand U1351 (N_1351,N_635,N_740);
nand U1352 (N_1352,N_1192,N_1027);
xnor U1353 (N_1353,N_858,N_853);
nor U1354 (N_1354,N_621,N_721);
and U1355 (N_1355,N_1023,N_1040);
nor U1356 (N_1356,N_1096,N_830);
nor U1357 (N_1357,N_1074,N_1101);
nand U1358 (N_1358,N_970,N_1103);
and U1359 (N_1359,N_763,N_1132);
nand U1360 (N_1360,N_624,N_851);
nor U1361 (N_1361,N_1041,N_1068);
and U1362 (N_1362,N_1148,N_1140);
nor U1363 (N_1363,N_874,N_961);
nor U1364 (N_1364,N_697,N_757);
and U1365 (N_1365,N_620,N_962);
nor U1366 (N_1366,N_1021,N_692);
nor U1367 (N_1367,N_653,N_613);
nor U1368 (N_1368,N_798,N_847);
nor U1369 (N_1369,N_822,N_806);
nand U1370 (N_1370,N_1010,N_1108);
xnor U1371 (N_1371,N_1093,N_1124);
or U1372 (N_1372,N_1188,N_923);
nor U1373 (N_1373,N_738,N_801);
nand U1374 (N_1374,N_836,N_840);
and U1375 (N_1375,N_873,N_777);
xor U1376 (N_1376,N_695,N_1097);
and U1377 (N_1377,N_946,N_1184);
and U1378 (N_1378,N_639,N_733);
or U1379 (N_1379,N_1151,N_766);
nor U1380 (N_1380,N_1120,N_762);
nor U1381 (N_1381,N_767,N_790);
nor U1382 (N_1382,N_1028,N_626);
or U1383 (N_1383,N_973,N_939);
nor U1384 (N_1384,N_1022,N_1011);
nor U1385 (N_1385,N_800,N_730);
and U1386 (N_1386,N_708,N_693);
or U1387 (N_1387,N_936,N_784);
nand U1388 (N_1388,N_682,N_1115);
or U1389 (N_1389,N_1016,N_799);
and U1390 (N_1390,N_1087,N_739);
nor U1391 (N_1391,N_1080,N_811);
xor U1392 (N_1392,N_670,N_810);
and U1393 (N_1393,N_864,N_1070);
nand U1394 (N_1394,N_1018,N_954);
nand U1395 (N_1395,N_1145,N_913);
or U1396 (N_1396,N_657,N_945);
and U1397 (N_1397,N_636,N_759);
nor U1398 (N_1398,N_1147,N_932);
or U1399 (N_1399,N_716,N_729);
nor U1400 (N_1400,N_834,N_666);
and U1401 (N_1401,N_1063,N_1065);
nor U1402 (N_1402,N_1149,N_1029);
or U1403 (N_1403,N_748,N_781);
and U1404 (N_1404,N_1156,N_968);
nor U1405 (N_1405,N_1058,N_709);
or U1406 (N_1406,N_686,N_612);
and U1407 (N_1407,N_673,N_1072);
and U1408 (N_1408,N_856,N_687);
nor U1409 (N_1409,N_967,N_720);
or U1410 (N_1410,N_605,N_1141);
and U1411 (N_1411,N_665,N_679);
nand U1412 (N_1412,N_616,N_1032);
nand U1413 (N_1413,N_1082,N_924);
nor U1414 (N_1414,N_601,N_1006);
and U1415 (N_1415,N_641,N_1073);
and U1416 (N_1416,N_906,N_909);
nand U1417 (N_1417,N_956,N_889);
and U1418 (N_1418,N_688,N_761);
nor U1419 (N_1419,N_646,N_1009);
nand U1420 (N_1420,N_1089,N_867);
nor U1421 (N_1421,N_1092,N_663);
nor U1422 (N_1422,N_1125,N_756);
nor U1423 (N_1423,N_792,N_938);
nand U1424 (N_1424,N_655,N_1050);
nor U1425 (N_1425,N_600,N_794);
nand U1426 (N_1426,N_629,N_651);
or U1427 (N_1427,N_703,N_1146);
or U1428 (N_1428,N_770,N_778);
nand U1429 (N_1429,N_1014,N_895);
xnor U1430 (N_1430,N_625,N_1112);
and U1431 (N_1431,N_948,N_1133);
nor U1432 (N_1432,N_1043,N_816);
nor U1433 (N_1433,N_791,N_664);
nand U1434 (N_1434,N_658,N_660);
nand U1435 (N_1435,N_1083,N_746);
nor U1436 (N_1436,N_1131,N_986);
nand U1437 (N_1437,N_700,N_680);
or U1438 (N_1438,N_1044,N_838);
or U1439 (N_1439,N_985,N_966);
nand U1440 (N_1440,N_701,N_955);
and U1441 (N_1441,N_944,N_1055);
or U1442 (N_1442,N_1144,N_1095);
nor U1443 (N_1443,N_920,N_776);
or U1444 (N_1444,N_914,N_831);
nor U1445 (N_1445,N_793,N_919);
nor U1446 (N_1446,N_779,N_1000);
nand U1447 (N_1447,N_1163,N_1176);
or U1448 (N_1448,N_749,N_1113);
nand U1449 (N_1449,N_674,N_854);
or U1450 (N_1450,N_606,N_1139);
nor U1451 (N_1451,N_832,N_805);
and U1452 (N_1452,N_719,N_1178);
and U1453 (N_1453,N_850,N_722);
or U1454 (N_1454,N_989,N_1019);
or U1455 (N_1455,N_689,N_828);
xor U1456 (N_1456,N_642,N_1085);
and U1457 (N_1457,N_702,N_1005);
or U1458 (N_1458,N_987,N_929);
nand U1459 (N_1459,N_839,N_647);
nand U1460 (N_1460,N_676,N_1180);
and U1461 (N_1461,N_908,N_1002);
or U1462 (N_1462,N_789,N_678);
or U1463 (N_1463,N_694,N_1166);
and U1464 (N_1464,N_1077,N_632);
nand U1465 (N_1465,N_975,N_1048);
or U1466 (N_1466,N_943,N_852);
nor U1467 (N_1467,N_976,N_928);
nor U1468 (N_1468,N_1117,N_725);
or U1469 (N_1469,N_1102,N_622);
nand U1470 (N_1470,N_958,N_681);
and U1471 (N_1471,N_623,N_992);
or U1472 (N_1472,N_751,N_1038);
or U1473 (N_1473,N_833,N_1194);
and U1474 (N_1474,N_859,N_711);
nand U1475 (N_1475,N_837,N_758);
nor U1476 (N_1476,N_1049,N_824);
nor U1477 (N_1477,N_1099,N_1017);
and U1478 (N_1478,N_969,N_857);
nor U1479 (N_1479,N_849,N_1170);
nand U1480 (N_1480,N_971,N_869);
or U1481 (N_1481,N_991,N_710);
nor U1482 (N_1482,N_953,N_627);
and U1483 (N_1483,N_731,N_736);
and U1484 (N_1484,N_1045,N_752);
nand U1485 (N_1485,N_912,N_880);
or U1486 (N_1486,N_891,N_1118);
or U1487 (N_1487,N_705,N_706);
nor U1488 (N_1488,N_774,N_1094);
nand U1489 (N_1489,N_787,N_994);
nor U1490 (N_1490,N_744,N_933);
and U1491 (N_1491,N_1105,N_644);
nand U1492 (N_1492,N_1061,N_1177);
nor U1493 (N_1493,N_875,N_1051);
nor U1494 (N_1494,N_1136,N_813);
or U1495 (N_1495,N_648,N_1190);
nor U1496 (N_1496,N_827,N_896);
nand U1497 (N_1497,N_1033,N_887);
nand U1498 (N_1498,N_633,N_769);
nand U1499 (N_1499,N_915,N_1162);
and U1500 (N_1500,N_748,N_734);
or U1501 (N_1501,N_1140,N_659);
nor U1502 (N_1502,N_1091,N_796);
nor U1503 (N_1503,N_724,N_888);
nor U1504 (N_1504,N_986,N_956);
nor U1505 (N_1505,N_1190,N_1004);
or U1506 (N_1506,N_651,N_647);
nand U1507 (N_1507,N_1199,N_736);
nor U1508 (N_1508,N_1189,N_778);
and U1509 (N_1509,N_726,N_1094);
nand U1510 (N_1510,N_719,N_779);
and U1511 (N_1511,N_907,N_1196);
nor U1512 (N_1512,N_815,N_672);
nor U1513 (N_1513,N_955,N_1039);
and U1514 (N_1514,N_884,N_1050);
and U1515 (N_1515,N_766,N_1139);
nand U1516 (N_1516,N_750,N_1179);
nand U1517 (N_1517,N_753,N_1064);
nor U1518 (N_1518,N_930,N_922);
nor U1519 (N_1519,N_958,N_995);
or U1520 (N_1520,N_647,N_851);
and U1521 (N_1521,N_717,N_847);
nor U1522 (N_1522,N_682,N_1051);
or U1523 (N_1523,N_1160,N_968);
or U1524 (N_1524,N_1026,N_888);
xor U1525 (N_1525,N_1054,N_739);
nor U1526 (N_1526,N_1079,N_963);
and U1527 (N_1527,N_774,N_1110);
nor U1528 (N_1528,N_1025,N_1000);
and U1529 (N_1529,N_1125,N_1139);
nand U1530 (N_1530,N_987,N_1146);
nand U1531 (N_1531,N_808,N_960);
and U1532 (N_1532,N_1152,N_714);
nand U1533 (N_1533,N_789,N_628);
or U1534 (N_1534,N_957,N_922);
and U1535 (N_1535,N_739,N_952);
nor U1536 (N_1536,N_1117,N_624);
nor U1537 (N_1537,N_895,N_870);
xnor U1538 (N_1538,N_1121,N_945);
or U1539 (N_1539,N_924,N_805);
nor U1540 (N_1540,N_1062,N_950);
or U1541 (N_1541,N_1163,N_785);
xnor U1542 (N_1542,N_960,N_730);
nor U1543 (N_1543,N_791,N_981);
or U1544 (N_1544,N_1125,N_1022);
or U1545 (N_1545,N_853,N_868);
or U1546 (N_1546,N_1086,N_1074);
or U1547 (N_1547,N_964,N_745);
and U1548 (N_1548,N_900,N_749);
or U1549 (N_1549,N_790,N_1024);
nand U1550 (N_1550,N_986,N_1180);
xnor U1551 (N_1551,N_1046,N_743);
or U1552 (N_1552,N_1015,N_899);
nor U1553 (N_1553,N_801,N_1046);
nand U1554 (N_1554,N_616,N_1052);
or U1555 (N_1555,N_1190,N_809);
nor U1556 (N_1556,N_688,N_874);
and U1557 (N_1557,N_674,N_1087);
nand U1558 (N_1558,N_877,N_965);
nand U1559 (N_1559,N_783,N_694);
nor U1560 (N_1560,N_667,N_1102);
nor U1561 (N_1561,N_1101,N_608);
or U1562 (N_1562,N_790,N_891);
and U1563 (N_1563,N_894,N_745);
nand U1564 (N_1564,N_1066,N_1113);
nor U1565 (N_1565,N_904,N_1178);
nor U1566 (N_1566,N_1011,N_1157);
nand U1567 (N_1567,N_768,N_729);
nand U1568 (N_1568,N_621,N_821);
or U1569 (N_1569,N_915,N_765);
or U1570 (N_1570,N_712,N_875);
and U1571 (N_1571,N_721,N_649);
nor U1572 (N_1572,N_1061,N_1168);
nor U1573 (N_1573,N_883,N_604);
or U1574 (N_1574,N_1129,N_1136);
or U1575 (N_1575,N_693,N_617);
or U1576 (N_1576,N_1053,N_732);
nor U1577 (N_1577,N_657,N_775);
nor U1578 (N_1578,N_619,N_789);
nor U1579 (N_1579,N_635,N_902);
or U1580 (N_1580,N_758,N_951);
nand U1581 (N_1581,N_779,N_628);
nand U1582 (N_1582,N_800,N_1071);
and U1583 (N_1583,N_924,N_933);
nor U1584 (N_1584,N_666,N_698);
xor U1585 (N_1585,N_881,N_836);
nand U1586 (N_1586,N_632,N_975);
and U1587 (N_1587,N_800,N_1026);
or U1588 (N_1588,N_904,N_844);
or U1589 (N_1589,N_1156,N_1128);
nand U1590 (N_1590,N_1173,N_952);
nor U1591 (N_1591,N_1162,N_1159);
nand U1592 (N_1592,N_819,N_870);
and U1593 (N_1593,N_834,N_616);
or U1594 (N_1594,N_1184,N_739);
and U1595 (N_1595,N_1062,N_997);
nor U1596 (N_1596,N_1168,N_909);
or U1597 (N_1597,N_770,N_1135);
and U1598 (N_1598,N_1026,N_661);
and U1599 (N_1599,N_714,N_1062);
or U1600 (N_1600,N_670,N_1143);
or U1601 (N_1601,N_705,N_640);
and U1602 (N_1602,N_805,N_647);
and U1603 (N_1603,N_1024,N_1058);
nor U1604 (N_1604,N_1154,N_982);
and U1605 (N_1605,N_772,N_1198);
or U1606 (N_1606,N_1068,N_763);
nand U1607 (N_1607,N_714,N_1068);
and U1608 (N_1608,N_622,N_814);
nand U1609 (N_1609,N_807,N_618);
or U1610 (N_1610,N_716,N_708);
nor U1611 (N_1611,N_1029,N_1046);
or U1612 (N_1612,N_998,N_752);
or U1613 (N_1613,N_789,N_998);
or U1614 (N_1614,N_980,N_1099);
and U1615 (N_1615,N_1017,N_1133);
or U1616 (N_1616,N_798,N_685);
and U1617 (N_1617,N_768,N_644);
nand U1618 (N_1618,N_1078,N_691);
nor U1619 (N_1619,N_742,N_999);
and U1620 (N_1620,N_732,N_1148);
nor U1621 (N_1621,N_719,N_926);
nor U1622 (N_1622,N_748,N_886);
or U1623 (N_1623,N_1084,N_1130);
xnor U1624 (N_1624,N_721,N_1004);
nand U1625 (N_1625,N_974,N_1004);
nand U1626 (N_1626,N_719,N_1029);
nand U1627 (N_1627,N_723,N_754);
nor U1628 (N_1628,N_1050,N_1192);
and U1629 (N_1629,N_1047,N_618);
or U1630 (N_1630,N_1106,N_661);
nand U1631 (N_1631,N_1121,N_904);
nand U1632 (N_1632,N_853,N_758);
and U1633 (N_1633,N_1108,N_660);
and U1634 (N_1634,N_821,N_725);
xnor U1635 (N_1635,N_600,N_1124);
or U1636 (N_1636,N_1168,N_830);
nor U1637 (N_1637,N_883,N_611);
or U1638 (N_1638,N_891,N_1000);
or U1639 (N_1639,N_943,N_823);
nand U1640 (N_1640,N_1087,N_812);
xor U1641 (N_1641,N_1199,N_765);
nor U1642 (N_1642,N_685,N_674);
nand U1643 (N_1643,N_1023,N_870);
nand U1644 (N_1644,N_933,N_671);
and U1645 (N_1645,N_872,N_829);
and U1646 (N_1646,N_770,N_1172);
and U1647 (N_1647,N_935,N_1133);
and U1648 (N_1648,N_701,N_887);
or U1649 (N_1649,N_665,N_699);
or U1650 (N_1650,N_794,N_1040);
or U1651 (N_1651,N_896,N_826);
or U1652 (N_1652,N_620,N_1002);
nor U1653 (N_1653,N_678,N_1018);
nand U1654 (N_1654,N_1147,N_679);
or U1655 (N_1655,N_723,N_600);
nor U1656 (N_1656,N_655,N_1162);
or U1657 (N_1657,N_1045,N_953);
and U1658 (N_1658,N_976,N_962);
nor U1659 (N_1659,N_790,N_759);
nand U1660 (N_1660,N_639,N_1008);
nand U1661 (N_1661,N_1164,N_878);
xnor U1662 (N_1662,N_1199,N_710);
nor U1663 (N_1663,N_680,N_769);
and U1664 (N_1664,N_861,N_710);
and U1665 (N_1665,N_814,N_1070);
nand U1666 (N_1666,N_682,N_755);
or U1667 (N_1667,N_907,N_1151);
nand U1668 (N_1668,N_629,N_1147);
nand U1669 (N_1669,N_1144,N_1010);
nand U1670 (N_1670,N_667,N_962);
nor U1671 (N_1671,N_1125,N_943);
and U1672 (N_1672,N_821,N_1013);
nor U1673 (N_1673,N_856,N_1045);
and U1674 (N_1674,N_1019,N_837);
and U1675 (N_1675,N_781,N_953);
nor U1676 (N_1676,N_741,N_725);
xor U1677 (N_1677,N_782,N_914);
nand U1678 (N_1678,N_1046,N_843);
and U1679 (N_1679,N_1160,N_764);
nor U1680 (N_1680,N_1150,N_775);
xor U1681 (N_1681,N_1027,N_750);
or U1682 (N_1682,N_1042,N_1031);
or U1683 (N_1683,N_690,N_727);
nand U1684 (N_1684,N_937,N_601);
and U1685 (N_1685,N_892,N_943);
and U1686 (N_1686,N_1034,N_1063);
nor U1687 (N_1687,N_884,N_785);
nor U1688 (N_1688,N_1183,N_1079);
or U1689 (N_1689,N_780,N_710);
or U1690 (N_1690,N_1015,N_1020);
nand U1691 (N_1691,N_632,N_723);
nand U1692 (N_1692,N_652,N_891);
nand U1693 (N_1693,N_674,N_747);
nand U1694 (N_1694,N_892,N_975);
nand U1695 (N_1695,N_849,N_933);
or U1696 (N_1696,N_667,N_713);
or U1697 (N_1697,N_1155,N_805);
nor U1698 (N_1698,N_1186,N_1158);
or U1699 (N_1699,N_746,N_1111);
nand U1700 (N_1700,N_1063,N_1188);
or U1701 (N_1701,N_846,N_643);
nor U1702 (N_1702,N_961,N_771);
and U1703 (N_1703,N_905,N_768);
and U1704 (N_1704,N_1131,N_905);
nand U1705 (N_1705,N_626,N_981);
or U1706 (N_1706,N_954,N_1146);
nand U1707 (N_1707,N_1037,N_659);
xor U1708 (N_1708,N_1121,N_1104);
and U1709 (N_1709,N_706,N_893);
nor U1710 (N_1710,N_863,N_644);
and U1711 (N_1711,N_1042,N_832);
or U1712 (N_1712,N_622,N_980);
nand U1713 (N_1713,N_669,N_876);
or U1714 (N_1714,N_936,N_901);
nand U1715 (N_1715,N_1129,N_627);
nand U1716 (N_1716,N_1080,N_1048);
nand U1717 (N_1717,N_877,N_1156);
and U1718 (N_1718,N_732,N_626);
or U1719 (N_1719,N_725,N_954);
and U1720 (N_1720,N_1178,N_911);
or U1721 (N_1721,N_647,N_879);
or U1722 (N_1722,N_829,N_779);
nor U1723 (N_1723,N_1145,N_1180);
nand U1724 (N_1724,N_628,N_1108);
or U1725 (N_1725,N_870,N_973);
or U1726 (N_1726,N_840,N_868);
or U1727 (N_1727,N_936,N_975);
or U1728 (N_1728,N_1144,N_648);
or U1729 (N_1729,N_1055,N_1069);
nand U1730 (N_1730,N_693,N_989);
nor U1731 (N_1731,N_869,N_740);
nor U1732 (N_1732,N_759,N_675);
or U1733 (N_1733,N_1151,N_1111);
nand U1734 (N_1734,N_788,N_1094);
nor U1735 (N_1735,N_1039,N_1016);
and U1736 (N_1736,N_1045,N_728);
nor U1737 (N_1737,N_807,N_916);
nor U1738 (N_1738,N_875,N_658);
nand U1739 (N_1739,N_684,N_993);
or U1740 (N_1740,N_1152,N_853);
nor U1741 (N_1741,N_1148,N_710);
nor U1742 (N_1742,N_726,N_1157);
or U1743 (N_1743,N_674,N_1178);
or U1744 (N_1744,N_635,N_727);
or U1745 (N_1745,N_782,N_1055);
nor U1746 (N_1746,N_685,N_1075);
and U1747 (N_1747,N_1059,N_794);
or U1748 (N_1748,N_1178,N_829);
nand U1749 (N_1749,N_1018,N_1187);
nand U1750 (N_1750,N_830,N_615);
nor U1751 (N_1751,N_688,N_973);
nor U1752 (N_1752,N_649,N_631);
or U1753 (N_1753,N_958,N_658);
and U1754 (N_1754,N_762,N_1141);
and U1755 (N_1755,N_1123,N_680);
nand U1756 (N_1756,N_722,N_1143);
nor U1757 (N_1757,N_792,N_1011);
nand U1758 (N_1758,N_816,N_622);
and U1759 (N_1759,N_1101,N_765);
nand U1760 (N_1760,N_731,N_613);
nand U1761 (N_1761,N_886,N_852);
and U1762 (N_1762,N_1138,N_996);
or U1763 (N_1763,N_624,N_636);
nand U1764 (N_1764,N_639,N_1104);
nor U1765 (N_1765,N_935,N_1069);
nor U1766 (N_1766,N_699,N_1011);
or U1767 (N_1767,N_808,N_838);
nor U1768 (N_1768,N_936,N_1192);
nor U1769 (N_1769,N_1045,N_797);
nor U1770 (N_1770,N_1145,N_1138);
nand U1771 (N_1771,N_816,N_964);
or U1772 (N_1772,N_1081,N_1018);
or U1773 (N_1773,N_1096,N_706);
and U1774 (N_1774,N_1131,N_987);
or U1775 (N_1775,N_729,N_1008);
nand U1776 (N_1776,N_1167,N_952);
nand U1777 (N_1777,N_935,N_987);
nand U1778 (N_1778,N_790,N_749);
nand U1779 (N_1779,N_641,N_659);
or U1780 (N_1780,N_605,N_718);
or U1781 (N_1781,N_770,N_1025);
and U1782 (N_1782,N_748,N_918);
or U1783 (N_1783,N_1172,N_870);
nand U1784 (N_1784,N_639,N_991);
and U1785 (N_1785,N_834,N_1007);
and U1786 (N_1786,N_786,N_968);
nor U1787 (N_1787,N_654,N_936);
nor U1788 (N_1788,N_1008,N_813);
or U1789 (N_1789,N_1169,N_890);
xnor U1790 (N_1790,N_665,N_1013);
nor U1791 (N_1791,N_806,N_1049);
nand U1792 (N_1792,N_1008,N_1137);
nor U1793 (N_1793,N_852,N_1182);
nor U1794 (N_1794,N_1008,N_948);
nand U1795 (N_1795,N_1154,N_994);
and U1796 (N_1796,N_712,N_704);
nor U1797 (N_1797,N_984,N_872);
and U1798 (N_1798,N_911,N_830);
or U1799 (N_1799,N_1194,N_1003);
nor U1800 (N_1800,N_1304,N_1515);
or U1801 (N_1801,N_1337,N_1480);
or U1802 (N_1802,N_1421,N_1722);
nor U1803 (N_1803,N_1547,N_1615);
or U1804 (N_1804,N_1567,N_1368);
and U1805 (N_1805,N_1593,N_1591);
nand U1806 (N_1806,N_1339,N_1393);
nor U1807 (N_1807,N_1281,N_1796);
nand U1808 (N_1808,N_1469,N_1303);
nand U1809 (N_1809,N_1442,N_1579);
nand U1810 (N_1810,N_1344,N_1295);
nand U1811 (N_1811,N_1521,N_1320);
nor U1812 (N_1812,N_1632,N_1355);
nand U1813 (N_1813,N_1730,N_1535);
nor U1814 (N_1814,N_1504,N_1653);
nand U1815 (N_1815,N_1500,N_1331);
nor U1816 (N_1816,N_1416,N_1525);
and U1817 (N_1817,N_1392,N_1422);
nor U1818 (N_1818,N_1738,N_1540);
or U1819 (N_1819,N_1300,N_1353);
and U1820 (N_1820,N_1232,N_1340);
and U1821 (N_1821,N_1265,N_1296);
nor U1822 (N_1822,N_1670,N_1621);
and U1823 (N_1823,N_1214,N_1276);
nor U1824 (N_1824,N_1267,N_1542);
xnor U1825 (N_1825,N_1473,N_1305);
nand U1826 (N_1826,N_1466,N_1546);
nand U1827 (N_1827,N_1586,N_1465);
and U1828 (N_1828,N_1260,N_1585);
nor U1829 (N_1829,N_1543,N_1612);
xor U1830 (N_1830,N_1629,N_1693);
or U1831 (N_1831,N_1522,N_1576);
nand U1832 (N_1832,N_1666,N_1775);
or U1833 (N_1833,N_1335,N_1311);
nor U1834 (N_1834,N_1204,N_1222);
and U1835 (N_1835,N_1258,N_1205);
and U1836 (N_1836,N_1408,N_1397);
nor U1837 (N_1837,N_1657,N_1380);
or U1838 (N_1838,N_1507,N_1505);
and U1839 (N_1839,N_1484,N_1235);
or U1840 (N_1840,N_1414,N_1766);
nor U1841 (N_1841,N_1524,N_1789);
nor U1842 (N_1842,N_1782,N_1274);
nor U1843 (N_1843,N_1487,N_1423);
nor U1844 (N_1844,N_1566,N_1695);
and U1845 (N_1845,N_1644,N_1426);
and U1846 (N_1846,N_1491,N_1602);
nor U1847 (N_1847,N_1709,N_1213);
and U1848 (N_1848,N_1681,N_1209);
and U1849 (N_1849,N_1747,N_1312);
nor U1850 (N_1850,N_1432,N_1221);
or U1851 (N_1851,N_1288,N_1248);
and U1852 (N_1852,N_1669,N_1269);
or U1853 (N_1853,N_1479,N_1429);
and U1854 (N_1854,N_1379,N_1637);
and U1855 (N_1855,N_1529,N_1253);
nor U1856 (N_1856,N_1278,N_1697);
nand U1857 (N_1857,N_1779,N_1444);
or U1858 (N_1858,N_1490,N_1301);
and U1859 (N_1859,N_1528,N_1275);
nor U1860 (N_1860,N_1388,N_1233);
and U1861 (N_1861,N_1715,N_1351);
nor U1862 (N_1862,N_1562,N_1451);
nor U1863 (N_1863,N_1284,N_1461);
nor U1864 (N_1864,N_1742,N_1406);
nor U1865 (N_1865,N_1718,N_1571);
or U1866 (N_1866,N_1506,N_1783);
or U1867 (N_1867,N_1371,N_1623);
and U1868 (N_1868,N_1446,N_1272);
or U1869 (N_1869,N_1399,N_1625);
xor U1870 (N_1870,N_1329,N_1592);
or U1871 (N_1871,N_1707,N_1332);
or U1872 (N_1872,N_1552,N_1387);
nor U1873 (N_1873,N_1494,N_1780);
and U1874 (N_1874,N_1223,N_1383);
nor U1875 (N_1875,N_1264,N_1784);
or U1876 (N_1876,N_1425,N_1785);
and U1877 (N_1877,N_1293,N_1533);
nor U1878 (N_1878,N_1765,N_1658);
nand U1879 (N_1879,N_1440,N_1729);
and U1880 (N_1880,N_1651,N_1268);
or U1881 (N_1881,N_1532,N_1362);
nand U1882 (N_1882,N_1788,N_1659);
nand U1883 (N_1883,N_1514,N_1714);
and U1884 (N_1884,N_1476,N_1231);
or U1885 (N_1885,N_1472,N_1550);
nand U1886 (N_1886,N_1431,N_1776);
or U1887 (N_1887,N_1676,N_1726);
xnor U1888 (N_1888,N_1672,N_1492);
nand U1889 (N_1889,N_1212,N_1544);
and U1890 (N_1890,N_1460,N_1698);
or U1891 (N_1891,N_1445,N_1555);
nand U1892 (N_1892,N_1786,N_1639);
or U1893 (N_1893,N_1563,N_1502);
nand U1894 (N_1894,N_1413,N_1367);
or U1895 (N_1895,N_1321,N_1675);
nand U1896 (N_1896,N_1583,N_1475);
or U1897 (N_1897,N_1554,N_1449);
or U1898 (N_1898,N_1725,N_1510);
nor U1899 (N_1899,N_1370,N_1617);
and U1900 (N_1900,N_1516,N_1758);
and U1901 (N_1901,N_1680,N_1358);
and U1902 (N_1902,N_1298,N_1418);
nand U1903 (N_1903,N_1702,N_1290);
nor U1904 (N_1904,N_1609,N_1503);
xor U1905 (N_1905,N_1318,N_1292);
and U1906 (N_1906,N_1790,N_1673);
nor U1907 (N_1907,N_1727,N_1630);
nand U1908 (N_1908,N_1589,N_1237);
and U1909 (N_1909,N_1316,N_1624);
or U1910 (N_1910,N_1417,N_1671);
nand U1911 (N_1911,N_1508,N_1744);
and U1912 (N_1912,N_1313,N_1220);
or U1913 (N_1913,N_1315,N_1511);
nand U1914 (N_1914,N_1610,N_1463);
or U1915 (N_1915,N_1343,N_1415);
nand U1916 (N_1916,N_1564,N_1336);
nor U1917 (N_1917,N_1603,N_1536);
nor U1918 (N_1918,N_1706,N_1635);
nand U1919 (N_1919,N_1489,N_1330);
or U1920 (N_1920,N_1763,N_1595);
nand U1921 (N_1921,N_1456,N_1654);
nand U1922 (N_1922,N_1403,N_1682);
or U1923 (N_1923,N_1787,N_1636);
xnor U1924 (N_1924,N_1410,N_1338);
nor U1925 (N_1925,N_1211,N_1798);
nor U1926 (N_1926,N_1381,N_1679);
or U1927 (N_1927,N_1495,N_1647);
or U1928 (N_1928,N_1286,N_1369);
nor U1929 (N_1929,N_1247,N_1732);
and U1930 (N_1930,N_1450,N_1478);
or U1931 (N_1931,N_1597,N_1354);
nor U1932 (N_1932,N_1459,N_1750);
and U1933 (N_1933,N_1594,N_1513);
nor U1934 (N_1934,N_1457,N_1447);
or U1935 (N_1935,N_1700,N_1322);
and U1936 (N_1936,N_1745,N_1793);
or U1937 (N_1937,N_1386,N_1759);
and U1938 (N_1938,N_1470,N_1501);
and U1939 (N_1939,N_1225,N_1723);
nor U1940 (N_1940,N_1645,N_1572);
and U1941 (N_1941,N_1349,N_1746);
nor U1942 (N_1942,N_1665,N_1606);
and U1943 (N_1943,N_1259,N_1646);
nand U1944 (N_1944,N_1441,N_1769);
and U1945 (N_1945,N_1662,N_1739);
nor U1946 (N_1946,N_1207,N_1708);
xnor U1947 (N_1947,N_1334,N_1584);
nor U1948 (N_1948,N_1791,N_1748);
or U1949 (N_1949,N_1254,N_1346);
nand U1950 (N_1950,N_1498,N_1217);
nand U1951 (N_1951,N_1438,N_1283);
nand U1952 (N_1952,N_1587,N_1424);
and U1953 (N_1953,N_1310,N_1545);
xor U1954 (N_1954,N_1740,N_1361);
nor U1955 (N_1955,N_1768,N_1620);
nor U1956 (N_1956,N_1716,N_1448);
or U1957 (N_1957,N_1240,N_1282);
and U1958 (N_1958,N_1384,N_1691);
nor U1959 (N_1959,N_1685,N_1777);
and U1960 (N_1960,N_1569,N_1236);
and U1961 (N_1961,N_1711,N_1402);
and U1962 (N_1962,N_1683,N_1356);
or U1963 (N_1963,N_1385,N_1704);
xor U1964 (N_1964,N_1611,N_1694);
nand U1965 (N_1965,N_1266,N_1359);
nor U1966 (N_1966,N_1604,N_1557);
and U1967 (N_1967,N_1720,N_1641);
and U1968 (N_1968,N_1756,N_1795);
or U1969 (N_1969,N_1599,N_1526);
nor U1970 (N_1970,N_1497,N_1434);
and U1971 (N_1971,N_1252,N_1411);
nand U1972 (N_1972,N_1761,N_1216);
nor U1973 (N_1973,N_1622,N_1559);
nor U1974 (N_1974,N_1203,N_1537);
and U1975 (N_1975,N_1664,N_1364);
nor U1976 (N_1976,N_1737,N_1229);
nor U1977 (N_1977,N_1616,N_1674);
nor U1978 (N_1978,N_1781,N_1327);
nor U1979 (N_1979,N_1751,N_1394);
and U1980 (N_1980,N_1660,N_1270);
nor U1981 (N_1981,N_1684,N_1201);
nand U1982 (N_1982,N_1255,N_1430);
or U1983 (N_1983,N_1294,N_1439);
and U1984 (N_1984,N_1243,N_1696);
nand U1985 (N_1985,N_1482,N_1299);
nand U1986 (N_1986,N_1376,N_1578);
nor U1987 (N_1987,N_1226,N_1754);
and U1988 (N_1988,N_1655,N_1558);
or U1989 (N_1989,N_1391,N_1573);
nand U1990 (N_1990,N_1518,N_1519);
and U1991 (N_1991,N_1230,N_1468);
nor U1992 (N_1992,N_1378,N_1712);
nor U1993 (N_1993,N_1208,N_1263);
and U1994 (N_1994,N_1297,N_1347);
nand U1995 (N_1995,N_1633,N_1608);
and U1996 (N_1996,N_1319,N_1360);
nor U1997 (N_1997,N_1256,N_1242);
or U1998 (N_1998,N_1488,N_1582);
nor U1999 (N_1999,N_1549,N_1428);
or U2000 (N_2000,N_1588,N_1462);
nand U2001 (N_2001,N_1333,N_1580);
or U2002 (N_2002,N_1631,N_1435);
and U2003 (N_2003,N_1753,N_1395);
and U2004 (N_2004,N_1607,N_1755);
or U2005 (N_2005,N_1713,N_1250);
xor U2006 (N_2006,N_1251,N_1724);
and U2007 (N_2007,N_1574,N_1496);
nand U2008 (N_2008,N_1643,N_1663);
or U2009 (N_2009,N_1271,N_1794);
or U2010 (N_2010,N_1733,N_1493);
and U2011 (N_2011,N_1734,N_1605);
or U2012 (N_2012,N_1512,N_1570);
nor U2013 (N_2013,N_1443,N_1317);
or U2014 (N_2014,N_1539,N_1757);
and U2015 (N_2015,N_1365,N_1596);
nor U2016 (N_2016,N_1614,N_1499);
or U2017 (N_2017,N_1308,N_1273);
or U2018 (N_2018,N_1771,N_1257);
and U2019 (N_2019,N_1530,N_1531);
nor U2020 (N_2020,N_1731,N_1400);
nor U2021 (N_2021,N_1401,N_1749);
nor U2022 (N_2022,N_1244,N_1736);
and U2023 (N_2023,N_1228,N_1686);
nor U2024 (N_2024,N_1458,N_1390);
or U2025 (N_2025,N_1398,N_1486);
or U2026 (N_2026,N_1467,N_1710);
nand U2027 (N_2027,N_1420,N_1728);
and U2028 (N_2028,N_1452,N_1309);
nor U2029 (N_2029,N_1372,N_1581);
or U2030 (N_2030,N_1561,N_1436);
and U2031 (N_2031,N_1262,N_1455);
nor U2032 (N_2032,N_1404,N_1634);
and U2033 (N_2033,N_1261,N_1743);
xor U2034 (N_2034,N_1481,N_1705);
and U2035 (N_2035,N_1721,N_1289);
nand U2036 (N_2036,N_1453,N_1206);
or U2037 (N_2037,N_1227,N_1419);
and U2038 (N_2038,N_1619,N_1661);
nand U2039 (N_2039,N_1668,N_1363);
and U2040 (N_2040,N_1389,N_1701);
nand U2041 (N_2041,N_1239,N_1677);
nor U2042 (N_2042,N_1433,N_1437);
nand U2043 (N_2043,N_1764,N_1760);
nand U2044 (N_2044,N_1277,N_1210);
or U2045 (N_2045,N_1246,N_1409);
and U2046 (N_2046,N_1534,N_1717);
or U2047 (N_2047,N_1352,N_1314);
nor U2048 (N_2048,N_1373,N_1374);
nor U2049 (N_2049,N_1770,N_1306);
nor U2050 (N_2050,N_1202,N_1454);
and U2051 (N_2051,N_1350,N_1412);
nor U2052 (N_2052,N_1553,N_1649);
or U2053 (N_2053,N_1640,N_1618);
and U2054 (N_2054,N_1326,N_1200);
and U2055 (N_2055,N_1407,N_1735);
and U2056 (N_2056,N_1767,N_1601);
xor U2057 (N_2057,N_1405,N_1541);
or U2058 (N_2058,N_1692,N_1642);
nor U2059 (N_2059,N_1538,N_1678);
or U2060 (N_2060,N_1762,N_1568);
and U2061 (N_2061,N_1628,N_1577);
and U2062 (N_2062,N_1650,N_1772);
nand U2063 (N_2063,N_1377,N_1799);
nor U2064 (N_2064,N_1792,N_1548);
and U2065 (N_2065,N_1638,N_1302);
nor U2066 (N_2066,N_1556,N_1648);
nand U2067 (N_2067,N_1797,N_1427);
or U2068 (N_2068,N_1575,N_1613);
and U2069 (N_2069,N_1241,N_1509);
nand U2070 (N_2070,N_1752,N_1249);
nand U2071 (N_2071,N_1325,N_1652);
or U2072 (N_2072,N_1474,N_1690);
and U2073 (N_2073,N_1345,N_1699);
and U2074 (N_2074,N_1323,N_1719);
nor U2075 (N_2075,N_1285,N_1774);
or U2076 (N_2076,N_1375,N_1600);
nor U2077 (N_2077,N_1689,N_1477);
nor U2078 (N_2078,N_1741,N_1590);
nand U2079 (N_2079,N_1219,N_1627);
nand U2080 (N_2080,N_1342,N_1773);
or U2081 (N_2081,N_1520,N_1626);
and U2082 (N_2082,N_1279,N_1341);
nand U2083 (N_2083,N_1224,N_1517);
or U2084 (N_2084,N_1324,N_1287);
nor U2085 (N_2085,N_1667,N_1560);
nor U2086 (N_2086,N_1703,N_1656);
nand U2087 (N_2087,N_1464,N_1688);
or U2088 (N_2088,N_1396,N_1382);
and U2089 (N_2089,N_1598,N_1328);
nor U2090 (N_2090,N_1238,N_1234);
xnor U2091 (N_2091,N_1280,N_1687);
nor U2092 (N_2092,N_1357,N_1348);
and U2093 (N_2093,N_1565,N_1483);
nand U2094 (N_2094,N_1471,N_1778);
nor U2095 (N_2095,N_1218,N_1551);
xnor U2096 (N_2096,N_1215,N_1523);
nand U2097 (N_2097,N_1245,N_1366);
or U2098 (N_2098,N_1485,N_1527);
nor U2099 (N_2099,N_1291,N_1307);
nor U2100 (N_2100,N_1272,N_1623);
or U2101 (N_2101,N_1494,N_1545);
nand U2102 (N_2102,N_1647,N_1760);
nand U2103 (N_2103,N_1478,N_1511);
nand U2104 (N_2104,N_1436,N_1322);
nor U2105 (N_2105,N_1258,N_1452);
and U2106 (N_2106,N_1749,N_1574);
or U2107 (N_2107,N_1477,N_1514);
and U2108 (N_2108,N_1639,N_1319);
nand U2109 (N_2109,N_1334,N_1351);
or U2110 (N_2110,N_1584,N_1548);
nor U2111 (N_2111,N_1553,N_1358);
nand U2112 (N_2112,N_1404,N_1772);
and U2113 (N_2113,N_1580,N_1278);
and U2114 (N_2114,N_1400,N_1468);
nor U2115 (N_2115,N_1464,N_1488);
or U2116 (N_2116,N_1383,N_1518);
and U2117 (N_2117,N_1209,N_1268);
nor U2118 (N_2118,N_1561,N_1656);
nand U2119 (N_2119,N_1511,N_1679);
nand U2120 (N_2120,N_1718,N_1554);
and U2121 (N_2121,N_1498,N_1403);
nor U2122 (N_2122,N_1411,N_1572);
nand U2123 (N_2123,N_1701,N_1268);
or U2124 (N_2124,N_1738,N_1788);
and U2125 (N_2125,N_1352,N_1484);
and U2126 (N_2126,N_1454,N_1785);
nand U2127 (N_2127,N_1781,N_1590);
nor U2128 (N_2128,N_1373,N_1322);
or U2129 (N_2129,N_1356,N_1634);
and U2130 (N_2130,N_1514,N_1761);
and U2131 (N_2131,N_1786,N_1448);
and U2132 (N_2132,N_1715,N_1298);
nor U2133 (N_2133,N_1344,N_1403);
and U2134 (N_2134,N_1691,N_1749);
nor U2135 (N_2135,N_1662,N_1417);
nand U2136 (N_2136,N_1236,N_1266);
nand U2137 (N_2137,N_1532,N_1584);
or U2138 (N_2138,N_1360,N_1558);
nand U2139 (N_2139,N_1356,N_1281);
nor U2140 (N_2140,N_1287,N_1753);
nor U2141 (N_2141,N_1250,N_1514);
nand U2142 (N_2142,N_1629,N_1460);
or U2143 (N_2143,N_1773,N_1619);
or U2144 (N_2144,N_1351,N_1283);
or U2145 (N_2145,N_1494,N_1235);
nand U2146 (N_2146,N_1264,N_1566);
nand U2147 (N_2147,N_1633,N_1220);
or U2148 (N_2148,N_1568,N_1316);
or U2149 (N_2149,N_1689,N_1582);
and U2150 (N_2150,N_1341,N_1702);
or U2151 (N_2151,N_1766,N_1265);
and U2152 (N_2152,N_1599,N_1453);
nor U2153 (N_2153,N_1243,N_1405);
and U2154 (N_2154,N_1376,N_1288);
and U2155 (N_2155,N_1572,N_1579);
nor U2156 (N_2156,N_1688,N_1546);
or U2157 (N_2157,N_1384,N_1696);
nor U2158 (N_2158,N_1268,N_1670);
nor U2159 (N_2159,N_1638,N_1623);
or U2160 (N_2160,N_1566,N_1731);
and U2161 (N_2161,N_1664,N_1383);
or U2162 (N_2162,N_1291,N_1797);
and U2163 (N_2163,N_1608,N_1509);
nor U2164 (N_2164,N_1614,N_1403);
nor U2165 (N_2165,N_1446,N_1250);
nor U2166 (N_2166,N_1768,N_1305);
or U2167 (N_2167,N_1347,N_1352);
nor U2168 (N_2168,N_1634,N_1548);
or U2169 (N_2169,N_1565,N_1488);
nand U2170 (N_2170,N_1606,N_1733);
nor U2171 (N_2171,N_1317,N_1357);
nand U2172 (N_2172,N_1551,N_1606);
and U2173 (N_2173,N_1295,N_1710);
and U2174 (N_2174,N_1321,N_1722);
nand U2175 (N_2175,N_1692,N_1757);
and U2176 (N_2176,N_1662,N_1692);
nand U2177 (N_2177,N_1615,N_1466);
or U2178 (N_2178,N_1672,N_1651);
nand U2179 (N_2179,N_1225,N_1687);
nand U2180 (N_2180,N_1739,N_1589);
nor U2181 (N_2181,N_1518,N_1536);
nor U2182 (N_2182,N_1332,N_1627);
nand U2183 (N_2183,N_1508,N_1580);
nor U2184 (N_2184,N_1438,N_1771);
nand U2185 (N_2185,N_1275,N_1692);
or U2186 (N_2186,N_1790,N_1203);
xnor U2187 (N_2187,N_1693,N_1475);
nor U2188 (N_2188,N_1463,N_1301);
and U2189 (N_2189,N_1457,N_1571);
nand U2190 (N_2190,N_1799,N_1288);
or U2191 (N_2191,N_1298,N_1505);
and U2192 (N_2192,N_1205,N_1452);
nor U2193 (N_2193,N_1520,N_1214);
nand U2194 (N_2194,N_1629,N_1434);
nor U2195 (N_2195,N_1205,N_1730);
and U2196 (N_2196,N_1328,N_1294);
nand U2197 (N_2197,N_1664,N_1281);
nor U2198 (N_2198,N_1691,N_1587);
and U2199 (N_2199,N_1728,N_1774);
nor U2200 (N_2200,N_1711,N_1536);
nand U2201 (N_2201,N_1394,N_1402);
nor U2202 (N_2202,N_1412,N_1690);
or U2203 (N_2203,N_1429,N_1725);
nand U2204 (N_2204,N_1270,N_1601);
nor U2205 (N_2205,N_1305,N_1781);
nand U2206 (N_2206,N_1408,N_1308);
and U2207 (N_2207,N_1367,N_1226);
or U2208 (N_2208,N_1424,N_1776);
nor U2209 (N_2209,N_1202,N_1262);
nor U2210 (N_2210,N_1367,N_1434);
or U2211 (N_2211,N_1725,N_1478);
and U2212 (N_2212,N_1475,N_1210);
or U2213 (N_2213,N_1333,N_1788);
nand U2214 (N_2214,N_1735,N_1676);
nand U2215 (N_2215,N_1595,N_1551);
and U2216 (N_2216,N_1378,N_1387);
and U2217 (N_2217,N_1380,N_1704);
or U2218 (N_2218,N_1613,N_1563);
or U2219 (N_2219,N_1458,N_1524);
nor U2220 (N_2220,N_1783,N_1266);
nand U2221 (N_2221,N_1431,N_1531);
and U2222 (N_2222,N_1281,N_1698);
nand U2223 (N_2223,N_1766,N_1408);
nand U2224 (N_2224,N_1605,N_1356);
nand U2225 (N_2225,N_1568,N_1269);
nor U2226 (N_2226,N_1412,N_1430);
and U2227 (N_2227,N_1450,N_1576);
nand U2228 (N_2228,N_1400,N_1356);
nand U2229 (N_2229,N_1204,N_1359);
and U2230 (N_2230,N_1266,N_1475);
nor U2231 (N_2231,N_1647,N_1532);
xnor U2232 (N_2232,N_1393,N_1587);
nand U2233 (N_2233,N_1204,N_1424);
nor U2234 (N_2234,N_1505,N_1495);
or U2235 (N_2235,N_1405,N_1482);
nor U2236 (N_2236,N_1517,N_1577);
and U2237 (N_2237,N_1798,N_1401);
nand U2238 (N_2238,N_1691,N_1400);
and U2239 (N_2239,N_1638,N_1393);
and U2240 (N_2240,N_1676,N_1641);
xor U2241 (N_2241,N_1554,N_1461);
nand U2242 (N_2242,N_1384,N_1200);
and U2243 (N_2243,N_1567,N_1751);
nand U2244 (N_2244,N_1500,N_1364);
and U2245 (N_2245,N_1454,N_1609);
or U2246 (N_2246,N_1790,N_1378);
or U2247 (N_2247,N_1715,N_1229);
or U2248 (N_2248,N_1592,N_1632);
nand U2249 (N_2249,N_1273,N_1310);
and U2250 (N_2250,N_1585,N_1515);
nor U2251 (N_2251,N_1616,N_1610);
and U2252 (N_2252,N_1796,N_1351);
nand U2253 (N_2253,N_1658,N_1424);
nand U2254 (N_2254,N_1216,N_1266);
nand U2255 (N_2255,N_1201,N_1218);
nor U2256 (N_2256,N_1455,N_1659);
or U2257 (N_2257,N_1345,N_1245);
or U2258 (N_2258,N_1237,N_1383);
or U2259 (N_2259,N_1682,N_1604);
or U2260 (N_2260,N_1686,N_1218);
and U2261 (N_2261,N_1611,N_1330);
and U2262 (N_2262,N_1677,N_1554);
nand U2263 (N_2263,N_1321,N_1567);
and U2264 (N_2264,N_1637,N_1691);
nand U2265 (N_2265,N_1754,N_1773);
nand U2266 (N_2266,N_1597,N_1447);
or U2267 (N_2267,N_1409,N_1608);
nor U2268 (N_2268,N_1480,N_1375);
and U2269 (N_2269,N_1799,N_1505);
nand U2270 (N_2270,N_1615,N_1541);
xnor U2271 (N_2271,N_1644,N_1710);
or U2272 (N_2272,N_1215,N_1438);
or U2273 (N_2273,N_1219,N_1276);
or U2274 (N_2274,N_1231,N_1246);
nand U2275 (N_2275,N_1478,N_1633);
nor U2276 (N_2276,N_1544,N_1471);
or U2277 (N_2277,N_1756,N_1769);
or U2278 (N_2278,N_1267,N_1706);
and U2279 (N_2279,N_1692,N_1725);
nor U2280 (N_2280,N_1664,N_1460);
or U2281 (N_2281,N_1325,N_1301);
and U2282 (N_2282,N_1225,N_1677);
and U2283 (N_2283,N_1780,N_1469);
nand U2284 (N_2284,N_1450,N_1647);
or U2285 (N_2285,N_1693,N_1593);
and U2286 (N_2286,N_1626,N_1616);
nand U2287 (N_2287,N_1735,N_1470);
nand U2288 (N_2288,N_1676,N_1308);
and U2289 (N_2289,N_1692,N_1412);
or U2290 (N_2290,N_1726,N_1402);
nor U2291 (N_2291,N_1271,N_1777);
and U2292 (N_2292,N_1352,N_1715);
xor U2293 (N_2293,N_1291,N_1521);
or U2294 (N_2294,N_1703,N_1604);
nor U2295 (N_2295,N_1511,N_1651);
nand U2296 (N_2296,N_1620,N_1798);
nand U2297 (N_2297,N_1281,N_1793);
nand U2298 (N_2298,N_1469,N_1683);
or U2299 (N_2299,N_1238,N_1410);
or U2300 (N_2300,N_1302,N_1287);
or U2301 (N_2301,N_1497,N_1455);
or U2302 (N_2302,N_1256,N_1547);
nor U2303 (N_2303,N_1272,N_1569);
and U2304 (N_2304,N_1400,N_1749);
and U2305 (N_2305,N_1413,N_1744);
and U2306 (N_2306,N_1328,N_1339);
and U2307 (N_2307,N_1358,N_1309);
nand U2308 (N_2308,N_1772,N_1204);
nand U2309 (N_2309,N_1346,N_1572);
and U2310 (N_2310,N_1606,N_1796);
or U2311 (N_2311,N_1744,N_1617);
nand U2312 (N_2312,N_1590,N_1514);
nand U2313 (N_2313,N_1445,N_1588);
nor U2314 (N_2314,N_1497,N_1703);
and U2315 (N_2315,N_1504,N_1796);
or U2316 (N_2316,N_1352,N_1501);
nand U2317 (N_2317,N_1304,N_1481);
nand U2318 (N_2318,N_1528,N_1599);
nand U2319 (N_2319,N_1431,N_1299);
nor U2320 (N_2320,N_1680,N_1679);
and U2321 (N_2321,N_1506,N_1306);
and U2322 (N_2322,N_1556,N_1299);
nand U2323 (N_2323,N_1526,N_1586);
nor U2324 (N_2324,N_1518,N_1768);
or U2325 (N_2325,N_1712,N_1501);
nor U2326 (N_2326,N_1603,N_1676);
nor U2327 (N_2327,N_1298,N_1221);
nor U2328 (N_2328,N_1549,N_1554);
nor U2329 (N_2329,N_1484,N_1631);
or U2330 (N_2330,N_1393,N_1788);
or U2331 (N_2331,N_1698,N_1247);
nand U2332 (N_2332,N_1348,N_1349);
and U2333 (N_2333,N_1581,N_1392);
nor U2334 (N_2334,N_1299,N_1589);
and U2335 (N_2335,N_1744,N_1784);
nand U2336 (N_2336,N_1579,N_1530);
nand U2337 (N_2337,N_1332,N_1226);
or U2338 (N_2338,N_1399,N_1659);
xnor U2339 (N_2339,N_1441,N_1572);
and U2340 (N_2340,N_1759,N_1219);
xor U2341 (N_2341,N_1501,N_1255);
nor U2342 (N_2342,N_1251,N_1766);
nor U2343 (N_2343,N_1275,N_1543);
nor U2344 (N_2344,N_1619,N_1417);
nor U2345 (N_2345,N_1666,N_1207);
and U2346 (N_2346,N_1732,N_1735);
nor U2347 (N_2347,N_1535,N_1592);
xor U2348 (N_2348,N_1751,N_1488);
xnor U2349 (N_2349,N_1315,N_1301);
and U2350 (N_2350,N_1679,N_1379);
nor U2351 (N_2351,N_1491,N_1342);
nor U2352 (N_2352,N_1747,N_1750);
nor U2353 (N_2353,N_1749,N_1521);
nand U2354 (N_2354,N_1203,N_1590);
nand U2355 (N_2355,N_1230,N_1673);
nor U2356 (N_2356,N_1442,N_1740);
and U2357 (N_2357,N_1730,N_1635);
nand U2358 (N_2358,N_1624,N_1602);
or U2359 (N_2359,N_1643,N_1337);
or U2360 (N_2360,N_1392,N_1202);
nand U2361 (N_2361,N_1740,N_1222);
nor U2362 (N_2362,N_1646,N_1657);
and U2363 (N_2363,N_1561,N_1539);
or U2364 (N_2364,N_1403,N_1373);
and U2365 (N_2365,N_1453,N_1729);
nor U2366 (N_2366,N_1690,N_1573);
or U2367 (N_2367,N_1634,N_1559);
nand U2368 (N_2368,N_1415,N_1693);
nand U2369 (N_2369,N_1461,N_1678);
and U2370 (N_2370,N_1682,N_1350);
or U2371 (N_2371,N_1527,N_1375);
nand U2372 (N_2372,N_1348,N_1641);
nand U2373 (N_2373,N_1499,N_1262);
xor U2374 (N_2374,N_1532,N_1316);
nor U2375 (N_2375,N_1565,N_1780);
nand U2376 (N_2376,N_1508,N_1251);
nor U2377 (N_2377,N_1318,N_1784);
or U2378 (N_2378,N_1359,N_1757);
nor U2379 (N_2379,N_1788,N_1203);
and U2380 (N_2380,N_1614,N_1760);
nand U2381 (N_2381,N_1603,N_1654);
and U2382 (N_2382,N_1393,N_1711);
nand U2383 (N_2383,N_1508,N_1765);
nand U2384 (N_2384,N_1542,N_1501);
or U2385 (N_2385,N_1324,N_1719);
nor U2386 (N_2386,N_1689,N_1273);
nor U2387 (N_2387,N_1659,N_1648);
and U2388 (N_2388,N_1381,N_1299);
nand U2389 (N_2389,N_1280,N_1402);
nand U2390 (N_2390,N_1437,N_1412);
nand U2391 (N_2391,N_1461,N_1736);
nand U2392 (N_2392,N_1683,N_1715);
or U2393 (N_2393,N_1216,N_1666);
nand U2394 (N_2394,N_1695,N_1706);
nor U2395 (N_2395,N_1765,N_1654);
nor U2396 (N_2396,N_1500,N_1629);
or U2397 (N_2397,N_1647,N_1208);
nor U2398 (N_2398,N_1726,N_1693);
nor U2399 (N_2399,N_1478,N_1593);
nand U2400 (N_2400,N_1893,N_2373);
or U2401 (N_2401,N_2326,N_2266);
nor U2402 (N_2402,N_2301,N_1833);
and U2403 (N_2403,N_1950,N_2319);
nor U2404 (N_2404,N_1851,N_1954);
and U2405 (N_2405,N_2192,N_1968);
nor U2406 (N_2406,N_2377,N_1808);
or U2407 (N_2407,N_2020,N_2360);
and U2408 (N_2408,N_2072,N_2103);
and U2409 (N_2409,N_2245,N_1809);
and U2410 (N_2410,N_2043,N_2311);
nand U2411 (N_2411,N_2285,N_2068);
or U2412 (N_2412,N_1897,N_2287);
and U2413 (N_2413,N_2108,N_2034);
nor U2414 (N_2414,N_2016,N_2293);
or U2415 (N_2415,N_2008,N_1824);
or U2416 (N_2416,N_2084,N_2075);
nor U2417 (N_2417,N_2169,N_2397);
or U2418 (N_2418,N_2310,N_1818);
nand U2419 (N_2419,N_1982,N_1991);
nand U2420 (N_2420,N_2249,N_1821);
nand U2421 (N_2421,N_1877,N_2339);
nand U2422 (N_2422,N_1935,N_1956);
or U2423 (N_2423,N_2231,N_2063);
and U2424 (N_2424,N_1998,N_2296);
and U2425 (N_2425,N_2226,N_1942);
nor U2426 (N_2426,N_2195,N_1858);
or U2427 (N_2427,N_1928,N_2346);
and U2428 (N_2428,N_1911,N_2253);
nand U2429 (N_2429,N_1879,N_1919);
and U2430 (N_2430,N_2205,N_2041);
nor U2431 (N_2431,N_2292,N_2357);
nand U2432 (N_2432,N_2307,N_2269);
nand U2433 (N_2433,N_2222,N_2003);
nor U2434 (N_2434,N_2191,N_2190);
and U2435 (N_2435,N_1841,N_1984);
nor U2436 (N_2436,N_2382,N_2198);
and U2437 (N_2437,N_2267,N_1864);
and U2438 (N_2438,N_1848,N_2188);
nand U2439 (N_2439,N_2265,N_2044);
and U2440 (N_2440,N_1936,N_1921);
nand U2441 (N_2441,N_1817,N_1983);
nand U2442 (N_2442,N_1845,N_1804);
nand U2443 (N_2443,N_1907,N_2129);
nand U2444 (N_2444,N_1957,N_2013);
nand U2445 (N_2445,N_2217,N_1912);
and U2446 (N_2446,N_1898,N_2300);
nand U2447 (N_2447,N_2137,N_2365);
and U2448 (N_2448,N_1924,N_2393);
nor U2449 (N_2449,N_2256,N_2193);
or U2450 (N_2450,N_2141,N_1948);
nand U2451 (N_2451,N_1926,N_1944);
or U2452 (N_2452,N_2240,N_2261);
nor U2453 (N_2453,N_2302,N_2270);
nand U2454 (N_2454,N_2229,N_2381);
nor U2455 (N_2455,N_2209,N_1860);
nor U2456 (N_2456,N_2395,N_2100);
nor U2457 (N_2457,N_1994,N_1806);
nand U2458 (N_2458,N_2160,N_2105);
and U2459 (N_2459,N_1857,N_2203);
or U2460 (N_2460,N_2021,N_2047);
and U2461 (N_2461,N_2180,N_1871);
nor U2462 (N_2462,N_1838,N_2220);
nand U2463 (N_2463,N_2370,N_1902);
or U2464 (N_2464,N_2276,N_2336);
or U2465 (N_2465,N_2278,N_2116);
nor U2466 (N_2466,N_1930,N_1803);
nor U2467 (N_2467,N_2128,N_2046);
and U2468 (N_2468,N_2207,N_2183);
or U2469 (N_2469,N_1843,N_2272);
and U2470 (N_2470,N_2288,N_2102);
nor U2471 (N_2471,N_2051,N_1958);
nand U2472 (N_2472,N_2338,N_2158);
nor U2473 (N_2473,N_2390,N_1829);
and U2474 (N_2474,N_2036,N_1993);
nand U2475 (N_2475,N_2219,N_1888);
nand U2476 (N_2476,N_1955,N_2282);
nor U2477 (N_2477,N_1947,N_2080);
and U2478 (N_2478,N_2242,N_2258);
nor U2479 (N_2479,N_2283,N_1802);
xnor U2480 (N_2480,N_1887,N_2175);
xnor U2481 (N_2481,N_2216,N_2061);
and U2482 (N_2482,N_2074,N_1929);
nor U2483 (N_2483,N_1883,N_1961);
or U2484 (N_2484,N_1977,N_2130);
nand U2485 (N_2485,N_2165,N_1820);
and U2486 (N_2486,N_1856,N_2264);
nor U2487 (N_2487,N_1995,N_2306);
and U2488 (N_2488,N_1932,N_2241);
and U2489 (N_2489,N_2015,N_1884);
nand U2490 (N_2490,N_2082,N_1960);
nor U2491 (N_2491,N_2070,N_2153);
or U2492 (N_2492,N_2095,N_1896);
nor U2493 (N_2493,N_2386,N_1839);
or U2494 (N_2494,N_2383,N_2259);
or U2495 (N_2495,N_2040,N_1966);
nor U2496 (N_2496,N_1816,N_1840);
nand U2497 (N_2497,N_1901,N_2340);
xnor U2498 (N_2498,N_1850,N_2343);
nand U2499 (N_2499,N_2098,N_2056);
nand U2500 (N_2500,N_2014,N_2361);
nand U2501 (N_2501,N_2247,N_2161);
and U2502 (N_2502,N_2274,N_1985);
nor U2503 (N_2503,N_1874,N_2035);
nor U2504 (N_2504,N_2398,N_2384);
or U2505 (N_2505,N_1910,N_2236);
and U2506 (N_2506,N_1801,N_2050);
or U2507 (N_2507,N_2322,N_1959);
and U2508 (N_2508,N_2369,N_2138);
nor U2509 (N_2509,N_2107,N_2054);
xnor U2510 (N_2510,N_2006,N_1825);
or U2511 (N_2511,N_2151,N_2359);
and U2512 (N_2512,N_1952,N_2001);
nor U2513 (N_2513,N_1940,N_2234);
and U2514 (N_2514,N_2115,N_2118);
nor U2515 (N_2515,N_2134,N_1811);
or U2516 (N_2516,N_2064,N_2255);
nand U2517 (N_2517,N_2355,N_1885);
and U2518 (N_2518,N_2168,N_1971);
nand U2519 (N_2519,N_2167,N_2148);
nor U2520 (N_2520,N_2000,N_1873);
nor U2521 (N_2521,N_1867,N_2176);
and U2522 (N_2522,N_1927,N_1831);
and U2523 (N_2523,N_2097,N_2388);
nand U2524 (N_2524,N_2055,N_2092);
or U2525 (N_2525,N_1810,N_2387);
nor U2526 (N_2526,N_1931,N_2351);
nand U2527 (N_2527,N_1844,N_2279);
and U2528 (N_2528,N_2017,N_1836);
and U2529 (N_2529,N_2251,N_2156);
and U2530 (N_2530,N_1909,N_1812);
and U2531 (N_2531,N_2045,N_2335);
nor U2532 (N_2532,N_2225,N_2091);
nor U2533 (N_2533,N_1925,N_1855);
or U2534 (N_2534,N_2121,N_2159);
nor U2535 (N_2535,N_2099,N_2037);
or U2536 (N_2536,N_2132,N_2010);
and U2537 (N_2537,N_2120,N_2111);
and U2538 (N_2538,N_2362,N_1837);
or U2539 (N_2539,N_2083,N_2366);
and U2540 (N_2540,N_1830,N_2039);
and U2541 (N_2541,N_2356,N_1918);
and U2542 (N_2542,N_1964,N_2331);
or U2543 (N_2543,N_2002,N_2350);
or U2544 (N_2544,N_2178,N_2106);
and U2545 (N_2545,N_1875,N_2181);
nand U2546 (N_2546,N_1915,N_2227);
nand U2547 (N_2547,N_2260,N_1807);
or U2548 (N_2548,N_2060,N_1939);
and U2549 (N_2549,N_2009,N_2136);
nand U2550 (N_2550,N_2329,N_2157);
or U2551 (N_2551,N_2076,N_2396);
or U2552 (N_2552,N_2368,N_2312);
and U2553 (N_2553,N_2011,N_1819);
nor U2554 (N_2554,N_2252,N_2170);
or U2555 (N_2555,N_2109,N_1834);
nand U2556 (N_2556,N_2114,N_2349);
and U2557 (N_2557,N_1814,N_2257);
nand U2558 (N_2558,N_2337,N_2277);
or U2559 (N_2559,N_2280,N_2210);
or U2560 (N_2560,N_2328,N_2110);
nor U2561 (N_2561,N_2078,N_1869);
nand U2562 (N_2562,N_2135,N_2024);
nand U2563 (N_2563,N_2348,N_2235);
or U2564 (N_2564,N_2246,N_2172);
nor U2565 (N_2565,N_1905,N_1989);
nand U2566 (N_2566,N_2318,N_2149);
or U2567 (N_2567,N_2023,N_2150);
and U2568 (N_2568,N_2254,N_2087);
and U2569 (N_2569,N_2372,N_2309);
and U2570 (N_2570,N_1962,N_1996);
nand U2571 (N_2571,N_1943,N_2012);
and U2572 (N_2572,N_1846,N_2353);
nor U2573 (N_2573,N_2347,N_2239);
nor U2574 (N_2574,N_1920,N_2367);
nor U2575 (N_2575,N_1862,N_1866);
and U2576 (N_2576,N_1953,N_2031);
and U2577 (N_2577,N_2320,N_2038);
and U2578 (N_2578,N_2086,N_2004);
nand U2579 (N_2579,N_1813,N_1886);
nand U2580 (N_2580,N_2224,N_2022);
or U2581 (N_2581,N_1889,N_2019);
nand U2582 (N_2582,N_1852,N_1882);
and U2583 (N_2583,N_1974,N_1999);
and U2584 (N_2584,N_1872,N_2295);
or U2585 (N_2585,N_1969,N_1973);
and U2586 (N_2586,N_1890,N_2299);
or U2587 (N_2587,N_1832,N_2273);
and U2588 (N_2588,N_2354,N_1988);
nand U2589 (N_2589,N_2263,N_2248);
and U2590 (N_2590,N_2088,N_1891);
or U2591 (N_2591,N_1899,N_1827);
xor U2592 (N_2592,N_2139,N_2321);
and U2593 (N_2593,N_2237,N_1870);
and U2594 (N_2594,N_2094,N_1876);
nor U2595 (N_2595,N_2385,N_2303);
nand U2596 (N_2596,N_2030,N_2332);
or U2597 (N_2597,N_2112,N_2152);
or U2598 (N_2598,N_2345,N_2155);
nand U2599 (N_2599,N_2334,N_2018);
nor U2600 (N_2600,N_1900,N_2342);
nand U2601 (N_2601,N_2223,N_2375);
or U2602 (N_2602,N_2052,N_2113);
and U2603 (N_2603,N_2163,N_2268);
or U2604 (N_2604,N_2212,N_1847);
nor U2605 (N_2605,N_1805,N_2142);
nand U2606 (N_2606,N_1868,N_1822);
nand U2607 (N_2607,N_2308,N_2380);
nand U2608 (N_2608,N_2154,N_2090);
and U2609 (N_2609,N_2316,N_2297);
nand U2610 (N_2610,N_2048,N_2077);
or U2611 (N_2611,N_2049,N_1895);
nor U2612 (N_2612,N_1976,N_1933);
nand U2613 (N_2613,N_1946,N_2284);
nand U2614 (N_2614,N_2218,N_2123);
nor U2615 (N_2615,N_1941,N_2202);
nor U2616 (N_2616,N_2032,N_2005);
and U2617 (N_2617,N_2291,N_2315);
nor U2618 (N_2618,N_1937,N_2262);
nor U2619 (N_2619,N_2327,N_1903);
nor U2620 (N_2620,N_2117,N_1979);
and U2621 (N_2621,N_2325,N_1949);
nand U2622 (N_2622,N_2162,N_1938);
or U2623 (N_2623,N_2394,N_1967);
and U2624 (N_2624,N_2174,N_2096);
nor U2625 (N_2625,N_1865,N_2281);
and U2626 (N_2626,N_2029,N_2101);
nand U2627 (N_2627,N_2204,N_2062);
nand U2628 (N_2628,N_2069,N_1906);
and U2629 (N_2629,N_2314,N_2333);
nand U2630 (N_2630,N_2131,N_1965);
or U2631 (N_2631,N_1987,N_1951);
or U2632 (N_2632,N_2125,N_1849);
nor U2633 (N_2633,N_2208,N_2066);
nor U2634 (N_2634,N_2294,N_2271);
and U2635 (N_2635,N_2140,N_2007);
nand U2636 (N_2636,N_1970,N_2173);
nor U2637 (N_2637,N_2027,N_1922);
and U2638 (N_2638,N_2275,N_2215);
xor U2639 (N_2639,N_2025,N_2244);
and U2640 (N_2640,N_2391,N_1828);
and U2641 (N_2641,N_2363,N_2243);
nor U2642 (N_2642,N_1978,N_2399);
and U2643 (N_2643,N_2378,N_2389);
or U2644 (N_2644,N_2177,N_2073);
nor U2645 (N_2645,N_2119,N_2144);
and U2646 (N_2646,N_2344,N_2194);
and U2647 (N_2647,N_1800,N_2200);
nand U2648 (N_2648,N_1980,N_2182);
nor U2649 (N_2649,N_2079,N_2290);
nor U2650 (N_2650,N_1863,N_2313);
and U2651 (N_2651,N_2057,N_2067);
or U2652 (N_2652,N_1853,N_1861);
or U2653 (N_2653,N_2058,N_2164);
nand U2654 (N_2654,N_1908,N_2199);
nand U2655 (N_2655,N_2379,N_2352);
or U2656 (N_2656,N_1892,N_2085);
and U2657 (N_2657,N_2147,N_2185);
or U2658 (N_2658,N_1854,N_2341);
or U2659 (N_2659,N_2289,N_1990);
nor U2660 (N_2660,N_1963,N_2026);
and U2661 (N_2661,N_2042,N_2081);
and U2662 (N_2662,N_2324,N_2146);
and U2663 (N_2663,N_1934,N_2376);
nand U2664 (N_2664,N_1894,N_2179);
nand U2665 (N_2665,N_2358,N_2323);
nor U2666 (N_2666,N_2211,N_2189);
or U2667 (N_2667,N_2392,N_1917);
nor U2668 (N_2668,N_1975,N_2033);
and U2669 (N_2669,N_2171,N_2065);
and U2670 (N_2670,N_1945,N_1881);
or U2671 (N_2671,N_1916,N_2286);
or U2672 (N_2672,N_2071,N_2143);
nand U2673 (N_2673,N_2145,N_1859);
nor U2674 (N_2674,N_2201,N_1823);
and U2675 (N_2675,N_2197,N_2133);
nor U2676 (N_2676,N_2124,N_1878);
nand U2677 (N_2677,N_2374,N_1981);
and U2678 (N_2678,N_2093,N_2238);
nand U2679 (N_2679,N_2330,N_2232);
nand U2680 (N_2680,N_2196,N_1815);
or U2681 (N_2681,N_2250,N_2230);
nor U2682 (N_2682,N_2298,N_2228);
nor U2683 (N_2683,N_1835,N_1923);
nand U2684 (N_2684,N_1904,N_2304);
or U2685 (N_2685,N_1913,N_2166);
nand U2686 (N_2686,N_2187,N_1826);
nand U2687 (N_2687,N_2233,N_2317);
and U2688 (N_2688,N_2186,N_2213);
nor U2689 (N_2689,N_2028,N_1914);
nand U2690 (N_2690,N_2127,N_2122);
and U2691 (N_2691,N_2214,N_1972);
nor U2692 (N_2692,N_2089,N_2206);
nor U2693 (N_2693,N_2305,N_1997);
nor U2694 (N_2694,N_1992,N_2059);
nor U2695 (N_2695,N_2104,N_2221);
nor U2696 (N_2696,N_2184,N_1880);
or U2697 (N_2697,N_2126,N_2364);
nand U2698 (N_2698,N_2371,N_1986);
nand U2699 (N_2699,N_2053,N_1842);
or U2700 (N_2700,N_2108,N_1939);
nand U2701 (N_2701,N_2160,N_2279);
nor U2702 (N_2702,N_2299,N_2236);
nand U2703 (N_2703,N_2030,N_2017);
or U2704 (N_2704,N_2101,N_2311);
nor U2705 (N_2705,N_2096,N_2059);
or U2706 (N_2706,N_2091,N_2037);
nor U2707 (N_2707,N_1894,N_2268);
nor U2708 (N_2708,N_1878,N_2204);
nor U2709 (N_2709,N_1994,N_2351);
and U2710 (N_2710,N_2195,N_2027);
nand U2711 (N_2711,N_2322,N_2270);
nor U2712 (N_2712,N_1818,N_2085);
and U2713 (N_2713,N_2286,N_1896);
nand U2714 (N_2714,N_2334,N_2027);
nand U2715 (N_2715,N_1978,N_2057);
or U2716 (N_2716,N_1853,N_2380);
or U2717 (N_2717,N_2320,N_2173);
xnor U2718 (N_2718,N_1901,N_2360);
and U2719 (N_2719,N_2330,N_2362);
nand U2720 (N_2720,N_1957,N_2271);
nand U2721 (N_2721,N_1887,N_2232);
nor U2722 (N_2722,N_2178,N_1995);
nand U2723 (N_2723,N_2028,N_1982);
or U2724 (N_2724,N_1813,N_1881);
and U2725 (N_2725,N_1875,N_2227);
xor U2726 (N_2726,N_2395,N_2388);
nand U2727 (N_2727,N_2181,N_2378);
and U2728 (N_2728,N_1985,N_2323);
nand U2729 (N_2729,N_2343,N_1881);
or U2730 (N_2730,N_2028,N_2311);
and U2731 (N_2731,N_2343,N_2315);
nand U2732 (N_2732,N_2087,N_1862);
nor U2733 (N_2733,N_1897,N_1986);
nand U2734 (N_2734,N_1873,N_2022);
nand U2735 (N_2735,N_1964,N_1832);
nand U2736 (N_2736,N_1813,N_2000);
nor U2737 (N_2737,N_1807,N_2358);
or U2738 (N_2738,N_2275,N_2394);
or U2739 (N_2739,N_2347,N_1918);
nand U2740 (N_2740,N_2195,N_2236);
nor U2741 (N_2741,N_2180,N_1996);
and U2742 (N_2742,N_2070,N_1860);
or U2743 (N_2743,N_2128,N_2387);
and U2744 (N_2744,N_1830,N_2192);
or U2745 (N_2745,N_2198,N_1821);
and U2746 (N_2746,N_1950,N_2184);
or U2747 (N_2747,N_2070,N_2051);
nand U2748 (N_2748,N_2204,N_1928);
nand U2749 (N_2749,N_2256,N_1915);
or U2750 (N_2750,N_1981,N_2255);
nand U2751 (N_2751,N_1846,N_1873);
nor U2752 (N_2752,N_1832,N_2062);
nor U2753 (N_2753,N_2105,N_1864);
or U2754 (N_2754,N_1865,N_1861);
nand U2755 (N_2755,N_1938,N_1805);
and U2756 (N_2756,N_1868,N_2178);
or U2757 (N_2757,N_2234,N_2250);
or U2758 (N_2758,N_2229,N_1983);
nor U2759 (N_2759,N_2041,N_2193);
and U2760 (N_2760,N_1952,N_2204);
nor U2761 (N_2761,N_2232,N_2137);
nor U2762 (N_2762,N_1968,N_2244);
and U2763 (N_2763,N_2085,N_2154);
or U2764 (N_2764,N_2194,N_2169);
and U2765 (N_2765,N_2268,N_2245);
or U2766 (N_2766,N_2028,N_1889);
nor U2767 (N_2767,N_1924,N_1874);
or U2768 (N_2768,N_2018,N_1905);
or U2769 (N_2769,N_2059,N_1893);
nand U2770 (N_2770,N_2036,N_2263);
or U2771 (N_2771,N_1951,N_2259);
nor U2772 (N_2772,N_2356,N_1880);
nand U2773 (N_2773,N_1945,N_2341);
nand U2774 (N_2774,N_2295,N_2331);
nand U2775 (N_2775,N_2305,N_2042);
and U2776 (N_2776,N_2286,N_1876);
or U2777 (N_2777,N_2369,N_2092);
nor U2778 (N_2778,N_2328,N_2010);
and U2779 (N_2779,N_1870,N_1997);
or U2780 (N_2780,N_2328,N_2341);
nor U2781 (N_2781,N_1949,N_1885);
nor U2782 (N_2782,N_2397,N_1992);
or U2783 (N_2783,N_2111,N_2028);
or U2784 (N_2784,N_2174,N_1976);
nor U2785 (N_2785,N_2172,N_1982);
nand U2786 (N_2786,N_2353,N_1981);
or U2787 (N_2787,N_2034,N_2291);
xor U2788 (N_2788,N_2366,N_2160);
and U2789 (N_2789,N_2018,N_2111);
nand U2790 (N_2790,N_2043,N_2180);
or U2791 (N_2791,N_2001,N_2000);
and U2792 (N_2792,N_2295,N_2025);
nand U2793 (N_2793,N_2228,N_2198);
nand U2794 (N_2794,N_2243,N_1988);
nor U2795 (N_2795,N_2267,N_2211);
or U2796 (N_2796,N_1881,N_2132);
and U2797 (N_2797,N_2377,N_2232);
and U2798 (N_2798,N_2100,N_2173);
nor U2799 (N_2799,N_1832,N_2032);
or U2800 (N_2800,N_2279,N_1928);
and U2801 (N_2801,N_1931,N_2191);
nand U2802 (N_2802,N_2058,N_2344);
or U2803 (N_2803,N_2011,N_1850);
nor U2804 (N_2804,N_1899,N_1854);
or U2805 (N_2805,N_2073,N_1806);
nor U2806 (N_2806,N_1984,N_1948);
nor U2807 (N_2807,N_2274,N_2052);
and U2808 (N_2808,N_2041,N_2039);
nand U2809 (N_2809,N_2054,N_2389);
nand U2810 (N_2810,N_2103,N_1884);
or U2811 (N_2811,N_2218,N_2297);
or U2812 (N_2812,N_2196,N_2363);
xnor U2813 (N_2813,N_1887,N_2129);
nor U2814 (N_2814,N_2163,N_2172);
nor U2815 (N_2815,N_2262,N_2334);
nand U2816 (N_2816,N_2320,N_1986);
or U2817 (N_2817,N_2082,N_1985);
nor U2818 (N_2818,N_1829,N_1880);
or U2819 (N_2819,N_2208,N_2270);
nand U2820 (N_2820,N_1942,N_2261);
or U2821 (N_2821,N_1844,N_2090);
nor U2822 (N_2822,N_2399,N_2306);
or U2823 (N_2823,N_2073,N_1983);
nor U2824 (N_2824,N_2002,N_2189);
nand U2825 (N_2825,N_2256,N_2235);
and U2826 (N_2826,N_2308,N_1866);
and U2827 (N_2827,N_2327,N_2382);
nand U2828 (N_2828,N_1861,N_1859);
and U2829 (N_2829,N_2080,N_2050);
and U2830 (N_2830,N_2093,N_2124);
and U2831 (N_2831,N_2340,N_2317);
nor U2832 (N_2832,N_2239,N_2228);
nand U2833 (N_2833,N_1961,N_2087);
nor U2834 (N_2834,N_2008,N_2215);
nor U2835 (N_2835,N_2317,N_2343);
or U2836 (N_2836,N_1809,N_2112);
and U2837 (N_2837,N_2205,N_2162);
or U2838 (N_2838,N_2355,N_1856);
and U2839 (N_2839,N_2036,N_1930);
nand U2840 (N_2840,N_2077,N_1875);
or U2841 (N_2841,N_1992,N_2206);
nand U2842 (N_2842,N_1972,N_1872);
nor U2843 (N_2843,N_2283,N_1970);
and U2844 (N_2844,N_1918,N_1855);
nor U2845 (N_2845,N_2381,N_2247);
or U2846 (N_2846,N_1913,N_2304);
nor U2847 (N_2847,N_2068,N_2321);
nand U2848 (N_2848,N_1810,N_1885);
and U2849 (N_2849,N_1870,N_1963);
nand U2850 (N_2850,N_2210,N_2034);
nor U2851 (N_2851,N_2389,N_1821);
and U2852 (N_2852,N_1949,N_2322);
xor U2853 (N_2853,N_2155,N_2131);
nor U2854 (N_2854,N_2097,N_1841);
or U2855 (N_2855,N_1998,N_2165);
nor U2856 (N_2856,N_2236,N_2210);
or U2857 (N_2857,N_1820,N_2352);
nor U2858 (N_2858,N_1927,N_1955);
and U2859 (N_2859,N_2269,N_1925);
or U2860 (N_2860,N_1885,N_2012);
nand U2861 (N_2861,N_1913,N_2042);
nand U2862 (N_2862,N_2207,N_2192);
nand U2863 (N_2863,N_2157,N_2051);
or U2864 (N_2864,N_2380,N_1813);
nand U2865 (N_2865,N_2325,N_2207);
and U2866 (N_2866,N_2279,N_2139);
nor U2867 (N_2867,N_2207,N_2126);
or U2868 (N_2868,N_2077,N_2166);
and U2869 (N_2869,N_2156,N_2074);
or U2870 (N_2870,N_2106,N_2179);
or U2871 (N_2871,N_2149,N_2074);
or U2872 (N_2872,N_2272,N_2228);
or U2873 (N_2873,N_1968,N_2143);
and U2874 (N_2874,N_1905,N_2110);
and U2875 (N_2875,N_1947,N_1891);
and U2876 (N_2876,N_1885,N_1973);
xnor U2877 (N_2877,N_1901,N_2066);
or U2878 (N_2878,N_2235,N_2134);
nand U2879 (N_2879,N_2222,N_1927);
xnor U2880 (N_2880,N_2106,N_1858);
nor U2881 (N_2881,N_1927,N_2130);
and U2882 (N_2882,N_2304,N_2367);
nor U2883 (N_2883,N_2325,N_2261);
and U2884 (N_2884,N_1837,N_2072);
and U2885 (N_2885,N_2357,N_2213);
or U2886 (N_2886,N_2300,N_1988);
and U2887 (N_2887,N_1882,N_1932);
nor U2888 (N_2888,N_2104,N_2078);
nor U2889 (N_2889,N_1976,N_2154);
nand U2890 (N_2890,N_2077,N_2148);
nor U2891 (N_2891,N_2105,N_2180);
and U2892 (N_2892,N_2129,N_2211);
nand U2893 (N_2893,N_1916,N_1822);
nand U2894 (N_2894,N_1801,N_2282);
and U2895 (N_2895,N_1828,N_2369);
and U2896 (N_2896,N_1926,N_1939);
nor U2897 (N_2897,N_2319,N_2207);
nor U2898 (N_2898,N_1881,N_2013);
nor U2899 (N_2899,N_2233,N_1979);
or U2900 (N_2900,N_2286,N_2142);
or U2901 (N_2901,N_2019,N_2286);
and U2902 (N_2902,N_2068,N_1957);
and U2903 (N_2903,N_2360,N_1833);
and U2904 (N_2904,N_2210,N_2039);
nor U2905 (N_2905,N_2350,N_1803);
nor U2906 (N_2906,N_2323,N_1869);
or U2907 (N_2907,N_1878,N_2049);
nand U2908 (N_2908,N_2076,N_1875);
nor U2909 (N_2909,N_2242,N_2275);
nor U2910 (N_2910,N_1841,N_2318);
and U2911 (N_2911,N_2239,N_2391);
and U2912 (N_2912,N_2201,N_2009);
nand U2913 (N_2913,N_2227,N_2355);
nor U2914 (N_2914,N_2185,N_2346);
or U2915 (N_2915,N_2320,N_2260);
nand U2916 (N_2916,N_1828,N_1939);
and U2917 (N_2917,N_2365,N_2142);
or U2918 (N_2918,N_2066,N_2023);
nor U2919 (N_2919,N_2018,N_2104);
nand U2920 (N_2920,N_1878,N_2031);
nand U2921 (N_2921,N_2367,N_2198);
nor U2922 (N_2922,N_2237,N_2337);
or U2923 (N_2923,N_1939,N_2375);
and U2924 (N_2924,N_2211,N_2387);
or U2925 (N_2925,N_1851,N_1921);
nand U2926 (N_2926,N_1877,N_2207);
nand U2927 (N_2927,N_1809,N_2363);
or U2928 (N_2928,N_2240,N_1870);
nor U2929 (N_2929,N_2153,N_1895);
or U2930 (N_2930,N_2302,N_2038);
and U2931 (N_2931,N_2391,N_2199);
and U2932 (N_2932,N_2187,N_1899);
and U2933 (N_2933,N_2253,N_2174);
or U2934 (N_2934,N_1992,N_2101);
or U2935 (N_2935,N_2259,N_2147);
or U2936 (N_2936,N_2009,N_2343);
and U2937 (N_2937,N_1963,N_2109);
or U2938 (N_2938,N_2304,N_2016);
and U2939 (N_2939,N_2144,N_1930);
nand U2940 (N_2940,N_1850,N_2162);
xor U2941 (N_2941,N_2399,N_1841);
or U2942 (N_2942,N_1895,N_1924);
nor U2943 (N_2943,N_2014,N_2139);
nand U2944 (N_2944,N_2023,N_1957);
and U2945 (N_2945,N_2019,N_2089);
or U2946 (N_2946,N_1965,N_2291);
nand U2947 (N_2947,N_2112,N_2354);
and U2948 (N_2948,N_2055,N_2392);
nand U2949 (N_2949,N_2377,N_2370);
nor U2950 (N_2950,N_1902,N_1871);
or U2951 (N_2951,N_2140,N_1854);
and U2952 (N_2952,N_2164,N_2197);
nor U2953 (N_2953,N_2178,N_2348);
nor U2954 (N_2954,N_2143,N_1844);
and U2955 (N_2955,N_1952,N_1853);
nor U2956 (N_2956,N_2079,N_2155);
and U2957 (N_2957,N_2366,N_2146);
nand U2958 (N_2958,N_2305,N_2252);
nor U2959 (N_2959,N_2369,N_1990);
nor U2960 (N_2960,N_2302,N_2135);
nand U2961 (N_2961,N_1804,N_1950);
xor U2962 (N_2962,N_2179,N_1838);
nand U2963 (N_2963,N_1832,N_2095);
nand U2964 (N_2964,N_2150,N_2114);
and U2965 (N_2965,N_2171,N_2086);
and U2966 (N_2966,N_1887,N_1960);
nor U2967 (N_2967,N_2366,N_2333);
nand U2968 (N_2968,N_2344,N_2139);
nand U2969 (N_2969,N_2008,N_1862);
and U2970 (N_2970,N_2180,N_2349);
nand U2971 (N_2971,N_1858,N_2364);
or U2972 (N_2972,N_2037,N_2305);
and U2973 (N_2973,N_2176,N_2056);
nor U2974 (N_2974,N_2157,N_2317);
or U2975 (N_2975,N_2114,N_1915);
nand U2976 (N_2976,N_1905,N_2373);
nor U2977 (N_2977,N_2195,N_2158);
and U2978 (N_2978,N_1975,N_2187);
nand U2979 (N_2979,N_1827,N_2352);
nor U2980 (N_2980,N_2184,N_2377);
or U2981 (N_2981,N_2261,N_1923);
and U2982 (N_2982,N_2224,N_1833);
or U2983 (N_2983,N_2075,N_1999);
or U2984 (N_2984,N_2149,N_2097);
nor U2985 (N_2985,N_2075,N_1993);
or U2986 (N_2986,N_1862,N_1825);
and U2987 (N_2987,N_1990,N_2001);
or U2988 (N_2988,N_2378,N_1982);
nand U2989 (N_2989,N_2210,N_2309);
nor U2990 (N_2990,N_1874,N_2116);
nand U2991 (N_2991,N_1911,N_1895);
and U2992 (N_2992,N_2153,N_2076);
nor U2993 (N_2993,N_2161,N_2342);
nand U2994 (N_2994,N_2153,N_2030);
nand U2995 (N_2995,N_2126,N_2135);
xnor U2996 (N_2996,N_2246,N_2039);
nand U2997 (N_2997,N_1874,N_2244);
or U2998 (N_2998,N_2111,N_2348);
nand U2999 (N_2999,N_2142,N_1911);
or UO_0 (O_0,N_2629,N_2423);
and UO_1 (O_1,N_2532,N_2542);
nand UO_2 (O_2,N_2992,N_2968);
and UO_3 (O_3,N_2639,N_2678);
and UO_4 (O_4,N_2619,N_2624);
nand UO_5 (O_5,N_2617,N_2779);
or UO_6 (O_6,N_2812,N_2965);
nor UO_7 (O_7,N_2508,N_2738);
nor UO_8 (O_8,N_2455,N_2649);
nor UO_9 (O_9,N_2940,N_2748);
nand UO_10 (O_10,N_2895,N_2635);
nor UO_11 (O_11,N_2687,N_2874);
nor UO_12 (O_12,N_2887,N_2730);
nor UO_13 (O_13,N_2973,N_2995);
or UO_14 (O_14,N_2837,N_2596);
or UO_15 (O_15,N_2510,N_2789);
or UO_16 (O_16,N_2760,N_2964);
or UO_17 (O_17,N_2491,N_2918);
and UO_18 (O_18,N_2770,N_2605);
nand UO_19 (O_19,N_2483,N_2453);
nor UO_20 (O_20,N_2728,N_2817);
and UO_21 (O_21,N_2660,N_2886);
xor UO_22 (O_22,N_2425,N_2801);
and UO_23 (O_23,N_2791,N_2990);
or UO_24 (O_24,N_2869,N_2939);
nand UO_25 (O_25,N_2559,N_2420);
nand UO_26 (O_26,N_2818,N_2433);
and UO_27 (O_27,N_2419,N_2948);
and UO_28 (O_28,N_2668,N_2470);
and UO_29 (O_29,N_2488,N_2442);
and UO_30 (O_30,N_2766,N_2829);
nand UO_31 (O_31,N_2552,N_2839);
or UO_32 (O_32,N_2636,N_2997);
and UO_33 (O_33,N_2686,N_2896);
nor UO_34 (O_34,N_2947,N_2473);
nor UO_35 (O_35,N_2880,N_2611);
xnor UO_36 (O_36,N_2480,N_2569);
or UO_37 (O_37,N_2894,N_2441);
nor UO_38 (O_38,N_2661,N_2720);
or UO_39 (O_39,N_2590,N_2615);
and UO_40 (O_40,N_2755,N_2924);
and UO_41 (O_41,N_2716,N_2603);
and UO_42 (O_42,N_2969,N_2852);
and UO_43 (O_43,N_2489,N_2452);
nor UO_44 (O_44,N_2910,N_2937);
nor UO_45 (O_45,N_2953,N_2681);
nor UO_46 (O_46,N_2875,N_2855);
nor UO_47 (O_47,N_2505,N_2921);
nor UO_48 (O_48,N_2461,N_2666);
or UO_49 (O_49,N_2761,N_2550);
or UO_50 (O_50,N_2980,N_2827);
or UO_51 (O_51,N_2691,N_2466);
and UO_52 (O_52,N_2702,N_2606);
nor UO_53 (O_53,N_2906,N_2447);
or UO_54 (O_54,N_2417,N_2664);
and UO_55 (O_55,N_2946,N_2640);
nand UO_56 (O_56,N_2733,N_2723);
or UO_57 (O_57,N_2774,N_2721);
and UO_58 (O_58,N_2509,N_2979);
nand UO_59 (O_59,N_2669,N_2991);
and UO_60 (O_60,N_2469,N_2614);
nor UO_61 (O_61,N_2872,N_2983);
and UO_62 (O_62,N_2955,N_2485);
nor UO_63 (O_63,N_2741,N_2777);
nor UO_64 (O_64,N_2904,N_2727);
and UO_65 (O_65,N_2667,N_2902);
nor UO_66 (O_66,N_2870,N_2807);
and UO_67 (O_67,N_2600,N_2739);
nor UO_68 (O_68,N_2683,N_2934);
or UO_69 (O_69,N_2927,N_2407);
and UO_70 (O_70,N_2451,N_2695);
and UO_71 (O_71,N_2864,N_2633);
and UO_72 (O_72,N_2487,N_2712);
or UO_73 (O_73,N_2731,N_2850);
nor UO_74 (O_74,N_2725,N_2450);
nor UO_75 (O_75,N_2699,N_2623);
or UO_76 (O_76,N_2457,N_2634);
and UO_77 (O_77,N_2612,N_2520);
nor UO_78 (O_78,N_2462,N_2555);
xor UO_79 (O_79,N_2402,N_2949);
or UO_80 (O_80,N_2482,N_2860);
nor UO_81 (O_81,N_2601,N_2471);
xor UO_82 (O_82,N_2662,N_2657);
xor UO_83 (O_83,N_2942,N_2638);
nand UO_84 (O_84,N_2688,N_2684);
or UO_85 (O_85,N_2710,N_2539);
nand UO_86 (O_86,N_2517,N_2844);
and UO_87 (O_87,N_2982,N_2900);
nand UO_88 (O_88,N_2805,N_2588);
nand UO_89 (O_89,N_2602,N_2868);
and UO_90 (O_90,N_2808,N_2907);
or UO_91 (O_91,N_2888,N_2680);
nand UO_92 (O_92,N_2828,N_2785);
or UO_93 (O_93,N_2515,N_2565);
nor UO_94 (O_94,N_2556,N_2796);
nor UO_95 (O_95,N_2573,N_2406);
or UO_96 (O_96,N_2412,N_2424);
nor UO_97 (O_97,N_2432,N_2707);
and UO_98 (O_98,N_2563,N_2804);
and UO_99 (O_99,N_2853,N_2987);
nand UO_100 (O_100,N_2978,N_2715);
nor UO_101 (O_101,N_2831,N_2551);
nor UO_102 (O_102,N_2421,N_2445);
and UO_103 (O_103,N_2977,N_2673);
and UO_104 (O_104,N_2644,N_2865);
and UO_105 (O_105,N_2490,N_2714);
nor UO_106 (O_106,N_2535,N_2759);
nor UO_107 (O_107,N_2786,N_2816);
and UO_108 (O_108,N_2444,N_2959);
or UO_109 (O_109,N_2586,N_2652);
nor UO_110 (O_110,N_2478,N_2866);
or UO_111 (O_111,N_2694,N_2911);
nor UO_112 (O_112,N_2988,N_2996);
nand UO_113 (O_113,N_2670,N_2460);
and UO_114 (O_114,N_2527,N_2599);
nor UO_115 (O_115,N_2632,N_2467);
or UO_116 (O_116,N_2754,N_2861);
nand UO_117 (O_117,N_2437,N_2431);
and UO_118 (O_118,N_2521,N_2859);
nor UO_119 (O_119,N_2833,N_2957);
and UO_120 (O_120,N_2583,N_2971);
or UO_121 (O_121,N_2597,N_2967);
xnor UO_122 (O_122,N_2506,N_2576);
nand UO_123 (O_123,N_2595,N_2905);
and UO_124 (O_124,N_2798,N_2713);
or UO_125 (O_125,N_2908,N_2788);
or UO_126 (O_126,N_2848,N_2647);
nor UO_127 (O_127,N_2851,N_2562);
nor UO_128 (O_128,N_2836,N_2993);
and UO_129 (O_129,N_2709,N_2708);
nor UO_130 (O_130,N_2845,N_2915);
or UO_131 (O_131,N_2416,N_2726);
nor UO_132 (O_132,N_2404,N_2526);
nor UO_133 (O_133,N_2581,N_2484);
nand UO_134 (O_134,N_2566,N_2497);
nor UO_135 (O_135,N_2516,N_2734);
or UO_136 (O_136,N_2514,N_2703);
or UO_137 (O_137,N_2449,N_2544);
or UO_138 (O_138,N_2543,N_2752);
and UO_139 (O_139,N_2758,N_2568);
and UO_140 (O_140,N_2950,N_2405);
or UO_141 (O_141,N_2513,N_2692);
or UO_142 (O_142,N_2945,N_2878);
or UO_143 (O_143,N_2890,N_2418);
nor UO_144 (O_144,N_2787,N_2511);
nor UO_145 (O_145,N_2561,N_2830);
or UO_146 (O_146,N_2577,N_2742);
or UO_147 (O_147,N_2572,N_2504);
nand UO_148 (O_148,N_2881,N_2503);
or UO_149 (O_149,N_2524,N_2591);
xor UO_150 (O_150,N_2975,N_2486);
nor UO_151 (O_151,N_2456,N_2919);
nor UO_152 (O_152,N_2622,N_2832);
and UO_153 (O_153,N_2536,N_2693);
or UO_154 (O_154,N_2523,N_2954);
nand UO_155 (O_155,N_2826,N_2665);
or UO_156 (O_156,N_2522,N_2928);
or UO_157 (O_157,N_2682,N_2659);
and UO_158 (O_158,N_2443,N_2757);
nor UO_159 (O_159,N_2815,N_2642);
nand UO_160 (O_160,N_2820,N_2529);
and UO_161 (O_161,N_2744,N_2960);
or UO_162 (O_162,N_2841,N_2414);
and UO_163 (O_163,N_2898,N_2540);
or UO_164 (O_164,N_2884,N_2737);
nand UO_165 (O_165,N_2458,N_2962);
xor UO_166 (O_166,N_2704,N_2956);
and UO_167 (O_167,N_2912,N_2970);
and UO_168 (O_168,N_2794,N_2637);
nand UO_169 (O_169,N_2630,N_2803);
nor UO_170 (O_170,N_2897,N_2784);
or UO_171 (O_171,N_2674,N_2711);
nand UO_172 (O_172,N_2775,N_2613);
nor UO_173 (O_173,N_2646,N_2580);
nand UO_174 (O_174,N_2475,N_2534);
nor UO_175 (O_175,N_2554,N_2879);
and UO_176 (O_176,N_2771,N_2916);
and UO_177 (O_177,N_2935,N_2790);
or UO_178 (O_178,N_2889,N_2654);
nor UO_179 (O_179,N_2474,N_2476);
nor UO_180 (O_180,N_2658,N_2920);
or UO_181 (O_181,N_2593,N_2876);
xnor UO_182 (O_182,N_2925,N_2428);
nor UO_183 (O_183,N_2675,N_2840);
nand UO_184 (O_184,N_2732,N_2999);
and UO_185 (O_185,N_2834,N_2843);
nand UO_186 (O_186,N_2722,N_2951);
and UO_187 (O_187,N_2594,N_2972);
or UO_188 (O_188,N_2974,N_2729);
and UO_189 (O_189,N_2944,N_2767);
or UO_190 (O_190,N_2923,N_2496);
nor UO_191 (O_191,N_2985,N_2762);
nand UO_192 (O_192,N_2824,N_2809);
nor UO_193 (O_193,N_2795,N_2835);
nand UO_194 (O_194,N_2701,N_2413);
nor UO_195 (O_195,N_2679,N_2763);
nor UO_196 (O_196,N_2984,N_2574);
nand UO_197 (O_197,N_2538,N_2847);
or UO_198 (O_198,N_2427,N_2604);
and UO_199 (O_199,N_2782,N_2650);
nand UO_200 (O_200,N_2592,N_2438);
or UO_201 (O_201,N_2531,N_2740);
nor UO_202 (O_202,N_2823,N_2854);
nand UO_203 (O_203,N_2751,N_2717);
or UO_204 (O_204,N_2400,N_2799);
and UO_205 (O_205,N_2891,N_2648);
and UO_206 (O_206,N_2549,N_2893);
and UO_207 (O_207,N_2645,N_2797);
or UO_208 (O_208,N_2537,N_2641);
and UO_209 (O_209,N_2696,N_2819);
nand UO_210 (O_210,N_2541,N_2938);
and UO_211 (O_211,N_2736,N_2403);
or UO_212 (O_212,N_2415,N_2961);
nand UO_213 (O_213,N_2952,N_2976);
or UO_214 (O_214,N_2587,N_2883);
or UO_215 (O_215,N_2436,N_2718);
or UO_216 (O_216,N_2772,N_2813);
or UO_217 (O_217,N_2477,N_2719);
or UO_218 (O_218,N_2871,N_2663);
and UO_219 (O_219,N_2863,N_2745);
and UO_220 (O_220,N_2931,N_2685);
nor UO_221 (O_221,N_2493,N_2747);
and UO_222 (O_222,N_2689,N_2507);
nor UO_223 (O_223,N_2800,N_2671);
nor UO_224 (O_224,N_2429,N_2705);
nand UO_225 (O_225,N_2627,N_2917);
or UO_226 (O_226,N_2756,N_2560);
and UO_227 (O_227,N_2643,N_2778);
nand UO_228 (O_228,N_2481,N_2783);
nand UO_229 (O_229,N_2582,N_2810);
or UO_230 (O_230,N_2409,N_2571);
or UO_231 (O_231,N_2700,N_2410);
and UO_232 (O_232,N_2621,N_2903);
nand UO_233 (O_233,N_2530,N_2858);
xor UO_234 (O_234,N_2439,N_2856);
nor UO_235 (O_235,N_2567,N_2926);
nand UO_236 (O_236,N_2846,N_2877);
or UO_237 (O_237,N_2780,N_2557);
nand UO_238 (O_238,N_2608,N_2873);
nand UO_239 (O_239,N_2929,N_2966);
nand UO_240 (O_240,N_2401,N_2806);
nor UO_241 (O_241,N_2610,N_2909);
or UO_242 (O_242,N_2564,N_2465);
nor UO_243 (O_243,N_2677,N_2913);
or UO_244 (O_244,N_2764,N_2579);
and UO_245 (O_245,N_2628,N_2446);
nand UO_246 (O_246,N_2598,N_2479);
nand UO_247 (O_247,N_2620,N_2697);
or UO_248 (O_248,N_2570,N_2494);
and UO_249 (O_249,N_2857,N_2989);
and UO_250 (O_250,N_2558,N_2495);
nor UO_251 (O_251,N_2578,N_2842);
and UO_252 (O_252,N_2618,N_2459);
or UO_253 (O_253,N_2548,N_2655);
nor UO_254 (O_254,N_2792,N_2464);
or UO_255 (O_255,N_2472,N_2768);
or UO_256 (O_256,N_2430,N_2882);
and UO_257 (O_257,N_2941,N_2781);
nand UO_258 (O_258,N_2943,N_2653);
or UO_259 (O_259,N_2492,N_2811);
nor UO_260 (O_260,N_2434,N_2616);
or UO_261 (O_261,N_2930,N_2631);
and UO_262 (O_262,N_2498,N_2584);
nand UO_263 (O_263,N_2547,N_2849);
xor UO_264 (O_264,N_2862,N_2892);
nor UO_265 (O_265,N_2440,N_2776);
or UO_266 (O_266,N_2518,N_2724);
and UO_267 (O_267,N_2994,N_2502);
nand UO_268 (O_268,N_2793,N_2899);
nor UO_269 (O_269,N_2981,N_2625);
or UO_270 (O_270,N_2914,N_2512);
and UO_271 (O_271,N_2821,N_2468);
or UO_272 (O_272,N_2769,N_2519);
and UO_273 (O_273,N_2932,N_2533);
or UO_274 (O_274,N_2545,N_2422);
or UO_275 (O_275,N_2838,N_2867);
or UO_276 (O_276,N_2500,N_2656);
or UO_277 (O_277,N_2676,N_2986);
nand UO_278 (O_278,N_2607,N_2463);
nor UO_279 (O_279,N_2553,N_2753);
nor UO_280 (O_280,N_2749,N_2922);
and UO_281 (O_281,N_2609,N_2958);
nand UO_282 (O_282,N_2743,N_2933);
or UO_283 (O_283,N_2589,N_2626);
or UO_284 (O_284,N_2528,N_2575);
and UO_285 (O_285,N_2690,N_2408);
nand UO_286 (O_286,N_2825,N_2651);
nand UO_287 (O_287,N_2963,N_2773);
nand UO_288 (O_288,N_2546,N_2454);
nand UO_289 (O_289,N_2765,N_2750);
or UO_290 (O_290,N_2585,N_2735);
nand UO_291 (O_291,N_2525,N_2802);
or UO_292 (O_292,N_2672,N_2998);
and UO_293 (O_293,N_2746,N_2885);
nand UO_294 (O_294,N_2426,N_2698);
and UO_295 (O_295,N_2936,N_2499);
and UO_296 (O_296,N_2706,N_2901);
nand UO_297 (O_297,N_2448,N_2814);
or UO_298 (O_298,N_2501,N_2411);
or UO_299 (O_299,N_2822,N_2435);
nor UO_300 (O_300,N_2540,N_2965);
and UO_301 (O_301,N_2951,N_2636);
nor UO_302 (O_302,N_2597,N_2846);
nor UO_303 (O_303,N_2942,N_2541);
and UO_304 (O_304,N_2795,N_2645);
and UO_305 (O_305,N_2459,N_2763);
or UO_306 (O_306,N_2763,N_2674);
nand UO_307 (O_307,N_2615,N_2606);
xor UO_308 (O_308,N_2923,N_2472);
and UO_309 (O_309,N_2497,N_2805);
and UO_310 (O_310,N_2768,N_2835);
or UO_311 (O_311,N_2651,N_2800);
nor UO_312 (O_312,N_2689,N_2692);
nor UO_313 (O_313,N_2440,N_2572);
nand UO_314 (O_314,N_2407,N_2494);
or UO_315 (O_315,N_2758,N_2925);
and UO_316 (O_316,N_2876,N_2727);
nand UO_317 (O_317,N_2865,N_2670);
nand UO_318 (O_318,N_2595,N_2749);
or UO_319 (O_319,N_2903,N_2417);
nand UO_320 (O_320,N_2896,N_2913);
nand UO_321 (O_321,N_2533,N_2816);
or UO_322 (O_322,N_2583,N_2547);
and UO_323 (O_323,N_2423,N_2443);
and UO_324 (O_324,N_2469,N_2861);
and UO_325 (O_325,N_2806,N_2849);
nand UO_326 (O_326,N_2818,N_2584);
nor UO_327 (O_327,N_2584,N_2869);
or UO_328 (O_328,N_2963,N_2644);
xor UO_329 (O_329,N_2920,N_2774);
or UO_330 (O_330,N_2833,N_2735);
nor UO_331 (O_331,N_2607,N_2434);
nor UO_332 (O_332,N_2909,N_2908);
nor UO_333 (O_333,N_2409,N_2989);
nand UO_334 (O_334,N_2965,N_2559);
nor UO_335 (O_335,N_2657,N_2900);
nor UO_336 (O_336,N_2586,N_2748);
or UO_337 (O_337,N_2868,N_2881);
or UO_338 (O_338,N_2878,N_2708);
or UO_339 (O_339,N_2826,N_2661);
and UO_340 (O_340,N_2768,N_2774);
and UO_341 (O_341,N_2584,N_2552);
nand UO_342 (O_342,N_2947,N_2428);
and UO_343 (O_343,N_2935,N_2748);
nand UO_344 (O_344,N_2448,N_2773);
or UO_345 (O_345,N_2541,N_2820);
nand UO_346 (O_346,N_2400,N_2479);
and UO_347 (O_347,N_2976,N_2794);
nand UO_348 (O_348,N_2868,N_2943);
and UO_349 (O_349,N_2729,N_2501);
nor UO_350 (O_350,N_2564,N_2598);
nand UO_351 (O_351,N_2401,N_2429);
and UO_352 (O_352,N_2840,N_2625);
xnor UO_353 (O_353,N_2957,N_2519);
nand UO_354 (O_354,N_2410,N_2916);
nor UO_355 (O_355,N_2418,N_2704);
nor UO_356 (O_356,N_2609,N_2917);
or UO_357 (O_357,N_2575,N_2576);
or UO_358 (O_358,N_2619,N_2491);
nand UO_359 (O_359,N_2745,N_2750);
and UO_360 (O_360,N_2834,N_2988);
nand UO_361 (O_361,N_2513,N_2830);
or UO_362 (O_362,N_2480,N_2460);
nor UO_363 (O_363,N_2971,N_2446);
or UO_364 (O_364,N_2965,N_2513);
nand UO_365 (O_365,N_2797,N_2711);
nand UO_366 (O_366,N_2628,N_2490);
or UO_367 (O_367,N_2414,N_2842);
nor UO_368 (O_368,N_2822,N_2754);
nor UO_369 (O_369,N_2711,N_2471);
or UO_370 (O_370,N_2726,N_2638);
or UO_371 (O_371,N_2790,N_2877);
nand UO_372 (O_372,N_2805,N_2542);
nand UO_373 (O_373,N_2506,N_2730);
nor UO_374 (O_374,N_2586,N_2734);
or UO_375 (O_375,N_2888,N_2784);
or UO_376 (O_376,N_2970,N_2989);
nand UO_377 (O_377,N_2433,N_2998);
and UO_378 (O_378,N_2862,N_2514);
nand UO_379 (O_379,N_2852,N_2974);
or UO_380 (O_380,N_2817,N_2678);
nand UO_381 (O_381,N_2849,N_2645);
nand UO_382 (O_382,N_2769,N_2459);
nor UO_383 (O_383,N_2738,N_2754);
nor UO_384 (O_384,N_2897,N_2546);
or UO_385 (O_385,N_2974,N_2677);
nor UO_386 (O_386,N_2789,N_2981);
and UO_387 (O_387,N_2511,N_2911);
nand UO_388 (O_388,N_2695,N_2486);
and UO_389 (O_389,N_2691,N_2493);
or UO_390 (O_390,N_2442,N_2710);
nor UO_391 (O_391,N_2603,N_2574);
or UO_392 (O_392,N_2596,N_2875);
nor UO_393 (O_393,N_2417,N_2502);
nor UO_394 (O_394,N_2418,N_2977);
or UO_395 (O_395,N_2860,N_2640);
and UO_396 (O_396,N_2516,N_2977);
or UO_397 (O_397,N_2427,N_2502);
xnor UO_398 (O_398,N_2624,N_2998);
nor UO_399 (O_399,N_2941,N_2951);
nand UO_400 (O_400,N_2850,N_2896);
and UO_401 (O_401,N_2763,N_2911);
nand UO_402 (O_402,N_2565,N_2837);
and UO_403 (O_403,N_2824,N_2658);
or UO_404 (O_404,N_2786,N_2604);
nor UO_405 (O_405,N_2944,N_2718);
or UO_406 (O_406,N_2595,N_2881);
and UO_407 (O_407,N_2577,N_2528);
nand UO_408 (O_408,N_2661,N_2923);
and UO_409 (O_409,N_2990,N_2820);
and UO_410 (O_410,N_2948,N_2460);
and UO_411 (O_411,N_2923,N_2981);
and UO_412 (O_412,N_2401,N_2997);
nor UO_413 (O_413,N_2682,N_2635);
or UO_414 (O_414,N_2649,N_2976);
or UO_415 (O_415,N_2625,N_2841);
nand UO_416 (O_416,N_2552,N_2948);
nand UO_417 (O_417,N_2925,N_2571);
nor UO_418 (O_418,N_2716,N_2452);
nand UO_419 (O_419,N_2726,N_2430);
nand UO_420 (O_420,N_2893,N_2407);
and UO_421 (O_421,N_2540,N_2731);
and UO_422 (O_422,N_2493,N_2779);
nor UO_423 (O_423,N_2892,N_2651);
nand UO_424 (O_424,N_2621,N_2518);
xnor UO_425 (O_425,N_2405,N_2670);
xor UO_426 (O_426,N_2664,N_2718);
nor UO_427 (O_427,N_2661,N_2516);
nor UO_428 (O_428,N_2913,N_2488);
or UO_429 (O_429,N_2581,N_2496);
nor UO_430 (O_430,N_2880,N_2953);
or UO_431 (O_431,N_2476,N_2654);
nand UO_432 (O_432,N_2951,N_2864);
nand UO_433 (O_433,N_2441,N_2709);
and UO_434 (O_434,N_2990,N_2829);
nor UO_435 (O_435,N_2781,N_2401);
and UO_436 (O_436,N_2919,N_2410);
or UO_437 (O_437,N_2585,N_2661);
and UO_438 (O_438,N_2630,N_2845);
nand UO_439 (O_439,N_2567,N_2697);
nand UO_440 (O_440,N_2847,N_2415);
or UO_441 (O_441,N_2878,N_2579);
nand UO_442 (O_442,N_2455,N_2814);
nand UO_443 (O_443,N_2893,N_2759);
and UO_444 (O_444,N_2741,N_2419);
nor UO_445 (O_445,N_2483,N_2403);
or UO_446 (O_446,N_2508,N_2443);
nor UO_447 (O_447,N_2716,N_2766);
nor UO_448 (O_448,N_2692,N_2638);
nand UO_449 (O_449,N_2898,N_2463);
and UO_450 (O_450,N_2495,N_2896);
nand UO_451 (O_451,N_2462,N_2677);
and UO_452 (O_452,N_2566,N_2866);
and UO_453 (O_453,N_2995,N_2657);
nand UO_454 (O_454,N_2953,N_2892);
nand UO_455 (O_455,N_2414,N_2558);
or UO_456 (O_456,N_2743,N_2588);
and UO_457 (O_457,N_2945,N_2952);
nor UO_458 (O_458,N_2448,N_2649);
nand UO_459 (O_459,N_2846,N_2732);
nand UO_460 (O_460,N_2611,N_2690);
nand UO_461 (O_461,N_2817,N_2998);
nor UO_462 (O_462,N_2524,N_2668);
nor UO_463 (O_463,N_2438,N_2610);
nand UO_464 (O_464,N_2890,N_2793);
or UO_465 (O_465,N_2431,N_2535);
nand UO_466 (O_466,N_2674,N_2601);
nand UO_467 (O_467,N_2907,N_2763);
or UO_468 (O_468,N_2696,N_2890);
nor UO_469 (O_469,N_2734,N_2730);
nand UO_470 (O_470,N_2960,N_2443);
nand UO_471 (O_471,N_2732,N_2451);
and UO_472 (O_472,N_2555,N_2706);
nor UO_473 (O_473,N_2785,N_2882);
or UO_474 (O_474,N_2715,N_2412);
nand UO_475 (O_475,N_2711,N_2724);
or UO_476 (O_476,N_2615,N_2738);
nand UO_477 (O_477,N_2720,N_2970);
or UO_478 (O_478,N_2619,N_2644);
or UO_479 (O_479,N_2569,N_2630);
nand UO_480 (O_480,N_2792,N_2798);
nand UO_481 (O_481,N_2649,N_2814);
and UO_482 (O_482,N_2663,N_2498);
and UO_483 (O_483,N_2577,N_2965);
or UO_484 (O_484,N_2704,N_2718);
nor UO_485 (O_485,N_2886,N_2642);
nor UO_486 (O_486,N_2406,N_2692);
nand UO_487 (O_487,N_2676,N_2446);
or UO_488 (O_488,N_2462,N_2601);
nor UO_489 (O_489,N_2459,N_2803);
or UO_490 (O_490,N_2484,N_2533);
nand UO_491 (O_491,N_2986,N_2660);
and UO_492 (O_492,N_2948,N_2626);
or UO_493 (O_493,N_2754,N_2770);
and UO_494 (O_494,N_2625,N_2684);
or UO_495 (O_495,N_2881,N_2668);
nand UO_496 (O_496,N_2997,N_2610);
nor UO_497 (O_497,N_2895,N_2694);
or UO_498 (O_498,N_2454,N_2592);
nor UO_499 (O_499,N_2838,N_2995);
endmodule