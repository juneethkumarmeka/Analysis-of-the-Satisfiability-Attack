module basic_1000_10000_1500_20_levels_2xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nor U0 (N_0,In_703,In_314);
nor U1 (N_1,In_460,In_173);
or U2 (N_2,In_382,In_108);
nor U3 (N_3,In_685,In_562);
or U4 (N_4,In_144,In_780);
xor U5 (N_5,In_284,In_588);
and U6 (N_6,In_696,In_304);
nand U7 (N_7,In_156,In_140);
and U8 (N_8,In_514,In_46);
nand U9 (N_9,In_798,In_99);
or U10 (N_10,In_700,In_848);
nor U11 (N_11,In_982,In_879);
nand U12 (N_12,In_821,In_312);
nand U13 (N_13,In_319,In_956);
and U14 (N_14,In_711,In_836);
or U15 (N_15,In_357,In_142);
and U16 (N_16,In_378,In_496);
or U17 (N_17,In_568,In_465);
or U18 (N_18,In_648,In_98);
or U19 (N_19,In_490,In_82);
nand U20 (N_20,In_387,In_784);
and U21 (N_21,In_972,In_772);
nor U22 (N_22,In_522,In_47);
nor U23 (N_23,In_572,In_179);
nand U24 (N_24,In_883,In_812);
nor U25 (N_25,In_469,In_379);
and U26 (N_26,In_27,In_782);
or U27 (N_27,In_199,In_310);
and U28 (N_28,In_421,In_801);
or U29 (N_29,In_191,In_654);
nand U30 (N_30,In_251,In_946);
nor U31 (N_31,In_369,In_130);
and U32 (N_32,In_534,In_886);
or U33 (N_33,In_32,In_560);
and U34 (N_34,In_487,In_442);
nor U35 (N_35,In_234,In_26);
or U36 (N_36,In_210,In_826);
nor U37 (N_37,In_204,In_827);
nand U38 (N_38,In_841,In_190);
nand U39 (N_39,In_352,In_75);
nand U40 (N_40,In_898,In_719);
or U41 (N_41,In_705,In_28);
nand U42 (N_42,In_775,In_736);
nand U43 (N_43,In_66,In_596);
and U44 (N_44,In_61,In_530);
nand U45 (N_45,In_417,In_609);
or U46 (N_46,In_335,In_748);
or U47 (N_47,In_383,In_164);
nor U48 (N_48,In_712,In_891);
or U49 (N_49,In_74,In_63);
and U50 (N_50,In_296,In_934);
nand U51 (N_51,In_542,In_59);
nand U52 (N_52,In_511,In_458);
and U53 (N_53,In_292,In_329);
nand U54 (N_54,In_363,In_797);
or U55 (N_55,In_96,In_20);
nor U56 (N_56,In_139,In_664);
nand U57 (N_57,In_136,In_92);
and U58 (N_58,In_731,In_850);
nand U59 (N_59,In_630,In_611);
or U60 (N_60,In_790,In_155);
and U61 (N_61,In_236,In_709);
or U62 (N_62,In_656,In_792);
and U63 (N_63,In_464,In_181);
nand U64 (N_64,In_247,In_275);
nor U65 (N_65,In_541,In_300);
or U66 (N_66,In_629,In_260);
and U67 (N_67,In_160,In_881);
and U68 (N_68,In_437,In_803);
or U69 (N_69,In_713,In_264);
nor U70 (N_70,In_874,In_777);
and U71 (N_71,In_904,In_622);
xnor U72 (N_72,In_192,In_925);
and U73 (N_73,In_870,In_407);
and U74 (N_74,In_852,In_5);
nand U75 (N_75,In_259,In_395);
nand U76 (N_76,In_763,In_261);
or U77 (N_77,In_809,In_185);
and U78 (N_78,In_452,In_390);
nor U79 (N_79,In_76,In_635);
and U80 (N_80,In_678,In_166);
and U81 (N_81,In_740,In_184);
and U82 (N_82,In_582,In_19);
or U83 (N_83,In_770,In_4);
nand U84 (N_84,In_698,In_707);
or U85 (N_85,In_810,In_476);
nand U86 (N_86,In_752,In_340);
and U87 (N_87,In_24,In_599);
nand U88 (N_88,In_644,In_570);
or U89 (N_89,In_571,In_478);
nor U90 (N_90,In_773,In_295);
nor U91 (N_91,In_360,In_124);
nor U92 (N_92,In_877,In_433);
and U93 (N_93,In_17,In_970);
nor U94 (N_94,In_616,In_332);
nor U95 (N_95,In_449,In_226);
or U96 (N_96,In_482,In_765);
nor U97 (N_97,In_294,In_756);
nor U98 (N_98,In_987,In_961);
nand U99 (N_99,In_154,In_313);
or U100 (N_100,In_758,In_281);
or U101 (N_101,In_301,In_646);
nand U102 (N_102,In_868,In_903);
or U103 (N_103,In_855,In_808);
or U104 (N_104,In_681,In_574);
nor U105 (N_105,In_815,In_196);
or U106 (N_106,In_849,In_730);
nand U107 (N_107,In_44,In_806);
nand U108 (N_108,In_254,In_893);
nand U109 (N_109,In_687,In_639);
and U110 (N_110,In_388,In_101);
and U111 (N_111,In_392,In_3);
or U112 (N_112,In_649,In_58);
nand U113 (N_113,In_983,In_172);
and U114 (N_114,In_643,In_919);
nand U115 (N_115,In_869,In_962);
nor U116 (N_116,In_483,In_271);
nor U117 (N_117,In_999,In_125);
nand U118 (N_118,In_370,In_677);
or U119 (N_119,In_2,In_12);
nor U120 (N_120,In_710,In_412);
nor U121 (N_121,In_218,In_342);
nor U122 (N_122,In_104,In_331);
nor U123 (N_123,In_624,In_913);
nor U124 (N_124,In_188,In_822);
nor U125 (N_125,In_978,In_384);
or U126 (N_126,In_580,In_969);
nand U127 (N_127,In_170,In_265);
nand U128 (N_128,In_800,In_908);
xor U129 (N_129,In_863,In_964);
and U130 (N_130,In_735,In_660);
and U131 (N_131,In_591,In_641);
and U132 (N_132,In_725,In_198);
nor U133 (N_133,In_1,In_244);
or U134 (N_134,In_195,In_910);
or U135 (N_135,In_739,In_148);
nand U136 (N_136,In_508,In_86);
nand U137 (N_137,In_814,In_512);
or U138 (N_138,In_285,In_381);
or U139 (N_139,In_317,In_977);
nand U140 (N_140,In_431,In_912);
or U141 (N_141,In_427,In_280);
nand U142 (N_142,In_330,In_459);
nor U143 (N_143,In_842,In_959);
nor U144 (N_144,In_344,In_804);
or U145 (N_145,In_269,In_273);
nand U146 (N_146,In_846,In_759);
nand U147 (N_147,In_322,In_688);
nor U148 (N_148,In_102,In_230);
nand U149 (N_149,In_921,In_121);
nor U150 (N_150,In_422,In_944);
or U151 (N_151,In_666,In_35);
xor U152 (N_152,In_889,In_145);
and U153 (N_153,In_537,In_267);
nand U154 (N_154,In_36,In_386);
or U155 (N_155,In_405,In_277);
nor U156 (N_156,In_31,In_657);
or U157 (N_157,In_747,In_434);
nor U158 (N_158,In_345,In_856);
nand U159 (N_159,In_43,In_684);
nor U160 (N_160,In_992,In_486);
nor U161 (N_161,In_262,In_410);
nand U162 (N_162,In_746,In_607);
or U163 (N_163,In_732,In_761);
and U164 (N_164,In_443,In_691);
nand U165 (N_165,In_150,In_828);
and U166 (N_166,In_857,In_127);
or U167 (N_167,In_603,In_966);
nor U168 (N_168,In_11,In_291);
nor U169 (N_169,In_403,In_667);
nand U170 (N_170,In_887,In_468);
nor U171 (N_171,In_741,In_393);
nor U172 (N_172,In_222,In_536);
nand U173 (N_173,In_167,In_492);
or U174 (N_174,In_94,In_93);
nor U175 (N_175,In_787,In_751);
and U176 (N_176,In_785,In_621);
or U177 (N_177,In_618,In_767);
and U178 (N_178,In_137,In_860);
nor U179 (N_179,In_202,In_477);
nor U180 (N_180,In_565,In_149);
or U181 (N_181,In_22,In_882);
and U182 (N_182,In_343,In_385);
and U183 (N_183,In_817,In_445);
and U184 (N_184,In_30,In_432);
or U185 (N_185,In_73,In_766);
nand U186 (N_186,In_62,In_8);
nor U187 (N_187,In_152,In_897);
nor U188 (N_188,In_628,In_847);
and U189 (N_189,In_915,In_548);
nand U190 (N_190,In_51,In_209);
nor U191 (N_191,In_544,In_608);
and U192 (N_192,In_636,In_626);
and U193 (N_193,In_105,In_968);
nand U194 (N_194,In_858,In_500);
or U195 (N_195,In_581,In_521);
and U196 (N_196,In_779,In_690);
and U197 (N_197,In_693,In_819);
xor U198 (N_198,In_945,In_7);
and U199 (N_199,In_920,In_578);
and U200 (N_200,In_447,In_871);
nand U201 (N_201,In_778,In_161);
or U202 (N_202,In_951,In_940);
nor U203 (N_203,In_876,In_408);
nor U204 (N_204,In_561,In_930);
nand U205 (N_205,In_186,In_470);
xor U206 (N_206,In_287,In_337);
or U207 (N_207,In_106,In_699);
nor U208 (N_208,In_771,In_223);
or U209 (N_209,In_795,In_120);
nor U210 (N_210,In_435,In_286);
nand U211 (N_211,In_0,In_135);
xnor U212 (N_212,In_757,In_400);
nor U213 (N_213,In_256,In_948);
or U214 (N_214,In_429,In_231);
and U215 (N_215,In_351,In_967);
and U216 (N_216,In_653,In_131);
or U217 (N_217,In_927,In_553);
nor U218 (N_218,In_613,In_601);
nor U219 (N_219,In_529,In_123);
nand U220 (N_220,In_455,In_444);
nor U221 (N_221,In_531,In_993);
or U222 (N_222,In_723,In_602);
or U223 (N_223,In_200,In_620);
nor U224 (N_224,In_60,In_554);
nor U225 (N_225,In_840,In_67);
nand U226 (N_226,In_960,In_504);
or U227 (N_227,In_734,In_923);
nor U228 (N_228,In_745,In_952);
nor U229 (N_229,In_738,In_834);
or U230 (N_230,In_462,In_37);
xnor U231 (N_231,In_979,In_320);
or U232 (N_232,In_854,In_631);
nand U233 (N_233,In_900,In_559);
nor U234 (N_234,In_479,In_851);
or U235 (N_235,In_651,In_957);
or U236 (N_236,In_650,In_526);
and U237 (N_237,In_34,In_107);
nor U238 (N_238,In_714,In_614);
or U239 (N_239,In_776,In_371);
or U240 (N_240,In_566,In_532);
xor U241 (N_241,In_380,In_211);
and U242 (N_242,In_176,In_576);
nor U243 (N_243,In_91,In_818);
or U244 (N_244,In_55,In_917);
nor U245 (N_245,In_706,In_126);
nand U246 (N_246,In_974,In_971);
or U247 (N_247,In_843,In_663);
and U248 (N_248,In_717,In_513);
nor U249 (N_249,In_193,In_708);
or U250 (N_250,In_556,In_53);
or U251 (N_251,In_84,In_884);
nor U252 (N_252,In_353,In_503);
nand U253 (N_253,In_14,In_327);
and U254 (N_254,In_895,In_610);
and U255 (N_255,In_438,In_764);
nor U256 (N_256,In_662,In_103);
nor U257 (N_257,In_615,In_88);
or U258 (N_258,In_165,In_197);
nor U259 (N_259,In_268,In_111);
xnor U260 (N_260,In_791,In_178);
nand U261 (N_261,In_348,In_816);
and U262 (N_262,In_228,In_10);
nand U263 (N_263,In_282,In_689);
nand U264 (N_264,In_682,In_416);
nand U265 (N_265,In_563,In_880);
nor U266 (N_266,In_546,In_425);
nand U267 (N_267,In_668,In_697);
nor U268 (N_268,In_888,In_45);
nand U269 (N_269,In_375,In_151);
and U270 (N_270,In_377,In_303);
nor U271 (N_271,In_141,In_965);
or U272 (N_272,In_594,In_307);
nand U273 (N_273,In_68,In_481);
nand U274 (N_274,In_215,In_749);
nor U275 (N_275,In_875,In_658);
or U276 (N_276,In_402,In_769);
nand U277 (N_277,In_448,In_569);
and U278 (N_278,In_950,In_220);
xor U279 (N_279,In_590,In_293);
or U280 (N_280,In_859,In_661);
nand U281 (N_281,In_305,In_253);
nor U282 (N_282,In_949,In_939);
nand U283 (N_283,In_902,In_391);
nand U284 (N_284,In_805,In_864);
nand U285 (N_285,In_175,In_133);
nor U286 (N_286,In_309,In_973);
nand U287 (N_287,In_592,In_593);
or U288 (N_288,In_867,In_750);
nor U289 (N_289,In_837,In_6);
nand U290 (N_290,In_577,In_80);
or U291 (N_291,In_450,In_938);
nand U292 (N_292,In_288,In_339);
nor U293 (N_293,In_523,In_214);
or U294 (N_294,In_638,In_985);
nand U295 (N_295,In_905,In_575);
nand U296 (N_296,In_844,In_652);
nand U297 (N_297,In_516,In_242);
xor U298 (N_298,In_354,In_411);
nand U299 (N_299,In_182,In_224);
nor U300 (N_300,In_206,In_225);
nor U301 (N_301,In_954,In_311);
or U302 (N_302,In_365,In_783);
or U303 (N_303,In_52,In_499);
and U304 (N_304,In_168,In_835);
nand U305 (N_305,In_238,In_832);
nor U306 (N_306,In_676,In_694);
or U307 (N_307,In_398,In_722);
nor U308 (N_308,In_216,In_501);
and U309 (N_309,In_116,In_372);
or U310 (N_310,In_799,In_742);
nand U311 (N_311,In_958,In_341);
or U312 (N_312,In_896,In_509);
or U313 (N_313,In_926,In_349);
xor U314 (N_314,In_794,In_79);
nor U315 (N_315,In_551,In_143);
and U316 (N_316,In_647,In_505);
or U317 (N_317,In_793,In_23);
or U318 (N_318,In_540,In_467);
nor U319 (N_319,In_823,In_389);
nor U320 (N_320,In_361,In_642);
nor U321 (N_321,In_334,In_922);
nor U322 (N_322,In_446,In_941);
nand U323 (N_323,In_42,In_786);
and U324 (N_324,In_283,In_475);
nand U325 (N_325,In_419,In_302);
nor U326 (N_326,In_159,In_85);
xnor U327 (N_327,In_413,In_171);
nand U328 (N_328,In_990,In_78);
nor U329 (N_329,In_246,In_57);
nor U330 (N_330,In_894,In_659);
and U331 (N_331,In_328,In_781);
nor U332 (N_332,In_489,In_48);
or U333 (N_333,In_87,In_39);
and U334 (N_334,In_906,In_38);
or U335 (N_335,In_916,In_89);
or U336 (N_336,In_169,In_279);
and U337 (N_337,In_257,In_671);
xor U338 (N_338,In_811,In_440);
nor U339 (N_339,In_480,In_704);
and U340 (N_340,In_623,In_789);
and U341 (N_341,In_515,In_441);
nand U342 (N_342,In_457,In_232);
nor U343 (N_343,In_366,In_180);
or U344 (N_344,In_632,In_484);
xnor U345 (N_345,In_720,In_240);
nor U346 (N_346,In_605,In_679);
nand U347 (N_347,In_907,In_16);
or U348 (N_348,In_396,In_9);
or U349 (N_349,In_13,In_862);
or U350 (N_350,In_989,In_373);
nor U351 (N_351,In_947,In_584);
nor U352 (N_352,In_909,In_90);
and U353 (N_353,In_737,In_221);
nand U354 (N_354,In_81,In_217);
or U355 (N_355,In_297,In_463);
or U356 (N_356,In_65,In_118);
nor U357 (N_357,In_557,In_524);
nand U358 (N_358,In_729,In_70);
nor U359 (N_359,In_71,In_243);
nand U360 (N_360,In_64,In_507);
and U361 (N_361,In_25,In_885);
and U362 (N_362,In_640,In_115);
or U363 (N_363,In_203,In_237);
and U364 (N_364,In_493,In_692);
or U365 (N_365,In_645,In_350);
and U366 (N_366,In_252,In_336);
or U367 (N_367,In_550,In_18);
nand U368 (N_368,In_270,In_401);
nor U369 (N_369,In_995,In_937);
nor U370 (N_370,In_669,In_368);
and U371 (N_371,In_420,In_290);
or U372 (N_372,In_519,In_975);
nor U373 (N_373,In_845,In_266);
nand U374 (N_374,In_113,In_397);
nor U375 (N_375,In_589,In_963);
nand U376 (N_376,In_986,In_890);
nand U377 (N_377,In_918,In_241);
or U378 (N_378,In_718,In_77);
and U379 (N_379,In_472,In_829);
nand U380 (N_380,In_587,In_753);
or U381 (N_381,In_715,In_943);
and U382 (N_382,In_606,In_461);
nor U383 (N_383,In_488,In_436);
or U384 (N_384,In_866,In_306);
and U385 (N_385,In_675,In_213);
or U386 (N_386,In_597,In_356);
nor U387 (N_387,In_333,In_549);
or U388 (N_388,In_128,In_453);
or U389 (N_389,In_600,In_726);
nor U390 (N_390,In_83,In_298);
nor U391 (N_391,In_485,In_69);
or U392 (N_392,In_683,In_755);
and U393 (N_393,In_670,In_338);
nand U394 (N_394,In_158,In_743);
nor U395 (N_395,In_153,In_355);
nand U396 (N_396,In_617,In_673);
nand U397 (N_397,In_899,In_535);
and U398 (N_398,In_612,In_558);
nand U399 (N_399,In_762,In_122);
or U400 (N_400,In_474,In_316);
or U401 (N_401,In_768,In_40);
and U402 (N_402,In_498,In_49);
nand U403 (N_403,In_163,In_456);
nor U404 (N_404,In_984,In_29);
and U405 (N_405,In_911,In_976);
or U406 (N_406,In_323,In_929);
nor U407 (N_407,In_21,In_861);
nor U408 (N_408,In_518,In_716);
nand U409 (N_409,In_994,In_833);
nand U410 (N_410,In_598,In_585);
nor U411 (N_411,In_539,In_194);
and U412 (N_412,In_56,In_831);
or U413 (N_413,In_996,In_796);
and U414 (N_414,In_728,In_528);
nand U415 (N_415,In_665,In_533);
or U416 (N_416,In_187,In_207);
xnor U417 (N_417,In_672,In_998);
and U418 (N_418,In_318,In_41);
xnor U419 (N_419,In_701,In_324);
or U420 (N_420,In_655,In_399);
nand U421 (N_421,In_935,In_555);
nor U422 (N_422,In_936,In_276);
or U423 (N_423,In_547,In_724);
nor U424 (N_424,In_212,In_162);
xnor U425 (N_425,In_358,In_695);
nor U426 (N_426,In_579,In_418);
nor U427 (N_427,In_674,In_633);
nand U428 (N_428,In_825,In_991);
nor U429 (N_429,In_423,In_586);
or U430 (N_430,In_543,In_278);
nor U431 (N_431,In_272,In_733);
nor U432 (N_432,In_15,In_404);
or U433 (N_433,In_129,In_788);
and U434 (N_434,In_564,In_50);
and U435 (N_435,In_227,In_409);
or U436 (N_436,In_157,In_495);
nand U437 (N_437,In_72,In_525);
nor U438 (N_438,In_112,In_321);
and U439 (N_439,In_177,In_119);
nor U440 (N_440,In_117,In_567);
or U441 (N_441,In_394,In_219);
nand U442 (N_442,In_208,In_744);
and U443 (N_443,In_174,In_604);
or U444 (N_444,In_229,In_325);
nor U445 (N_445,In_721,In_263);
nand U446 (N_446,In_430,In_878);
xor U447 (N_447,In_502,In_595);
and U448 (N_448,In_573,In_754);
or U449 (N_449,In_838,In_258);
nand U450 (N_450,In_473,In_510);
and U451 (N_451,In_97,In_583);
and U452 (N_452,In_109,In_686);
nor U453 (N_453,In_988,In_820);
nor U454 (N_454,In_406,In_326);
or U455 (N_455,In_942,In_245);
or U456 (N_456,In_824,In_892);
or U457 (N_457,In_538,In_527);
and U458 (N_458,In_552,In_931);
or U459 (N_459,In_471,In_637);
or U460 (N_460,In_839,In_189);
nand U461 (N_461,In_374,In_619);
nor U462 (N_462,In_506,In_138);
and U463 (N_463,In_239,In_439);
or U464 (N_464,In_201,In_95);
nor U465 (N_465,In_517,In_924);
nor U466 (N_466,In_134,In_359);
and U467 (N_467,In_955,In_414);
or U468 (N_468,In_997,In_953);
nor U469 (N_469,In_233,In_727);
and U470 (N_470,In_376,In_634);
or U471 (N_471,In_853,In_428);
or U472 (N_472,In_33,In_255);
and U473 (N_473,In_830,In_362);
nand U474 (N_474,In_289,In_54);
nand U475 (N_475,In_110,In_451);
and U476 (N_476,In_183,In_146);
nor U477 (N_477,In_625,In_114);
and U478 (N_478,In_980,In_249);
and U479 (N_479,In_520,In_760);
or U480 (N_480,In_454,In_347);
and U481 (N_481,In_813,In_132);
nand U482 (N_482,In_491,In_250);
and U483 (N_483,In_100,In_299);
nand U484 (N_484,In_865,In_627);
nand U485 (N_485,In_494,In_774);
nand U486 (N_486,In_367,In_932);
nand U487 (N_487,In_308,In_981);
or U488 (N_488,In_807,In_424);
nor U489 (N_489,In_364,In_346);
nor U490 (N_490,In_466,In_248);
nand U491 (N_491,In_933,In_901);
and U492 (N_492,In_802,In_205);
or U493 (N_493,In_545,In_147);
and U494 (N_494,In_415,In_315);
nor U495 (N_495,In_426,In_702);
and U496 (N_496,In_274,In_873);
nand U497 (N_497,In_914,In_680);
or U498 (N_498,In_235,In_497);
nor U499 (N_499,In_872,In_928);
nor U500 (N_500,N_110,N_263);
and U501 (N_501,N_393,N_406);
or U502 (N_502,N_220,N_135);
and U503 (N_503,N_371,N_390);
nand U504 (N_504,N_212,N_280);
and U505 (N_505,N_158,N_317);
and U506 (N_506,N_41,N_247);
nand U507 (N_507,N_315,N_11);
and U508 (N_508,N_300,N_350);
nor U509 (N_509,N_471,N_114);
or U510 (N_510,N_225,N_454);
and U511 (N_511,N_161,N_203);
nor U512 (N_512,N_194,N_446);
and U513 (N_513,N_99,N_362);
and U514 (N_514,N_483,N_229);
or U515 (N_515,N_58,N_40);
and U516 (N_516,N_0,N_163);
or U517 (N_517,N_324,N_344);
nor U518 (N_518,N_155,N_217);
or U519 (N_519,N_295,N_189);
and U520 (N_520,N_17,N_477);
nor U521 (N_521,N_474,N_461);
nor U522 (N_522,N_417,N_166);
or U523 (N_523,N_224,N_485);
and U524 (N_524,N_381,N_146);
and U525 (N_525,N_90,N_338);
nand U526 (N_526,N_35,N_377);
nor U527 (N_527,N_388,N_195);
nand U528 (N_528,N_401,N_491);
nor U529 (N_529,N_25,N_479);
and U530 (N_530,N_379,N_361);
nand U531 (N_531,N_48,N_349);
nor U532 (N_532,N_380,N_43);
and U533 (N_533,N_357,N_70);
nand U534 (N_534,N_126,N_200);
nand U535 (N_535,N_34,N_116);
nand U536 (N_536,N_269,N_20);
nor U537 (N_537,N_258,N_308);
and U538 (N_538,N_392,N_244);
nor U539 (N_539,N_487,N_193);
and U540 (N_540,N_480,N_372);
or U541 (N_541,N_292,N_469);
or U542 (N_542,N_498,N_455);
and U543 (N_543,N_274,N_55);
nor U544 (N_544,N_142,N_249);
nand U545 (N_545,N_51,N_436);
or U546 (N_546,N_137,N_118);
or U547 (N_547,N_374,N_191);
nand U548 (N_548,N_496,N_27);
and U549 (N_549,N_10,N_196);
nand U550 (N_550,N_464,N_445);
and U551 (N_551,N_108,N_318);
nand U552 (N_552,N_78,N_298);
and U553 (N_553,N_105,N_341);
nor U554 (N_554,N_242,N_299);
nand U555 (N_555,N_138,N_275);
nand U556 (N_556,N_467,N_28);
nand U557 (N_557,N_103,N_228);
nor U558 (N_558,N_383,N_38);
nor U559 (N_559,N_345,N_325);
nor U560 (N_560,N_160,N_81);
nand U561 (N_561,N_124,N_168);
or U562 (N_562,N_321,N_53);
xnor U563 (N_563,N_184,N_231);
nand U564 (N_564,N_199,N_169);
and U565 (N_565,N_96,N_210);
nand U566 (N_566,N_227,N_452);
or U567 (N_567,N_93,N_451);
or U568 (N_568,N_470,N_165);
or U569 (N_569,N_140,N_113);
or U570 (N_570,N_282,N_171);
or U571 (N_571,N_141,N_133);
or U572 (N_572,N_433,N_444);
nand U573 (N_573,N_358,N_403);
nor U574 (N_574,N_495,N_386);
or U575 (N_575,N_475,N_230);
or U576 (N_576,N_185,N_351);
nor U577 (N_577,N_177,N_159);
nand U578 (N_578,N_6,N_175);
and U579 (N_579,N_339,N_443);
or U580 (N_580,N_164,N_482);
xor U581 (N_581,N_373,N_248);
nand U582 (N_582,N_405,N_214);
or U583 (N_583,N_156,N_281);
and U584 (N_584,N_369,N_36);
and U585 (N_585,N_77,N_296);
nand U586 (N_586,N_302,N_208);
nor U587 (N_587,N_394,N_100);
nand U588 (N_588,N_435,N_431);
nor U589 (N_589,N_422,N_365);
or U590 (N_590,N_432,N_376);
or U591 (N_591,N_347,N_205);
nor U592 (N_592,N_273,N_327);
nor U593 (N_593,N_79,N_364);
nand U594 (N_594,N_131,N_484);
nor U595 (N_595,N_162,N_62);
or U596 (N_596,N_102,N_87);
xnor U597 (N_597,N_419,N_180);
nand U598 (N_598,N_382,N_1);
nor U599 (N_599,N_286,N_490);
nand U600 (N_600,N_387,N_29);
and U601 (N_601,N_3,N_411);
nor U602 (N_602,N_219,N_143);
and U603 (N_603,N_329,N_399);
or U604 (N_604,N_288,N_328);
and U605 (N_605,N_92,N_277);
nor U606 (N_606,N_54,N_186);
or U607 (N_607,N_438,N_201);
nand U608 (N_608,N_408,N_353);
or U609 (N_609,N_427,N_215);
nor U610 (N_610,N_235,N_223);
and U611 (N_611,N_128,N_101);
nand U612 (N_612,N_190,N_416);
or U613 (N_613,N_354,N_202);
or U614 (N_614,N_398,N_64);
and U615 (N_615,N_226,N_278);
and U616 (N_616,N_197,N_154);
or U617 (N_617,N_14,N_72);
and U618 (N_618,N_236,N_303);
or U619 (N_619,N_49,N_314);
nor U620 (N_620,N_47,N_449);
nor U621 (N_621,N_346,N_237);
nor U622 (N_622,N_4,N_262);
nor U623 (N_623,N_415,N_331);
nor U624 (N_624,N_30,N_473);
and U625 (N_625,N_24,N_460);
xnor U626 (N_626,N_337,N_352);
or U627 (N_627,N_356,N_342);
nand U628 (N_628,N_333,N_499);
and U629 (N_629,N_316,N_69);
nor U630 (N_630,N_462,N_332);
or U631 (N_631,N_74,N_409);
nand U632 (N_632,N_253,N_494);
nor U633 (N_633,N_183,N_7);
nand U634 (N_634,N_111,N_82);
nand U635 (N_635,N_149,N_33);
or U636 (N_636,N_410,N_97);
nor U637 (N_637,N_239,N_213);
nor U638 (N_638,N_414,N_89);
nor U639 (N_639,N_95,N_268);
or U640 (N_640,N_57,N_170);
nor U641 (N_641,N_265,N_52);
nand U642 (N_642,N_389,N_271);
and U643 (N_643,N_366,N_463);
nor U644 (N_644,N_400,N_343);
nor U645 (N_645,N_238,N_45);
nand U646 (N_646,N_442,N_181);
and U647 (N_647,N_279,N_391);
nor U648 (N_648,N_294,N_150);
nor U649 (N_649,N_246,N_66);
nor U650 (N_650,N_39,N_428);
or U651 (N_651,N_283,N_153);
nand U652 (N_652,N_407,N_148);
nor U653 (N_653,N_285,N_234);
nand U654 (N_654,N_453,N_335);
or U655 (N_655,N_104,N_67);
nor U656 (N_656,N_221,N_91);
or U657 (N_657,N_425,N_241);
nand U658 (N_658,N_413,N_420);
and U659 (N_659,N_423,N_240);
nand U660 (N_660,N_188,N_492);
nor U661 (N_661,N_173,N_85);
nand U662 (N_662,N_59,N_172);
or U663 (N_663,N_402,N_75);
or U664 (N_664,N_115,N_9);
nand U665 (N_665,N_8,N_187);
nor U666 (N_666,N_251,N_206);
and U667 (N_667,N_478,N_472);
nand U668 (N_668,N_123,N_359);
nand U669 (N_669,N_15,N_305);
nand U670 (N_670,N_439,N_421);
nor U671 (N_671,N_145,N_290);
nor U672 (N_672,N_370,N_493);
and U673 (N_673,N_174,N_465);
nand U674 (N_674,N_243,N_254);
and U675 (N_675,N_65,N_310);
nand U676 (N_676,N_476,N_488);
nor U677 (N_677,N_264,N_232);
nor U678 (N_678,N_396,N_384);
or U679 (N_679,N_204,N_130);
or U680 (N_680,N_16,N_125);
nor U681 (N_681,N_83,N_468);
or U682 (N_682,N_157,N_21);
or U683 (N_683,N_434,N_73);
nor U684 (N_684,N_355,N_378);
and U685 (N_685,N_19,N_289);
or U686 (N_686,N_367,N_12);
nand U687 (N_687,N_129,N_151);
nand U688 (N_688,N_222,N_481);
nor U689 (N_689,N_457,N_330);
and U690 (N_690,N_192,N_5);
nor U691 (N_691,N_336,N_412);
nand U692 (N_692,N_120,N_256);
and U693 (N_693,N_31,N_80);
nand U694 (N_694,N_313,N_182);
or U695 (N_695,N_22,N_233);
nor U696 (N_696,N_56,N_136);
or U697 (N_697,N_309,N_458);
or U698 (N_698,N_257,N_301);
xor U699 (N_699,N_88,N_291);
and U700 (N_700,N_297,N_348);
xor U701 (N_701,N_84,N_178);
nand U702 (N_702,N_360,N_430);
nand U703 (N_703,N_63,N_284);
nand U704 (N_704,N_307,N_46);
nor U705 (N_705,N_429,N_447);
and U706 (N_706,N_144,N_61);
nor U707 (N_707,N_37,N_13);
nor U708 (N_708,N_385,N_76);
and U709 (N_709,N_418,N_179);
nor U710 (N_710,N_397,N_441);
or U711 (N_711,N_86,N_266);
and U712 (N_712,N_320,N_440);
nand U713 (N_713,N_198,N_147);
nand U714 (N_714,N_437,N_121);
nor U715 (N_715,N_245,N_368);
nand U716 (N_716,N_60,N_98);
or U717 (N_717,N_139,N_323);
nor U718 (N_718,N_218,N_404);
nand U719 (N_719,N_334,N_112);
nand U720 (N_720,N_255,N_132);
nor U721 (N_721,N_426,N_272);
nand U722 (N_722,N_267,N_276);
and U723 (N_723,N_107,N_32);
or U724 (N_724,N_152,N_326);
or U725 (N_725,N_71,N_68);
nor U726 (N_726,N_287,N_340);
and U727 (N_727,N_270,N_134);
nor U728 (N_728,N_119,N_306);
or U729 (N_729,N_250,N_261);
nand U730 (N_730,N_312,N_311);
nand U731 (N_731,N_18,N_94);
nand U732 (N_732,N_304,N_176);
nor U733 (N_733,N_127,N_26);
nor U734 (N_734,N_117,N_322);
nand U735 (N_735,N_209,N_216);
nand U736 (N_736,N_319,N_207);
nand U737 (N_737,N_167,N_2);
nor U738 (N_738,N_122,N_489);
nor U739 (N_739,N_260,N_375);
or U740 (N_740,N_450,N_486);
nand U741 (N_741,N_466,N_293);
nand U742 (N_742,N_44,N_363);
xor U743 (N_743,N_259,N_456);
and U744 (N_744,N_424,N_50);
nand U745 (N_745,N_497,N_23);
or U746 (N_746,N_211,N_106);
or U747 (N_747,N_109,N_459);
nand U748 (N_748,N_252,N_42);
and U749 (N_749,N_395,N_448);
or U750 (N_750,N_421,N_394);
nand U751 (N_751,N_160,N_16);
and U752 (N_752,N_207,N_64);
or U753 (N_753,N_359,N_384);
and U754 (N_754,N_374,N_168);
nor U755 (N_755,N_406,N_326);
nor U756 (N_756,N_228,N_464);
nand U757 (N_757,N_69,N_493);
and U758 (N_758,N_26,N_70);
or U759 (N_759,N_477,N_250);
nor U760 (N_760,N_318,N_485);
or U761 (N_761,N_247,N_6);
or U762 (N_762,N_130,N_485);
nand U763 (N_763,N_467,N_412);
and U764 (N_764,N_263,N_264);
or U765 (N_765,N_477,N_367);
and U766 (N_766,N_324,N_320);
or U767 (N_767,N_336,N_99);
nand U768 (N_768,N_338,N_494);
and U769 (N_769,N_391,N_39);
nor U770 (N_770,N_274,N_5);
and U771 (N_771,N_450,N_325);
nand U772 (N_772,N_337,N_213);
nor U773 (N_773,N_262,N_116);
nor U774 (N_774,N_317,N_119);
and U775 (N_775,N_383,N_309);
and U776 (N_776,N_5,N_239);
or U777 (N_777,N_28,N_299);
nand U778 (N_778,N_451,N_155);
and U779 (N_779,N_20,N_282);
or U780 (N_780,N_468,N_298);
or U781 (N_781,N_76,N_371);
nor U782 (N_782,N_186,N_235);
and U783 (N_783,N_174,N_127);
nor U784 (N_784,N_327,N_114);
and U785 (N_785,N_215,N_46);
nor U786 (N_786,N_191,N_321);
or U787 (N_787,N_122,N_312);
nor U788 (N_788,N_98,N_432);
or U789 (N_789,N_84,N_276);
xnor U790 (N_790,N_312,N_241);
and U791 (N_791,N_448,N_141);
and U792 (N_792,N_122,N_462);
nand U793 (N_793,N_39,N_443);
and U794 (N_794,N_314,N_453);
and U795 (N_795,N_409,N_298);
nor U796 (N_796,N_201,N_207);
and U797 (N_797,N_214,N_254);
or U798 (N_798,N_315,N_44);
xnor U799 (N_799,N_101,N_215);
xor U800 (N_800,N_199,N_419);
or U801 (N_801,N_449,N_124);
nand U802 (N_802,N_415,N_337);
or U803 (N_803,N_329,N_125);
nand U804 (N_804,N_322,N_343);
and U805 (N_805,N_8,N_209);
or U806 (N_806,N_438,N_46);
xor U807 (N_807,N_425,N_41);
and U808 (N_808,N_279,N_185);
and U809 (N_809,N_21,N_97);
and U810 (N_810,N_148,N_279);
or U811 (N_811,N_385,N_382);
and U812 (N_812,N_160,N_318);
nor U813 (N_813,N_316,N_363);
nor U814 (N_814,N_52,N_264);
or U815 (N_815,N_313,N_473);
or U816 (N_816,N_4,N_177);
or U817 (N_817,N_367,N_38);
nand U818 (N_818,N_26,N_47);
or U819 (N_819,N_154,N_44);
nand U820 (N_820,N_201,N_23);
nor U821 (N_821,N_135,N_496);
nor U822 (N_822,N_146,N_370);
nor U823 (N_823,N_251,N_394);
and U824 (N_824,N_147,N_312);
nand U825 (N_825,N_496,N_15);
and U826 (N_826,N_467,N_284);
nand U827 (N_827,N_107,N_24);
nand U828 (N_828,N_230,N_80);
nor U829 (N_829,N_293,N_8);
or U830 (N_830,N_146,N_136);
and U831 (N_831,N_176,N_113);
and U832 (N_832,N_169,N_88);
or U833 (N_833,N_438,N_450);
nand U834 (N_834,N_396,N_198);
and U835 (N_835,N_240,N_108);
nor U836 (N_836,N_0,N_124);
or U837 (N_837,N_436,N_83);
and U838 (N_838,N_166,N_368);
nor U839 (N_839,N_467,N_483);
nand U840 (N_840,N_315,N_161);
or U841 (N_841,N_269,N_315);
and U842 (N_842,N_204,N_416);
nand U843 (N_843,N_129,N_431);
or U844 (N_844,N_206,N_333);
nor U845 (N_845,N_443,N_86);
nand U846 (N_846,N_343,N_334);
or U847 (N_847,N_367,N_242);
nor U848 (N_848,N_344,N_71);
nor U849 (N_849,N_41,N_335);
nand U850 (N_850,N_372,N_469);
or U851 (N_851,N_142,N_364);
nor U852 (N_852,N_298,N_151);
nand U853 (N_853,N_399,N_491);
nand U854 (N_854,N_378,N_332);
and U855 (N_855,N_74,N_135);
nor U856 (N_856,N_216,N_135);
or U857 (N_857,N_89,N_126);
and U858 (N_858,N_345,N_202);
nand U859 (N_859,N_336,N_288);
nand U860 (N_860,N_432,N_195);
nor U861 (N_861,N_433,N_187);
nand U862 (N_862,N_259,N_166);
and U863 (N_863,N_89,N_152);
or U864 (N_864,N_178,N_173);
nand U865 (N_865,N_102,N_136);
nor U866 (N_866,N_67,N_309);
nor U867 (N_867,N_363,N_308);
and U868 (N_868,N_157,N_297);
or U869 (N_869,N_161,N_479);
nand U870 (N_870,N_265,N_425);
and U871 (N_871,N_179,N_72);
nor U872 (N_872,N_8,N_91);
and U873 (N_873,N_395,N_475);
or U874 (N_874,N_494,N_448);
nand U875 (N_875,N_51,N_29);
and U876 (N_876,N_116,N_305);
or U877 (N_877,N_471,N_246);
and U878 (N_878,N_25,N_214);
and U879 (N_879,N_206,N_369);
xor U880 (N_880,N_116,N_146);
nand U881 (N_881,N_119,N_49);
and U882 (N_882,N_486,N_395);
and U883 (N_883,N_360,N_453);
and U884 (N_884,N_173,N_129);
and U885 (N_885,N_411,N_368);
or U886 (N_886,N_208,N_261);
and U887 (N_887,N_221,N_151);
nand U888 (N_888,N_352,N_320);
and U889 (N_889,N_211,N_486);
nand U890 (N_890,N_60,N_141);
and U891 (N_891,N_48,N_43);
and U892 (N_892,N_89,N_83);
nand U893 (N_893,N_13,N_87);
and U894 (N_894,N_472,N_188);
nor U895 (N_895,N_214,N_383);
and U896 (N_896,N_305,N_197);
nand U897 (N_897,N_161,N_478);
nor U898 (N_898,N_357,N_225);
nor U899 (N_899,N_381,N_135);
nand U900 (N_900,N_113,N_149);
or U901 (N_901,N_303,N_154);
nor U902 (N_902,N_455,N_275);
and U903 (N_903,N_149,N_360);
or U904 (N_904,N_222,N_400);
nor U905 (N_905,N_437,N_419);
nor U906 (N_906,N_166,N_209);
and U907 (N_907,N_84,N_498);
nand U908 (N_908,N_152,N_223);
or U909 (N_909,N_209,N_147);
and U910 (N_910,N_460,N_465);
and U911 (N_911,N_337,N_229);
nand U912 (N_912,N_52,N_18);
or U913 (N_913,N_337,N_268);
nand U914 (N_914,N_480,N_22);
nor U915 (N_915,N_32,N_454);
or U916 (N_916,N_484,N_94);
nand U917 (N_917,N_419,N_189);
and U918 (N_918,N_31,N_67);
nor U919 (N_919,N_364,N_245);
or U920 (N_920,N_460,N_436);
nor U921 (N_921,N_160,N_287);
and U922 (N_922,N_370,N_347);
and U923 (N_923,N_475,N_370);
or U924 (N_924,N_396,N_481);
and U925 (N_925,N_250,N_119);
nand U926 (N_926,N_77,N_316);
or U927 (N_927,N_70,N_258);
or U928 (N_928,N_61,N_276);
nor U929 (N_929,N_31,N_468);
nor U930 (N_930,N_63,N_385);
or U931 (N_931,N_386,N_385);
or U932 (N_932,N_379,N_125);
or U933 (N_933,N_436,N_47);
nor U934 (N_934,N_197,N_461);
or U935 (N_935,N_369,N_300);
nand U936 (N_936,N_82,N_91);
or U937 (N_937,N_273,N_22);
nand U938 (N_938,N_183,N_225);
nand U939 (N_939,N_105,N_136);
and U940 (N_940,N_57,N_18);
or U941 (N_941,N_364,N_499);
nand U942 (N_942,N_455,N_8);
and U943 (N_943,N_404,N_278);
and U944 (N_944,N_81,N_47);
nor U945 (N_945,N_41,N_314);
or U946 (N_946,N_117,N_318);
and U947 (N_947,N_192,N_373);
nor U948 (N_948,N_401,N_136);
nor U949 (N_949,N_283,N_373);
nor U950 (N_950,N_7,N_61);
nor U951 (N_951,N_108,N_301);
nor U952 (N_952,N_345,N_391);
and U953 (N_953,N_336,N_436);
nand U954 (N_954,N_475,N_25);
nor U955 (N_955,N_128,N_397);
nand U956 (N_956,N_427,N_327);
or U957 (N_957,N_353,N_283);
nand U958 (N_958,N_437,N_476);
or U959 (N_959,N_316,N_72);
nand U960 (N_960,N_0,N_491);
or U961 (N_961,N_400,N_14);
and U962 (N_962,N_386,N_212);
or U963 (N_963,N_172,N_492);
xnor U964 (N_964,N_494,N_190);
or U965 (N_965,N_128,N_163);
and U966 (N_966,N_18,N_346);
nand U967 (N_967,N_374,N_156);
or U968 (N_968,N_153,N_246);
nor U969 (N_969,N_113,N_75);
or U970 (N_970,N_24,N_66);
or U971 (N_971,N_184,N_1);
nor U972 (N_972,N_258,N_140);
and U973 (N_973,N_123,N_68);
nor U974 (N_974,N_228,N_318);
nor U975 (N_975,N_174,N_34);
nand U976 (N_976,N_5,N_20);
or U977 (N_977,N_266,N_295);
nand U978 (N_978,N_134,N_316);
or U979 (N_979,N_281,N_430);
or U980 (N_980,N_189,N_223);
nor U981 (N_981,N_403,N_79);
nand U982 (N_982,N_28,N_56);
xor U983 (N_983,N_44,N_146);
and U984 (N_984,N_54,N_266);
and U985 (N_985,N_172,N_115);
and U986 (N_986,N_421,N_216);
or U987 (N_987,N_63,N_467);
nand U988 (N_988,N_355,N_351);
or U989 (N_989,N_93,N_329);
or U990 (N_990,N_51,N_371);
or U991 (N_991,N_429,N_1);
nor U992 (N_992,N_329,N_3);
nand U993 (N_993,N_371,N_55);
or U994 (N_994,N_223,N_234);
nand U995 (N_995,N_82,N_2);
nand U996 (N_996,N_466,N_194);
or U997 (N_997,N_89,N_66);
or U998 (N_998,N_239,N_82);
and U999 (N_999,N_348,N_272);
or U1000 (N_1000,N_861,N_868);
nand U1001 (N_1001,N_804,N_892);
nor U1002 (N_1002,N_936,N_932);
nor U1003 (N_1003,N_866,N_622);
nor U1004 (N_1004,N_755,N_831);
nand U1005 (N_1005,N_604,N_748);
nand U1006 (N_1006,N_606,N_642);
nand U1007 (N_1007,N_577,N_949);
or U1008 (N_1008,N_505,N_741);
nor U1009 (N_1009,N_980,N_625);
nand U1010 (N_1010,N_933,N_615);
and U1011 (N_1011,N_994,N_517);
nand U1012 (N_1012,N_734,N_706);
nor U1013 (N_1013,N_504,N_679);
or U1014 (N_1014,N_830,N_926);
nor U1015 (N_1015,N_954,N_847);
nand U1016 (N_1016,N_930,N_668);
nand U1017 (N_1017,N_662,N_888);
and U1018 (N_1018,N_685,N_514);
nand U1019 (N_1019,N_582,N_855);
and U1020 (N_1020,N_844,N_590);
nor U1021 (N_1021,N_968,N_784);
or U1022 (N_1022,N_914,N_873);
and U1023 (N_1023,N_686,N_787);
and U1024 (N_1024,N_691,N_939);
and U1025 (N_1025,N_982,N_707);
and U1026 (N_1026,N_569,N_717);
nor U1027 (N_1027,N_526,N_924);
nor U1028 (N_1028,N_780,N_798);
nor U1029 (N_1029,N_714,N_829);
and U1030 (N_1030,N_728,N_506);
and U1031 (N_1031,N_836,N_631);
nand U1032 (N_1032,N_637,N_681);
or U1033 (N_1033,N_712,N_987);
and U1034 (N_1034,N_843,N_901);
nand U1035 (N_1035,N_589,N_785);
and U1036 (N_1036,N_752,N_731);
nor U1037 (N_1037,N_733,N_689);
nand U1038 (N_1038,N_635,N_815);
and U1039 (N_1039,N_702,N_549);
nor U1040 (N_1040,N_767,N_556);
and U1041 (N_1041,N_587,N_923);
nand U1042 (N_1042,N_957,N_557);
or U1043 (N_1043,N_682,N_940);
and U1044 (N_1044,N_596,N_666);
nand U1045 (N_1045,N_769,N_974);
or U1046 (N_1046,N_793,N_657);
nand U1047 (N_1047,N_763,N_947);
nand U1048 (N_1048,N_902,N_956);
nand U1049 (N_1049,N_764,N_611);
nand U1050 (N_1050,N_634,N_906);
or U1051 (N_1051,N_789,N_975);
and U1052 (N_1052,N_656,N_953);
and U1053 (N_1053,N_903,N_768);
nand U1054 (N_1054,N_601,N_799);
nor U1055 (N_1055,N_825,N_508);
nand U1056 (N_1056,N_883,N_729);
nand U1057 (N_1057,N_701,N_553);
or U1058 (N_1058,N_951,N_651);
nand U1059 (N_1059,N_623,N_573);
or U1060 (N_1060,N_619,N_792);
nand U1061 (N_1061,N_791,N_568);
xnor U1062 (N_1062,N_925,N_661);
nand U1063 (N_1063,N_915,N_562);
nand U1064 (N_1064,N_858,N_528);
nor U1065 (N_1065,N_993,N_870);
nand U1066 (N_1066,N_718,N_943);
nor U1067 (N_1067,N_745,N_995);
and U1068 (N_1068,N_897,N_966);
or U1069 (N_1069,N_840,N_907);
nor U1070 (N_1070,N_778,N_960);
or U1071 (N_1071,N_913,N_709);
and U1072 (N_1072,N_570,N_972);
or U1073 (N_1073,N_877,N_558);
nor U1074 (N_1074,N_786,N_602);
xnor U1075 (N_1075,N_564,N_610);
and U1076 (N_1076,N_800,N_713);
and U1077 (N_1077,N_853,N_614);
nand U1078 (N_1078,N_796,N_579);
or U1079 (N_1079,N_757,N_534);
and U1080 (N_1080,N_751,N_929);
and U1081 (N_1081,N_571,N_970);
nor U1082 (N_1082,N_600,N_598);
nor U1083 (N_1083,N_979,N_884);
nor U1084 (N_1084,N_754,N_576);
and U1085 (N_1085,N_819,N_538);
nor U1086 (N_1086,N_833,N_613);
and U1087 (N_1087,N_852,N_574);
or U1088 (N_1088,N_874,N_667);
nand U1089 (N_1089,N_705,N_889);
nand U1090 (N_1090,N_524,N_758);
nor U1091 (N_1091,N_511,N_585);
nor U1092 (N_1092,N_698,N_885);
nand U1093 (N_1093,N_626,N_826);
or U1094 (N_1094,N_969,N_967);
and U1095 (N_1095,N_674,N_650);
nand U1096 (N_1096,N_919,N_802);
and U1097 (N_1097,N_869,N_854);
or U1098 (N_1098,N_981,N_565);
nand U1099 (N_1099,N_898,N_997);
nor U1100 (N_1100,N_896,N_950);
or U1101 (N_1101,N_917,N_864);
and U1102 (N_1102,N_886,N_856);
nor U1103 (N_1103,N_618,N_654);
nand U1104 (N_1104,N_964,N_620);
or U1105 (N_1105,N_921,N_990);
and U1106 (N_1106,N_742,N_737);
nand U1107 (N_1107,N_770,N_597);
nor U1108 (N_1108,N_605,N_759);
or U1109 (N_1109,N_920,N_744);
or U1110 (N_1110,N_849,N_910);
nor U1111 (N_1111,N_848,N_941);
and U1112 (N_1112,N_937,N_973);
nand U1113 (N_1113,N_665,N_663);
nor U1114 (N_1114,N_653,N_760);
nor U1115 (N_1115,N_581,N_599);
nor U1116 (N_1116,N_776,N_520);
and U1117 (N_1117,N_801,N_984);
nand U1118 (N_1118,N_961,N_648);
nand U1119 (N_1119,N_958,N_945);
nor U1120 (N_1120,N_540,N_659);
nand U1121 (N_1121,N_513,N_895);
nand U1122 (N_1122,N_697,N_783);
nor U1123 (N_1123,N_749,N_664);
nand U1124 (N_1124,N_992,N_779);
or U1125 (N_1125,N_525,N_746);
nor U1126 (N_1126,N_724,N_551);
nor U1127 (N_1127,N_814,N_880);
nor U1128 (N_1128,N_838,N_998);
nand U1129 (N_1129,N_629,N_580);
nand U1130 (N_1130,N_607,N_879);
nand U1131 (N_1131,N_908,N_593);
nand U1132 (N_1132,N_773,N_545);
nand U1133 (N_1133,N_771,N_750);
nand U1134 (N_1134,N_890,N_775);
nand U1135 (N_1135,N_916,N_716);
nor U1136 (N_1136,N_859,N_554);
nand U1137 (N_1137,N_660,N_671);
or U1138 (N_1138,N_546,N_676);
or U1139 (N_1139,N_875,N_743);
and U1140 (N_1140,N_703,N_708);
nand U1141 (N_1141,N_837,N_882);
and U1142 (N_1142,N_766,N_948);
and U1143 (N_1143,N_753,N_983);
and U1144 (N_1144,N_928,N_552);
or U1145 (N_1145,N_616,N_756);
nor U1146 (N_1146,N_516,N_946);
xor U1147 (N_1147,N_938,N_523);
nor U1148 (N_1148,N_696,N_560);
and U1149 (N_1149,N_693,N_777);
nor U1150 (N_1150,N_810,N_850);
nand U1151 (N_1151,N_730,N_677);
or U1152 (N_1152,N_872,N_539);
and U1153 (N_1153,N_781,N_699);
or U1154 (N_1154,N_911,N_658);
nand U1155 (N_1155,N_927,N_512);
nor U1156 (N_1156,N_561,N_971);
nand U1157 (N_1157,N_851,N_672);
or U1158 (N_1158,N_976,N_641);
nand U1159 (N_1159,N_559,N_627);
nand U1160 (N_1160,N_739,N_963);
nand U1161 (N_1161,N_509,N_624);
or U1162 (N_1162,N_965,N_740);
and U1163 (N_1163,N_899,N_772);
nand U1164 (N_1164,N_944,N_541);
nor U1165 (N_1165,N_846,N_527);
nor U1166 (N_1166,N_694,N_811);
or U1167 (N_1167,N_867,N_692);
or U1168 (N_1168,N_592,N_537);
nor U1169 (N_1169,N_722,N_871);
and U1170 (N_1170,N_894,N_547);
or U1171 (N_1171,N_715,N_909);
nor U1172 (N_1172,N_647,N_905);
and U1173 (N_1173,N_865,N_639);
or U1174 (N_1174,N_794,N_736);
or U1175 (N_1175,N_555,N_803);
or U1176 (N_1176,N_621,N_507);
nand U1177 (N_1177,N_841,N_824);
nor U1178 (N_1178,N_567,N_931);
nor U1179 (N_1179,N_578,N_881);
or U1180 (N_1180,N_809,N_735);
nand U1181 (N_1181,N_518,N_644);
and U1182 (N_1182,N_532,N_986);
or U1183 (N_1183,N_821,N_918);
nand U1184 (N_1184,N_649,N_529);
nand U1185 (N_1185,N_887,N_584);
nor U1186 (N_1186,N_630,N_823);
or U1187 (N_1187,N_738,N_575);
nor U1188 (N_1188,N_989,N_991);
or U1189 (N_1189,N_603,N_684);
and U1190 (N_1190,N_669,N_536);
nand U1191 (N_1191,N_594,N_727);
nand U1192 (N_1192,N_788,N_959);
nor U1193 (N_1193,N_822,N_591);
and U1194 (N_1194,N_519,N_812);
xor U1195 (N_1195,N_687,N_904);
and U1196 (N_1196,N_827,N_655);
and U1197 (N_1197,N_543,N_782);
nor U1198 (N_1198,N_863,N_818);
nand U1199 (N_1199,N_761,N_996);
or U1200 (N_1200,N_632,N_790);
nand U1201 (N_1201,N_962,N_544);
and U1202 (N_1202,N_640,N_645);
nor U1203 (N_1203,N_515,N_550);
and U1204 (N_1204,N_817,N_985);
and U1205 (N_1205,N_942,N_500);
nand U1206 (N_1206,N_617,N_900);
nand U1207 (N_1207,N_683,N_795);
xor U1208 (N_1208,N_633,N_566);
nor U1209 (N_1209,N_690,N_542);
nor U1210 (N_1210,N_502,N_710);
nand U1211 (N_1211,N_732,N_893);
or U1212 (N_1212,N_721,N_711);
nor U1213 (N_1213,N_678,N_636);
or U1214 (N_1214,N_762,N_726);
or U1215 (N_1215,N_988,N_834);
or U1216 (N_1216,N_797,N_680);
nand U1217 (N_1217,N_807,N_839);
nor U1218 (N_1218,N_588,N_832);
or U1219 (N_1219,N_548,N_719);
or U1220 (N_1220,N_934,N_595);
and U1221 (N_1221,N_725,N_586);
nand U1222 (N_1222,N_860,N_922);
and U1223 (N_1223,N_530,N_638);
nand U1224 (N_1224,N_695,N_531);
xor U1225 (N_1225,N_522,N_643);
or U1226 (N_1226,N_628,N_952);
xor U1227 (N_1227,N_572,N_955);
nand U1228 (N_1228,N_533,N_999);
nand U1229 (N_1229,N_912,N_978);
or U1230 (N_1230,N_608,N_813);
or U1231 (N_1231,N_501,N_670);
nand U1232 (N_1232,N_563,N_646);
or U1233 (N_1233,N_806,N_857);
and U1234 (N_1234,N_535,N_845);
nand U1235 (N_1235,N_935,N_688);
nand U1236 (N_1236,N_583,N_675);
nor U1237 (N_1237,N_816,N_765);
nor U1238 (N_1238,N_805,N_842);
or U1239 (N_1239,N_652,N_723);
or U1240 (N_1240,N_808,N_876);
nand U1241 (N_1241,N_835,N_891);
nand U1242 (N_1242,N_878,N_521);
nand U1243 (N_1243,N_720,N_609);
nand U1244 (N_1244,N_828,N_747);
nand U1245 (N_1245,N_673,N_704);
nor U1246 (N_1246,N_862,N_700);
nor U1247 (N_1247,N_977,N_503);
nand U1248 (N_1248,N_612,N_774);
or U1249 (N_1249,N_510,N_820);
nand U1250 (N_1250,N_911,N_590);
nand U1251 (N_1251,N_811,N_599);
nor U1252 (N_1252,N_576,N_538);
nand U1253 (N_1253,N_689,N_627);
and U1254 (N_1254,N_520,N_548);
nand U1255 (N_1255,N_811,N_981);
nor U1256 (N_1256,N_539,N_747);
nor U1257 (N_1257,N_817,N_833);
and U1258 (N_1258,N_643,N_662);
nor U1259 (N_1259,N_670,N_887);
and U1260 (N_1260,N_829,N_827);
nor U1261 (N_1261,N_545,N_795);
nand U1262 (N_1262,N_792,N_909);
and U1263 (N_1263,N_589,N_691);
nor U1264 (N_1264,N_647,N_979);
nor U1265 (N_1265,N_843,N_771);
nor U1266 (N_1266,N_580,N_916);
or U1267 (N_1267,N_761,N_681);
nand U1268 (N_1268,N_648,N_549);
nand U1269 (N_1269,N_520,N_950);
and U1270 (N_1270,N_793,N_804);
nand U1271 (N_1271,N_973,N_946);
xor U1272 (N_1272,N_507,N_642);
and U1273 (N_1273,N_565,N_838);
and U1274 (N_1274,N_936,N_955);
nor U1275 (N_1275,N_627,N_821);
or U1276 (N_1276,N_971,N_650);
and U1277 (N_1277,N_760,N_744);
nand U1278 (N_1278,N_950,N_745);
or U1279 (N_1279,N_842,N_884);
xnor U1280 (N_1280,N_855,N_780);
nand U1281 (N_1281,N_629,N_941);
or U1282 (N_1282,N_682,N_576);
and U1283 (N_1283,N_574,N_804);
or U1284 (N_1284,N_560,N_648);
nand U1285 (N_1285,N_565,N_857);
nand U1286 (N_1286,N_894,N_720);
nor U1287 (N_1287,N_588,N_720);
or U1288 (N_1288,N_547,N_983);
and U1289 (N_1289,N_682,N_772);
and U1290 (N_1290,N_681,N_858);
nor U1291 (N_1291,N_680,N_589);
or U1292 (N_1292,N_646,N_709);
nor U1293 (N_1293,N_670,N_859);
nand U1294 (N_1294,N_789,N_933);
and U1295 (N_1295,N_794,N_767);
or U1296 (N_1296,N_948,N_649);
nor U1297 (N_1297,N_816,N_661);
nand U1298 (N_1298,N_867,N_759);
nand U1299 (N_1299,N_513,N_647);
or U1300 (N_1300,N_535,N_558);
or U1301 (N_1301,N_899,N_663);
and U1302 (N_1302,N_703,N_917);
and U1303 (N_1303,N_722,N_900);
nor U1304 (N_1304,N_755,N_774);
nor U1305 (N_1305,N_701,N_759);
nand U1306 (N_1306,N_859,N_961);
or U1307 (N_1307,N_589,N_504);
or U1308 (N_1308,N_649,N_508);
nand U1309 (N_1309,N_538,N_703);
xnor U1310 (N_1310,N_666,N_765);
nor U1311 (N_1311,N_982,N_727);
or U1312 (N_1312,N_530,N_939);
or U1313 (N_1313,N_667,N_788);
nor U1314 (N_1314,N_751,N_737);
and U1315 (N_1315,N_687,N_820);
and U1316 (N_1316,N_970,N_792);
nor U1317 (N_1317,N_914,N_607);
nor U1318 (N_1318,N_970,N_889);
nor U1319 (N_1319,N_803,N_764);
and U1320 (N_1320,N_570,N_698);
nand U1321 (N_1321,N_813,N_533);
and U1322 (N_1322,N_560,N_786);
nor U1323 (N_1323,N_607,N_565);
nor U1324 (N_1324,N_982,N_731);
nor U1325 (N_1325,N_822,N_630);
or U1326 (N_1326,N_585,N_756);
and U1327 (N_1327,N_510,N_503);
nand U1328 (N_1328,N_961,N_955);
or U1329 (N_1329,N_798,N_714);
nor U1330 (N_1330,N_531,N_992);
or U1331 (N_1331,N_884,N_835);
or U1332 (N_1332,N_646,N_507);
or U1333 (N_1333,N_936,N_773);
and U1334 (N_1334,N_863,N_774);
or U1335 (N_1335,N_926,N_944);
xnor U1336 (N_1336,N_691,N_957);
and U1337 (N_1337,N_887,N_770);
and U1338 (N_1338,N_581,N_959);
nor U1339 (N_1339,N_967,N_829);
nor U1340 (N_1340,N_767,N_883);
or U1341 (N_1341,N_557,N_995);
and U1342 (N_1342,N_646,N_602);
or U1343 (N_1343,N_937,N_681);
nor U1344 (N_1344,N_952,N_937);
nor U1345 (N_1345,N_793,N_717);
and U1346 (N_1346,N_803,N_607);
nor U1347 (N_1347,N_893,N_690);
xor U1348 (N_1348,N_934,N_670);
and U1349 (N_1349,N_658,N_892);
nor U1350 (N_1350,N_713,N_513);
nor U1351 (N_1351,N_774,N_903);
and U1352 (N_1352,N_784,N_710);
nor U1353 (N_1353,N_974,N_738);
nand U1354 (N_1354,N_971,N_873);
nor U1355 (N_1355,N_996,N_833);
nand U1356 (N_1356,N_537,N_956);
or U1357 (N_1357,N_637,N_662);
nand U1358 (N_1358,N_705,N_997);
and U1359 (N_1359,N_943,N_702);
nand U1360 (N_1360,N_676,N_563);
nand U1361 (N_1361,N_567,N_661);
nand U1362 (N_1362,N_561,N_533);
and U1363 (N_1363,N_948,N_897);
or U1364 (N_1364,N_584,N_515);
nor U1365 (N_1365,N_659,N_703);
nand U1366 (N_1366,N_973,N_746);
nor U1367 (N_1367,N_675,N_733);
or U1368 (N_1368,N_572,N_616);
nor U1369 (N_1369,N_825,N_975);
and U1370 (N_1370,N_916,N_612);
nor U1371 (N_1371,N_539,N_587);
nor U1372 (N_1372,N_547,N_549);
or U1373 (N_1373,N_593,N_551);
nor U1374 (N_1374,N_626,N_778);
nand U1375 (N_1375,N_745,N_533);
and U1376 (N_1376,N_557,N_969);
or U1377 (N_1377,N_883,N_525);
nand U1378 (N_1378,N_517,N_930);
nand U1379 (N_1379,N_976,N_807);
nand U1380 (N_1380,N_949,N_897);
and U1381 (N_1381,N_575,N_860);
or U1382 (N_1382,N_937,N_903);
or U1383 (N_1383,N_912,N_907);
or U1384 (N_1384,N_672,N_981);
or U1385 (N_1385,N_693,N_947);
and U1386 (N_1386,N_870,N_689);
and U1387 (N_1387,N_825,N_941);
and U1388 (N_1388,N_500,N_512);
or U1389 (N_1389,N_526,N_832);
or U1390 (N_1390,N_723,N_977);
nor U1391 (N_1391,N_814,N_796);
or U1392 (N_1392,N_818,N_671);
nor U1393 (N_1393,N_906,N_840);
and U1394 (N_1394,N_735,N_588);
nand U1395 (N_1395,N_515,N_733);
or U1396 (N_1396,N_876,N_868);
and U1397 (N_1397,N_583,N_666);
and U1398 (N_1398,N_738,N_740);
and U1399 (N_1399,N_850,N_642);
nor U1400 (N_1400,N_946,N_559);
nand U1401 (N_1401,N_760,N_745);
xor U1402 (N_1402,N_774,N_748);
or U1403 (N_1403,N_628,N_919);
and U1404 (N_1404,N_596,N_866);
or U1405 (N_1405,N_813,N_517);
and U1406 (N_1406,N_755,N_515);
nor U1407 (N_1407,N_599,N_638);
nand U1408 (N_1408,N_760,N_896);
nand U1409 (N_1409,N_953,N_610);
nand U1410 (N_1410,N_607,N_572);
nor U1411 (N_1411,N_698,N_656);
nor U1412 (N_1412,N_758,N_777);
nor U1413 (N_1413,N_892,N_521);
or U1414 (N_1414,N_953,N_957);
nand U1415 (N_1415,N_896,N_759);
nor U1416 (N_1416,N_735,N_857);
xor U1417 (N_1417,N_926,N_920);
or U1418 (N_1418,N_670,N_879);
nor U1419 (N_1419,N_800,N_636);
xor U1420 (N_1420,N_767,N_810);
nor U1421 (N_1421,N_887,N_922);
nand U1422 (N_1422,N_907,N_660);
nor U1423 (N_1423,N_661,N_700);
or U1424 (N_1424,N_987,N_993);
nand U1425 (N_1425,N_874,N_634);
nand U1426 (N_1426,N_589,N_987);
nand U1427 (N_1427,N_525,N_796);
nand U1428 (N_1428,N_955,N_622);
and U1429 (N_1429,N_741,N_700);
nor U1430 (N_1430,N_524,N_737);
and U1431 (N_1431,N_581,N_660);
and U1432 (N_1432,N_675,N_989);
nand U1433 (N_1433,N_820,N_945);
nand U1434 (N_1434,N_983,N_597);
nor U1435 (N_1435,N_503,N_812);
nor U1436 (N_1436,N_933,N_978);
and U1437 (N_1437,N_936,N_798);
nand U1438 (N_1438,N_731,N_577);
or U1439 (N_1439,N_618,N_525);
nand U1440 (N_1440,N_797,N_508);
nor U1441 (N_1441,N_712,N_524);
xnor U1442 (N_1442,N_960,N_551);
nor U1443 (N_1443,N_972,N_669);
nand U1444 (N_1444,N_952,N_935);
nor U1445 (N_1445,N_586,N_954);
or U1446 (N_1446,N_501,N_755);
and U1447 (N_1447,N_525,N_876);
or U1448 (N_1448,N_522,N_888);
nor U1449 (N_1449,N_646,N_505);
nor U1450 (N_1450,N_650,N_788);
nor U1451 (N_1451,N_744,N_921);
or U1452 (N_1452,N_511,N_843);
nand U1453 (N_1453,N_533,N_833);
nand U1454 (N_1454,N_815,N_927);
nor U1455 (N_1455,N_778,N_794);
nor U1456 (N_1456,N_751,N_809);
nor U1457 (N_1457,N_985,N_940);
nand U1458 (N_1458,N_945,N_768);
nand U1459 (N_1459,N_813,N_996);
nor U1460 (N_1460,N_708,N_531);
nand U1461 (N_1461,N_749,N_815);
xor U1462 (N_1462,N_765,N_616);
or U1463 (N_1463,N_586,N_560);
or U1464 (N_1464,N_772,N_850);
or U1465 (N_1465,N_794,N_833);
and U1466 (N_1466,N_843,N_665);
nand U1467 (N_1467,N_733,N_905);
nand U1468 (N_1468,N_680,N_543);
or U1469 (N_1469,N_971,N_781);
nand U1470 (N_1470,N_542,N_731);
xnor U1471 (N_1471,N_672,N_989);
or U1472 (N_1472,N_869,N_510);
or U1473 (N_1473,N_662,N_920);
nand U1474 (N_1474,N_667,N_953);
nand U1475 (N_1475,N_711,N_547);
nor U1476 (N_1476,N_984,N_918);
nand U1477 (N_1477,N_526,N_862);
or U1478 (N_1478,N_847,N_553);
nor U1479 (N_1479,N_789,N_596);
nor U1480 (N_1480,N_920,N_869);
or U1481 (N_1481,N_959,N_835);
and U1482 (N_1482,N_685,N_733);
nor U1483 (N_1483,N_941,N_716);
and U1484 (N_1484,N_857,N_815);
nor U1485 (N_1485,N_925,N_667);
nor U1486 (N_1486,N_747,N_533);
and U1487 (N_1487,N_660,N_566);
nor U1488 (N_1488,N_500,N_984);
or U1489 (N_1489,N_635,N_708);
nor U1490 (N_1490,N_841,N_726);
nor U1491 (N_1491,N_526,N_704);
nand U1492 (N_1492,N_726,N_883);
nor U1493 (N_1493,N_869,N_845);
nand U1494 (N_1494,N_853,N_655);
nor U1495 (N_1495,N_833,N_749);
or U1496 (N_1496,N_562,N_894);
and U1497 (N_1497,N_700,N_888);
nor U1498 (N_1498,N_796,N_878);
or U1499 (N_1499,N_896,N_621);
nor U1500 (N_1500,N_1126,N_1215);
nor U1501 (N_1501,N_1248,N_1097);
or U1502 (N_1502,N_1310,N_1120);
or U1503 (N_1503,N_1375,N_1205);
and U1504 (N_1504,N_1137,N_1077);
or U1505 (N_1505,N_1407,N_1256);
or U1506 (N_1506,N_1087,N_1368);
and U1507 (N_1507,N_1003,N_1498);
nand U1508 (N_1508,N_1315,N_1391);
nor U1509 (N_1509,N_1383,N_1442);
and U1510 (N_1510,N_1450,N_1245);
nor U1511 (N_1511,N_1489,N_1354);
or U1512 (N_1512,N_1389,N_1240);
nand U1513 (N_1513,N_1209,N_1467);
nand U1514 (N_1514,N_1221,N_1312);
and U1515 (N_1515,N_1082,N_1365);
or U1516 (N_1516,N_1364,N_1358);
nor U1517 (N_1517,N_1011,N_1136);
nand U1518 (N_1518,N_1348,N_1193);
and U1519 (N_1519,N_1323,N_1061);
or U1520 (N_1520,N_1017,N_1283);
or U1521 (N_1521,N_1410,N_1040);
nor U1522 (N_1522,N_1438,N_1239);
and U1523 (N_1523,N_1455,N_1255);
nor U1524 (N_1524,N_1388,N_1101);
nand U1525 (N_1525,N_1491,N_1010);
nand U1526 (N_1526,N_1191,N_1385);
nor U1527 (N_1527,N_1124,N_1189);
and U1528 (N_1528,N_1357,N_1242);
nand U1529 (N_1529,N_1280,N_1028);
and U1530 (N_1530,N_1369,N_1402);
and U1531 (N_1531,N_1143,N_1400);
and U1532 (N_1532,N_1018,N_1490);
nand U1533 (N_1533,N_1133,N_1261);
nand U1534 (N_1534,N_1163,N_1452);
and U1535 (N_1535,N_1084,N_1482);
or U1536 (N_1536,N_1339,N_1381);
nand U1537 (N_1537,N_1481,N_1337);
and U1538 (N_1538,N_1433,N_1131);
or U1539 (N_1539,N_1463,N_1155);
nor U1540 (N_1540,N_1278,N_1122);
or U1541 (N_1541,N_1472,N_1457);
nor U1542 (N_1542,N_1477,N_1019);
or U1543 (N_1543,N_1401,N_1423);
nor U1544 (N_1544,N_1065,N_1178);
and U1545 (N_1545,N_1479,N_1378);
nand U1546 (N_1546,N_1192,N_1076);
nand U1547 (N_1547,N_1068,N_1217);
nand U1548 (N_1548,N_1026,N_1016);
nor U1549 (N_1549,N_1487,N_1355);
and U1550 (N_1550,N_1132,N_1092);
nor U1551 (N_1551,N_1333,N_1230);
and U1552 (N_1552,N_1259,N_1308);
nor U1553 (N_1553,N_1380,N_1089);
or U1554 (N_1554,N_1458,N_1233);
nand U1555 (N_1555,N_1246,N_1225);
or U1556 (N_1556,N_1033,N_1392);
nor U1557 (N_1557,N_1188,N_1125);
nand U1558 (N_1558,N_1220,N_1166);
or U1559 (N_1559,N_1396,N_1462);
and U1560 (N_1560,N_1000,N_1444);
nor U1561 (N_1561,N_1258,N_1447);
nand U1562 (N_1562,N_1134,N_1107);
nor U1563 (N_1563,N_1359,N_1332);
nand U1564 (N_1564,N_1446,N_1231);
nor U1565 (N_1565,N_1173,N_1409);
nor U1566 (N_1566,N_1476,N_1045);
nor U1567 (N_1567,N_1440,N_1336);
nor U1568 (N_1568,N_1063,N_1064);
nand U1569 (N_1569,N_1007,N_1275);
nand U1570 (N_1570,N_1135,N_1443);
and U1571 (N_1571,N_1198,N_1439);
nor U1572 (N_1572,N_1321,N_1214);
nand U1573 (N_1573,N_1437,N_1090);
nand U1574 (N_1574,N_1372,N_1282);
nand U1575 (N_1575,N_1024,N_1478);
and U1576 (N_1576,N_1327,N_1116);
and U1577 (N_1577,N_1432,N_1361);
and U1578 (N_1578,N_1300,N_1006);
or U1579 (N_1579,N_1460,N_1497);
or U1580 (N_1580,N_1352,N_1085);
and U1581 (N_1581,N_1121,N_1080);
or U1582 (N_1582,N_1397,N_1168);
nor U1583 (N_1583,N_1167,N_1265);
nand U1584 (N_1584,N_1043,N_1032);
nand U1585 (N_1585,N_1422,N_1203);
nand U1586 (N_1586,N_1324,N_1164);
nor U1587 (N_1587,N_1316,N_1109);
nand U1588 (N_1588,N_1334,N_1330);
nand U1589 (N_1589,N_1050,N_1022);
nand U1590 (N_1590,N_1170,N_1023);
and U1591 (N_1591,N_1343,N_1196);
or U1592 (N_1592,N_1128,N_1252);
and U1593 (N_1593,N_1474,N_1066);
nor U1594 (N_1594,N_1150,N_1073);
nor U1595 (N_1595,N_1218,N_1235);
nor U1596 (N_1596,N_1340,N_1318);
or U1597 (N_1597,N_1042,N_1495);
or U1598 (N_1598,N_1075,N_1480);
and U1599 (N_1599,N_1374,N_1186);
nor U1600 (N_1600,N_1176,N_1031);
nor U1601 (N_1601,N_1453,N_1306);
nand U1602 (N_1602,N_1058,N_1296);
nand U1603 (N_1603,N_1399,N_1053);
nand U1604 (N_1604,N_1144,N_1162);
and U1605 (N_1605,N_1456,N_1421);
or U1606 (N_1606,N_1366,N_1147);
nand U1607 (N_1607,N_1347,N_1273);
or U1608 (N_1608,N_1370,N_1108);
nand U1609 (N_1609,N_1473,N_1102);
nor U1610 (N_1610,N_1005,N_1408);
nor U1611 (N_1611,N_1349,N_1213);
nor U1612 (N_1612,N_1431,N_1057);
and U1613 (N_1613,N_1054,N_1413);
nand U1614 (N_1614,N_1140,N_1394);
and U1615 (N_1615,N_1448,N_1153);
nand U1616 (N_1616,N_1141,N_1486);
xnor U1617 (N_1617,N_1086,N_1226);
nand U1618 (N_1618,N_1160,N_1288);
nand U1619 (N_1619,N_1430,N_1158);
and U1620 (N_1620,N_1243,N_1441);
and U1621 (N_1621,N_1403,N_1048);
nor U1622 (N_1622,N_1350,N_1237);
nor U1623 (N_1623,N_1382,N_1384);
nor U1624 (N_1624,N_1184,N_1004);
nor U1625 (N_1625,N_1244,N_1099);
nand U1626 (N_1626,N_1113,N_1279);
and U1627 (N_1627,N_1103,N_1216);
nand U1628 (N_1628,N_1056,N_1062);
and U1629 (N_1629,N_1014,N_1311);
or U1630 (N_1630,N_1157,N_1183);
nand U1631 (N_1631,N_1302,N_1039);
nand U1632 (N_1632,N_1331,N_1201);
and U1633 (N_1633,N_1105,N_1274);
or U1634 (N_1634,N_1286,N_1229);
and U1635 (N_1635,N_1204,N_1284);
nor U1636 (N_1636,N_1129,N_1001);
nor U1637 (N_1637,N_1294,N_1346);
nor U1638 (N_1638,N_1414,N_1098);
and U1639 (N_1639,N_1224,N_1276);
xnor U1640 (N_1640,N_1376,N_1207);
and U1641 (N_1641,N_1379,N_1345);
or U1642 (N_1642,N_1436,N_1494);
nor U1643 (N_1643,N_1013,N_1069);
nand U1644 (N_1644,N_1094,N_1353);
or U1645 (N_1645,N_1029,N_1470);
nand U1646 (N_1646,N_1373,N_1088);
nand U1647 (N_1647,N_1325,N_1272);
nor U1648 (N_1648,N_1145,N_1428);
and U1649 (N_1649,N_1138,N_1449);
xnor U1650 (N_1650,N_1222,N_1303);
or U1651 (N_1651,N_1236,N_1371);
nor U1652 (N_1652,N_1263,N_1281);
or U1653 (N_1653,N_1367,N_1046);
or U1654 (N_1654,N_1036,N_1002);
or U1655 (N_1655,N_1172,N_1344);
nor U1656 (N_1656,N_1475,N_1074);
nor U1657 (N_1657,N_1251,N_1299);
xnor U1658 (N_1658,N_1257,N_1290);
nand U1659 (N_1659,N_1177,N_1021);
nor U1660 (N_1660,N_1268,N_1362);
or U1661 (N_1661,N_1289,N_1307);
and U1662 (N_1662,N_1484,N_1119);
and U1663 (N_1663,N_1466,N_1180);
nand U1664 (N_1664,N_1154,N_1200);
nor U1665 (N_1665,N_1227,N_1386);
and U1666 (N_1666,N_1412,N_1118);
nand U1667 (N_1667,N_1037,N_1151);
nand U1668 (N_1668,N_1406,N_1055);
xor U1669 (N_1669,N_1293,N_1052);
or U1670 (N_1670,N_1493,N_1038);
or U1671 (N_1671,N_1174,N_1059);
xnor U1672 (N_1672,N_1093,N_1020);
and U1673 (N_1673,N_1329,N_1072);
and U1674 (N_1674,N_1405,N_1291);
or U1675 (N_1675,N_1060,N_1496);
nand U1676 (N_1676,N_1030,N_1304);
and U1677 (N_1677,N_1165,N_1404);
and U1678 (N_1678,N_1210,N_1451);
and U1679 (N_1679,N_1338,N_1320);
or U1680 (N_1680,N_1335,N_1175);
and U1681 (N_1681,N_1197,N_1426);
xnor U1682 (N_1682,N_1488,N_1313);
and U1683 (N_1683,N_1083,N_1115);
or U1684 (N_1684,N_1127,N_1309);
xor U1685 (N_1685,N_1341,N_1459);
or U1686 (N_1686,N_1202,N_1418);
and U1687 (N_1687,N_1269,N_1260);
nand U1688 (N_1688,N_1499,N_1398);
nand U1689 (N_1689,N_1429,N_1254);
nor U1690 (N_1690,N_1071,N_1253);
nand U1691 (N_1691,N_1182,N_1395);
and U1692 (N_1692,N_1148,N_1195);
nand U1693 (N_1693,N_1208,N_1419);
or U1694 (N_1694,N_1425,N_1228);
nand U1695 (N_1695,N_1416,N_1483);
nand U1696 (N_1696,N_1044,N_1078);
and U1697 (N_1697,N_1305,N_1149);
nand U1698 (N_1698,N_1356,N_1110);
nor U1699 (N_1699,N_1123,N_1009);
nor U1700 (N_1700,N_1106,N_1424);
and U1701 (N_1701,N_1034,N_1464);
and U1702 (N_1702,N_1264,N_1211);
or U1703 (N_1703,N_1411,N_1100);
nor U1704 (N_1704,N_1190,N_1096);
nor U1705 (N_1705,N_1223,N_1271);
and U1706 (N_1706,N_1156,N_1298);
nor U1707 (N_1707,N_1161,N_1301);
and U1708 (N_1708,N_1465,N_1035);
nor U1709 (N_1709,N_1095,N_1212);
xor U1710 (N_1710,N_1461,N_1266);
nor U1711 (N_1711,N_1169,N_1270);
and U1712 (N_1712,N_1387,N_1250);
or U1713 (N_1713,N_1319,N_1492);
and U1714 (N_1714,N_1417,N_1130);
and U1715 (N_1715,N_1111,N_1117);
and U1716 (N_1716,N_1008,N_1326);
xor U1717 (N_1717,N_1390,N_1199);
or U1718 (N_1718,N_1393,N_1206);
nand U1719 (N_1719,N_1314,N_1171);
nand U1720 (N_1720,N_1295,N_1027);
nor U1721 (N_1721,N_1241,N_1091);
nor U1722 (N_1722,N_1360,N_1238);
nand U1723 (N_1723,N_1139,N_1179);
nand U1724 (N_1724,N_1104,N_1415);
nand U1725 (N_1725,N_1277,N_1152);
and U1726 (N_1726,N_1351,N_1469);
or U1727 (N_1727,N_1079,N_1081);
or U1728 (N_1728,N_1297,N_1445);
nor U1729 (N_1729,N_1194,N_1049);
and U1730 (N_1730,N_1485,N_1363);
nand U1731 (N_1731,N_1232,N_1051);
nor U1732 (N_1732,N_1317,N_1025);
and U1733 (N_1733,N_1187,N_1041);
nor U1734 (N_1734,N_1247,N_1287);
and U1735 (N_1735,N_1146,N_1112);
and U1736 (N_1736,N_1015,N_1219);
xnor U1737 (N_1737,N_1285,N_1471);
nor U1738 (N_1738,N_1070,N_1267);
or U1739 (N_1739,N_1047,N_1420);
nor U1740 (N_1740,N_1142,N_1377);
or U1741 (N_1741,N_1434,N_1159);
and U1742 (N_1742,N_1185,N_1435);
nor U1743 (N_1743,N_1234,N_1012);
or U1744 (N_1744,N_1181,N_1342);
nor U1745 (N_1745,N_1427,N_1454);
and U1746 (N_1746,N_1328,N_1114);
nand U1747 (N_1747,N_1067,N_1262);
xor U1748 (N_1748,N_1322,N_1249);
or U1749 (N_1749,N_1292,N_1468);
and U1750 (N_1750,N_1287,N_1421);
nand U1751 (N_1751,N_1190,N_1380);
and U1752 (N_1752,N_1179,N_1003);
or U1753 (N_1753,N_1354,N_1265);
nand U1754 (N_1754,N_1295,N_1312);
nor U1755 (N_1755,N_1427,N_1253);
nor U1756 (N_1756,N_1134,N_1498);
and U1757 (N_1757,N_1201,N_1130);
and U1758 (N_1758,N_1351,N_1385);
nand U1759 (N_1759,N_1494,N_1310);
nor U1760 (N_1760,N_1092,N_1425);
or U1761 (N_1761,N_1014,N_1135);
and U1762 (N_1762,N_1359,N_1387);
nor U1763 (N_1763,N_1461,N_1119);
xor U1764 (N_1764,N_1236,N_1493);
nand U1765 (N_1765,N_1389,N_1373);
nor U1766 (N_1766,N_1476,N_1100);
or U1767 (N_1767,N_1077,N_1189);
or U1768 (N_1768,N_1203,N_1180);
and U1769 (N_1769,N_1344,N_1434);
nor U1770 (N_1770,N_1365,N_1330);
or U1771 (N_1771,N_1465,N_1267);
and U1772 (N_1772,N_1275,N_1207);
or U1773 (N_1773,N_1411,N_1343);
nand U1774 (N_1774,N_1470,N_1348);
or U1775 (N_1775,N_1191,N_1158);
nand U1776 (N_1776,N_1395,N_1163);
nand U1777 (N_1777,N_1110,N_1111);
or U1778 (N_1778,N_1162,N_1169);
nor U1779 (N_1779,N_1384,N_1073);
or U1780 (N_1780,N_1142,N_1435);
nand U1781 (N_1781,N_1052,N_1386);
nand U1782 (N_1782,N_1258,N_1095);
or U1783 (N_1783,N_1453,N_1330);
or U1784 (N_1784,N_1066,N_1273);
nand U1785 (N_1785,N_1040,N_1394);
nand U1786 (N_1786,N_1377,N_1380);
nand U1787 (N_1787,N_1044,N_1111);
xor U1788 (N_1788,N_1443,N_1253);
nand U1789 (N_1789,N_1157,N_1258);
nand U1790 (N_1790,N_1297,N_1394);
nand U1791 (N_1791,N_1384,N_1219);
and U1792 (N_1792,N_1016,N_1462);
nor U1793 (N_1793,N_1370,N_1291);
or U1794 (N_1794,N_1188,N_1142);
and U1795 (N_1795,N_1333,N_1004);
nand U1796 (N_1796,N_1298,N_1040);
nand U1797 (N_1797,N_1056,N_1389);
and U1798 (N_1798,N_1275,N_1204);
and U1799 (N_1799,N_1477,N_1319);
or U1800 (N_1800,N_1458,N_1032);
nand U1801 (N_1801,N_1219,N_1001);
and U1802 (N_1802,N_1035,N_1349);
nand U1803 (N_1803,N_1137,N_1092);
nand U1804 (N_1804,N_1041,N_1481);
nor U1805 (N_1805,N_1394,N_1447);
nand U1806 (N_1806,N_1311,N_1312);
or U1807 (N_1807,N_1342,N_1187);
nand U1808 (N_1808,N_1346,N_1359);
or U1809 (N_1809,N_1103,N_1235);
or U1810 (N_1810,N_1436,N_1272);
or U1811 (N_1811,N_1024,N_1017);
xnor U1812 (N_1812,N_1215,N_1347);
nand U1813 (N_1813,N_1235,N_1387);
nor U1814 (N_1814,N_1419,N_1375);
nand U1815 (N_1815,N_1057,N_1213);
nand U1816 (N_1816,N_1083,N_1350);
and U1817 (N_1817,N_1450,N_1066);
nand U1818 (N_1818,N_1442,N_1021);
and U1819 (N_1819,N_1379,N_1019);
nand U1820 (N_1820,N_1366,N_1271);
nor U1821 (N_1821,N_1356,N_1369);
or U1822 (N_1822,N_1416,N_1053);
and U1823 (N_1823,N_1488,N_1449);
or U1824 (N_1824,N_1134,N_1296);
and U1825 (N_1825,N_1126,N_1314);
or U1826 (N_1826,N_1347,N_1341);
and U1827 (N_1827,N_1138,N_1108);
nand U1828 (N_1828,N_1346,N_1456);
nand U1829 (N_1829,N_1244,N_1357);
nand U1830 (N_1830,N_1210,N_1149);
nand U1831 (N_1831,N_1019,N_1060);
nand U1832 (N_1832,N_1358,N_1206);
or U1833 (N_1833,N_1291,N_1162);
or U1834 (N_1834,N_1392,N_1051);
nand U1835 (N_1835,N_1123,N_1440);
or U1836 (N_1836,N_1070,N_1355);
or U1837 (N_1837,N_1165,N_1337);
or U1838 (N_1838,N_1248,N_1032);
nand U1839 (N_1839,N_1429,N_1104);
nand U1840 (N_1840,N_1376,N_1173);
or U1841 (N_1841,N_1366,N_1426);
or U1842 (N_1842,N_1381,N_1008);
or U1843 (N_1843,N_1302,N_1219);
nand U1844 (N_1844,N_1130,N_1129);
and U1845 (N_1845,N_1460,N_1353);
nand U1846 (N_1846,N_1182,N_1269);
nand U1847 (N_1847,N_1186,N_1167);
nor U1848 (N_1848,N_1000,N_1375);
nand U1849 (N_1849,N_1043,N_1063);
nor U1850 (N_1850,N_1295,N_1066);
nor U1851 (N_1851,N_1291,N_1358);
or U1852 (N_1852,N_1355,N_1245);
or U1853 (N_1853,N_1052,N_1241);
nor U1854 (N_1854,N_1181,N_1091);
nor U1855 (N_1855,N_1171,N_1305);
or U1856 (N_1856,N_1249,N_1031);
or U1857 (N_1857,N_1071,N_1082);
nor U1858 (N_1858,N_1235,N_1211);
nor U1859 (N_1859,N_1229,N_1432);
or U1860 (N_1860,N_1273,N_1477);
and U1861 (N_1861,N_1439,N_1024);
or U1862 (N_1862,N_1379,N_1435);
nand U1863 (N_1863,N_1398,N_1482);
or U1864 (N_1864,N_1195,N_1354);
and U1865 (N_1865,N_1409,N_1040);
nand U1866 (N_1866,N_1093,N_1428);
nor U1867 (N_1867,N_1100,N_1382);
xnor U1868 (N_1868,N_1111,N_1446);
nor U1869 (N_1869,N_1212,N_1143);
and U1870 (N_1870,N_1274,N_1460);
and U1871 (N_1871,N_1114,N_1322);
nand U1872 (N_1872,N_1140,N_1465);
nand U1873 (N_1873,N_1375,N_1036);
nand U1874 (N_1874,N_1058,N_1307);
nand U1875 (N_1875,N_1473,N_1095);
and U1876 (N_1876,N_1188,N_1369);
nand U1877 (N_1877,N_1225,N_1028);
or U1878 (N_1878,N_1415,N_1010);
nand U1879 (N_1879,N_1478,N_1129);
nor U1880 (N_1880,N_1293,N_1054);
nor U1881 (N_1881,N_1479,N_1056);
or U1882 (N_1882,N_1316,N_1343);
nand U1883 (N_1883,N_1000,N_1396);
nand U1884 (N_1884,N_1458,N_1230);
nor U1885 (N_1885,N_1162,N_1053);
xnor U1886 (N_1886,N_1137,N_1091);
and U1887 (N_1887,N_1416,N_1277);
and U1888 (N_1888,N_1318,N_1358);
nand U1889 (N_1889,N_1319,N_1378);
nand U1890 (N_1890,N_1068,N_1082);
or U1891 (N_1891,N_1348,N_1011);
or U1892 (N_1892,N_1174,N_1332);
nor U1893 (N_1893,N_1189,N_1393);
and U1894 (N_1894,N_1389,N_1459);
nor U1895 (N_1895,N_1405,N_1184);
nor U1896 (N_1896,N_1354,N_1073);
nand U1897 (N_1897,N_1058,N_1295);
nand U1898 (N_1898,N_1241,N_1409);
nand U1899 (N_1899,N_1369,N_1270);
nor U1900 (N_1900,N_1280,N_1404);
nand U1901 (N_1901,N_1159,N_1096);
nand U1902 (N_1902,N_1402,N_1006);
or U1903 (N_1903,N_1443,N_1435);
or U1904 (N_1904,N_1120,N_1112);
nor U1905 (N_1905,N_1302,N_1325);
and U1906 (N_1906,N_1292,N_1236);
or U1907 (N_1907,N_1013,N_1459);
nand U1908 (N_1908,N_1397,N_1003);
and U1909 (N_1909,N_1495,N_1118);
nand U1910 (N_1910,N_1440,N_1286);
and U1911 (N_1911,N_1262,N_1109);
nand U1912 (N_1912,N_1483,N_1460);
or U1913 (N_1913,N_1289,N_1081);
and U1914 (N_1914,N_1022,N_1409);
and U1915 (N_1915,N_1421,N_1005);
nor U1916 (N_1916,N_1484,N_1476);
or U1917 (N_1917,N_1412,N_1345);
or U1918 (N_1918,N_1394,N_1465);
or U1919 (N_1919,N_1477,N_1499);
nor U1920 (N_1920,N_1336,N_1124);
and U1921 (N_1921,N_1059,N_1484);
or U1922 (N_1922,N_1110,N_1380);
or U1923 (N_1923,N_1347,N_1390);
nor U1924 (N_1924,N_1057,N_1095);
or U1925 (N_1925,N_1388,N_1389);
or U1926 (N_1926,N_1265,N_1388);
and U1927 (N_1927,N_1221,N_1030);
or U1928 (N_1928,N_1033,N_1363);
nand U1929 (N_1929,N_1298,N_1013);
and U1930 (N_1930,N_1248,N_1219);
nand U1931 (N_1931,N_1445,N_1494);
or U1932 (N_1932,N_1118,N_1434);
xnor U1933 (N_1933,N_1147,N_1238);
nor U1934 (N_1934,N_1163,N_1336);
nor U1935 (N_1935,N_1071,N_1320);
nand U1936 (N_1936,N_1461,N_1138);
nor U1937 (N_1937,N_1487,N_1310);
and U1938 (N_1938,N_1300,N_1067);
and U1939 (N_1939,N_1482,N_1473);
nor U1940 (N_1940,N_1145,N_1017);
and U1941 (N_1941,N_1374,N_1453);
nand U1942 (N_1942,N_1419,N_1418);
or U1943 (N_1943,N_1259,N_1254);
and U1944 (N_1944,N_1024,N_1259);
nand U1945 (N_1945,N_1144,N_1368);
or U1946 (N_1946,N_1336,N_1000);
nor U1947 (N_1947,N_1268,N_1020);
or U1948 (N_1948,N_1318,N_1105);
nor U1949 (N_1949,N_1349,N_1443);
or U1950 (N_1950,N_1177,N_1248);
nor U1951 (N_1951,N_1254,N_1077);
or U1952 (N_1952,N_1168,N_1013);
nor U1953 (N_1953,N_1276,N_1140);
or U1954 (N_1954,N_1069,N_1407);
and U1955 (N_1955,N_1197,N_1488);
nand U1956 (N_1956,N_1476,N_1498);
or U1957 (N_1957,N_1147,N_1241);
nand U1958 (N_1958,N_1154,N_1314);
and U1959 (N_1959,N_1035,N_1267);
and U1960 (N_1960,N_1012,N_1277);
nand U1961 (N_1961,N_1026,N_1137);
nor U1962 (N_1962,N_1024,N_1070);
nor U1963 (N_1963,N_1464,N_1297);
and U1964 (N_1964,N_1067,N_1220);
nor U1965 (N_1965,N_1258,N_1036);
nand U1966 (N_1966,N_1184,N_1303);
or U1967 (N_1967,N_1248,N_1066);
nor U1968 (N_1968,N_1267,N_1216);
nor U1969 (N_1969,N_1066,N_1349);
nand U1970 (N_1970,N_1418,N_1046);
or U1971 (N_1971,N_1407,N_1116);
or U1972 (N_1972,N_1357,N_1389);
nor U1973 (N_1973,N_1282,N_1103);
or U1974 (N_1974,N_1265,N_1427);
or U1975 (N_1975,N_1298,N_1286);
nand U1976 (N_1976,N_1319,N_1427);
or U1977 (N_1977,N_1234,N_1423);
nor U1978 (N_1978,N_1297,N_1258);
or U1979 (N_1979,N_1144,N_1495);
and U1980 (N_1980,N_1259,N_1059);
nor U1981 (N_1981,N_1105,N_1494);
nor U1982 (N_1982,N_1479,N_1055);
and U1983 (N_1983,N_1437,N_1171);
and U1984 (N_1984,N_1001,N_1007);
or U1985 (N_1985,N_1067,N_1431);
nor U1986 (N_1986,N_1472,N_1355);
nor U1987 (N_1987,N_1329,N_1057);
or U1988 (N_1988,N_1007,N_1321);
or U1989 (N_1989,N_1251,N_1375);
and U1990 (N_1990,N_1186,N_1201);
and U1991 (N_1991,N_1264,N_1145);
or U1992 (N_1992,N_1444,N_1355);
and U1993 (N_1993,N_1066,N_1151);
and U1994 (N_1994,N_1461,N_1349);
or U1995 (N_1995,N_1144,N_1203);
nand U1996 (N_1996,N_1296,N_1261);
and U1997 (N_1997,N_1037,N_1053);
xnor U1998 (N_1998,N_1426,N_1388);
or U1999 (N_1999,N_1413,N_1192);
or U2000 (N_2000,N_1643,N_1733);
or U2001 (N_2001,N_1908,N_1925);
and U2002 (N_2002,N_1566,N_1957);
or U2003 (N_2003,N_1800,N_1633);
nor U2004 (N_2004,N_1543,N_1847);
or U2005 (N_2005,N_1831,N_1690);
or U2006 (N_2006,N_1639,N_1801);
or U2007 (N_2007,N_1828,N_1877);
nor U2008 (N_2008,N_1568,N_1616);
nor U2009 (N_2009,N_1506,N_1587);
nor U2010 (N_2010,N_1897,N_1960);
nand U2011 (N_2011,N_1588,N_1868);
or U2012 (N_2012,N_1597,N_1786);
or U2013 (N_2013,N_1958,N_1904);
or U2014 (N_2014,N_1551,N_1905);
xnor U2015 (N_2015,N_1559,N_1640);
nor U2016 (N_2016,N_1554,N_1522);
and U2017 (N_2017,N_1656,N_1624);
nand U2018 (N_2018,N_1818,N_1862);
nor U2019 (N_2019,N_1684,N_1758);
and U2020 (N_2020,N_1713,N_1557);
or U2021 (N_2021,N_1726,N_1714);
or U2022 (N_2022,N_1542,N_1707);
and U2023 (N_2023,N_1916,N_1553);
and U2024 (N_2024,N_1832,N_1665);
or U2025 (N_2025,N_1621,N_1744);
and U2026 (N_2026,N_1547,N_1924);
nand U2027 (N_2027,N_1914,N_1545);
nor U2028 (N_2028,N_1569,N_1702);
and U2029 (N_2029,N_1515,N_1693);
nand U2030 (N_2030,N_1647,N_1892);
nand U2031 (N_2031,N_1798,N_1792);
nand U2032 (N_2032,N_1748,N_1951);
nor U2033 (N_2033,N_1963,N_1876);
nand U2034 (N_2034,N_1563,N_1606);
nor U2035 (N_2035,N_1909,N_1926);
nand U2036 (N_2036,N_1592,N_1980);
and U2037 (N_2037,N_1612,N_1580);
or U2038 (N_2038,N_1516,N_1885);
and U2039 (N_2039,N_1536,N_1835);
or U2040 (N_2040,N_1986,N_1583);
nor U2041 (N_2041,N_1556,N_1803);
and U2042 (N_2042,N_1742,N_1760);
or U2043 (N_2043,N_1562,N_1988);
nand U2044 (N_2044,N_1799,N_1692);
nor U2045 (N_2045,N_1768,N_1864);
and U2046 (N_2046,N_1593,N_1519);
xnor U2047 (N_2047,N_1991,N_1802);
and U2048 (N_2048,N_1823,N_1763);
and U2049 (N_2049,N_1718,N_1765);
nor U2050 (N_2050,N_1687,N_1791);
nor U2051 (N_2051,N_1699,N_1708);
nor U2052 (N_2052,N_1977,N_1810);
or U2053 (N_2053,N_1975,N_1852);
nand U2054 (N_2054,N_1788,N_1603);
or U2055 (N_2055,N_1922,N_1691);
nand U2056 (N_2056,N_1739,N_1659);
and U2057 (N_2057,N_1648,N_1664);
nor U2058 (N_2058,N_1895,N_1590);
or U2059 (N_2059,N_1777,N_1900);
and U2060 (N_2060,N_1564,N_1584);
or U2061 (N_2061,N_1613,N_1837);
nor U2062 (N_2062,N_1710,N_1813);
or U2063 (N_2063,N_1513,N_1928);
and U2064 (N_2064,N_1662,N_1622);
and U2065 (N_2065,N_1582,N_1577);
or U2066 (N_2066,N_1842,N_1652);
and U2067 (N_2067,N_1517,N_1682);
nand U2068 (N_2068,N_1673,N_1887);
nand U2069 (N_2069,N_1504,N_1911);
xnor U2070 (N_2070,N_1781,N_1761);
and U2071 (N_2071,N_1934,N_1981);
nor U2072 (N_2072,N_1598,N_1944);
or U2073 (N_2073,N_1734,N_1697);
or U2074 (N_2074,N_1610,N_1931);
and U2075 (N_2075,N_1759,N_1881);
and U2076 (N_2076,N_1782,N_1848);
and U2077 (N_2077,N_1548,N_1851);
or U2078 (N_2078,N_1555,N_1970);
and U2079 (N_2079,N_1880,N_1669);
nand U2080 (N_2080,N_1956,N_1722);
xnor U2081 (N_2081,N_1838,N_1634);
and U2082 (N_2082,N_1965,N_1663);
nor U2083 (N_2083,N_1997,N_1626);
or U2084 (N_2084,N_1749,N_1844);
nand U2085 (N_2085,N_1537,N_1780);
and U2086 (N_2086,N_1968,N_1787);
or U2087 (N_2087,N_1561,N_1821);
and U2088 (N_2088,N_1833,N_1525);
or U2089 (N_2089,N_1755,N_1503);
nor U2090 (N_2090,N_1609,N_1694);
nor U2091 (N_2091,N_1632,N_1841);
nand U2092 (N_2092,N_1771,N_1716);
nor U2093 (N_2093,N_1910,N_1962);
nand U2094 (N_2094,N_1972,N_1620);
nor U2095 (N_2095,N_1964,N_1989);
xor U2096 (N_2096,N_1874,N_1945);
or U2097 (N_2097,N_1888,N_1933);
nand U2098 (N_2098,N_1521,N_1510);
nand U2099 (N_2099,N_1701,N_1614);
or U2100 (N_2100,N_1839,N_1549);
and U2101 (N_2101,N_1501,N_1947);
xnor U2102 (N_2102,N_1608,N_1820);
or U2103 (N_2103,N_1657,N_1976);
nand U2104 (N_2104,N_1974,N_1658);
nand U2105 (N_2105,N_1856,N_1853);
nor U2106 (N_2106,N_1756,N_1752);
nand U2107 (N_2107,N_1539,N_1567);
or U2108 (N_2108,N_1688,N_1811);
nor U2109 (N_2109,N_1967,N_1732);
nor U2110 (N_2110,N_1772,N_1825);
nor U2111 (N_2111,N_1937,N_1990);
or U2112 (N_2112,N_1731,N_1611);
and U2113 (N_2113,N_1923,N_1952);
nor U2114 (N_2114,N_1858,N_1953);
and U2115 (N_2115,N_1829,N_1578);
or U2116 (N_2116,N_1660,N_1630);
or U2117 (N_2117,N_1637,N_1779);
nand U2118 (N_2118,N_1942,N_1689);
nor U2119 (N_2119,N_1894,N_1747);
and U2120 (N_2120,N_1999,N_1604);
nor U2121 (N_2121,N_1720,N_1745);
nor U2122 (N_2122,N_1625,N_1729);
nor U2123 (N_2123,N_1954,N_1532);
and U2124 (N_2124,N_1783,N_1629);
nor U2125 (N_2125,N_1906,N_1985);
or U2126 (N_2126,N_1635,N_1861);
nand U2127 (N_2127,N_1645,N_1959);
nor U2128 (N_2128,N_1676,N_1873);
or U2129 (N_2129,N_1882,N_1715);
nand U2130 (N_2130,N_1601,N_1751);
nand U2131 (N_2131,N_1767,N_1793);
nand U2132 (N_2132,N_1642,N_1631);
nor U2133 (N_2133,N_1845,N_1875);
nor U2134 (N_2134,N_1785,N_1995);
and U2135 (N_2135,N_1889,N_1675);
nand U2136 (N_2136,N_1698,N_1728);
nor U2137 (N_2137,N_1738,N_1737);
or U2138 (N_2138,N_1773,N_1512);
nor U2139 (N_2139,N_1753,N_1508);
nor U2140 (N_2140,N_1654,N_1600);
nor U2141 (N_2141,N_1514,N_1843);
nor U2142 (N_2142,N_1903,N_1819);
and U2143 (N_2143,N_1533,N_1619);
or U2144 (N_2144,N_1769,N_1849);
or U2145 (N_2145,N_1860,N_1949);
and U2146 (N_2146,N_1774,N_1917);
or U2147 (N_2147,N_1727,N_1719);
or U2148 (N_2148,N_1794,N_1840);
nor U2149 (N_2149,N_1824,N_1526);
or U2150 (N_2150,N_1850,N_1796);
nand U2151 (N_2151,N_1834,N_1987);
nand U2152 (N_2152,N_1636,N_1594);
nand U2153 (N_2153,N_1581,N_1700);
or U2154 (N_2154,N_1816,N_1921);
or U2155 (N_2155,N_1983,N_1805);
or U2156 (N_2156,N_1721,N_1867);
nand U2157 (N_2157,N_1929,N_1705);
nor U2158 (N_2158,N_1570,N_1685);
and U2159 (N_2159,N_1735,N_1961);
and U2160 (N_2160,N_1898,N_1878);
or U2161 (N_2161,N_1661,N_1674);
or U2162 (N_2162,N_1886,N_1530);
nor U2163 (N_2163,N_1671,N_1871);
nand U2164 (N_2164,N_1940,N_1695);
nor U2165 (N_2165,N_1591,N_1511);
nand U2166 (N_2166,N_1969,N_1935);
nand U2167 (N_2167,N_1529,N_1520);
and U2168 (N_2168,N_1883,N_1984);
nand U2169 (N_2169,N_1650,N_1724);
or U2170 (N_2170,N_1750,N_1681);
and U2171 (N_2171,N_1507,N_1891);
nand U2172 (N_2172,N_1927,N_1994);
nand U2173 (N_2173,N_1730,N_1915);
or U2174 (N_2174,N_1740,N_1943);
or U2175 (N_2175,N_1797,N_1854);
or U2176 (N_2176,N_1950,N_1572);
or U2177 (N_2177,N_1743,N_1599);
nand U2178 (N_2178,N_1778,N_1930);
nor U2179 (N_2179,N_1683,N_1736);
and U2180 (N_2180,N_1919,N_1766);
nor U2181 (N_2181,N_1540,N_1560);
or U2182 (N_2182,N_1941,N_1884);
or U2183 (N_2183,N_1527,N_1576);
or U2184 (N_2184,N_1672,N_1955);
or U2185 (N_2185,N_1741,N_1509);
or U2186 (N_2186,N_1920,N_1998);
nand U2187 (N_2187,N_1649,N_1896);
nor U2188 (N_2188,N_1535,N_1806);
nor U2189 (N_2189,N_1706,N_1946);
or U2190 (N_2190,N_1971,N_1826);
nor U2191 (N_2191,N_1901,N_1615);
nor U2192 (N_2192,N_1596,N_1807);
or U2193 (N_2193,N_1565,N_1523);
nand U2194 (N_2194,N_1531,N_1541);
or U2195 (N_2195,N_1809,N_1872);
and U2196 (N_2196,N_1667,N_1812);
nor U2197 (N_2197,N_1836,N_1764);
nor U2198 (N_2198,N_1703,N_1680);
and U2199 (N_2199,N_1717,N_1973);
nor U2200 (N_2200,N_1817,N_1846);
and U2201 (N_2201,N_1770,N_1863);
and U2202 (N_2202,N_1754,N_1666);
nand U2203 (N_2203,N_1586,N_1938);
and U2204 (N_2204,N_1879,N_1538);
xor U2205 (N_2205,N_1651,N_1890);
nor U2206 (N_2206,N_1869,N_1932);
and U2207 (N_2207,N_1762,N_1679);
or U2208 (N_2208,N_1912,N_1830);
and U2209 (N_2209,N_1776,N_1804);
or U2210 (N_2210,N_1712,N_1678);
or U2211 (N_2211,N_1709,N_1544);
nor U2212 (N_2212,N_1696,N_1686);
or U2213 (N_2213,N_1618,N_1757);
nor U2214 (N_2214,N_1996,N_1589);
or U2215 (N_2215,N_1870,N_1505);
nor U2216 (N_2216,N_1902,N_1628);
or U2217 (N_2217,N_1670,N_1574);
nand U2218 (N_2218,N_1808,N_1641);
nand U2219 (N_2219,N_1502,N_1907);
nand U2220 (N_2220,N_1585,N_1605);
or U2221 (N_2221,N_1865,N_1866);
nor U2222 (N_2222,N_1795,N_1575);
nor U2223 (N_2223,N_1855,N_1723);
nand U2224 (N_2224,N_1982,N_1775);
or U2225 (N_2225,N_1534,N_1993);
nand U2226 (N_2226,N_1859,N_1966);
and U2227 (N_2227,N_1579,N_1725);
or U2228 (N_2228,N_1827,N_1711);
nand U2229 (N_2229,N_1546,N_1668);
nand U2230 (N_2230,N_1815,N_1913);
or U2231 (N_2231,N_1638,N_1992);
and U2232 (N_2232,N_1518,N_1746);
or U2233 (N_2233,N_1500,N_1644);
nor U2234 (N_2234,N_1573,N_1571);
nand U2235 (N_2235,N_1978,N_1939);
or U2236 (N_2236,N_1948,N_1789);
nand U2237 (N_2237,N_1524,N_1784);
nand U2238 (N_2238,N_1558,N_1655);
or U2239 (N_2239,N_1646,N_1528);
nor U2240 (N_2240,N_1822,N_1653);
or U2241 (N_2241,N_1595,N_1857);
xor U2242 (N_2242,N_1623,N_1550);
nand U2243 (N_2243,N_1704,N_1677);
or U2244 (N_2244,N_1607,N_1617);
or U2245 (N_2245,N_1602,N_1814);
nor U2246 (N_2246,N_1936,N_1627);
nor U2247 (N_2247,N_1918,N_1979);
and U2248 (N_2248,N_1552,N_1893);
nor U2249 (N_2249,N_1899,N_1790);
and U2250 (N_2250,N_1714,N_1772);
or U2251 (N_2251,N_1683,N_1794);
and U2252 (N_2252,N_1627,N_1923);
nor U2253 (N_2253,N_1700,N_1800);
nor U2254 (N_2254,N_1780,N_1504);
and U2255 (N_2255,N_1768,N_1665);
or U2256 (N_2256,N_1698,N_1765);
and U2257 (N_2257,N_1763,N_1717);
or U2258 (N_2258,N_1804,N_1702);
nand U2259 (N_2259,N_1723,N_1563);
nand U2260 (N_2260,N_1826,N_1633);
nor U2261 (N_2261,N_1673,N_1821);
xor U2262 (N_2262,N_1667,N_1879);
nand U2263 (N_2263,N_1654,N_1918);
xor U2264 (N_2264,N_1512,N_1827);
nor U2265 (N_2265,N_1918,N_1949);
or U2266 (N_2266,N_1643,N_1716);
nor U2267 (N_2267,N_1615,N_1720);
nor U2268 (N_2268,N_1921,N_1866);
or U2269 (N_2269,N_1800,N_1942);
and U2270 (N_2270,N_1789,N_1816);
and U2271 (N_2271,N_1547,N_1669);
or U2272 (N_2272,N_1581,N_1863);
and U2273 (N_2273,N_1658,N_1828);
nor U2274 (N_2274,N_1880,N_1842);
or U2275 (N_2275,N_1717,N_1693);
or U2276 (N_2276,N_1853,N_1898);
nand U2277 (N_2277,N_1618,N_1522);
nor U2278 (N_2278,N_1541,N_1589);
and U2279 (N_2279,N_1712,N_1689);
nand U2280 (N_2280,N_1622,N_1817);
or U2281 (N_2281,N_1736,N_1805);
nor U2282 (N_2282,N_1805,N_1952);
or U2283 (N_2283,N_1805,N_1786);
and U2284 (N_2284,N_1652,N_1597);
nor U2285 (N_2285,N_1773,N_1582);
nand U2286 (N_2286,N_1962,N_1500);
and U2287 (N_2287,N_1582,N_1526);
or U2288 (N_2288,N_1909,N_1617);
nor U2289 (N_2289,N_1926,N_1696);
and U2290 (N_2290,N_1680,N_1985);
xor U2291 (N_2291,N_1967,N_1573);
and U2292 (N_2292,N_1831,N_1898);
nand U2293 (N_2293,N_1815,N_1923);
nand U2294 (N_2294,N_1942,N_1982);
xor U2295 (N_2295,N_1669,N_1876);
nand U2296 (N_2296,N_1717,N_1729);
xor U2297 (N_2297,N_1941,N_1953);
nor U2298 (N_2298,N_1595,N_1911);
nor U2299 (N_2299,N_1875,N_1634);
and U2300 (N_2300,N_1655,N_1724);
nor U2301 (N_2301,N_1572,N_1978);
nor U2302 (N_2302,N_1801,N_1539);
xnor U2303 (N_2303,N_1887,N_1798);
nand U2304 (N_2304,N_1928,N_1559);
nand U2305 (N_2305,N_1941,N_1513);
or U2306 (N_2306,N_1632,N_1963);
and U2307 (N_2307,N_1609,N_1783);
and U2308 (N_2308,N_1707,N_1888);
xnor U2309 (N_2309,N_1719,N_1588);
xnor U2310 (N_2310,N_1832,N_1827);
nand U2311 (N_2311,N_1935,N_1743);
nand U2312 (N_2312,N_1718,N_1850);
nand U2313 (N_2313,N_1675,N_1568);
and U2314 (N_2314,N_1911,N_1628);
or U2315 (N_2315,N_1700,N_1677);
and U2316 (N_2316,N_1592,N_1875);
nand U2317 (N_2317,N_1855,N_1825);
nand U2318 (N_2318,N_1954,N_1993);
nand U2319 (N_2319,N_1961,N_1746);
nor U2320 (N_2320,N_1596,N_1862);
nand U2321 (N_2321,N_1609,N_1644);
or U2322 (N_2322,N_1534,N_1919);
or U2323 (N_2323,N_1703,N_1927);
nor U2324 (N_2324,N_1664,N_1582);
and U2325 (N_2325,N_1523,N_1745);
or U2326 (N_2326,N_1938,N_1945);
nor U2327 (N_2327,N_1864,N_1533);
and U2328 (N_2328,N_1684,N_1736);
nor U2329 (N_2329,N_1768,N_1534);
nand U2330 (N_2330,N_1817,N_1891);
or U2331 (N_2331,N_1842,N_1506);
nor U2332 (N_2332,N_1592,N_1562);
and U2333 (N_2333,N_1681,N_1791);
or U2334 (N_2334,N_1768,N_1689);
or U2335 (N_2335,N_1965,N_1797);
or U2336 (N_2336,N_1758,N_1889);
and U2337 (N_2337,N_1790,N_1733);
and U2338 (N_2338,N_1871,N_1727);
or U2339 (N_2339,N_1941,N_1589);
and U2340 (N_2340,N_1845,N_1964);
nand U2341 (N_2341,N_1857,N_1923);
nand U2342 (N_2342,N_1824,N_1955);
nand U2343 (N_2343,N_1554,N_1824);
or U2344 (N_2344,N_1938,N_1725);
or U2345 (N_2345,N_1819,N_1892);
or U2346 (N_2346,N_1930,N_1588);
or U2347 (N_2347,N_1774,N_1578);
nand U2348 (N_2348,N_1812,N_1612);
nand U2349 (N_2349,N_1610,N_1555);
and U2350 (N_2350,N_1679,N_1825);
nor U2351 (N_2351,N_1611,N_1831);
nand U2352 (N_2352,N_1738,N_1688);
or U2353 (N_2353,N_1599,N_1574);
or U2354 (N_2354,N_1873,N_1847);
nand U2355 (N_2355,N_1815,N_1502);
nor U2356 (N_2356,N_1624,N_1730);
nand U2357 (N_2357,N_1515,N_1852);
and U2358 (N_2358,N_1677,N_1745);
nor U2359 (N_2359,N_1815,N_1915);
and U2360 (N_2360,N_1845,N_1973);
nand U2361 (N_2361,N_1768,N_1525);
nand U2362 (N_2362,N_1768,N_1666);
or U2363 (N_2363,N_1855,N_1949);
or U2364 (N_2364,N_1505,N_1540);
or U2365 (N_2365,N_1936,N_1578);
nand U2366 (N_2366,N_1516,N_1531);
and U2367 (N_2367,N_1704,N_1940);
nand U2368 (N_2368,N_1655,N_1625);
and U2369 (N_2369,N_1674,N_1921);
nand U2370 (N_2370,N_1788,N_1567);
and U2371 (N_2371,N_1987,N_1942);
and U2372 (N_2372,N_1760,N_1570);
or U2373 (N_2373,N_1685,N_1627);
nor U2374 (N_2374,N_1638,N_1625);
or U2375 (N_2375,N_1939,N_1949);
nor U2376 (N_2376,N_1994,N_1718);
nand U2377 (N_2377,N_1785,N_1725);
nand U2378 (N_2378,N_1909,N_1777);
nor U2379 (N_2379,N_1765,N_1974);
or U2380 (N_2380,N_1998,N_1841);
xor U2381 (N_2381,N_1778,N_1548);
or U2382 (N_2382,N_1812,N_1765);
or U2383 (N_2383,N_1581,N_1838);
or U2384 (N_2384,N_1787,N_1922);
nor U2385 (N_2385,N_1533,N_1898);
nor U2386 (N_2386,N_1978,N_1929);
nand U2387 (N_2387,N_1769,N_1695);
nor U2388 (N_2388,N_1902,N_1989);
nor U2389 (N_2389,N_1834,N_1951);
and U2390 (N_2390,N_1557,N_1769);
nand U2391 (N_2391,N_1773,N_1631);
nor U2392 (N_2392,N_1596,N_1743);
or U2393 (N_2393,N_1979,N_1682);
nand U2394 (N_2394,N_1699,N_1913);
nor U2395 (N_2395,N_1577,N_1693);
nor U2396 (N_2396,N_1834,N_1719);
nand U2397 (N_2397,N_1840,N_1508);
nor U2398 (N_2398,N_1913,N_1850);
and U2399 (N_2399,N_1877,N_1715);
nand U2400 (N_2400,N_1764,N_1866);
and U2401 (N_2401,N_1884,N_1686);
nand U2402 (N_2402,N_1617,N_1557);
nor U2403 (N_2403,N_1615,N_1882);
or U2404 (N_2404,N_1504,N_1520);
nor U2405 (N_2405,N_1938,N_1661);
nand U2406 (N_2406,N_1578,N_1543);
nor U2407 (N_2407,N_1926,N_1914);
or U2408 (N_2408,N_1968,N_1667);
or U2409 (N_2409,N_1553,N_1520);
nand U2410 (N_2410,N_1576,N_1904);
and U2411 (N_2411,N_1719,N_1966);
nand U2412 (N_2412,N_1639,N_1965);
nor U2413 (N_2413,N_1710,N_1854);
or U2414 (N_2414,N_1774,N_1664);
and U2415 (N_2415,N_1594,N_1684);
nor U2416 (N_2416,N_1860,N_1902);
nand U2417 (N_2417,N_1860,N_1723);
nor U2418 (N_2418,N_1528,N_1954);
or U2419 (N_2419,N_1958,N_1601);
or U2420 (N_2420,N_1833,N_1567);
xnor U2421 (N_2421,N_1811,N_1832);
or U2422 (N_2422,N_1830,N_1841);
nand U2423 (N_2423,N_1626,N_1908);
nand U2424 (N_2424,N_1793,N_1713);
xnor U2425 (N_2425,N_1628,N_1846);
and U2426 (N_2426,N_1961,N_1600);
or U2427 (N_2427,N_1548,N_1566);
or U2428 (N_2428,N_1738,N_1812);
and U2429 (N_2429,N_1824,N_1502);
and U2430 (N_2430,N_1654,N_1569);
or U2431 (N_2431,N_1688,N_1649);
nor U2432 (N_2432,N_1841,N_1733);
or U2433 (N_2433,N_1579,N_1665);
nand U2434 (N_2434,N_1789,N_1648);
and U2435 (N_2435,N_1666,N_1865);
nand U2436 (N_2436,N_1991,N_1759);
and U2437 (N_2437,N_1694,N_1870);
nor U2438 (N_2438,N_1845,N_1700);
nand U2439 (N_2439,N_1968,N_1802);
and U2440 (N_2440,N_1713,N_1976);
nor U2441 (N_2441,N_1578,N_1818);
or U2442 (N_2442,N_1817,N_1642);
nand U2443 (N_2443,N_1773,N_1608);
or U2444 (N_2444,N_1786,N_1977);
nand U2445 (N_2445,N_1525,N_1812);
nor U2446 (N_2446,N_1882,N_1583);
and U2447 (N_2447,N_1780,N_1787);
and U2448 (N_2448,N_1711,N_1801);
and U2449 (N_2449,N_1851,N_1508);
nor U2450 (N_2450,N_1534,N_1932);
or U2451 (N_2451,N_1770,N_1847);
and U2452 (N_2452,N_1976,N_1990);
nor U2453 (N_2453,N_1868,N_1614);
nor U2454 (N_2454,N_1968,N_1845);
nor U2455 (N_2455,N_1540,N_1744);
and U2456 (N_2456,N_1797,N_1760);
or U2457 (N_2457,N_1594,N_1731);
or U2458 (N_2458,N_1872,N_1848);
nor U2459 (N_2459,N_1952,N_1628);
nand U2460 (N_2460,N_1850,N_1933);
nor U2461 (N_2461,N_1659,N_1949);
nand U2462 (N_2462,N_1661,N_1769);
nand U2463 (N_2463,N_1712,N_1805);
and U2464 (N_2464,N_1785,N_1570);
nand U2465 (N_2465,N_1809,N_1585);
and U2466 (N_2466,N_1830,N_1990);
nor U2467 (N_2467,N_1838,N_1555);
nor U2468 (N_2468,N_1583,N_1543);
nand U2469 (N_2469,N_1785,N_1698);
or U2470 (N_2470,N_1687,N_1623);
and U2471 (N_2471,N_1960,N_1543);
nor U2472 (N_2472,N_1787,N_1649);
nor U2473 (N_2473,N_1890,N_1557);
or U2474 (N_2474,N_1588,N_1522);
or U2475 (N_2475,N_1942,N_1763);
nor U2476 (N_2476,N_1843,N_1973);
or U2477 (N_2477,N_1657,N_1711);
and U2478 (N_2478,N_1642,N_1896);
or U2479 (N_2479,N_1812,N_1664);
nand U2480 (N_2480,N_1690,N_1506);
nand U2481 (N_2481,N_1591,N_1814);
nand U2482 (N_2482,N_1653,N_1593);
nor U2483 (N_2483,N_1951,N_1593);
nor U2484 (N_2484,N_1783,N_1774);
nand U2485 (N_2485,N_1697,N_1799);
and U2486 (N_2486,N_1596,N_1867);
nand U2487 (N_2487,N_1770,N_1596);
or U2488 (N_2488,N_1938,N_1644);
and U2489 (N_2489,N_1713,N_1905);
nand U2490 (N_2490,N_1955,N_1624);
or U2491 (N_2491,N_1665,N_1551);
nand U2492 (N_2492,N_1766,N_1511);
and U2493 (N_2493,N_1660,N_1986);
nand U2494 (N_2494,N_1971,N_1954);
or U2495 (N_2495,N_1837,N_1707);
nor U2496 (N_2496,N_1669,N_1750);
nor U2497 (N_2497,N_1930,N_1541);
nand U2498 (N_2498,N_1676,N_1553);
or U2499 (N_2499,N_1630,N_1625);
or U2500 (N_2500,N_2344,N_2428);
and U2501 (N_2501,N_2369,N_2438);
and U2502 (N_2502,N_2487,N_2011);
nand U2503 (N_2503,N_2102,N_2051);
nor U2504 (N_2504,N_2057,N_2315);
nand U2505 (N_2505,N_2147,N_2424);
nor U2506 (N_2506,N_2292,N_2024);
nor U2507 (N_2507,N_2256,N_2193);
nand U2508 (N_2508,N_2139,N_2439);
nor U2509 (N_2509,N_2384,N_2341);
and U2510 (N_2510,N_2010,N_2278);
nand U2511 (N_2511,N_2155,N_2224);
and U2512 (N_2512,N_2423,N_2145);
and U2513 (N_2513,N_2414,N_2017);
nand U2514 (N_2514,N_2179,N_2127);
or U2515 (N_2515,N_2003,N_2436);
and U2516 (N_2516,N_2074,N_2406);
and U2517 (N_2517,N_2403,N_2449);
nor U2518 (N_2518,N_2036,N_2251);
nand U2519 (N_2519,N_2322,N_2112);
or U2520 (N_2520,N_2093,N_2343);
and U2521 (N_2521,N_2497,N_2265);
nand U2522 (N_2522,N_2018,N_2156);
or U2523 (N_2523,N_2433,N_2190);
nor U2524 (N_2524,N_2367,N_2081);
nor U2525 (N_2525,N_2159,N_2026);
nor U2526 (N_2526,N_2314,N_2482);
nor U2527 (N_2527,N_2498,N_2199);
or U2528 (N_2528,N_2393,N_2270);
and U2529 (N_2529,N_2073,N_2214);
nor U2530 (N_2530,N_2242,N_2039);
and U2531 (N_2531,N_2453,N_2308);
nand U2532 (N_2532,N_2217,N_2320);
nor U2533 (N_2533,N_2259,N_2437);
nor U2534 (N_2534,N_2106,N_2033);
or U2535 (N_2535,N_2022,N_2038);
or U2536 (N_2536,N_2178,N_2359);
nand U2537 (N_2537,N_2052,N_2196);
or U2538 (N_2538,N_2230,N_2146);
or U2539 (N_2539,N_2266,N_2426);
nand U2540 (N_2540,N_2338,N_2361);
nand U2541 (N_2541,N_2083,N_2056);
or U2542 (N_2542,N_2333,N_2336);
nand U2543 (N_2543,N_2268,N_2120);
or U2544 (N_2544,N_2180,N_2281);
and U2545 (N_2545,N_2138,N_2086);
nand U2546 (N_2546,N_2092,N_2477);
nor U2547 (N_2547,N_2280,N_2253);
or U2548 (N_2548,N_2401,N_2115);
nor U2549 (N_2549,N_2286,N_2069);
and U2550 (N_2550,N_2126,N_2412);
nor U2551 (N_2551,N_2442,N_2132);
nor U2552 (N_2552,N_2491,N_2284);
or U2553 (N_2553,N_2128,N_2096);
nand U2554 (N_2554,N_2109,N_2034);
nor U2555 (N_2555,N_2246,N_2450);
and U2556 (N_2556,N_2441,N_2060);
and U2557 (N_2557,N_2087,N_2030);
nor U2558 (N_2558,N_2249,N_2269);
or U2559 (N_2559,N_2160,N_2241);
and U2560 (N_2560,N_2407,N_2088);
and U2561 (N_2561,N_2296,N_2041);
xnor U2562 (N_2562,N_2481,N_2285);
or U2563 (N_2563,N_2025,N_2301);
xor U2564 (N_2564,N_2262,N_2062);
nand U2565 (N_2565,N_2451,N_2399);
nor U2566 (N_2566,N_2014,N_2172);
or U2567 (N_2567,N_2032,N_2144);
nand U2568 (N_2568,N_2045,N_2035);
and U2569 (N_2569,N_2304,N_2161);
nand U2570 (N_2570,N_2219,N_2028);
nor U2571 (N_2571,N_2125,N_2177);
or U2572 (N_2572,N_2388,N_2273);
or U2573 (N_2573,N_2104,N_2430);
or U2574 (N_2574,N_2371,N_2335);
or U2575 (N_2575,N_2287,N_2136);
or U2576 (N_2576,N_2100,N_2152);
and U2577 (N_2577,N_2049,N_2486);
nor U2578 (N_2578,N_2169,N_2306);
or U2579 (N_2579,N_2252,N_2229);
and U2580 (N_2580,N_2378,N_2085);
or U2581 (N_2581,N_2006,N_2002);
nand U2582 (N_2582,N_2429,N_2394);
nor U2583 (N_2583,N_2020,N_2303);
or U2584 (N_2584,N_2162,N_2282);
nor U2585 (N_2585,N_2148,N_2328);
nand U2586 (N_2586,N_2381,N_2077);
or U2587 (N_2587,N_2387,N_2211);
or U2588 (N_2588,N_2392,N_2360);
nand U2589 (N_2589,N_2205,N_2182);
nor U2590 (N_2590,N_2331,N_2483);
or U2591 (N_2591,N_2447,N_2225);
nor U2592 (N_2592,N_2363,N_2466);
nand U2593 (N_2593,N_2089,N_2133);
nand U2594 (N_2594,N_2302,N_2300);
and U2595 (N_2595,N_2295,N_2166);
nand U2596 (N_2596,N_2329,N_2472);
nor U2597 (N_2597,N_2065,N_2037);
nor U2598 (N_2598,N_2055,N_2345);
and U2599 (N_2599,N_2149,N_2379);
or U2600 (N_2600,N_2191,N_2048);
xnor U2601 (N_2601,N_2377,N_2061);
and U2602 (N_2602,N_2267,N_2337);
nand U2603 (N_2603,N_2461,N_2114);
xnor U2604 (N_2604,N_2194,N_2332);
or U2605 (N_2605,N_2317,N_2298);
nor U2606 (N_2606,N_2151,N_2290);
nor U2607 (N_2607,N_2170,N_2027);
nor U2608 (N_2608,N_2325,N_2464);
nor U2609 (N_2609,N_2352,N_2218);
nor U2610 (N_2610,N_2385,N_2163);
or U2611 (N_2611,N_2082,N_2473);
nor U2612 (N_2612,N_2054,N_2443);
nor U2613 (N_2613,N_2465,N_2124);
or U2614 (N_2614,N_2459,N_2351);
nor U2615 (N_2615,N_2174,N_2355);
and U2616 (N_2616,N_2228,N_2134);
or U2617 (N_2617,N_2123,N_2425);
and U2618 (N_2618,N_2066,N_2207);
nand U2619 (N_2619,N_2095,N_2130);
and U2620 (N_2620,N_2183,N_2356);
nor U2621 (N_2621,N_2140,N_2029);
or U2622 (N_2622,N_2213,N_2195);
or U2623 (N_2623,N_2410,N_2471);
and U2624 (N_2624,N_2390,N_2400);
and U2625 (N_2625,N_2008,N_2203);
and U2626 (N_2626,N_2236,N_2157);
nand U2627 (N_2627,N_2305,N_2454);
or U2628 (N_2628,N_2110,N_2475);
or U2629 (N_2629,N_2158,N_2150);
and U2630 (N_2630,N_2316,N_2283);
or U2631 (N_2631,N_2264,N_2495);
nand U2632 (N_2632,N_2181,N_2467);
nand U2633 (N_2633,N_2202,N_2274);
or U2634 (N_2634,N_2098,N_2007);
xor U2635 (N_2635,N_2142,N_2248);
and U2636 (N_2636,N_2116,N_2289);
or U2637 (N_2637,N_2012,N_2485);
or U2638 (N_2638,N_2489,N_2240);
or U2639 (N_2639,N_2413,N_2078);
nand U2640 (N_2640,N_2185,N_2044);
nor U2641 (N_2641,N_2323,N_2311);
nor U2642 (N_2642,N_2023,N_2452);
and U2643 (N_2643,N_2141,N_2309);
nor U2644 (N_2644,N_2097,N_2319);
nor U2645 (N_2645,N_2231,N_2245);
or U2646 (N_2646,N_2326,N_2226);
nand U2647 (N_2647,N_2434,N_2254);
and U2648 (N_2648,N_2094,N_2373);
and U2649 (N_2649,N_2067,N_2072);
xnor U2650 (N_2650,N_2001,N_2391);
nand U2651 (N_2651,N_2119,N_2470);
nor U2652 (N_2652,N_2247,N_2276);
xnor U2653 (N_2653,N_2350,N_2444);
and U2654 (N_2654,N_2164,N_2154);
and U2655 (N_2655,N_2382,N_2222);
and U2656 (N_2656,N_2448,N_2395);
nand U2657 (N_2657,N_2250,N_2118);
nand U2658 (N_2658,N_2063,N_2402);
and U2659 (N_2659,N_2405,N_2432);
nand U2660 (N_2660,N_2469,N_2076);
or U2661 (N_2661,N_2418,N_2111);
nor U2662 (N_2662,N_2212,N_2357);
nand U2663 (N_2663,N_2263,N_2313);
and U2664 (N_2664,N_2050,N_2108);
nor U2665 (N_2665,N_2009,N_2375);
nor U2666 (N_2666,N_2310,N_2376);
or U2667 (N_2667,N_2339,N_2365);
nand U2668 (N_2668,N_2137,N_2258);
nand U2669 (N_2669,N_2016,N_2197);
or U2670 (N_2670,N_2031,N_2496);
and U2671 (N_2671,N_2216,N_2291);
or U2672 (N_2672,N_2208,N_2422);
and U2673 (N_2673,N_2053,N_2321);
nand U2674 (N_2674,N_2348,N_2330);
or U2675 (N_2675,N_2223,N_2135);
and U2676 (N_2676,N_2084,N_2187);
nand U2677 (N_2677,N_2494,N_2200);
or U2678 (N_2678,N_2013,N_2171);
nor U2679 (N_2679,N_2455,N_2220);
nor U2680 (N_2680,N_2070,N_2404);
and U2681 (N_2681,N_2493,N_2421);
nor U2682 (N_2682,N_2420,N_2347);
or U2683 (N_2683,N_2293,N_2206);
nor U2684 (N_2684,N_2232,N_2215);
nand U2685 (N_2685,N_2233,N_2312);
or U2686 (N_2686,N_2046,N_2143);
xnor U2687 (N_2687,N_2271,N_2204);
or U2688 (N_2688,N_2015,N_2478);
nand U2689 (N_2689,N_2474,N_2349);
or U2690 (N_2690,N_2380,N_2440);
and U2691 (N_2691,N_2416,N_2080);
nand U2692 (N_2692,N_2383,N_2362);
nand U2693 (N_2693,N_2059,N_2173);
nand U2694 (N_2694,N_2468,N_2488);
or U2695 (N_2695,N_2103,N_2221);
and U2696 (N_2696,N_2275,N_2396);
or U2697 (N_2697,N_2353,N_2479);
nand U2698 (N_2698,N_2431,N_2091);
xor U2699 (N_2699,N_2090,N_2463);
or U2700 (N_2700,N_2188,N_2415);
nor U2701 (N_2701,N_2105,N_2368);
or U2702 (N_2702,N_2342,N_2327);
and U2703 (N_2703,N_2417,N_2005);
and U2704 (N_2704,N_2107,N_2113);
nand U2705 (N_2705,N_2307,N_2068);
and U2706 (N_2706,N_2457,N_2358);
nand U2707 (N_2707,N_2234,N_2043);
and U2708 (N_2708,N_2079,N_2040);
nand U2709 (N_2709,N_2318,N_2004);
xor U2710 (N_2710,N_2277,N_2435);
nand U2711 (N_2711,N_2255,N_2324);
xor U2712 (N_2712,N_2460,N_2480);
nor U2713 (N_2713,N_2257,N_2239);
nand U2714 (N_2714,N_2419,N_2184);
nand U2715 (N_2715,N_2490,N_2117);
nor U2716 (N_2716,N_2462,N_2260);
nand U2717 (N_2717,N_2192,N_2340);
or U2718 (N_2718,N_2058,N_2354);
and U2719 (N_2719,N_2075,N_2334);
and U2720 (N_2720,N_2189,N_2153);
or U2721 (N_2721,N_2243,N_2288);
or U2722 (N_2722,N_2201,N_2168);
nand U2723 (N_2723,N_2370,N_2209);
nor U2724 (N_2724,N_2021,N_2411);
and U2725 (N_2725,N_2446,N_2279);
or U2726 (N_2726,N_2374,N_2198);
or U2727 (N_2727,N_2131,N_2456);
nor U2728 (N_2728,N_2176,N_2398);
or U2729 (N_2729,N_2122,N_2047);
or U2730 (N_2730,N_2299,N_2042);
nor U2731 (N_2731,N_2121,N_2366);
or U2732 (N_2732,N_2227,N_2064);
and U2733 (N_2733,N_2397,N_2167);
nand U2734 (N_2734,N_2099,N_2427);
nand U2735 (N_2735,N_2386,N_2294);
or U2736 (N_2736,N_2372,N_2186);
nand U2737 (N_2737,N_2000,N_2165);
nor U2738 (N_2738,N_2484,N_2175);
or U2739 (N_2739,N_2408,N_2499);
nor U2740 (N_2740,N_2238,N_2101);
and U2741 (N_2741,N_2492,N_2235);
and U2742 (N_2742,N_2210,N_2409);
or U2743 (N_2743,N_2389,N_2364);
nand U2744 (N_2744,N_2244,N_2129);
and U2745 (N_2745,N_2297,N_2272);
nor U2746 (N_2746,N_2019,N_2445);
nor U2747 (N_2747,N_2071,N_2261);
and U2748 (N_2748,N_2237,N_2346);
nor U2749 (N_2749,N_2458,N_2476);
nor U2750 (N_2750,N_2163,N_2239);
nand U2751 (N_2751,N_2008,N_2038);
nor U2752 (N_2752,N_2163,N_2250);
or U2753 (N_2753,N_2224,N_2179);
nand U2754 (N_2754,N_2187,N_2050);
nor U2755 (N_2755,N_2215,N_2221);
nor U2756 (N_2756,N_2243,N_2169);
nor U2757 (N_2757,N_2216,N_2167);
or U2758 (N_2758,N_2095,N_2227);
or U2759 (N_2759,N_2492,N_2480);
and U2760 (N_2760,N_2254,N_2080);
nand U2761 (N_2761,N_2231,N_2033);
or U2762 (N_2762,N_2357,N_2142);
and U2763 (N_2763,N_2241,N_2176);
nor U2764 (N_2764,N_2194,N_2106);
nor U2765 (N_2765,N_2386,N_2196);
and U2766 (N_2766,N_2057,N_2287);
nor U2767 (N_2767,N_2026,N_2273);
and U2768 (N_2768,N_2487,N_2049);
nand U2769 (N_2769,N_2331,N_2342);
and U2770 (N_2770,N_2302,N_2116);
or U2771 (N_2771,N_2014,N_2279);
nand U2772 (N_2772,N_2260,N_2194);
nor U2773 (N_2773,N_2124,N_2488);
nor U2774 (N_2774,N_2478,N_2022);
or U2775 (N_2775,N_2150,N_2167);
or U2776 (N_2776,N_2289,N_2488);
and U2777 (N_2777,N_2417,N_2138);
nor U2778 (N_2778,N_2157,N_2489);
nor U2779 (N_2779,N_2496,N_2046);
or U2780 (N_2780,N_2084,N_2066);
nand U2781 (N_2781,N_2343,N_2248);
or U2782 (N_2782,N_2397,N_2045);
nor U2783 (N_2783,N_2447,N_2218);
nand U2784 (N_2784,N_2195,N_2043);
or U2785 (N_2785,N_2028,N_2256);
xnor U2786 (N_2786,N_2440,N_2318);
and U2787 (N_2787,N_2446,N_2098);
or U2788 (N_2788,N_2461,N_2278);
nor U2789 (N_2789,N_2294,N_2447);
and U2790 (N_2790,N_2003,N_2440);
nand U2791 (N_2791,N_2226,N_2491);
nor U2792 (N_2792,N_2161,N_2285);
or U2793 (N_2793,N_2330,N_2494);
or U2794 (N_2794,N_2157,N_2378);
nand U2795 (N_2795,N_2332,N_2342);
and U2796 (N_2796,N_2304,N_2095);
and U2797 (N_2797,N_2002,N_2125);
and U2798 (N_2798,N_2142,N_2330);
nand U2799 (N_2799,N_2427,N_2287);
or U2800 (N_2800,N_2351,N_2365);
nor U2801 (N_2801,N_2449,N_2122);
and U2802 (N_2802,N_2277,N_2451);
and U2803 (N_2803,N_2427,N_2258);
and U2804 (N_2804,N_2168,N_2347);
nand U2805 (N_2805,N_2195,N_2309);
and U2806 (N_2806,N_2383,N_2451);
nand U2807 (N_2807,N_2426,N_2413);
and U2808 (N_2808,N_2397,N_2011);
nor U2809 (N_2809,N_2257,N_2475);
and U2810 (N_2810,N_2367,N_2045);
or U2811 (N_2811,N_2197,N_2467);
or U2812 (N_2812,N_2370,N_2122);
nand U2813 (N_2813,N_2109,N_2011);
and U2814 (N_2814,N_2414,N_2025);
nor U2815 (N_2815,N_2342,N_2024);
or U2816 (N_2816,N_2294,N_2126);
and U2817 (N_2817,N_2209,N_2095);
or U2818 (N_2818,N_2449,N_2150);
nor U2819 (N_2819,N_2458,N_2180);
nand U2820 (N_2820,N_2064,N_2133);
and U2821 (N_2821,N_2234,N_2423);
nand U2822 (N_2822,N_2279,N_2307);
and U2823 (N_2823,N_2246,N_2178);
and U2824 (N_2824,N_2174,N_2153);
and U2825 (N_2825,N_2331,N_2328);
and U2826 (N_2826,N_2143,N_2455);
nand U2827 (N_2827,N_2107,N_2082);
nand U2828 (N_2828,N_2493,N_2293);
and U2829 (N_2829,N_2356,N_2351);
nor U2830 (N_2830,N_2273,N_2113);
nor U2831 (N_2831,N_2385,N_2411);
nand U2832 (N_2832,N_2206,N_2001);
nand U2833 (N_2833,N_2098,N_2267);
or U2834 (N_2834,N_2284,N_2018);
and U2835 (N_2835,N_2288,N_2433);
and U2836 (N_2836,N_2474,N_2414);
or U2837 (N_2837,N_2049,N_2150);
or U2838 (N_2838,N_2308,N_2032);
or U2839 (N_2839,N_2010,N_2263);
or U2840 (N_2840,N_2221,N_2326);
xor U2841 (N_2841,N_2170,N_2237);
nand U2842 (N_2842,N_2471,N_2095);
or U2843 (N_2843,N_2412,N_2436);
and U2844 (N_2844,N_2010,N_2209);
nor U2845 (N_2845,N_2136,N_2002);
nand U2846 (N_2846,N_2317,N_2117);
nand U2847 (N_2847,N_2147,N_2247);
nor U2848 (N_2848,N_2075,N_2222);
and U2849 (N_2849,N_2286,N_2207);
or U2850 (N_2850,N_2340,N_2462);
and U2851 (N_2851,N_2409,N_2235);
nand U2852 (N_2852,N_2022,N_2204);
or U2853 (N_2853,N_2330,N_2064);
and U2854 (N_2854,N_2052,N_2282);
nor U2855 (N_2855,N_2035,N_2031);
and U2856 (N_2856,N_2044,N_2372);
or U2857 (N_2857,N_2046,N_2325);
or U2858 (N_2858,N_2494,N_2290);
and U2859 (N_2859,N_2418,N_2213);
or U2860 (N_2860,N_2034,N_2087);
or U2861 (N_2861,N_2175,N_2091);
nor U2862 (N_2862,N_2262,N_2106);
and U2863 (N_2863,N_2303,N_2322);
nand U2864 (N_2864,N_2212,N_2118);
nand U2865 (N_2865,N_2361,N_2296);
or U2866 (N_2866,N_2458,N_2375);
nand U2867 (N_2867,N_2239,N_2193);
nand U2868 (N_2868,N_2066,N_2402);
nand U2869 (N_2869,N_2296,N_2213);
and U2870 (N_2870,N_2433,N_2233);
and U2871 (N_2871,N_2242,N_2012);
or U2872 (N_2872,N_2239,N_2017);
xnor U2873 (N_2873,N_2220,N_2073);
or U2874 (N_2874,N_2101,N_2379);
xnor U2875 (N_2875,N_2421,N_2243);
nand U2876 (N_2876,N_2005,N_2377);
and U2877 (N_2877,N_2009,N_2468);
nor U2878 (N_2878,N_2494,N_2108);
nand U2879 (N_2879,N_2065,N_2011);
nor U2880 (N_2880,N_2183,N_2265);
nand U2881 (N_2881,N_2451,N_2344);
and U2882 (N_2882,N_2105,N_2091);
or U2883 (N_2883,N_2269,N_2457);
or U2884 (N_2884,N_2105,N_2352);
or U2885 (N_2885,N_2053,N_2162);
nand U2886 (N_2886,N_2475,N_2305);
nand U2887 (N_2887,N_2127,N_2393);
nor U2888 (N_2888,N_2488,N_2154);
nand U2889 (N_2889,N_2034,N_2131);
nor U2890 (N_2890,N_2393,N_2028);
and U2891 (N_2891,N_2448,N_2109);
nor U2892 (N_2892,N_2372,N_2101);
nor U2893 (N_2893,N_2288,N_2065);
nor U2894 (N_2894,N_2214,N_2173);
or U2895 (N_2895,N_2109,N_2360);
nand U2896 (N_2896,N_2297,N_2388);
and U2897 (N_2897,N_2457,N_2268);
and U2898 (N_2898,N_2337,N_2198);
or U2899 (N_2899,N_2310,N_2091);
nor U2900 (N_2900,N_2202,N_2227);
and U2901 (N_2901,N_2346,N_2319);
nor U2902 (N_2902,N_2480,N_2434);
or U2903 (N_2903,N_2412,N_2417);
nand U2904 (N_2904,N_2380,N_2283);
or U2905 (N_2905,N_2084,N_2041);
nor U2906 (N_2906,N_2463,N_2168);
nor U2907 (N_2907,N_2114,N_2375);
nor U2908 (N_2908,N_2495,N_2330);
and U2909 (N_2909,N_2241,N_2142);
or U2910 (N_2910,N_2343,N_2259);
or U2911 (N_2911,N_2303,N_2281);
and U2912 (N_2912,N_2410,N_2113);
nand U2913 (N_2913,N_2169,N_2099);
nand U2914 (N_2914,N_2380,N_2272);
nand U2915 (N_2915,N_2015,N_2401);
nor U2916 (N_2916,N_2075,N_2165);
or U2917 (N_2917,N_2302,N_2258);
nor U2918 (N_2918,N_2273,N_2126);
nand U2919 (N_2919,N_2070,N_2090);
nor U2920 (N_2920,N_2086,N_2058);
or U2921 (N_2921,N_2200,N_2390);
and U2922 (N_2922,N_2074,N_2280);
nand U2923 (N_2923,N_2467,N_2338);
nor U2924 (N_2924,N_2110,N_2318);
nor U2925 (N_2925,N_2256,N_2353);
and U2926 (N_2926,N_2434,N_2075);
nor U2927 (N_2927,N_2467,N_2472);
nand U2928 (N_2928,N_2156,N_2015);
nor U2929 (N_2929,N_2091,N_2100);
and U2930 (N_2930,N_2224,N_2090);
and U2931 (N_2931,N_2001,N_2236);
xnor U2932 (N_2932,N_2073,N_2406);
nand U2933 (N_2933,N_2329,N_2337);
and U2934 (N_2934,N_2062,N_2186);
and U2935 (N_2935,N_2195,N_2206);
nand U2936 (N_2936,N_2135,N_2329);
nand U2937 (N_2937,N_2249,N_2128);
nor U2938 (N_2938,N_2256,N_2142);
or U2939 (N_2939,N_2040,N_2226);
and U2940 (N_2940,N_2204,N_2393);
nand U2941 (N_2941,N_2356,N_2242);
nand U2942 (N_2942,N_2046,N_2164);
nor U2943 (N_2943,N_2462,N_2202);
nand U2944 (N_2944,N_2405,N_2059);
nor U2945 (N_2945,N_2449,N_2024);
nand U2946 (N_2946,N_2148,N_2313);
nor U2947 (N_2947,N_2295,N_2139);
nor U2948 (N_2948,N_2381,N_2097);
or U2949 (N_2949,N_2307,N_2120);
nor U2950 (N_2950,N_2226,N_2036);
nand U2951 (N_2951,N_2143,N_2047);
nand U2952 (N_2952,N_2338,N_2292);
and U2953 (N_2953,N_2191,N_2104);
nor U2954 (N_2954,N_2040,N_2124);
nand U2955 (N_2955,N_2335,N_2486);
nor U2956 (N_2956,N_2404,N_2061);
and U2957 (N_2957,N_2302,N_2235);
and U2958 (N_2958,N_2396,N_2036);
nand U2959 (N_2959,N_2128,N_2078);
nand U2960 (N_2960,N_2120,N_2313);
nor U2961 (N_2961,N_2111,N_2450);
and U2962 (N_2962,N_2448,N_2299);
and U2963 (N_2963,N_2225,N_2253);
and U2964 (N_2964,N_2318,N_2187);
or U2965 (N_2965,N_2169,N_2291);
and U2966 (N_2966,N_2084,N_2230);
or U2967 (N_2967,N_2222,N_2040);
nor U2968 (N_2968,N_2099,N_2151);
or U2969 (N_2969,N_2479,N_2186);
and U2970 (N_2970,N_2058,N_2009);
nand U2971 (N_2971,N_2034,N_2110);
nand U2972 (N_2972,N_2190,N_2477);
nand U2973 (N_2973,N_2122,N_2191);
or U2974 (N_2974,N_2298,N_2079);
or U2975 (N_2975,N_2333,N_2149);
or U2976 (N_2976,N_2413,N_2110);
nand U2977 (N_2977,N_2392,N_2171);
nand U2978 (N_2978,N_2341,N_2439);
nand U2979 (N_2979,N_2382,N_2170);
and U2980 (N_2980,N_2099,N_2358);
nor U2981 (N_2981,N_2197,N_2240);
and U2982 (N_2982,N_2458,N_2486);
nor U2983 (N_2983,N_2271,N_2220);
and U2984 (N_2984,N_2191,N_2004);
nor U2985 (N_2985,N_2423,N_2494);
nor U2986 (N_2986,N_2326,N_2418);
nand U2987 (N_2987,N_2188,N_2257);
nand U2988 (N_2988,N_2437,N_2151);
nor U2989 (N_2989,N_2113,N_2258);
nor U2990 (N_2990,N_2162,N_2348);
and U2991 (N_2991,N_2301,N_2409);
xnor U2992 (N_2992,N_2387,N_2308);
and U2993 (N_2993,N_2311,N_2426);
nor U2994 (N_2994,N_2107,N_2218);
and U2995 (N_2995,N_2394,N_2178);
nand U2996 (N_2996,N_2169,N_2196);
or U2997 (N_2997,N_2154,N_2493);
nor U2998 (N_2998,N_2204,N_2058);
and U2999 (N_2999,N_2184,N_2307);
or U3000 (N_3000,N_2660,N_2622);
nor U3001 (N_3001,N_2697,N_2820);
or U3002 (N_3002,N_2706,N_2857);
nor U3003 (N_3003,N_2804,N_2604);
nand U3004 (N_3004,N_2687,N_2765);
and U3005 (N_3005,N_2731,N_2954);
nor U3006 (N_3006,N_2542,N_2789);
or U3007 (N_3007,N_2716,N_2669);
and U3008 (N_3008,N_2574,N_2988);
or U3009 (N_3009,N_2578,N_2708);
nand U3010 (N_3010,N_2942,N_2720);
nand U3011 (N_3011,N_2576,N_2762);
nor U3012 (N_3012,N_2545,N_2650);
and U3013 (N_3013,N_2569,N_2616);
xnor U3014 (N_3014,N_2785,N_2620);
nor U3015 (N_3015,N_2749,N_2537);
nand U3016 (N_3016,N_2631,N_2568);
and U3017 (N_3017,N_2584,N_2596);
nand U3018 (N_3018,N_2725,N_2922);
nor U3019 (N_3019,N_2863,N_2573);
and U3020 (N_3020,N_2906,N_2860);
and U3021 (N_3021,N_2675,N_2872);
or U3022 (N_3022,N_2972,N_2796);
nand U3023 (N_3023,N_2674,N_2558);
or U3024 (N_3024,N_2665,N_2531);
nor U3025 (N_3025,N_2614,N_2962);
or U3026 (N_3026,N_2866,N_2781);
or U3027 (N_3027,N_2905,N_2734);
nor U3028 (N_3028,N_2953,N_2521);
xnor U3029 (N_3029,N_2759,N_2703);
or U3030 (N_3030,N_2694,N_2814);
nor U3031 (N_3031,N_2858,N_2770);
nor U3032 (N_3032,N_2812,N_2806);
or U3033 (N_3033,N_2721,N_2935);
nor U3034 (N_3034,N_2733,N_2549);
nor U3035 (N_3035,N_2657,N_2979);
and U3036 (N_3036,N_2779,N_2994);
nand U3037 (N_3037,N_2617,N_2647);
nand U3038 (N_3038,N_2559,N_2798);
xor U3039 (N_3039,N_2534,N_2685);
nor U3040 (N_3040,N_2634,N_2713);
nand U3041 (N_3041,N_2740,N_2523);
or U3042 (N_3042,N_2773,N_2655);
or U3043 (N_3043,N_2817,N_2777);
and U3044 (N_3044,N_2567,N_2892);
nand U3045 (N_3045,N_2824,N_2724);
nor U3046 (N_3046,N_2654,N_2856);
nand U3047 (N_3047,N_2799,N_2591);
nor U3048 (N_3048,N_2566,N_2852);
nor U3049 (N_3049,N_2950,N_2801);
nand U3050 (N_3050,N_2964,N_2682);
or U3051 (N_3051,N_2512,N_2934);
nor U3052 (N_3052,N_2931,N_2618);
nand U3053 (N_3053,N_2587,N_2589);
and U3054 (N_3054,N_2921,N_2513);
nor U3055 (N_3055,N_2896,N_2890);
and U3056 (N_3056,N_2711,N_2973);
xor U3057 (N_3057,N_2782,N_2901);
nor U3058 (N_3058,N_2848,N_2751);
nand U3059 (N_3059,N_2585,N_2730);
xor U3060 (N_3060,N_2956,N_2967);
nand U3061 (N_3061,N_2514,N_2989);
or U3062 (N_3062,N_2547,N_2705);
nor U3063 (N_3063,N_2530,N_2895);
and U3064 (N_3064,N_2875,N_2902);
nand U3065 (N_3065,N_2509,N_2912);
or U3066 (N_3066,N_2946,N_2690);
nand U3067 (N_3067,N_2851,N_2949);
xor U3068 (N_3068,N_2686,N_2610);
or U3069 (N_3069,N_2517,N_2987);
nand U3070 (N_3070,N_2554,N_2739);
nand U3071 (N_3071,N_2638,N_2511);
or U3072 (N_3072,N_2715,N_2900);
nand U3073 (N_3073,N_2528,N_2503);
nand U3074 (N_3074,N_2570,N_2698);
nand U3075 (N_3075,N_2577,N_2790);
and U3076 (N_3076,N_2599,N_2560);
or U3077 (N_3077,N_2649,N_2668);
and U3078 (N_3078,N_2629,N_2784);
nand U3079 (N_3079,N_2502,N_2842);
xor U3080 (N_3080,N_2924,N_2709);
and U3081 (N_3081,N_2609,N_2677);
or U3082 (N_3082,N_2932,N_2944);
or U3083 (N_3083,N_2766,N_2681);
and U3084 (N_3084,N_2786,N_2691);
nor U3085 (N_3085,N_2689,N_2822);
nand U3086 (N_3086,N_2844,N_2507);
nor U3087 (N_3087,N_2775,N_2532);
nand U3088 (N_3088,N_2742,N_2877);
nand U3089 (N_3089,N_2952,N_2718);
nand U3090 (N_3090,N_2809,N_2791);
nor U3091 (N_3091,N_2993,N_2612);
or U3092 (N_3092,N_2772,N_2926);
and U3093 (N_3093,N_2623,N_2633);
nand U3094 (N_3094,N_2640,N_2893);
nor U3095 (N_3095,N_2868,N_2834);
and U3096 (N_3096,N_2529,N_2678);
and U3097 (N_3097,N_2891,N_2811);
nor U3098 (N_3098,N_2983,N_2627);
or U3099 (N_3099,N_2832,N_2522);
or U3100 (N_3100,N_2957,N_2644);
and U3101 (N_3101,N_2908,N_2847);
and U3102 (N_3102,N_2712,N_2586);
or U3103 (N_3103,N_2605,N_2758);
xnor U3104 (N_3104,N_2608,N_2619);
nand U3105 (N_3105,N_2659,N_2816);
nand U3106 (N_3106,N_2639,N_2774);
or U3107 (N_3107,N_2776,N_2524);
nor U3108 (N_3108,N_2563,N_2854);
and U3109 (N_3109,N_2548,N_2688);
nand U3110 (N_3110,N_2984,N_2861);
or U3111 (N_3111,N_2592,N_2969);
and U3112 (N_3112,N_2990,N_2898);
and U3113 (N_3113,N_2825,N_2710);
and U3114 (N_3114,N_2920,N_2505);
nor U3115 (N_3115,N_2601,N_2741);
or U3116 (N_3116,N_2571,N_2719);
nand U3117 (N_3117,N_2819,N_2632);
nor U3118 (N_3118,N_2837,N_2500);
nor U3119 (N_3119,N_2556,N_2607);
nand U3120 (N_3120,N_2539,N_2879);
and U3121 (N_3121,N_2978,N_2646);
and U3122 (N_3122,N_2611,N_2966);
or U3123 (N_3123,N_2696,N_2981);
and U3124 (N_3124,N_2746,N_2971);
and U3125 (N_3125,N_2828,N_2519);
and U3126 (N_3126,N_2830,N_2602);
nor U3127 (N_3127,N_2810,N_2752);
and U3128 (N_3128,N_2778,N_2840);
and U3129 (N_3129,N_2907,N_2636);
nor U3130 (N_3130,N_2645,N_2918);
or U3131 (N_3131,N_2870,N_2579);
nor U3132 (N_3132,N_2695,N_2794);
and U3133 (N_3133,N_2624,N_2525);
nor U3134 (N_3134,N_2729,N_2541);
nor U3135 (N_3135,N_2864,N_2831);
or U3136 (N_3136,N_2986,N_2927);
or U3137 (N_3137,N_2963,N_2862);
or U3138 (N_3138,N_2771,N_2916);
or U3139 (N_3139,N_2780,N_2662);
and U3140 (N_3140,N_2606,N_2580);
nor U3141 (N_3141,N_2876,N_2700);
and U3142 (N_3142,N_2663,N_2643);
nand U3143 (N_3143,N_2991,N_2551);
or U3144 (N_3144,N_2938,N_2980);
nand U3145 (N_3145,N_2818,N_2527);
nor U3146 (N_3146,N_2651,N_2727);
nor U3147 (N_3147,N_2835,N_2995);
nand U3148 (N_3148,N_2672,N_2555);
nand U3149 (N_3149,N_2676,N_2714);
or U3150 (N_3150,N_2594,N_2970);
and U3151 (N_3151,N_2894,N_2951);
nand U3152 (N_3152,N_2679,N_2557);
nand U3153 (N_3153,N_2515,N_2565);
or U3154 (N_3154,N_2526,N_2873);
and U3155 (N_3155,N_2745,N_2702);
or U3156 (N_3156,N_2726,N_2992);
nor U3157 (N_3157,N_2520,N_2881);
and U3158 (N_3158,N_2583,N_2915);
nand U3159 (N_3159,N_2546,N_2865);
nand U3160 (N_3160,N_2788,N_2823);
or U3161 (N_3161,N_2955,N_2805);
or U3162 (N_3162,N_2598,N_2976);
or U3163 (N_3163,N_2977,N_2968);
or U3164 (N_3164,N_2761,N_2518);
or U3165 (N_3165,N_2628,N_2913);
and U3166 (N_3166,N_2998,N_2763);
and U3167 (N_3167,N_2630,N_2878);
nor U3168 (N_3168,N_2648,N_2795);
or U3169 (N_3169,N_2826,N_2961);
and U3170 (N_3170,N_2827,N_2516);
nor U3171 (N_3171,N_2888,N_2664);
nor U3172 (N_3172,N_2670,N_2757);
nand U3173 (N_3173,N_2843,N_2635);
and U3174 (N_3174,N_2750,N_2754);
or U3175 (N_3175,N_2930,N_2945);
nor U3176 (N_3176,N_2874,N_2717);
nor U3177 (N_3177,N_2923,N_2936);
nor U3178 (N_3178,N_2748,N_2723);
nand U3179 (N_3179,N_2552,N_2732);
nand U3180 (N_3180,N_2550,N_2885);
nor U3181 (N_3181,N_2593,N_2783);
and U3182 (N_3182,N_2760,N_2886);
and U3183 (N_3183,N_2928,N_2974);
nand U3184 (N_3184,N_2575,N_2501);
and U3185 (N_3185,N_2919,N_2965);
nor U3186 (N_3186,N_2767,N_2807);
or U3187 (N_3187,N_2661,N_2510);
nand U3188 (N_3188,N_2543,N_2884);
nor U3189 (N_3189,N_2684,N_2735);
nor U3190 (N_3190,N_2590,N_2744);
or U3191 (N_3191,N_2508,N_2903);
nor U3192 (N_3192,N_2793,N_2850);
or U3193 (N_3193,N_2985,N_2813);
and U3194 (N_3194,N_2889,N_2937);
and U3195 (N_3195,N_2536,N_2588);
nand U3196 (N_3196,N_2656,N_2597);
xor U3197 (N_3197,N_2561,N_2603);
and U3198 (N_3198,N_2666,N_2768);
nor U3199 (N_3199,N_2582,N_2859);
nand U3200 (N_3200,N_2803,N_2871);
nand U3201 (N_3201,N_2941,N_2960);
nor U3202 (N_3202,N_2911,N_2821);
nor U3203 (N_3203,N_2887,N_2738);
nand U3204 (N_3204,N_2506,N_2613);
nor U3205 (N_3205,N_2836,N_2929);
or U3206 (N_3206,N_2769,N_2553);
and U3207 (N_3207,N_2917,N_2845);
nand U3208 (N_3208,N_2625,N_2736);
or U3209 (N_3209,N_2621,N_2667);
nor U3210 (N_3210,N_2910,N_2707);
nand U3211 (N_3211,N_2897,N_2939);
nor U3212 (N_3212,N_2699,N_2839);
and U3213 (N_3213,N_2704,N_2504);
and U3214 (N_3214,N_2572,N_2535);
or U3215 (N_3215,N_2947,N_2692);
nand U3216 (N_3216,N_2544,N_2600);
or U3217 (N_3217,N_2538,N_2846);
or U3218 (N_3218,N_2800,N_2637);
and U3219 (N_3219,N_2683,N_2722);
nor U3220 (N_3220,N_2652,N_2737);
nand U3221 (N_3221,N_2792,N_2743);
and U3222 (N_3222,N_2925,N_2653);
or U3223 (N_3223,N_2540,N_2867);
and U3224 (N_3224,N_2680,N_2909);
nand U3225 (N_3225,N_2802,N_2829);
nor U3226 (N_3226,N_2943,N_2904);
or U3227 (N_3227,N_2899,N_2671);
nand U3228 (N_3228,N_2853,N_2562);
nand U3229 (N_3229,N_2940,N_2914);
and U3230 (N_3230,N_2764,N_2595);
or U3231 (N_3231,N_2933,N_2693);
nor U3232 (N_3232,N_2787,N_2642);
nor U3233 (N_3233,N_2701,N_2581);
nor U3234 (N_3234,N_2959,N_2849);
or U3235 (N_3235,N_2728,N_2841);
and U3236 (N_3236,N_2880,N_2869);
or U3237 (N_3237,N_2996,N_2975);
nand U3238 (N_3238,N_2747,N_2658);
or U3239 (N_3239,N_2533,N_2997);
xnor U3240 (N_3240,N_2756,N_2883);
nor U3241 (N_3241,N_2797,N_2855);
and U3242 (N_3242,N_2815,N_2838);
nand U3243 (N_3243,N_2755,N_2641);
nor U3244 (N_3244,N_2808,N_2948);
and U3245 (N_3245,N_2882,N_2564);
nor U3246 (N_3246,N_2615,N_2958);
and U3247 (N_3247,N_2999,N_2753);
and U3248 (N_3248,N_2673,N_2626);
and U3249 (N_3249,N_2833,N_2982);
nor U3250 (N_3250,N_2977,N_2817);
and U3251 (N_3251,N_2685,N_2865);
and U3252 (N_3252,N_2625,N_2929);
nand U3253 (N_3253,N_2926,N_2555);
nand U3254 (N_3254,N_2683,N_2913);
xor U3255 (N_3255,N_2570,N_2851);
or U3256 (N_3256,N_2929,N_2638);
or U3257 (N_3257,N_2732,N_2736);
nand U3258 (N_3258,N_2600,N_2893);
and U3259 (N_3259,N_2681,N_2902);
nand U3260 (N_3260,N_2611,N_2975);
nor U3261 (N_3261,N_2720,N_2593);
or U3262 (N_3262,N_2653,N_2812);
or U3263 (N_3263,N_2931,N_2724);
nand U3264 (N_3264,N_2830,N_2978);
or U3265 (N_3265,N_2798,N_2599);
nand U3266 (N_3266,N_2638,N_2556);
and U3267 (N_3267,N_2788,N_2794);
or U3268 (N_3268,N_2830,N_2529);
xnor U3269 (N_3269,N_2722,N_2793);
and U3270 (N_3270,N_2988,N_2564);
nor U3271 (N_3271,N_2509,N_2949);
nand U3272 (N_3272,N_2878,N_2814);
and U3273 (N_3273,N_2729,N_2732);
and U3274 (N_3274,N_2788,N_2978);
or U3275 (N_3275,N_2905,N_2759);
nand U3276 (N_3276,N_2649,N_2963);
nand U3277 (N_3277,N_2645,N_2624);
or U3278 (N_3278,N_2948,N_2960);
xor U3279 (N_3279,N_2747,N_2592);
or U3280 (N_3280,N_2752,N_2589);
nand U3281 (N_3281,N_2818,N_2924);
or U3282 (N_3282,N_2695,N_2924);
nand U3283 (N_3283,N_2561,N_2862);
nand U3284 (N_3284,N_2524,N_2695);
xnor U3285 (N_3285,N_2614,N_2642);
or U3286 (N_3286,N_2860,N_2500);
nor U3287 (N_3287,N_2550,N_2772);
nand U3288 (N_3288,N_2902,N_2589);
or U3289 (N_3289,N_2921,N_2679);
nand U3290 (N_3290,N_2611,N_2541);
and U3291 (N_3291,N_2589,N_2553);
nor U3292 (N_3292,N_2919,N_2882);
and U3293 (N_3293,N_2996,N_2570);
nand U3294 (N_3294,N_2710,N_2937);
nor U3295 (N_3295,N_2814,N_2594);
nand U3296 (N_3296,N_2734,N_2567);
and U3297 (N_3297,N_2605,N_2977);
or U3298 (N_3298,N_2701,N_2924);
or U3299 (N_3299,N_2833,N_2647);
nor U3300 (N_3300,N_2580,N_2596);
or U3301 (N_3301,N_2708,N_2555);
xor U3302 (N_3302,N_2923,N_2773);
nor U3303 (N_3303,N_2745,N_2749);
nor U3304 (N_3304,N_2550,N_2879);
nor U3305 (N_3305,N_2648,N_2606);
nor U3306 (N_3306,N_2622,N_2734);
and U3307 (N_3307,N_2696,N_2707);
nand U3308 (N_3308,N_2798,N_2538);
nor U3309 (N_3309,N_2502,N_2819);
nor U3310 (N_3310,N_2850,N_2716);
nand U3311 (N_3311,N_2921,N_2998);
nor U3312 (N_3312,N_2713,N_2581);
or U3313 (N_3313,N_2915,N_2853);
nand U3314 (N_3314,N_2806,N_2863);
nand U3315 (N_3315,N_2663,N_2535);
or U3316 (N_3316,N_2856,N_2671);
and U3317 (N_3317,N_2776,N_2625);
or U3318 (N_3318,N_2631,N_2676);
nor U3319 (N_3319,N_2606,N_2826);
nand U3320 (N_3320,N_2663,N_2885);
and U3321 (N_3321,N_2909,N_2529);
or U3322 (N_3322,N_2773,N_2896);
nand U3323 (N_3323,N_2900,N_2780);
or U3324 (N_3324,N_2522,N_2503);
or U3325 (N_3325,N_2586,N_2538);
and U3326 (N_3326,N_2678,N_2554);
or U3327 (N_3327,N_2751,N_2723);
xor U3328 (N_3328,N_2762,N_2908);
nand U3329 (N_3329,N_2757,N_2686);
or U3330 (N_3330,N_2606,N_2636);
or U3331 (N_3331,N_2965,N_2806);
or U3332 (N_3332,N_2930,N_2861);
xnor U3333 (N_3333,N_2596,N_2808);
nor U3334 (N_3334,N_2825,N_2552);
or U3335 (N_3335,N_2657,N_2778);
nand U3336 (N_3336,N_2741,N_2859);
nand U3337 (N_3337,N_2677,N_2547);
and U3338 (N_3338,N_2768,N_2837);
nand U3339 (N_3339,N_2856,N_2784);
xor U3340 (N_3340,N_2544,N_2732);
and U3341 (N_3341,N_2802,N_2849);
nand U3342 (N_3342,N_2783,N_2655);
and U3343 (N_3343,N_2504,N_2835);
and U3344 (N_3344,N_2613,N_2899);
or U3345 (N_3345,N_2810,N_2888);
and U3346 (N_3346,N_2991,N_2589);
and U3347 (N_3347,N_2779,N_2795);
and U3348 (N_3348,N_2854,N_2783);
or U3349 (N_3349,N_2971,N_2630);
xor U3350 (N_3350,N_2999,N_2571);
or U3351 (N_3351,N_2855,N_2657);
and U3352 (N_3352,N_2739,N_2580);
nor U3353 (N_3353,N_2667,N_2605);
nor U3354 (N_3354,N_2636,N_2951);
nor U3355 (N_3355,N_2606,N_2697);
or U3356 (N_3356,N_2675,N_2958);
nor U3357 (N_3357,N_2881,N_2532);
or U3358 (N_3358,N_2836,N_2901);
and U3359 (N_3359,N_2628,N_2969);
or U3360 (N_3360,N_2563,N_2586);
or U3361 (N_3361,N_2646,N_2682);
or U3362 (N_3362,N_2860,N_2666);
nor U3363 (N_3363,N_2985,N_2895);
nand U3364 (N_3364,N_2929,N_2801);
nand U3365 (N_3365,N_2975,N_2819);
nor U3366 (N_3366,N_2932,N_2948);
or U3367 (N_3367,N_2907,N_2643);
and U3368 (N_3368,N_2717,N_2946);
nor U3369 (N_3369,N_2985,N_2834);
or U3370 (N_3370,N_2989,N_2682);
or U3371 (N_3371,N_2851,N_2542);
and U3372 (N_3372,N_2984,N_2970);
and U3373 (N_3373,N_2915,N_2636);
nor U3374 (N_3374,N_2814,N_2769);
nor U3375 (N_3375,N_2652,N_2804);
and U3376 (N_3376,N_2964,N_2991);
nand U3377 (N_3377,N_2796,N_2819);
nor U3378 (N_3378,N_2870,N_2857);
nor U3379 (N_3379,N_2641,N_2812);
nor U3380 (N_3380,N_2933,N_2866);
nand U3381 (N_3381,N_2526,N_2511);
nand U3382 (N_3382,N_2539,N_2798);
and U3383 (N_3383,N_2768,N_2681);
nor U3384 (N_3384,N_2893,N_2923);
and U3385 (N_3385,N_2732,N_2833);
xor U3386 (N_3386,N_2554,N_2506);
and U3387 (N_3387,N_2952,N_2894);
or U3388 (N_3388,N_2954,N_2534);
nand U3389 (N_3389,N_2760,N_2686);
nand U3390 (N_3390,N_2785,N_2536);
nand U3391 (N_3391,N_2750,N_2979);
or U3392 (N_3392,N_2871,N_2823);
and U3393 (N_3393,N_2542,N_2893);
and U3394 (N_3394,N_2990,N_2653);
and U3395 (N_3395,N_2534,N_2947);
and U3396 (N_3396,N_2827,N_2624);
and U3397 (N_3397,N_2740,N_2515);
and U3398 (N_3398,N_2977,N_2833);
and U3399 (N_3399,N_2827,N_2531);
nor U3400 (N_3400,N_2918,N_2951);
nand U3401 (N_3401,N_2946,N_2726);
nand U3402 (N_3402,N_2861,N_2828);
nand U3403 (N_3403,N_2666,N_2889);
nor U3404 (N_3404,N_2687,N_2822);
nand U3405 (N_3405,N_2533,N_2652);
nor U3406 (N_3406,N_2803,N_2747);
xor U3407 (N_3407,N_2541,N_2781);
or U3408 (N_3408,N_2987,N_2614);
nand U3409 (N_3409,N_2919,N_2688);
or U3410 (N_3410,N_2892,N_2517);
nor U3411 (N_3411,N_2761,N_2508);
or U3412 (N_3412,N_2818,N_2782);
and U3413 (N_3413,N_2832,N_2903);
or U3414 (N_3414,N_2873,N_2720);
nor U3415 (N_3415,N_2755,N_2522);
nand U3416 (N_3416,N_2926,N_2604);
nor U3417 (N_3417,N_2707,N_2892);
nor U3418 (N_3418,N_2870,N_2941);
nor U3419 (N_3419,N_2840,N_2884);
and U3420 (N_3420,N_2682,N_2844);
nor U3421 (N_3421,N_2847,N_2535);
and U3422 (N_3422,N_2750,N_2772);
nand U3423 (N_3423,N_2584,N_2812);
nand U3424 (N_3424,N_2703,N_2879);
nand U3425 (N_3425,N_2984,N_2986);
or U3426 (N_3426,N_2585,N_2635);
nand U3427 (N_3427,N_2975,N_2722);
nand U3428 (N_3428,N_2960,N_2903);
and U3429 (N_3429,N_2581,N_2594);
nand U3430 (N_3430,N_2650,N_2783);
nand U3431 (N_3431,N_2556,N_2666);
and U3432 (N_3432,N_2676,N_2982);
xnor U3433 (N_3433,N_2580,N_2694);
nor U3434 (N_3434,N_2525,N_2705);
or U3435 (N_3435,N_2758,N_2667);
or U3436 (N_3436,N_2619,N_2630);
nor U3437 (N_3437,N_2924,N_2844);
and U3438 (N_3438,N_2780,N_2740);
nor U3439 (N_3439,N_2538,N_2768);
nand U3440 (N_3440,N_2700,N_2505);
nor U3441 (N_3441,N_2720,N_2878);
or U3442 (N_3442,N_2544,N_2956);
or U3443 (N_3443,N_2507,N_2565);
and U3444 (N_3444,N_2526,N_2694);
or U3445 (N_3445,N_2631,N_2729);
and U3446 (N_3446,N_2791,N_2810);
and U3447 (N_3447,N_2573,N_2663);
or U3448 (N_3448,N_2918,N_2771);
and U3449 (N_3449,N_2909,N_2593);
nor U3450 (N_3450,N_2909,N_2695);
and U3451 (N_3451,N_2583,N_2869);
and U3452 (N_3452,N_2787,N_2633);
or U3453 (N_3453,N_2862,N_2549);
and U3454 (N_3454,N_2649,N_2746);
nand U3455 (N_3455,N_2810,N_2607);
and U3456 (N_3456,N_2559,N_2986);
or U3457 (N_3457,N_2726,N_2563);
or U3458 (N_3458,N_2829,N_2670);
nand U3459 (N_3459,N_2879,N_2807);
or U3460 (N_3460,N_2883,N_2618);
nand U3461 (N_3461,N_2903,N_2915);
or U3462 (N_3462,N_2504,N_2911);
nor U3463 (N_3463,N_2682,N_2834);
nor U3464 (N_3464,N_2818,N_2996);
xnor U3465 (N_3465,N_2675,N_2898);
xnor U3466 (N_3466,N_2594,N_2993);
nand U3467 (N_3467,N_2926,N_2986);
or U3468 (N_3468,N_2951,N_2748);
and U3469 (N_3469,N_2647,N_2810);
or U3470 (N_3470,N_2698,N_2539);
or U3471 (N_3471,N_2714,N_2830);
nor U3472 (N_3472,N_2562,N_2721);
nand U3473 (N_3473,N_2532,N_2505);
or U3474 (N_3474,N_2747,N_2721);
and U3475 (N_3475,N_2715,N_2786);
and U3476 (N_3476,N_2965,N_2633);
or U3477 (N_3477,N_2759,N_2765);
nand U3478 (N_3478,N_2732,N_2744);
and U3479 (N_3479,N_2501,N_2596);
nor U3480 (N_3480,N_2684,N_2804);
or U3481 (N_3481,N_2506,N_2594);
or U3482 (N_3482,N_2875,N_2583);
nand U3483 (N_3483,N_2829,N_2507);
nor U3484 (N_3484,N_2682,N_2808);
nand U3485 (N_3485,N_2869,N_2823);
or U3486 (N_3486,N_2714,N_2973);
nand U3487 (N_3487,N_2988,N_2655);
nor U3488 (N_3488,N_2912,N_2980);
and U3489 (N_3489,N_2673,N_2797);
or U3490 (N_3490,N_2708,N_2967);
nor U3491 (N_3491,N_2962,N_2815);
nor U3492 (N_3492,N_2622,N_2976);
or U3493 (N_3493,N_2864,N_2860);
or U3494 (N_3494,N_2591,N_2994);
nor U3495 (N_3495,N_2730,N_2766);
nand U3496 (N_3496,N_2819,N_2685);
or U3497 (N_3497,N_2791,N_2762);
nand U3498 (N_3498,N_2953,N_2543);
nand U3499 (N_3499,N_2739,N_2800);
or U3500 (N_3500,N_3246,N_3092);
nand U3501 (N_3501,N_3208,N_3167);
nor U3502 (N_3502,N_3027,N_3442);
nand U3503 (N_3503,N_3130,N_3286);
or U3504 (N_3504,N_3362,N_3188);
nand U3505 (N_3505,N_3408,N_3174);
or U3506 (N_3506,N_3338,N_3200);
and U3507 (N_3507,N_3432,N_3068);
nand U3508 (N_3508,N_3054,N_3019);
or U3509 (N_3509,N_3146,N_3205);
nor U3510 (N_3510,N_3170,N_3486);
nand U3511 (N_3511,N_3302,N_3458);
or U3512 (N_3512,N_3241,N_3242);
or U3513 (N_3513,N_3180,N_3292);
or U3514 (N_3514,N_3049,N_3428);
and U3515 (N_3515,N_3096,N_3214);
nor U3516 (N_3516,N_3100,N_3058);
or U3517 (N_3517,N_3011,N_3059);
nand U3518 (N_3518,N_3371,N_3122);
or U3519 (N_3519,N_3411,N_3175);
or U3520 (N_3520,N_3209,N_3183);
or U3521 (N_3521,N_3143,N_3189);
and U3522 (N_3522,N_3072,N_3494);
and U3523 (N_3523,N_3156,N_3171);
nand U3524 (N_3524,N_3406,N_3103);
nor U3525 (N_3525,N_3397,N_3368);
nor U3526 (N_3526,N_3472,N_3135);
nor U3527 (N_3527,N_3086,N_3028);
nand U3528 (N_3528,N_3001,N_3332);
or U3529 (N_3529,N_3261,N_3221);
nor U3530 (N_3530,N_3319,N_3352);
or U3531 (N_3531,N_3416,N_3311);
nor U3532 (N_3532,N_3206,N_3219);
or U3533 (N_3533,N_3373,N_3479);
nand U3534 (N_3534,N_3119,N_3109);
and U3535 (N_3535,N_3230,N_3112);
nor U3536 (N_3536,N_3013,N_3313);
nand U3537 (N_3537,N_3163,N_3347);
nand U3538 (N_3538,N_3181,N_3253);
nor U3539 (N_3539,N_3139,N_3184);
nand U3540 (N_3540,N_3034,N_3430);
or U3541 (N_3541,N_3069,N_3084);
xnor U3542 (N_3542,N_3421,N_3033);
and U3543 (N_3543,N_3290,N_3267);
nor U3544 (N_3544,N_3095,N_3173);
nor U3545 (N_3545,N_3482,N_3457);
nor U3546 (N_3546,N_3433,N_3104);
nand U3547 (N_3547,N_3210,N_3003);
nor U3548 (N_3548,N_3275,N_3030);
or U3549 (N_3549,N_3248,N_3446);
xnor U3550 (N_3550,N_3009,N_3070);
or U3551 (N_3551,N_3272,N_3158);
nand U3552 (N_3552,N_3407,N_3493);
and U3553 (N_3553,N_3452,N_3199);
or U3554 (N_3554,N_3330,N_3106);
nor U3555 (N_3555,N_3198,N_3172);
nand U3556 (N_3556,N_3496,N_3263);
and U3557 (N_3557,N_3366,N_3404);
and U3558 (N_3558,N_3481,N_3322);
or U3559 (N_3559,N_3422,N_3451);
nand U3560 (N_3560,N_3178,N_3409);
and U3561 (N_3561,N_3125,N_3165);
nor U3562 (N_3562,N_3145,N_3310);
nand U3563 (N_3563,N_3448,N_3115);
and U3564 (N_3564,N_3066,N_3207);
and U3565 (N_3565,N_3052,N_3385);
or U3566 (N_3566,N_3055,N_3064);
nand U3567 (N_3567,N_3259,N_3085);
and U3568 (N_3568,N_3025,N_3294);
and U3569 (N_3569,N_3254,N_3437);
nor U3570 (N_3570,N_3291,N_3403);
nand U3571 (N_3571,N_3485,N_3359);
and U3572 (N_3572,N_3335,N_3090);
or U3573 (N_3573,N_3223,N_3160);
nand U3574 (N_3574,N_3169,N_3193);
nand U3575 (N_3575,N_3418,N_3306);
or U3576 (N_3576,N_3401,N_3060);
xnor U3577 (N_3577,N_3043,N_3120);
or U3578 (N_3578,N_3320,N_3140);
nor U3579 (N_3579,N_3282,N_3462);
or U3580 (N_3580,N_3257,N_3232);
nand U3581 (N_3581,N_3234,N_3177);
and U3582 (N_3582,N_3328,N_3340);
or U3583 (N_3583,N_3293,N_3051);
or U3584 (N_3584,N_3354,N_3016);
nand U3585 (N_3585,N_3217,N_3439);
nand U3586 (N_3586,N_3400,N_3023);
and U3587 (N_3587,N_3154,N_3111);
or U3588 (N_3588,N_3110,N_3327);
and U3589 (N_3589,N_3073,N_3007);
or U3590 (N_3590,N_3269,N_3078);
nand U3591 (N_3591,N_3105,N_3337);
or U3592 (N_3592,N_3295,N_3460);
nor U3593 (N_3593,N_3079,N_3076);
nor U3594 (N_3594,N_3357,N_3179);
nand U3595 (N_3595,N_3168,N_3386);
nor U3596 (N_3596,N_3420,N_3392);
or U3597 (N_3597,N_3062,N_3464);
nand U3598 (N_3598,N_3358,N_3334);
and U3599 (N_3599,N_3393,N_3444);
and U3600 (N_3600,N_3326,N_3351);
and U3601 (N_3601,N_3114,N_3431);
or U3602 (N_3602,N_3255,N_3374);
xor U3603 (N_3603,N_3074,N_3245);
nor U3604 (N_3604,N_3376,N_3341);
or U3605 (N_3605,N_3343,N_3365);
or U3606 (N_3606,N_3037,N_3192);
nor U3607 (N_3607,N_3469,N_3318);
nor U3608 (N_3608,N_3002,N_3161);
and U3609 (N_3609,N_3273,N_3157);
nand U3610 (N_3610,N_3128,N_3006);
nor U3611 (N_3611,N_3329,N_3447);
nor U3612 (N_3612,N_3346,N_3412);
or U3613 (N_3613,N_3356,N_3131);
and U3614 (N_3614,N_3423,N_3091);
or U3615 (N_3615,N_3410,N_3378);
or U3616 (N_3616,N_3123,N_3339);
or U3617 (N_3617,N_3081,N_3271);
and U3618 (N_3618,N_3162,N_3265);
and U3619 (N_3619,N_3056,N_3389);
nor U3620 (N_3620,N_3202,N_3190);
and U3621 (N_3621,N_3299,N_3147);
and U3622 (N_3622,N_3164,N_3467);
and U3623 (N_3623,N_3414,N_3010);
and U3624 (N_3624,N_3020,N_3468);
or U3625 (N_3625,N_3465,N_3218);
nand U3626 (N_3626,N_3425,N_3440);
and U3627 (N_3627,N_3048,N_3116);
or U3628 (N_3628,N_3053,N_3071);
nand U3629 (N_3629,N_3137,N_3063);
nand U3630 (N_3630,N_3093,N_3361);
nand U3631 (N_3631,N_3314,N_3434);
or U3632 (N_3632,N_3129,N_3321);
and U3633 (N_3633,N_3307,N_3415);
xnor U3634 (N_3634,N_3495,N_3089);
and U3635 (N_3635,N_3088,N_3155);
nor U3636 (N_3636,N_3196,N_3476);
nor U3637 (N_3637,N_3350,N_3345);
nand U3638 (N_3638,N_3277,N_3197);
nand U3639 (N_3639,N_3398,N_3124);
nor U3640 (N_3640,N_3466,N_3040);
nor U3641 (N_3641,N_3405,N_3436);
nor U3642 (N_3642,N_3377,N_3031);
nand U3643 (N_3643,N_3153,N_3427);
or U3644 (N_3644,N_3099,N_3266);
nor U3645 (N_3645,N_3251,N_3166);
or U3646 (N_3646,N_3022,N_3220);
xnor U3647 (N_3647,N_3132,N_3276);
or U3648 (N_3648,N_3268,N_3283);
nand U3649 (N_3649,N_3237,N_3459);
and U3650 (N_3650,N_3355,N_3287);
nor U3651 (N_3651,N_3182,N_3498);
and U3652 (N_3652,N_3252,N_3270);
and U3653 (N_3653,N_3381,N_3113);
and U3654 (N_3654,N_3151,N_3008);
or U3655 (N_3655,N_3492,N_3454);
or U3656 (N_3656,N_3014,N_3222);
and U3657 (N_3657,N_3264,N_3142);
xor U3658 (N_3658,N_3235,N_3187);
or U3659 (N_3659,N_3331,N_3000);
and U3660 (N_3660,N_3296,N_3256);
nand U3661 (N_3661,N_3044,N_3364);
nand U3662 (N_3662,N_3301,N_3036);
and U3663 (N_3663,N_3024,N_3126);
and U3664 (N_3664,N_3399,N_3212);
and U3665 (N_3665,N_3285,N_3224);
nor U3666 (N_3666,N_3121,N_3236);
nand U3667 (N_3667,N_3225,N_3441);
or U3668 (N_3668,N_3461,N_3108);
and U3669 (N_3669,N_3050,N_3012);
nand U3670 (N_3670,N_3244,N_3041);
and U3671 (N_3671,N_3144,N_3367);
nor U3672 (N_3672,N_3185,N_3038);
and U3673 (N_3673,N_3233,N_3402);
nor U3674 (N_3674,N_3046,N_3315);
nor U3675 (N_3675,N_3491,N_3489);
or U3676 (N_3676,N_3015,N_3215);
or U3677 (N_3677,N_3300,N_3380);
or U3678 (N_3678,N_3017,N_3342);
or U3679 (N_3679,N_3455,N_3443);
or U3680 (N_3680,N_3445,N_3211);
nand U3681 (N_3681,N_3229,N_3195);
or U3682 (N_3682,N_3284,N_3384);
or U3683 (N_3683,N_3383,N_3435);
nand U3684 (N_3684,N_3304,N_3107);
nor U3685 (N_3685,N_3097,N_3470);
nor U3686 (N_3686,N_3149,N_3039);
nor U3687 (N_3687,N_3262,N_3333);
or U3688 (N_3688,N_3152,N_3274);
nand U3689 (N_3689,N_3449,N_3201);
or U3690 (N_3690,N_3298,N_3098);
and U3691 (N_3691,N_3474,N_3349);
nand U3692 (N_3692,N_3308,N_3203);
nor U3693 (N_3693,N_3288,N_3082);
nor U3694 (N_3694,N_3227,N_3136);
or U3695 (N_3695,N_3450,N_3369);
nand U3696 (N_3696,N_3372,N_3336);
nand U3697 (N_3697,N_3317,N_3473);
or U3698 (N_3698,N_3388,N_3191);
and U3699 (N_3699,N_3303,N_3249);
or U3700 (N_3700,N_3243,N_3363);
nor U3701 (N_3701,N_3353,N_3018);
or U3702 (N_3702,N_3413,N_3379);
nor U3703 (N_3703,N_3463,N_3148);
and U3704 (N_3704,N_3323,N_3480);
and U3705 (N_3705,N_3438,N_3490);
and U3706 (N_3706,N_3087,N_3478);
and U3707 (N_3707,N_3061,N_3247);
nor U3708 (N_3708,N_3471,N_3228);
nor U3709 (N_3709,N_3419,N_3297);
nor U3710 (N_3710,N_3309,N_3394);
nand U3711 (N_3711,N_3216,N_3117);
and U3712 (N_3712,N_3021,N_3456);
nand U3713 (N_3713,N_3325,N_3238);
nand U3714 (N_3714,N_3194,N_3141);
and U3715 (N_3715,N_3127,N_3484);
nor U3716 (N_3716,N_3057,N_3279);
or U3717 (N_3717,N_3390,N_3391);
nor U3718 (N_3718,N_3424,N_3005);
and U3719 (N_3719,N_3102,N_3133);
nor U3720 (N_3720,N_3231,N_3344);
or U3721 (N_3721,N_3429,N_3487);
and U3722 (N_3722,N_3258,N_3312);
or U3723 (N_3723,N_3426,N_3239);
nor U3724 (N_3724,N_3250,N_3159);
nand U3725 (N_3725,N_3067,N_3032);
or U3726 (N_3726,N_3278,N_3045);
nor U3727 (N_3727,N_3417,N_3150);
nand U3728 (N_3728,N_3360,N_3075);
and U3729 (N_3729,N_3324,N_3134);
and U3730 (N_3730,N_3240,N_3042);
nand U3731 (N_3731,N_3094,N_3035);
nand U3732 (N_3732,N_3453,N_3305);
nand U3733 (N_3733,N_3138,N_3488);
and U3734 (N_3734,N_3026,N_3204);
nor U3735 (N_3735,N_3289,N_3047);
nand U3736 (N_3736,N_3475,N_3176);
nor U3737 (N_3737,N_3395,N_3080);
nor U3738 (N_3738,N_3396,N_3280);
nand U3739 (N_3739,N_3077,N_3499);
nand U3740 (N_3740,N_3260,N_3213);
and U3741 (N_3741,N_3226,N_3065);
nand U3742 (N_3742,N_3477,N_3186);
or U3743 (N_3743,N_3118,N_3101);
or U3744 (N_3744,N_3029,N_3348);
nor U3745 (N_3745,N_3281,N_3004);
and U3746 (N_3746,N_3316,N_3375);
and U3747 (N_3747,N_3483,N_3382);
or U3748 (N_3748,N_3370,N_3497);
and U3749 (N_3749,N_3387,N_3083);
or U3750 (N_3750,N_3330,N_3381);
nor U3751 (N_3751,N_3124,N_3183);
and U3752 (N_3752,N_3171,N_3237);
nor U3753 (N_3753,N_3030,N_3155);
nand U3754 (N_3754,N_3297,N_3215);
or U3755 (N_3755,N_3445,N_3107);
nand U3756 (N_3756,N_3193,N_3320);
and U3757 (N_3757,N_3250,N_3287);
nand U3758 (N_3758,N_3162,N_3076);
nand U3759 (N_3759,N_3407,N_3175);
xnor U3760 (N_3760,N_3207,N_3104);
nand U3761 (N_3761,N_3321,N_3157);
nor U3762 (N_3762,N_3419,N_3328);
and U3763 (N_3763,N_3224,N_3263);
nand U3764 (N_3764,N_3266,N_3312);
nor U3765 (N_3765,N_3067,N_3166);
nor U3766 (N_3766,N_3059,N_3220);
nor U3767 (N_3767,N_3152,N_3353);
and U3768 (N_3768,N_3160,N_3364);
nand U3769 (N_3769,N_3368,N_3431);
or U3770 (N_3770,N_3324,N_3184);
or U3771 (N_3771,N_3449,N_3368);
and U3772 (N_3772,N_3111,N_3375);
xor U3773 (N_3773,N_3443,N_3040);
or U3774 (N_3774,N_3015,N_3232);
and U3775 (N_3775,N_3279,N_3327);
or U3776 (N_3776,N_3089,N_3313);
or U3777 (N_3777,N_3239,N_3289);
nand U3778 (N_3778,N_3233,N_3232);
nand U3779 (N_3779,N_3422,N_3041);
nor U3780 (N_3780,N_3242,N_3164);
or U3781 (N_3781,N_3117,N_3447);
or U3782 (N_3782,N_3181,N_3286);
nand U3783 (N_3783,N_3253,N_3175);
nand U3784 (N_3784,N_3351,N_3079);
or U3785 (N_3785,N_3188,N_3073);
nand U3786 (N_3786,N_3191,N_3261);
nor U3787 (N_3787,N_3004,N_3128);
nor U3788 (N_3788,N_3388,N_3151);
nor U3789 (N_3789,N_3134,N_3201);
nand U3790 (N_3790,N_3328,N_3489);
nand U3791 (N_3791,N_3312,N_3396);
and U3792 (N_3792,N_3284,N_3068);
and U3793 (N_3793,N_3030,N_3089);
xnor U3794 (N_3794,N_3027,N_3083);
nand U3795 (N_3795,N_3169,N_3463);
nor U3796 (N_3796,N_3232,N_3461);
and U3797 (N_3797,N_3177,N_3420);
and U3798 (N_3798,N_3247,N_3012);
or U3799 (N_3799,N_3180,N_3479);
or U3800 (N_3800,N_3051,N_3397);
and U3801 (N_3801,N_3217,N_3491);
and U3802 (N_3802,N_3319,N_3394);
and U3803 (N_3803,N_3278,N_3292);
and U3804 (N_3804,N_3077,N_3481);
nor U3805 (N_3805,N_3005,N_3139);
nand U3806 (N_3806,N_3268,N_3493);
and U3807 (N_3807,N_3155,N_3361);
nand U3808 (N_3808,N_3126,N_3188);
nand U3809 (N_3809,N_3251,N_3161);
and U3810 (N_3810,N_3201,N_3196);
nand U3811 (N_3811,N_3339,N_3385);
nand U3812 (N_3812,N_3378,N_3183);
nor U3813 (N_3813,N_3413,N_3279);
xnor U3814 (N_3814,N_3237,N_3220);
or U3815 (N_3815,N_3059,N_3458);
and U3816 (N_3816,N_3160,N_3136);
nand U3817 (N_3817,N_3216,N_3155);
or U3818 (N_3818,N_3027,N_3346);
or U3819 (N_3819,N_3065,N_3153);
and U3820 (N_3820,N_3407,N_3069);
nor U3821 (N_3821,N_3074,N_3029);
or U3822 (N_3822,N_3275,N_3058);
nand U3823 (N_3823,N_3407,N_3195);
or U3824 (N_3824,N_3060,N_3131);
and U3825 (N_3825,N_3210,N_3059);
or U3826 (N_3826,N_3104,N_3475);
or U3827 (N_3827,N_3030,N_3495);
or U3828 (N_3828,N_3478,N_3313);
and U3829 (N_3829,N_3336,N_3300);
and U3830 (N_3830,N_3411,N_3214);
nand U3831 (N_3831,N_3381,N_3422);
or U3832 (N_3832,N_3087,N_3011);
nor U3833 (N_3833,N_3151,N_3335);
nand U3834 (N_3834,N_3065,N_3416);
or U3835 (N_3835,N_3468,N_3325);
nor U3836 (N_3836,N_3270,N_3382);
or U3837 (N_3837,N_3357,N_3079);
or U3838 (N_3838,N_3366,N_3185);
nor U3839 (N_3839,N_3066,N_3030);
and U3840 (N_3840,N_3411,N_3291);
and U3841 (N_3841,N_3464,N_3359);
nor U3842 (N_3842,N_3258,N_3203);
and U3843 (N_3843,N_3472,N_3326);
and U3844 (N_3844,N_3446,N_3339);
and U3845 (N_3845,N_3418,N_3350);
xor U3846 (N_3846,N_3458,N_3403);
and U3847 (N_3847,N_3219,N_3227);
nand U3848 (N_3848,N_3051,N_3150);
nand U3849 (N_3849,N_3400,N_3154);
nor U3850 (N_3850,N_3390,N_3333);
nand U3851 (N_3851,N_3423,N_3130);
nor U3852 (N_3852,N_3359,N_3072);
nand U3853 (N_3853,N_3470,N_3210);
and U3854 (N_3854,N_3147,N_3344);
nor U3855 (N_3855,N_3417,N_3362);
nand U3856 (N_3856,N_3106,N_3005);
xor U3857 (N_3857,N_3363,N_3321);
and U3858 (N_3858,N_3156,N_3373);
or U3859 (N_3859,N_3114,N_3324);
or U3860 (N_3860,N_3383,N_3148);
nand U3861 (N_3861,N_3047,N_3375);
and U3862 (N_3862,N_3315,N_3405);
or U3863 (N_3863,N_3106,N_3268);
or U3864 (N_3864,N_3135,N_3067);
xnor U3865 (N_3865,N_3219,N_3156);
and U3866 (N_3866,N_3439,N_3053);
nor U3867 (N_3867,N_3379,N_3368);
nand U3868 (N_3868,N_3404,N_3057);
or U3869 (N_3869,N_3012,N_3143);
and U3870 (N_3870,N_3226,N_3350);
nor U3871 (N_3871,N_3477,N_3307);
xnor U3872 (N_3872,N_3086,N_3429);
nor U3873 (N_3873,N_3427,N_3290);
nand U3874 (N_3874,N_3174,N_3428);
or U3875 (N_3875,N_3443,N_3068);
nor U3876 (N_3876,N_3129,N_3023);
nand U3877 (N_3877,N_3153,N_3115);
or U3878 (N_3878,N_3150,N_3350);
nand U3879 (N_3879,N_3274,N_3359);
nand U3880 (N_3880,N_3229,N_3104);
nor U3881 (N_3881,N_3452,N_3431);
or U3882 (N_3882,N_3395,N_3228);
nand U3883 (N_3883,N_3317,N_3401);
nand U3884 (N_3884,N_3410,N_3389);
or U3885 (N_3885,N_3490,N_3063);
nor U3886 (N_3886,N_3008,N_3240);
or U3887 (N_3887,N_3123,N_3397);
nand U3888 (N_3888,N_3315,N_3139);
or U3889 (N_3889,N_3287,N_3056);
nor U3890 (N_3890,N_3397,N_3287);
or U3891 (N_3891,N_3121,N_3256);
or U3892 (N_3892,N_3110,N_3469);
or U3893 (N_3893,N_3068,N_3138);
nor U3894 (N_3894,N_3345,N_3205);
nor U3895 (N_3895,N_3122,N_3397);
and U3896 (N_3896,N_3467,N_3431);
or U3897 (N_3897,N_3093,N_3101);
and U3898 (N_3898,N_3142,N_3355);
or U3899 (N_3899,N_3211,N_3280);
nor U3900 (N_3900,N_3310,N_3398);
or U3901 (N_3901,N_3391,N_3059);
and U3902 (N_3902,N_3132,N_3120);
and U3903 (N_3903,N_3039,N_3199);
or U3904 (N_3904,N_3311,N_3045);
and U3905 (N_3905,N_3254,N_3456);
or U3906 (N_3906,N_3385,N_3048);
nor U3907 (N_3907,N_3018,N_3135);
nand U3908 (N_3908,N_3218,N_3292);
nor U3909 (N_3909,N_3037,N_3030);
nor U3910 (N_3910,N_3126,N_3341);
nand U3911 (N_3911,N_3482,N_3178);
nand U3912 (N_3912,N_3299,N_3166);
xor U3913 (N_3913,N_3331,N_3488);
nor U3914 (N_3914,N_3411,N_3289);
nor U3915 (N_3915,N_3408,N_3483);
and U3916 (N_3916,N_3258,N_3144);
and U3917 (N_3917,N_3007,N_3330);
or U3918 (N_3918,N_3111,N_3478);
or U3919 (N_3919,N_3494,N_3267);
nand U3920 (N_3920,N_3097,N_3300);
nor U3921 (N_3921,N_3173,N_3084);
or U3922 (N_3922,N_3309,N_3020);
nor U3923 (N_3923,N_3267,N_3247);
nand U3924 (N_3924,N_3110,N_3498);
nand U3925 (N_3925,N_3439,N_3038);
nand U3926 (N_3926,N_3063,N_3418);
and U3927 (N_3927,N_3235,N_3184);
xnor U3928 (N_3928,N_3194,N_3421);
nand U3929 (N_3929,N_3014,N_3421);
or U3930 (N_3930,N_3200,N_3181);
or U3931 (N_3931,N_3161,N_3017);
and U3932 (N_3932,N_3406,N_3256);
nor U3933 (N_3933,N_3491,N_3166);
nand U3934 (N_3934,N_3021,N_3259);
nand U3935 (N_3935,N_3077,N_3187);
or U3936 (N_3936,N_3404,N_3132);
nand U3937 (N_3937,N_3317,N_3256);
nor U3938 (N_3938,N_3279,N_3369);
nor U3939 (N_3939,N_3091,N_3359);
nand U3940 (N_3940,N_3222,N_3003);
nor U3941 (N_3941,N_3457,N_3064);
or U3942 (N_3942,N_3231,N_3128);
and U3943 (N_3943,N_3236,N_3021);
nand U3944 (N_3944,N_3308,N_3086);
or U3945 (N_3945,N_3480,N_3141);
nor U3946 (N_3946,N_3037,N_3365);
and U3947 (N_3947,N_3353,N_3404);
and U3948 (N_3948,N_3378,N_3233);
nor U3949 (N_3949,N_3191,N_3034);
nand U3950 (N_3950,N_3003,N_3304);
nand U3951 (N_3951,N_3078,N_3303);
nor U3952 (N_3952,N_3196,N_3351);
and U3953 (N_3953,N_3159,N_3160);
or U3954 (N_3954,N_3186,N_3373);
nand U3955 (N_3955,N_3378,N_3274);
nor U3956 (N_3956,N_3417,N_3166);
nand U3957 (N_3957,N_3165,N_3324);
nor U3958 (N_3958,N_3143,N_3465);
nand U3959 (N_3959,N_3452,N_3020);
and U3960 (N_3960,N_3015,N_3080);
nand U3961 (N_3961,N_3381,N_3375);
and U3962 (N_3962,N_3074,N_3488);
nor U3963 (N_3963,N_3277,N_3378);
nand U3964 (N_3964,N_3291,N_3461);
or U3965 (N_3965,N_3478,N_3416);
or U3966 (N_3966,N_3237,N_3309);
nor U3967 (N_3967,N_3299,N_3282);
or U3968 (N_3968,N_3105,N_3464);
nand U3969 (N_3969,N_3174,N_3020);
or U3970 (N_3970,N_3183,N_3280);
or U3971 (N_3971,N_3135,N_3253);
nand U3972 (N_3972,N_3268,N_3264);
and U3973 (N_3973,N_3357,N_3253);
or U3974 (N_3974,N_3123,N_3479);
or U3975 (N_3975,N_3474,N_3442);
and U3976 (N_3976,N_3497,N_3140);
nor U3977 (N_3977,N_3005,N_3157);
and U3978 (N_3978,N_3155,N_3068);
nand U3979 (N_3979,N_3496,N_3257);
xor U3980 (N_3980,N_3057,N_3479);
and U3981 (N_3981,N_3183,N_3144);
and U3982 (N_3982,N_3482,N_3365);
nand U3983 (N_3983,N_3392,N_3235);
and U3984 (N_3984,N_3408,N_3466);
nand U3985 (N_3985,N_3011,N_3435);
nand U3986 (N_3986,N_3216,N_3039);
nor U3987 (N_3987,N_3236,N_3326);
nand U3988 (N_3988,N_3470,N_3175);
or U3989 (N_3989,N_3400,N_3124);
or U3990 (N_3990,N_3429,N_3377);
nand U3991 (N_3991,N_3147,N_3006);
nor U3992 (N_3992,N_3461,N_3236);
nand U3993 (N_3993,N_3381,N_3275);
or U3994 (N_3994,N_3364,N_3230);
nor U3995 (N_3995,N_3278,N_3105);
or U3996 (N_3996,N_3222,N_3432);
xor U3997 (N_3997,N_3184,N_3050);
nand U3998 (N_3998,N_3137,N_3106);
or U3999 (N_3999,N_3083,N_3128);
and U4000 (N_4000,N_3874,N_3705);
and U4001 (N_4001,N_3582,N_3509);
nand U4002 (N_4002,N_3899,N_3568);
nor U4003 (N_4003,N_3867,N_3846);
nor U4004 (N_4004,N_3937,N_3974);
nor U4005 (N_4005,N_3826,N_3779);
and U4006 (N_4006,N_3812,N_3680);
or U4007 (N_4007,N_3518,N_3638);
or U4008 (N_4008,N_3947,N_3813);
and U4009 (N_4009,N_3612,N_3967);
nor U4010 (N_4010,N_3957,N_3527);
nor U4011 (N_4011,N_3965,N_3619);
nand U4012 (N_4012,N_3713,N_3584);
nor U4013 (N_4013,N_3766,N_3905);
nor U4014 (N_4014,N_3685,N_3927);
or U4015 (N_4015,N_3842,N_3629);
nand U4016 (N_4016,N_3697,N_3637);
or U4017 (N_4017,N_3662,N_3576);
and U4018 (N_4018,N_3581,N_3722);
nand U4019 (N_4019,N_3661,N_3636);
nand U4020 (N_4020,N_3740,N_3736);
or U4021 (N_4021,N_3550,N_3829);
nor U4022 (N_4022,N_3989,N_3700);
and U4023 (N_4023,N_3635,N_3792);
xnor U4024 (N_4024,N_3903,N_3843);
or U4025 (N_4025,N_3593,N_3839);
and U4026 (N_4026,N_3849,N_3693);
xor U4027 (N_4027,N_3799,N_3953);
or U4028 (N_4028,N_3923,N_3652);
or U4029 (N_4029,N_3746,N_3984);
and U4030 (N_4030,N_3978,N_3748);
nand U4031 (N_4031,N_3827,N_3528);
or U4032 (N_4032,N_3971,N_3726);
and U4033 (N_4033,N_3871,N_3882);
nand U4034 (N_4034,N_3515,N_3969);
nand U4035 (N_4035,N_3698,N_3963);
nor U4036 (N_4036,N_3993,N_3720);
or U4037 (N_4037,N_3920,N_3526);
or U4038 (N_4038,N_3870,N_3679);
or U4039 (N_4039,N_3998,N_3815);
or U4040 (N_4040,N_3500,N_3694);
nor U4041 (N_4041,N_3966,N_3621);
and U4042 (N_4042,N_3864,N_3541);
and U4043 (N_4043,N_3944,N_3702);
or U4044 (N_4044,N_3511,N_3837);
and U4045 (N_4045,N_3625,N_3530);
and U4046 (N_4046,N_3687,N_3883);
and U4047 (N_4047,N_3686,N_3996);
or U4048 (N_4048,N_3880,N_3602);
nor U4049 (N_4049,N_3639,N_3531);
or U4050 (N_4050,N_3761,N_3537);
nand U4051 (N_4051,N_3900,N_3768);
nor U4052 (N_4052,N_3804,N_3868);
nand U4053 (N_4053,N_3847,N_3943);
nor U4054 (N_4054,N_3630,N_3573);
nor U4055 (N_4055,N_3933,N_3520);
nand U4056 (N_4056,N_3838,N_3668);
or U4057 (N_4057,N_3818,N_3773);
nor U4058 (N_4058,N_3725,N_3563);
nor U4059 (N_4059,N_3708,N_3982);
or U4060 (N_4060,N_3854,N_3578);
and U4061 (N_4061,N_3795,N_3556);
and U4062 (N_4062,N_3850,N_3566);
nor U4063 (N_4063,N_3523,N_3809);
and U4064 (N_4064,N_3760,N_3559);
nand U4065 (N_4065,N_3605,N_3771);
nand U4066 (N_4066,N_3791,N_3912);
and U4067 (N_4067,N_3876,N_3924);
or U4068 (N_4068,N_3921,N_3750);
nor U4069 (N_4069,N_3613,N_3805);
and U4070 (N_4070,N_3904,N_3825);
and U4071 (N_4071,N_3606,N_3915);
or U4072 (N_4072,N_3911,N_3611);
and U4073 (N_4073,N_3819,N_3742);
or U4074 (N_4074,N_3930,N_3738);
or U4075 (N_4075,N_3782,N_3951);
nand U4076 (N_4076,N_3586,N_3767);
nor U4077 (N_4077,N_3683,N_3862);
and U4078 (N_4078,N_3517,N_3892);
nor U4079 (N_4079,N_3999,N_3536);
and U4080 (N_4080,N_3848,N_3735);
nor U4081 (N_4081,N_3522,N_3962);
nor U4082 (N_4082,N_3806,N_3657);
nand U4083 (N_4083,N_3567,N_3810);
or U4084 (N_4084,N_3589,N_3929);
nand U4085 (N_4085,N_3754,N_3734);
and U4086 (N_4086,N_3594,N_3591);
nor U4087 (N_4087,N_3908,N_3814);
and U4088 (N_4088,N_3666,N_3519);
nand U4089 (N_4089,N_3769,N_3684);
and U4090 (N_4090,N_3763,N_3615);
or U4091 (N_4091,N_3506,N_3762);
nand U4092 (N_4092,N_3873,N_3676);
nor U4093 (N_4093,N_3744,N_3587);
or U4094 (N_4094,N_3885,N_3745);
or U4095 (N_4095,N_3898,N_3564);
nor U4096 (N_4096,N_3709,N_3616);
nor U4097 (N_4097,N_3758,N_3626);
nand U4098 (N_4098,N_3831,N_3878);
and U4099 (N_4099,N_3865,N_3730);
or U4100 (N_4100,N_3647,N_3986);
and U4101 (N_4101,N_3835,N_3718);
xnor U4102 (N_4102,N_3764,N_3670);
nor U4103 (N_4103,N_3671,N_3942);
xor U4104 (N_4104,N_3816,N_3712);
nand U4105 (N_4105,N_3936,N_3757);
xor U4106 (N_4106,N_3858,N_3570);
nor U4107 (N_4107,N_3675,N_3560);
nand U4108 (N_4108,N_3981,N_3886);
and U4109 (N_4109,N_3514,N_3588);
and U4110 (N_4110,N_3704,N_3901);
nor U4111 (N_4111,N_3565,N_3884);
nor U4112 (N_4112,N_3893,N_3516);
nor U4113 (N_4113,N_3557,N_3706);
nor U4114 (N_4114,N_3549,N_3833);
and U4115 (N_4115,N_3583,N_3665);
nor U4116 (N_4116,N_3774,N_3751);
and U4117 (N_4117,N_3599,N_3717);
or U4118 (N_4118,N_3551,N_3945);
and U4119 (N_4119,N_3590,N_3729);
nand U4120 (N_4120,N_3501,N_3907);
or U4121 (N_4121,N_3617,N_3650);
and U4122 (N_4122,N_3658,N_3783);
and U4123 (N_4123,N_3949,N_3925);
or U4124 (N_4124,N_3562,N_3844);
nand U4125 (N_4125,N_3968,N_3983);
nor U4126 (N_4126,N_3571,N_3631);
or U4127 (N_4127,N_3985,N_3772);
nor U4128 (N_4128,N_3752,N_3765);
nand U4129 (N_4129,N_3926,N_3823);
or U4130 (N_4130,N_3906,N_3545);
nand U4131 (N_4131,N_3728,N_3741);
nor U4132 (N_4132,N_3866,N_3995);
or U4133 (N_4133,N_3990,N_3948);
nand U4134 (N_4134,N_3916,N_3524);
nand U4135 (N_4135,N_3723,N_3651);
or U4136 (N_4136,N_3778,N_3955);
nand U4137 (N_4137,N_3853,N_3505);
nand U4138 (N_4138,N_3879,N_3543);
and U4139 (N_4139,N_3950,N_3913);
and U4140 (N_4140,N_3610,N_3634);
or U4141 (N_4141,N_3707,N_3852);
nand U4142 (N_4142,N_3784,N_3747);
or U4143 (N_4143,N_3572,N_3733);
nor U4144 (N_4144,N_3688,N_3869);
nor U4145 (N_4145,N_3737,N_3644);
and U4146 (N_4146,N_3811,N_3859);
nand U4147 (N_4147,N_3664,N_3719);
nand U4148 (N_4148,N_3695,N_3622);
nor U4149 (N_4149,N_3932,N_3817);
or U4150 (N_4150,N_3624,N_3532);
nand U4151 (N_4151,N_3682,N_3787);
nand U4152 (N_4152,N_3609,N_3896);
or U4153 (N_4153,N_3958,N_3699);
xnor U4154 (N_4154,N_3632,N_3788);
nand U4155 (N_4155,N_3672,N_3863);
or U4156 (N_4156,N_3994,N_3979);
nand U4157 (N_4157,N_3830,N_3663);
and U4158 (N_4158,N_3739,N_3715);
nor U4159 (N_4159,N_3701,N_3753);
xor U4160 (N_4160,N_3759,N_3521);
nand U4161 (N_4161,N_3931,N_3976);
and U4162 (N_4162,N_3659,N_3939);
and U4163 (N_4163,N_3975,N_3535);
nor U4164 (N_4164,N_3653,N_3643);
nor U4165 (N_4165,N_3674,N_3832);
nor U4166 (N_4166,N_3775,N_3724);
or U4167 (N_4167,N_3561,N_3623);
and U4168 (N_4168,N_3614,N_3529);
and U4169 (N_4169,N_3889,N_3642);
and U4170 (N_4170,N_3840,N_3800);
and U4171 (N_4171,N_3618,N_3977);
and U4172 (N_4172,N_3881,N_3544);
nor U4173 (N_4173,N_3952,N_3956);
nand U4174 (N_4174,N_3628,N_3553);
nand U4175 (N_4175,N_3732,N_3770);
nor U4176 (N_4176,N_3510,N_3743);
and U4177 (N_4177,N_3992,N_3660);
nand U4178 (N_4178,N_3954,N_3872);
nand U4179 (N_4179,N_3959,N_3897);
nand U4180 (N_4180,N_3703,N_3710);
nor U4181 (N_4181,N_3888,N_3756);
xor U4182 (N_4182,N_3542,N_3558);
and U4183 (N_4183,N_3727,N_3857);
and U4184 (N_4184,N_3777,N_3714);
nand U4185 (N_4185,N_3692,N_3533);
nor U4186 (N_4186,N_3946,N_3538);
nor U4187 (N_4187,N_3780,N_3877);
xor U4188 (N_4188,N_3673,N_3796);
and U4189 (N_4189,N_3656,N_3716);
nand U4190 (N_4190,N_3861,N_3938);
nor U4191 (N_4191,N_3824,N_3860);
or U4192 (N_4192,N_3807,N_3547);
or U4193 (N_4193,N_3988,N_3513);
nor U4194 (N_4194,N_3790,N_3502);
and U4195 (N_4195,N_3855,N_3603);
and U4196 (N_4196,N_3934,N_3546);
nor U4197 (N_4197,N_3525,N_3940);
or U4198 (N_4198,N_3677,N_3534);
or U4199 (N_4199,N_3711,N_3890);
and U4200 (N_4200,N_3928,N_3834);
or U4201 (N_4201,N_3776,N_3555);
or U4202 (N_4202,N_3808,N_3902);
nand U4203 (N_4203,N_3972,N_3973);
nor U4204 (N_4204,N_3601,N_3935);
nor U4205 (N_4205,N_3633,N_3909);
xnor U4206 (N_4206,N_3580,N_3669);
or U4207 (N_4207,N_3991,N_3607);
and U4208 (N_4208,N_3895,N_3781);
or U4209 (N_4209,N_3941,N_3654);
nor U4210 (N_4210,N_3577,N_3786);
and U4211 (N_4211,N_3667,N_3851);
nand U4212 (N_4212,N_3845,N_3964);
and U4213 (N_4213,N_3887,N_3822);
and U4214 (N_4214,N_3919,N_3649);
and U4215 (N_4215,N_3678,N_3841);
or U4216 (N_4216,N_3596,N_3980);
nor U4217 (N_4217,N_3970,N_3689);
nor U4218 (N_4218,N_3585,N_3721);
or U4219 (N_4219,N_3548,N_3648);
nor U4220 (N_4220,N_3821,N_3828);
nand U4221 (N_4221,N_3856,N_3627);
nand U4222 (N_4222,N_3575,N_3798);
nor U4223 (N_4223,N_3655,N_3598);
and U4224 (N_4224,N_3503,N_3802);
or U4225 (N_4225,N_3987,N_3691);
and U4226 (N_4226,N_3641,N_3910);
nand U4227 (N_4227,N_3681,N_3597);
or U4228 (N_4228,N_3731,N_3640);
or U4229 (N_4229,N_3961,N_3917);
nor U4230 (N_4230,N_3574,N_3960);
nor U4231 (N_4231,N_3785,N_3793);
nand U4232 (N_4232,N_3755,N_3891);
and U4233 (N_4233,N_3600,N_3569);
nor U4234 (N_4234,N_3801,N_3997);
and U4235 (N_4235,N_3579,N_3789);
nor U4236 (N_4236,N_3592,N_3820);
or U4237 (N_4237,N_3539,N_3836);
or U4238 (N_4238,N_3646,N_3645);
and U4239 (N_4239,N_3914,N_3696);
or U4240 (N_4240,N_3554,N_3507);
xnor U4241 (N_4241,N_3894,N_3540);
nor U4242 (N_4242,N_3604,N_3794);
nand U4243 (N_4243,N_3803,N_3749);
and U4244 (N_4244,N_3620,N_3552);
and U4245 (N_4245,N_3508,N_3608);
or U4246 (N_4246,N_3875,N_3922);
xor U4247 (N_4247,N_3797,N_3690);
or U4248 (N_4248,N_3512,N_3595);
nor U4249 (N_4249,N_3504,N_3918);
or U4250 (N_4250,N_3846,N_3661);
nand U4251 (N_4251,N_3717,N_3694);
nand U4252 (N_4252,N_3632,N_3502);
and U4253 (N_4253,N_3522,N_3889);
or U4254 (N_4254,N_3616,N_3711);
and U4255 (N_4255,N_3971,N_3534);
nor U4256 (N_4256,N_3964,N_3953);
nor U4257 (N_4257,N_3741,N_3639);
or U4258 (N_4258,N_3808,N_3648);
nor U4259 (N_4259,N_3905,N_3808);
xor U4260 (N_4260,N_3998,N_3903);
or U4261 (N_4261,N_3998,N_3975);
nand U4262 (N_4262,N_3960,N_3533);
and U4263 (N_4263,N_3582,N_3652);
nor U4264 (N_4264,N_3728,N_3793);
nor U4265 (N_4265,N_3639,N_3923);
or U4266 (N_4266,N_3842,N_3724);
nand U4267 (N_4267,N_3826,N_3842);
or U4268 (N_4268,N_3555,N_3730);
and U4269 (N_4269,N_3658,N_3739);
nand U4270 (N_4270,N_3707,N_3727);
and U4271 (N_4271,N_3553,N_3731);
nor U4272 (N_4272,N_3935,N_3727);
and U4273 (N_4273,N_3942,N_3627);
nor U4274 (N_4274,N_3859,N_3770);
or U4275 (N_4275,N_3638,N_3642);
nand U4276 (N_4276,N_3657,N_3761);
or U4277 (N_4277,N_3856,N_3831);
nor U4278 (N_4278,N_3813,N_3550);
and U4279 (N_4279,N_3849,N_3610);
or U4280 (N_4280,N_3673,N_3794);
nor U4281 (N_4281,N_3873,N_3963);
and U4282 (N_4282,N_3921,N_3752);
and U4283 (N_4283,N_3650,N_3552);
xnor U4284 (N_4284,N_3503,N_3782);
nand U4285 (N_4285,N_3555,N_3821);
xor U4286 (N_4286,N_3864,N_3576);
nor U4287 (N_4287,N_3775,N_3783);
or U4288 (N_4288,N_3761,N_3662);
or U4289 (N_4289,N_3851,N_3732);
or U4290 (N_4290,N_3654,N_3980);
xor U4291 (N_4291,N_3987,N_3802);
nand U4292 (N_4292,N_3743,N_3873);
nand U4293 (N_4293,N_3570,N_3667);
nor U4294 (N_4294,N_3763,N_3717);
nor U4295 (N_4295,N_3680,N_3808);
and U4296 (N_4296,N_3825,N_3675);
or U4297 (N_4297,N_3967,N_3677);
or U4298 (N_4298,N_3597,N_3756);
nand U4299 (N_4299,N_3842,N_3542);
or U4300 (N_4300,N_3506,N_3722);
nand U4301 (N_4301,N_3714,N_3665);
nor U4302 (N_4302,N_3889,N_3634);
nand U4303 (N_4303,N_3898,N_3576);
or U4304 (N_4304,N_3939,N_3886);
and U4305 (N_4305,N_3792,N_3534);
nor U4306 (N_4306,N_3831,N_3673);
and U4307 (N_4307,N_3921,N_3815);
and U4308 (N_4308,N_3937,N_3522);
and U4309 (N_4309,N_3824,N_3937);
or U4310 (N_4310,N_3728,N_3779);
nand U4311 (N_4311,N_3588,N_3528);
or U4312 (N_4312,N_3789,N_3838);
or U4313 (N_4313,N_3864,N_3794);
and U4314 (N_4314,N_3919,N_3664);
or U4315 (N_4315,N_3985,N_3716);
nor U4316 (N_4316,N_3638,N_3607);
nand U4317 (N_4317,N_3656,N_3536);
nor U4318 (N_4318,N_3952,N_3736);
or U4319 (N_4319,N_3633,N_3591);
or U4320 (N_4320,N_3701,N_3970);
nand U4321 (N_4321,N_3918,N_3660);
and U4322 (N_4322,N_3551,N_3826);
or U4323 (N_4323,N_3890,N_3649);
or U4324 (N_4324,N_3576,N_3530);
nor U4325 (N_4325,N_3676,N_3976);
and U4326 (N_4326,N_3745,N_3667);
nand U4327 (N_4327,N_3840,N_3601);
and U4328 (N_4328,N_3673,N_3975);
nor U4329 (N_4329,N_3825,N_3740);
or U4330 (N_4330,N_3897,N_3739);
nand U4331 (N_4331,N_3714,N_3766);
nand U4332 (N_4332,N_3901,N_3665);
nor U4333 (N_4333,N_3869,N_3775);
nor U4334 (N_4334,N_3968,N_3678);
or U4335 (N_4335,N_3831,N_3678);
or U4336 (N_4336,N_3808,N_3735);
nand U4337 (N_4337,N_3539,N_3631);
and U4338 (N_4338,N_3942,N_3658);
nand U4339 (N_4339,N_3877,N_3798);
nand U4340 (N_4340,N_3592,N_3994);
nor U4341 (N_4341,N_3602,N_3888);
nor U4342 (N_4342,N_3512,N_3810);
nand U4343 (N_4343,N_3621,N_3914);
and U4344 (N_4344,N_3734,N_3697);
or U4345 (N_4345,N_3683,N_3979);
nor U4346 (N_4346,N_3840,N_3727);
and U4347 (N_4347,N_3875,N_3566);
or U4348 (N_4348,N_3889,N_3808);
nor U4349 (N_4349,N_3765,N_3530);
nor U4350 (N_4350,N_3958,N_3689);
nand U4351 (N_4351,N_3659,N_3623);
or U4352 (N_4352,N_3862,N_3607);
or U4353 (N_4353,N_3689,N_3624);
or U4354 (N_4354,N_3576,N_3690);
nor U4355 (N_4355,N_3834,N_3968);
nand U4356 (N_4356,N_3623,N_3874);
nor U4357 (N_4357,N_3509,N_3793);
and U4358 (N_4358,N_3705,N_3726);
or U4359 (N_4359,N_3641,N_3809);
or U4360 (N_4360,N_3720,N_3680);
nand U4361 (N_4361,N_3807,N_3769);
or U4362 (N_4362,N_3540,N_3520);
or U4363 (N_4363,N_3604,N_3702);
and U4364 (N_4364,N_3644,N_3845);
and U4365 (N_4365,N_3861,N_3740);
nand U4366 (N_4366,N_3706,N_3773);
or U4367 (N_4367,N_3642,N_3542);
and U4368 (N_4368,N_3880,N_3761);
nand U4369 (N_4369,N_3891,N_3783);
or U4370 (N_4370,N_3816,N_3619);
or U4371 (N_4371,N_3577,N_3518);
and U4372 (N_4372,N_3509,N_3660);
nor U4373 (N_4373,N_3922,N_3681);
nand U4374 (N_4374,N_3975,N_3656);
or U4375 (N_4375,N_3862,N_3557);
nand U4376 (N_4376,N_3892,N_3545);
and U4377 (N_4377,N_3555,N_3706);
or U4378 (N_4378,N_3876,N_3543);
or U4379 (N_4379,N_3694,N_3730);
and U4380 (N_4380,N_3813,N_3729);
or U4381 (N_4381,N_3986,N_3909);
nor U4382 (N_4382,N_3636,N_3563);
and U4383 (N_4383,N_3573,N_3827);
and U4384 (N_4384,N_3968,N_3926);
nor U4385 (N_4385,N_3722,N_3540);
nor U4386 (N_4386,N_3731,N_3915);
nor U4387 (N_4387,N_3846,N_3544);
and U4388 (N_4388,N_3586,N_3642);
nand U4389 (N_4389,N_3680,N_3741);
and U4390 (N_4390,N_3649,N_3664);
nand U4391 (N_4391,N_3992,N_3697);
nand U4392 (N_4392,N_3732,N_3947);
and U4393 (N_4393,N_3627,N_3758);
or U4394 (N_4394,N_3717,N_3509);
nor U4395 (N_4395,N_3586,N_3916);
nor U4396 (N_4396,N_3575,N_3572);
or U4397 (N_4397,N_3944,N_3530);
and U4398 (N_4398,N_3690,N_3782);
and U4399 (N_4399,N_3539,N_3681);
or U4400 (N_4400,N_3626,N_3885);
nand U4401 (N_4401,N_3896,N_3877);
nand U4402 (N_4402,N_3993,N_3918);
nand U4403 (N_4403,N_3995,N_3984);
nor U4404 (N_4404,N_3535,N_3549);
and U4405 (N_4405,N_3682,N_3899);
nor U4406 (N_4406,N_3584,N_3856);
and U4407 (N_4407,N_3514,N_3698);
or U4408 (N_4408,N_3588,N_3690);
nand U4409 (N_4409,N_3891,N_3823);
and U4410 (N_4410,N_3515,N_3595);
nor U4411 (N_4411,N_3536,N_3705);
and U4412 (N_4412,N_3597,N_3840);
nand U4413 (N_4413,N_3615,N_3978);
and U4414 (N_4414,N_3920,N_3852);
nand U4415 (N_4415,N_3884,N_3504);
nand U4416 (N_4416,N_3620,N_3652);
and U4417 (N_4417,N_3650,N_3786);
or U4418 (N_4418,N_3965,N_3606);
nand U4419 (N_4419,N_3830,N_3823);
and U4420 (N_4420,N_3661,N_3592);
nand U4421 (N_4421,N_3745,N_3829);
or U4422 (N_4422,N_3698,N_3526);
nor U4423 (N_4423,N_3999,N_3830);
nor U4424 (N_4424,N_3984,N_3700);
nor U4425 (N_4425,N_3935,N_3773);
and U4426 (N_4426,N_3746,N_3710);
nand U4427 (N_4427,N_3814,N_3975);
nor U4428 (N_4428,N_3532,N_3916);
nor U4429 (N_4429,N_3510,N_3540);
and U4430 (N_4430,N_3837,N_3784);
nor U4431 (N_4431,N_3654,N_3951);
nand U4432 (N_4432,N_3731,N_3892);
and U4433 (N_4433,N_3847,N_3554);
nand U4434 (N_4434,N_3730,N_3981);
and U4435 (N_4435,N_3809,N_3564);
and U4436 (N_4436,N_3821,N_3829);
or U4437 (N_4437,N_3656,N_3646);
and U4438 (N_4438,N_3500,N_3712);
nand U4439 (N_4439,N_3519,N_3802);
nor U4440 (N_4440,N_3772,N_3950);
nand U4441 (N_4441,N_3931,N_3537);
nand U4442 (N_4442,N_3606,N_3563);
or U4443 (N_4443,N_3594,N_3877);
nor U4444 (N_4444,N_3744,N_3809);
or U4445 (N_4445,N_3675,N_3885);
nor U4446 (N_4446,N_3813,N_3841);
and U4447 (N_4447,N_3716,N_3760);
or U4448 (N_4448,N_3788,N_3936);
and U4449 (N_4449,N_3922,N_3807);
nor U4450 (N_4450,N_3980,N_3684);
nand U4451 (N_4451,N_3683,N_3934);
and U4452 (N_4452,N_3941,N_3959);
nand U4453 (N_4453,N_3778,N_3571);
and U4454 (N_4454,N_3661,N_3812);
and U4455 (N_4455,N_3908,N_3866);
and U4456 (N_4456,N_3743,N_3920);
and U4457 (N_4457,N_3628,N_3964);
or U4458 (N_4458,N_3578,N_3590);
nor U4459 (N_4459,N_3946,N_3738);
or U4460 (N_4460,N_3808,N_3795);
nor U4461 (N_4461,N_3500,N_3737);
nand U4462 (N_4462,N_3799,N_3849);
nand U4463 (N_4463,N_3987,N_3684);
nor U4464 (N_4464,N_3787,N_3996);
and U4465 (N_4465,N_3796,N_3589);
nor U4466 (N_4466,N_3924,N_3665);
nand U4467 (N_4467,N_3842,N_3893);
nand U4468 (N_4468,N_3923,N_3771);
nand U4469 (N_4469,N_3762,N_3659);
or U4470 (N_4470,N_3666,N_3850);
xor U4471 (N_4471,N_3640,N_3550);
nand U4472 (N_4472,N_3750,N_3993);
or U4473 (N_4473,N_3522,N_3908);
and U4474 (N_4474,N_3550,N_3755);
nand U4475 (N_4475,N_3895,N_3692);
nor U4476 (N_4476,N_3527,N_3529);
nor U4477 (N_4477,N_3719,N_3721);
and U4478 (N_4478,N_3634,N_3867);
nand U4479 (N_4479,N_3803,N_3617);
nor U4480 (N_4480,N_3612,N_3540);
xor U4481 (N_4481,N_3751,N_3661);
nand U4482 (N_4482,N_3775,N_3549);
and U4483 (N_4483,N_3714,N_3823);
nand U4484 (N_4484,N_3928,N_3922);
and U4485 (N_4485,N_3922,N_3566);
nor U4486 (N_4486,N_3859,N_3661);
or U4487 (N_4487,N_3977,N_3749);
or U4488 (N_4488,N_3787,N_3889);
or U4489 (N_4489,N_3736,N_3923);
nand U4490 (N_4490,N_3691,N_3523);
nand U4491 (N_4491,N_3769,N_3850);
and U4492 (N_4492,N_3630,N_3709);
and U4493 (N_4493,N_3896,N_3663);
nor U4494 (N_4494,N_3756,N_3587);
nor U4495 (N_4495,N_3535,N_3629);
or U4496 (N_4496,N_3648,N_3636);
nand U4497 (N_4497,N_3644,N_3959);
or U4498 (N_4498,N_3676,N_3637);
nor U4499 (N_4499,N_3788,N_3961);
nand U4500 (N_4500,N_4019,N_4497);
nor U4501 (N_4501,N_4456,N_4040);
nor U4502 (N_4502,N_4293,N_4350);
nand U4503 (N_4503,N_4191,N_4383);
and U4504 (N_4504,N_4169,N_4227);
and U4505 (N_4505,N_4374,N_4206);
nor U4506 (N_4506,N_4335,N_4312);
nor U4507 (N_4507,N_4268,N_4309);
nand U4508 (N_4508,N_4449,N_4194);
nor U4509 (N_4509,N_4247,N_4379);
and U4510 (N_4510,N_4468,N_4278);
nor U4511 (N_4511,N_4317,N_4226);
nand U4512 (N_4512,N_4238,N_4001);
nand U4513 (N_4513,N_4286,N_4410);
nand U4514 (N_4514,N_4302,N_4065);
nand U4515 (N_4515,N_4400,N_4341);
nand U4516 (N_4516,N_4114,N_4057);
nand U4517 (N_4517,N_4061,N_4440);
nand U4518 (N_4518,N_4337,N_4181);
nor U4519 (N_4519,N_4241,N_4078);
nand U4520 (N_4520,N_4289,N_4467);
or U4521 (N_4521,N_4232,N_4305);
and U4522 (N_4522,N_4397,N_4420);
nor U4523 (N_4523,N_4474,N_4407);
nand U4524 (N_4524,N_4259,N_4127);
nand U4525 (N_4525,N_4217,N_4149);
nor U4526 (N_4526,N_4074,N_4415);
nand U4527 (N_4527,N_4130,N_4208);
nand U4528 (N_4528,N_4178,N_4366);
and U4529 (N_4529,N_4160,N_4129);
nand U4530 (N_4530,N_4154,N_4105);
nor U4531 (N_4531,N_4425,N_4116);
nand U4532 (N_4532,N_4324,N_4347);
and U4533 (N_4533,N_4359,N_4058);
and U4534 (N_4534,N_4257,N_4368);
and U4535 (N_4535,N_4325,N_4031);
xor U4536 (N_4536,N_4292,N_4024);
or U4537 (N_4537,N_4012,N_4071);
or U4538 (N_4538,N_4205,N_4180);
or U4539 (N_4539,N_4103,N_4321);
or U4540 (N_4540,N_4336,N_4492);
nor U4541 (N_4541,N_4250,N_4426);
or U4542 (N_4542,N_4150,N_4135);
nor U4543 (N_4543,N_4446,N_4291);
and U4544 (N_4544,N_4199,N_4326);
or U4545 (N_4545,N_4120,N_4053);
or U4546 (N_4546,N_4087,N_4331);
nor U4547 (N_4547,N_4046,N_4088);
nand U4548 (N_4548,N_4195,N_4263);
nand U4549 (N_4549,N_4436,N_4262);
or U4550 (N_4550,N_4008,N_4264);
or U4551 (N_4551,N_4138,N_4075);
or U4552 (N_4552,N_4281,N_4006);
and U4553 (N_4553,N_4295,N_4102);
or U4554 (N_4554,N_4387,N_4451);
nor U4555 (N_4555,N_4245,N_4280);
and U4556 (N_4556,N_4219,N_4340);
and U4557 (N_4557,N_4274,N_4435);
nand U4558 (N_4558,N_4363,N_4398);
or U4559 (N_4559,N_4030,N_4438);
nand U4560 (N_4560,N_4299,N_4026);
nand U4561 (N_4561,N_4485,N_4318);
or U4562 (N_4562,N_4266,N_4197);
nand U4563 (N_4563,N_4351,N_4002);
and U4564 (N_4564,N_4444,N_4142);
or U4565 (N_4565,N_4342,N_4077);
xor U4566 (N_4566,N_4352,N_4434);
nor U4567 (N_4567,N_4156,N_4308);
nand U4568 (N_4568,N_4210,N_4171);
or U4569 (N_4569,N_4399,N_4069);
and U4570 (N_4570,N_4055,N_4394);
or U4571 (N_4571,N_4240,N_4211);
or U4572 (N_4572,N_4223,N_4361);
nand U4573 (N_4573,N_4028,N_4025);
and U4574 (N_4574,N_4005,N_4424);
or U4575 (N_4575,N_4381,N_4465);
or U4576 (N_4576,N_4373,N_4237);
nor U4577 (N_4577,N_4107,N_4354);
or U4578 (N_4578,N_4477,N_4345);
and U4579 (N_4579,N_4148,N_4097);
or U4580 (N_4580,N_4496,N_4329);
nand U4581 (N_4581,N_4183,N_4125);
or U4582 (N_4582,N_4495,N_4165);
and U4583 (N_4583,N_4290,N_4306);
or U4584 (N_4584,N_4301,N_4121);
nor U4585 (N_4585,N_4411,N_4172);
or U4586 (N_4586,N_4020,N_4119);
nor U4587 (N_4587,N_4101,N_4060);
nand U4588 (N_4588,N_4460,N_4035);
or U4589 (N_4589,N_4146,N_4215);
nand U4590 (N_4590,N_4117,N_4041);
and U4591 (N_4591,N_4021,N_4083);
nand U4592 (N_4592,N_4419,N_4187);
nor U4593 (N_4593,N_4243,N_4311);
and U4594 (N_4594,N_4168,N_4304);
or U4595 (N_4595,N_4099,N_4010);
and U4596 (N_4596,N_4173,N_4430);
nor U4597 (N_4597,N_4182,N_4421);
nor U4598 (N_4598,N_4098,N_4360);
nand U4599 (N_4599,N_4086,N_4044);
or U4600 (N_4600,N_4249,N_4463);
nor U4601 (N_4601,N_4380,N_4470);
xor U4602 (N_4602,N_4313,N_4045);
and U4603 (N_4603,N_4155,N_4126);
xor U4604 (N_4604,N_4104,N_4170);
nor U4605 (N_4605,N_4386,N_4017);
nor U4606 (N_4606,N_4252,N_4242);
nand U4607 (N_4607,N_4151,N_4370);
nand U4608 (N_4608,N_4458,N_4490);
nor U4609 (N_4609,N_4275,N_4375);
nor U4610 (N_4610,N_4417,N_4000);
nor U4611 (N_4611,N_4433,N_4482);
xor U4612 (N_4612,N_4052,N_4073);
nor U4613 (N_4613,N_4174,N_4498);
and U4614 (N_4614,N_4461,N_4176);
and U4615 (N_4615,N_4315,N_4228);
and U4616 (N_4616,N_4473,N_4453);
and U4617 (N_4617,N_4332,N_4395);
nor U4618 (N_4618,N_4207,N_4486);
nand U4619 (N_4619,N_4251,N_4034);
nor U4620 (N_4620,N_4392,N_4239);
nor U4621 (N_4621,N_4036,N_4288);
nor U4622 (N_4622,N_4277,N_4344);
nand U4623 (N_4623,N_4287,N_4300);
and U4624 (N_4624,N_4488,N_4457);
nand U4625 (N_4625,N_4179,N_4016);
or U4626 (N_4626,N_4464,N_4070);
and U4627 (N_4627,N_4225,N_4202);
nor U4628 (N_4628,N_4011,N_4231);
nand U4629 (N_4629,N_4201,N_4050);
nor U4630 (N_4630,N_4455,N_4448);
and U4631 (N_4631,N_4106,N_4412);
or U4632 (N_4632,N_4362,N_4294);
and U4633 (N_4633,N_4100,N_4283);
or U4634 (N_4634,N_4066,N_4186);
and U4635 (N_4635,N_4144,N_4447);
and U4636 (N_4636,N_4188,N_4338);
nor U4637 (N_4637,N_4109,N_4385);
nand U4638 (N_4638,N_4391,N_4079);
nand U4639 (N_4639,N_4431,N_4054);
nand U4640 (N_4640,N_4153,N_4285);
and U4641 (N_4641,N_4082,N_4462);
and U4642 (N_4642,N_4246,N_4184);
nand U4643 (N_4643,N_4093,N_4364);
and U4644 (N_4644,N_4409,N_4235);
or U4645 (N_4645,N_4320,N_4175);
nor U4646 (N_4646,N_4037,N_4346);
nand U4647 (N_4647,N_4244,N_4218);
or U4648 (N_4648,N_4203,N_4084);
and U4649 (N_4649,N_4166,N_4200);
or U4650 (N_4650,N_4479,N_4229);
nor U4651 (N_4651,N_4159,N_4416);
nor U4652 (N_4652,N_4272,N_4112);
xor U4653 (N_4653,N_4377,N_4459);
and U4654 (N_4654,N_4115,N_4494);
or U4655 (N_4655,N_4389,N_4152);
and U4656 (N_4656,N_4039,N_4038);
and U4657 (N_4657,N_4167,N_4357);
nand U4658 (N_4658,N_4056,N_4406);
nor U4659 (N_4659,N_4224,N_4110);
and U4660 (N_4660,N_4404,N_4483);
nor U4661 (N_4661,N_4390,N_4253);
or U4662 (N_4662,N_4085,N_4233);
nand U4663 (N_4663,N_4469,N_4216);
nand U4664 (N_4664,N_4348,N_4096);
nor U4665 (N_4665,N_4185,N_4319);
nor U4666 (N_4666,N_4248,N_4282);
or U4667 (N_4667,N_4343,N_4284);
nor U4668 (N_4668,N_4261,N_4372);
and U4669 (N_4669,N_4090,N_4443);
and U4670 (N_4670,N_4450,N_4429);
nor U4671 (N_4671,N_4113,N_4297);
and U4672 (N_4672,N_4134,N_4439);
nand U4673 (N_4673,N_4478,N_4273);
or U4674 (N_4674,N_4234,N_4310);
and U4675 (N_4675,N_4396,N_4163);
and U4676 (N_4676,N_4256,N_4442);
and U4677 (N_4677,N_4047,N_4189);
or U4678 (N_4678,N_4128,N_4303);
and U4679 (N_4679,N_4314,N_4428);
nor U4680 (N_4680,N_4158,N_4371);
nor U4681 (N_4681,N_4405,N_4339);
and U4682 (N_4682,N_4132,N_4164);
and U4683 (N_4683,N_4489,N_4422);
or U4684 (N_4684,N_4269,N_4327);
or U4685 (N_4685,N_4236,N_4192);
nand U4686 (N_4686,N_4136,N_4062);
nor U4687 (N_4687,N_4221,N_4323);
and U4688 (N_4688,N_4427,N_4076);
and U4689 (N_4689,N_4418,N_4414);
nand U4690 (N_4690,N_4177,N_4145);
nor U4691 (N_4691,N_4003,N_4081);
and U4692 (N_4692,N_4437,N_4027);
or U4693 (N_4693,N_4255,N_4022);
nor U4694 (N_4694,N_4067,N_4118);
nand U4695 (N_4695,N_4059,N_4139);
nand U4696 (N_4696,N_4131,N_4029);
nor U4697 (N_4697,N_4193,N_4316);
and U4698 (N_4698,N_4403,N_4475);
nor U4699 (N_4699,N_4157,N_4367);
nand U4700 (N_4700,N_4384,N_4330);
or U4701 (N_4701,N_4413,N_4401);
nand U4702 (N_4702,N_4378,N_4322);
nor U4703 (N_4703,N_4481,N_4212);
nand U4704 (N_4704,N_4355,N_4196);
and U4705 (N_4705,N_4271,N_4147);
or U4706 (N_4706,N_4408,N_4094);
and U4707 (N_4707,N_4402,N_4137);
nand U4708 (N_4708,N_4072,N_4393);
or U4709 (N_4709,N_4049,N_4124);
nand U4710 (N_4710,N_4111,N_4007);
and U4711 (N_4711,N_4108,N_4484);
and U4712 (N_4712,N_4472,N_4441);
or U4713 (N_4713,N_4015,N_4064);
or U4714 (N_4714,N_4220,N_4213);
nand U4715 (N_4715,N_4141,N_4491);
nor U4716 (N_4716,N_4161,N_4013);
xnor U4717 (N_4717,N_4222,N_4254);
nand U4718 (N_4718,N_4204,N_4445);
nor U4719 (N_4719,N_4258,N_4209);
and U4720 (N_4720,N_4043,N_4487);
nor U4721 (N_4721,N_4140,N_4095);
and U4722 (N_4722,N_4298,N_4092);
and U4723 (N_4723,N_4004,N_4328);
nor U4724 (N_4724,N_4270,N_4267);
nor U4725 (N_4725,N_4133,N_4432);
nand U4726 (N_4726,N_4018,N_4296);
and U4727 (N_4727,N_4068,N_4123);
and U4728 (N_4728,N_4279,N_4480);
nand U4729 (N_4729,N_4143,N_4307);
and U4730 (N_4730,N_4349,N_4353);
nand U4731 (N_4731,N_4333,N_4230);
or U4732 (N_4732,N_4023,N_4376);
nand U4733 (N_4733,N_4063,N_4014);
and U4734 (N_4734,N_4382,N_4009);
nor U4735 (N_4735,N_4423,N_4356);
or U4736 (N_4736,N_4214,N_4198);
and U4737 (N_4737,N_4454,N_4365);
nand U4738 (N_4738,N_4476,N_4452);
nor U4739 (N_4739,N_4276,N_4369);
or U4740 (N_4740,N_4032,N_4051);
nor U4741 (N_4741,N_4471,N_4080);
and U4742 (N_4742,N_4091,N_4358);
and U4743 (N_4743,N_4042,N_4122);
nor U4744 (N_4744,N_4033,N_4260);
or U4745 (N_4745,N_4334,N_4499);
nand U4746 (N_4746,N_4048,N_4493);
and U4747 (N_4747,N_4388,N_4265);
nand U4748 (N_4748,N_4190,N_4162);
and U4749 (N_4749,N_4466,N_4089);
and U4750 (N_4750,N_4142,N_4353);
or U4751 (N_4751,N_4243,N_4213);
or U4752 (N_4752,N_4025,N_4386);
nor U4753 (N_4753,N_4399,N_4056);
or U4754 (N_4754,N_4154,N_4214);
and U4755 (N_4755,N_4046,N_4048);
and U4756 (N_4756,N_4331,N_4003);
and U4757 (N_4757,N_4166,N_4061);
nand U4758 (N_4758,N_4155,N_4495);
nand U4759 (N_4759,N_4117,N_4288);
nand U4760 (N_4760,N_4204,N_4184);
nand U4761 (N_4761,N_4469,N_4475);
nor U4762 (N_4762,N_4046,N_4030);
and U4763 (N_4763,N_4351,N_4427);
nor U4764 (N_4764,N_4195,N_4299);
or U4765 (N_4765,N_4162,N_4376);
and U4766 (N_4766,N_4361,N_4308);
nand U4767 (N_4767,N_4058,N_4325);
nor U4768 (N_4768,N_4339,N_4343);
and U4769 (N_4769,N_4264,N_4113);
or U4770 (N_4770,N_4479,N_4158);
or U4771 (N_4771,N_4498,N_4104);
nor U4772 (N_4772,N_4366,N_4125);
and U4773 (N_4773,N_4340,N_4456);
nor U4774 (N_4774,N_4116,N_4018);
nand U4775 (N_4775,N_4378,N_4215);
nor U4776 (N_4776,N_4219,N_4456);
nor U4777 (N_4777,N_4418,N_4072);
and U4778 (N_4778,N_4384,N_4218);
nand U4779 (N_4779,N_4447,N_4095);
nor U4780 (N_4780,N_4215,N_4050);
nand U4781 (N_4781,N_4094,N_4065);
and U4782 (N_4782,N_4437,N_4075);
and U4783 (N_4783,N_4084,N_4419);
and U4784 (N_4784,N_4212,N_4262);
xnor U4785 (N_4785,N_4172,N_4221);
nor U4786 (N_4786,N_4487,N_4411);
nor U4787 (N_4787,N_4085,N_4455);
nand U4788 (N_4788,N_4065,N_4284);
and U4789 (N_4789,N_4405,N_4302);
nor U4790 (N_4790,N_4452,N_4315);
nor U4791 (N_4791,N_4203,N_4366);
xnor U4792 (N_4792,N_4057,N_4006);
or U4793 (N_4793,N_4433,N_4364);
and U4794 (N_4794,N_4320,N_4268);
nand U4795 (N_4795,N_4195,N_4122);
nand U4796 (N_4796,N_4440,N_4125);
nand U4797 (N_4797,N_4336,N_4390);
nor U4798 (N_4798,N_4195,N_4436);
xor U4799 (N_4799,N_4032,N_4050);
and U4800 (N_4800,N_4325,N_4465);
or U4801 (N_4801,N_4110,N_4148);
nor U4802 (N_4802,N_4043,N_4311);
nor U4803 (N_4803,N_4057,N_4000);
and U4804 (N_4804,N_4138,N_4149);
and U4805 (N_4805,N_4005,N_4148);
nor U4806 (N_4806,N_4037,N_4119);
xnor U4807 (N_4807,N_4108,N_4401);
nand U4808 (N_4808,N_4202,N_4343);
nor U4809 (N_4809,N_4489,N_4119);
or U4810 (N_4810,N_4135,N_4193);
or U4811 (N_4811,N_4258,N_4057);
nor U4812 (N_4812,N_4215,N_4226);
and U4813 (N_4813,N_4251,N_4030);
or U4814 (N_4814,N_4187,N_4080);
and U4815 (N_4815,N_4352,N_4167);
or U4816 (N_4816,N_4292,N_4051);
nor U4817 (N_4817,N_4458,N_4159);
nor U4818 (N_4818,N_4188,N_4175);
or U4819 (N_4819,N_4494,N_4202);
or U4820 (N_4820,N_4217,N_4368);
nand U4821 (N_4821,N_4119,N_4159);
and U4822 (N_4822,N_4275,N_4193);
or U4823 (N_4823,N_4138,N_4104);
nand U4824 (N_4824,N_4126,N_4370);
nand U4825 (N_4825,N_4145,N_4403);
and U4826 (N_4826,N_4473,N_4089);
and U4827 (N_4827,N_4125,N_4263);
nand U4828 (N_4828,N_4473,N_4420);
nor U4829 (N_4829,N_4440,N_4092);
and U4830 (N_4830,N_4371,N_4488);
nor U4831 (N_4831,N_4307,N_4139);
nor U4832 (N_4832,N_4470,N_4238);
nand U4833 (N_4833,N_4016,N_4201);
and U4834 (N_4834,N_4131,N_4178);
nor U4835 (N_4835,N_4410,N_4432);
and U4836 (N_4836,N_4419,N_4476);
nand U4837 (N_4837,N_4087,N_4453);
or U4838 (N_4838,N_4310,N_4141);
or U4839 (N_4839,N_4194,N_4178);
nand U4840 (N_4840,N_4182,N_4440);
and U4841 (N_4841,N_4050,N_4289);
and U4842 (N_4842,N_4394,N_4350);
nand U4843 (N_4843,N_4451,N_4104);
nand U4844 (N_4844,N_4371,N_4199);
or U4845 (N_4845,N_4437,N_4233);
nor U4846 (N_4846,N_4490,N_4017);
nand U4847 (N_4847,N_4160,N_4212);
and U4848 (N_4848,N_4256,N_4466);
and U4849 (N_4849,N_4398,N_4266);
nor U4850 (N_4850,N_4440,N_4080);
nor U4851 (N_4851,N_4210,N_4064);
and U4852 (N_4852,N_4493,N_4465);
nor U4853 (N_4853,N_4056,N_4181);
and U4854 (N_4854,N_4387,N_4029);
and U4855 (N_4855,N_4349,N_4466);
or U4856 (N_4856,N_4438,N_4333);
nor U4857 (N_4857,N_4353,N_4157);
nor U4858 (N_4858,N_4169,N_4190);
nor U4859 (N_4859,N_4464,N_4332);
nand U4860 (N_4860,N_4057,N_4329);
and U4861 (N_4861,N_4060,N_4255);
and U4862 (N_4862,N_4073,N_4472);
nor U4863 (N_4863,N_4431,N_4498);
and U4864 (N_4864,N_4082,N_4370);
nand U4865 (N_4865,N_4274,N_4268);
nand U4866 (N_4866,N_4336,N_4029);
and U4867 (N_4867,N_4478,N_4258);
and U4868 (N_4868,N_4290,N_4124);
and U4869 (N_4869,N_4289,N_4334);
nand U4870 (N_4870,N_4264,N_4216);
nand U4871 (N_4871,N_4243,N_4048);
nor U4872 (N_4872,N_4029,N_4000);
xor U4873 (N_4873,N_4238,N_4274);
xnor U4874 (N_4874,N_4415,N_4200);
nand U4875 (N_4875,N_4350,N_4269);
or U4876 (N_4876,N_4208,N_4061);
or U4877 (N_4877,N_4114,N_4063);
nand U4878 (N_4878,N_4448,N_4288);
nor U4879 (N_4879,N_4172,N_4211);
or U4880 (N_4880,N_4053,N_4292);
nor U4881 (N_4881,N_4347,N_4362);
nand U4882 (N_4882,N_4080,N_4032);
nand U4883 (N_4883,N_4098,N_4053);
nor U4884 (N_4884,N_4378,N_4227);
or U4885 (N_4885,N_4371,N_4483);
and U4886 (N_4886,N_4308,N_4275);
nor U4887 (N_4887,N_4170,N_4124);
nor U4888 (N_4888,N_4121,N_4433);
nand U4889 (N_4889,N_4268,N_4391);
or U4890 (N_4890,N_4295,N_4166);
nand U4891 (N_4891,N_4445,N_4423);
or U4892 (N_4892,N_4041,N_4140);
nor U4893 (N_4893,N_4180,N_4092);
nor U4894 (N_4894,N_4467,N_4107);
nor U4895 (N_4895,N_4370,N_4101);
xnor U4896 (N_4896,N_4454,N_4045);
and U4897 (N_4897,N_4146,N_4475);
nand U4898 (N_4898,N_4182,N_4173);
nor U4899 (N_4899,N_4034,N_4119);
or U4900 (N_4900,N_4326,N_4036);
and U4901 (N_4901,N_4386,N_4194);
and U4902 (N_4902,N_4219,N_4481);
xor U4903 (N_4903,N_4120,N_4293);
or U4904 (N_4904,N_4119,N_4193);
nand U4905 (N_4905,N_4343,N_4407);
or U4906 (N_4906,N_4311,N_4298);
nand U4907 (N_4907,N_4321,N_4070);
or U4908 (N_4908,N_4292,N_4235);
nor U4909 (N_4909,N_4317,N_4299);
and U4910 (N_4910,N_4226,N_4308);
nor U4911 (N_4911,N_4331,N_4230);
nor U4912 (N_4912,N_4225,N_4239);
and U4913 (N_4913,N_4067,N_4222);
nor U4914 (N_4914,N_4418,N_4180);
nand U4915 (N_4915,N_4132,N_4042);
and U4916 (N_4916,N_4064,N_4296);
and U4917 (N_4917,N_4465,N_4175);
nand U4918 (N_4918,N_4026,N_4313);
or U4919 (N_4919,N_4196,N_4107);
or U4920 (N_4920,N_4335,N_4145);
nand U4921 (N_4921,N_4337,N_4078);
or U4922 (N_4922,N_4203,N_4217);
nor U4923 (N_4923,N_4253,N_4350);
nor U4924 (N_4924,N_4382,N_4272);
xor U4925 (N_4925,N_4448,N_4141);
or U4926 (N_4926,N_4340,N_4207);
nand U4927 (N_4927,N_4338,N_4386);
and U4928 (N_4928,N_4050,N_4400);
nand U4929 (N_4929,N_4092,N_4223);
or U4930 (N_4930,N_4442,N_4272);
nand U4931 (N_4931,N_4267,N_4343);
nand U4932 (N_4932,N_4195,N_4012);
or U4933 (N_4933,N_4360,N_4183);
and U4934 (N_4934,N_4387,N_4222);
and U4935 (N_4935,N_4453,N_4025);
and U4936 (N_4936,N_4313,N_4265);
nand U4937 (N_4937,N_4062,N_4361);
nor U4938 (N_4938,N_4008,N_4311);
or U4939 (N_4939,N_4065,N_4191);
nor U4940 (N_4940,N_4365,N_4088);
and U4941 (N_4941,N_4340,N_4357);
or U4942 (N_4942,N_4400,N_4363);
nor U4943 (N_4943,N_4439,N_4074);
or U4944 (N_4944,N_4263,N_4457);
nor U4945 (N_4945,N_4155,N_4489);
or U4946 (N_4946,N_4384,N_4314);
or U4947 (N_4947,N_4335,N_4184);
nand U4948 (N_4948,N_4171,N_4133);
nand U4949 (N_4949,N_4370,N_4178);
nor U4950 (N_4950,N_4003,N_4384);
nor U4951 (N_4951,N_4322,N_4470);
nor U4952 (N_4952,N_4290,N_4176);
nor U4953 (N_4953,N_4417,N_4394);
nor U4954 (N_4954,N_4132,N_4094);
or U4955 (N_4955,N_4120,N_4492);
nand U4956 (N_4956,N_4391,N_4366);
nand U4957 (N_4957,N_4292,N_4367);
and U4958 (N_4958,N_4320,N_4111);
or U4959 (N_4959,N_4226,N_4078);
xnor U4960 (N_4960,N_4260,N_4182);
and U4961 (N_4961,N_4459,N_4256);
or U4962 (N_4962,N_4329,N_4067);
nor U4963 (N_4963,N_4177,N_4199);
and U4964 (N_4964,N_4162,N_4497);
or U4965 (N_4965,N_4493,N_4372);
or U4966 (N_4966,N_4229,N_4081);
nand U4967 (N_4967,N_4048,N_4289);
and U4968 (N_4968,N_4052,N_4266);
and U4969 (N_4969,N_4202,N_4136);
and U4970 (N_4970,N_4179,N_4466);
and U4971 (N_4971,N_4494,N_4342);
and U4972 (N_4972,N_4205,N_4147);
and U4973 (N_4973,N_4492,N_4174);
nor U4974 (N_4974,N_4444,N_4197);
or U4975 (N_4975,N_4017,N_4459);
and U4976 (N_4976,N_4325,N_4232);
and U4977 (N_4977,N_4236,N_4260);
or U4978 (N_4978,N_4221,N_4134);
nor U4979 (N_4979,N_4140,N_4382);
nor U4980 (N_4980,N_4085,N_4383);
nor U4981 (N_4981,N_4393,N_4451);
and U4982 (N_4982,N_4089,N_4071);
nor U4983 (N_4983,N_4289,N_4045);
nor U4984 (N_4984,N_4439,N_4403);
or U4985 (N_4985,N_4304,N_4227);
and U4986 (N_4986,N_4184,N_4451);
nand U4987 (N_4987,N_4160,N_4029);
or U4988 (N_4988,N_4110,N_4396);
or U4989 (N_4989,N_4067,N_4163);
nand U4990 (N_4990,N_4234,N_4185);
or U4991 (N_4991,N_4023,N_4272);
nand U4992 (N_4992,N_4358,N_4274);
and U4993 (N_4993,N_4251,N_4151);
nand U4994 (N_4994,N_4027,N_4062);
or U4995 (N_4995,N_4321,N_4477);
nand U4996 (N_4996,N_4107,N_4410);
and U4997 (N_4997,N_4446,N_4276);
and U4998 (N_4998,N_4131,N_4321);
or U4999 (N_4999,N_4364,N_4006);
and U5000 (N_5000,N_4776,N_4647);
or U5001 (N_5001,N_4768,N_4556);
nor U5002 (N_5002,N_4989,N_4933);
and U5003 (N_5003,N_4701,N_4530);
nand U5004 (N_5004,N_4554,N_4801);
or U5005 (N_5005,N_4730,N_4631);
nor U5006 (N_5006,N_4905,N_4812);
nand U5007 (N_5007,N_4813,N_4802);
nand U5008 (N_5008,N_4599,N_4714);
nor U5009 (N_5009,N_4743,N_4996);
and U5010 (N_5010,N_4712,N_4513);
nor U5011 (N_5011,N_4962,N_4635);
nor U5012 (N_5012,N_4832,N_4693);
nand U5013 (N_5013,N_4843,N_4895);
or U5014 (N_5014,N_4940,N_4548);
nor U5015 (N_5015,N_4755,N_4660);
nand U5016 (N_5016,N_4613,N_4793);
nor U5017 (N_5017,N_4963,N_4952);
nor U5018 (N_5018,N_4600,N_4577);
nor U5019 (N_5019,N_4625,N_4935);
nand U5020 (N_5020,N_4509,N_4855);
and U5021 (N_5021,N_4686,N_4931);
nand U5022 (N_5022,N_4649,N_4956);
nor U5023 (N_5023,N_4610,N_4669);
nand U5024 (N_5024,N_4945,N_4856);
or U5025 (N_5025,N_4773,N_4850);
nand U5026 (N_5026,N_4917,N_4771);
or U5027 (N_5027,N_4946,N_4573);
nor U5028 (N_5028,N_4898,N_4708);
and U5029 (N_5029,N_4927,N_4572);
and U5030 (N_5030,N_4562,N_4545);
and U5031 (N_5031,N_4966,N_4503);
nand U5032 (N_5032,N_4919,N_4664);
or U5033 (N_5033,N_4950,N_4552);
or U5034 (N_5034,N_4980,N_4637);
and U5035 (N_5035,N_4522,N_4586);
and U5036 (N_5036,N_4512,N_4805);
nor U5037 (N_5037,N_4597,N_4506);
or U5038 (N_5038,N_4991,N_4590);
nand U5039 (N_5039,N_4544,N_4567);
or U5040 (N_5040,N_4844,N_4681);
nor U5041 (N_5041,N_4923,N_4883);
and U5042 (N_5042,N_4908,N_4783);
nand U5043 (N_5043,N_4827,N_4863);
or U5044 (N_5044,N_4523,N_4738);
nor U5045 (N_5045,N_4820,N_4520);
and U5046 (N_5046,N_4551,N_4742);
xor U5047 (N_5047,N_4864,N_4729);
nand U5048 (N_5048,N_4559,N_4619);
or U5049 (N_5049,N_4689,N_4973);
nor U5050 (N_5050,N_4723,N_4621);
and U5051 (N_5051,N_4673,N_4944);
and U5052 (N_5052,N_4876,N_4526);
nor U5053 (N_5053,N_4837,N_4711);
nor U5054 (N_5054,N_4588,N_4561);
nand U5055 (N_5055,N_4505,N_4648);
nand U5056 (N_5056,N_4624,N_4961);
nand U5057 (N_5057,N_4695,N_4872);
and U5058 (N_5058,N_4968,N_4779);
or U5059 (N_5059,N_4921,N_4748);
and U5060 (N_5060,N_4978,N_4675);
or U5061 (N_5061,N_4994,N_4926);
nand U5062 (N_5062,N_4728,N_4897);
nor U5063 (N_5063,N_4672,N_4605);
and U5064 (N_5064,N_4835,N_4854);
and U5065 (N_5065,N_4690,N_4964);
nand U5066 (N_5066,N_4774,N_4948);
nor U5067 (N_5067,N_4810,N_4767);
and U5068 (N_5068,N_4880,N_4787);
nor U5069 (N_5069,N_4869,N_4745);
nand U5070 (N_5070,N_4736,N_4951);
or U5071 (N_5071,N_4609,N_4724);
nand U5072 (N_5072,N_4899,N_4816);
and U5073 (N_5073,N_4868,N_4784);
nor U5074 (N_5074,N_4514,N_4758);
nand U5075 (N_5075,N_4725,N_4694);
nor U5076 (N_5076,N_4636,N_4700);
nand U5077 (N_5077,N_4502,N_4823);
nor U5078 (N_5078,N_4997,N_4715);
nor U5079 (N_5079,N_4985,N_4896);
and U5080 (N_5080,N_4853,N_4772);
nor U5081 (N_5081,N_4575,N_4953);
or U5082 (N_5082,N_4517,N_4798);
or U5083 (N_5083,N_4800,N_4670);
and U5084 (N_5084,N_4970,N_4587);
and U5085 (N_5085,N_4560,N_4873);
and U5086 (N_5086,N_4604,N_4778);
and U5087 (N_5087,N_4759,N_4751);
and U5088 (N_5088,N_4822,N_4914);
nor U5089 (N_5089,N_4763,N_4884);
or U5090 (N_5090,N_4665,N_4533);
nand U5091 (N_5091,N_4942,N_4756);
nor U5092 (N_5092,N_4703,N_4949);
nor U5093 (N_5093,N_4583,N_4829);
nand U5094 (N_5094,N_4537,N_4511);
nand U5095 (N_5095,N_4757,N_4982);
xnor U5096 (N_5096,N_4607,N_4571);
nor U5097 (N_5097,N_4593,N_4565);
nand U5098 (N_5098,N_4885,N_4570);
nor U5099 (N_5099,N_4930,N_4750);
and U5100 (N_5100,N_4815,N_4867);
nor U5101 (N_5101,N_4903,N_4925);
nor U5102 (N_5102,N_4857,N_4893);
nand U5103 (N_5103,N_4842,N_4764);
nor U5104 (N_5104,N_4529,N_4987);
or U5105 (N_5105,N_4814,N_4806);
or U5106 (N_5106,N_4795,N_4707);
or U5107 (N_5107,N_4706,N_4539);
xnor U5108 (N_5108,N_4910,N_4959);
nand U5109 (N_5109,N_4580,N_4702);
nand U5110 (N_5110,N_4983,N_4726);
nand U5111 (N_5111,N_4947,N_4840);
nor U5112 (N_5112,N_4770,N_4594);
nand U5113 (N_5113,N_4932,N_4993);
nand U5114 (N_5114,N_4941,N_4841);
and U5115 (N_5115,N_4866,N_4722);
and U5116 (N_5116,N_4639,N_4746);
nor U5117 (N_5117,N_4521,N_4938);
nand U5118 (N_5118,N_4769,N_4762);
nor U5119 (N_5119,N_4564,N_4633);
nor U5120 (N_5120,N_4965,N_4979);
nor U5121 (N_5121,N_4630,N_4591);
nand U5122 (N_5122,N_4734,N_4786);
or U5123 (N_5123,N_4906,N_4603);
nand U5124 (N_5124,N_4667,N_4662);
and U5125 (N_5125,N_4986,N_4501);
or U5126 (N_5126,N_4928,N_4620);
and U5127 (N_5127,N_4704,N_4626);
nor U5128 (N_5128,N_4555,N_4902);
nor U5129 (N_5129,N_4716,N_4821);
or U5130 (N_5130,N_4627,N_4638);
and U5131 (N_5131,N_4998,N_4538);
or U5132 (N_5132,N_4881,N_4984);
and U5133 (N_5133,N_4717,N_4671);
nand U5134 (N_5134,N_4849,N_4612);
nor U5135 (N_5135,N_4628,N_4737);
or U5136 (N_5136,N_4553,N_4687);
nand U5137 (N_5137,N_4592,N_4792);
or U5138 (N_5138,N_4804,N_4532);
and U5139 (N_5139,N_4696,N_4870);
nor U5140 (N_5140,N_4744,N_4568);
nand U5141 (N_5141,N_4657,N_4830);
nand U5142 (N_5142,N_4534,N_4888);
nand U5143 (N_5143,N_4516,N_4611);
or U5144 (N_5144,N_4524,N_4710);
nand U5145 (N_5145,N_4641,N_4871);
nor U5146 (N_5146,N_4918,N_4542);
nor U5147 (N_5147,N_4684,N_4692);
nand U5148 (N_5148,N_4713,N_4799);
or U5149 (N_5149,N_4601,N_4833);
and U5150 (N_5150,N_4861,N_4536);
or U5151 (N_5151,N_4622,N_4981);
and U5152 (N_5152,N_4992,N_4691);
nand U5153 (N_5153,N_4683,N_4907);
and U5154 (N_5154,N_4685,N_4582);
xor U5155 (N_5155,N_4652,N_4845);
or U5156 (N_5156,N_4990,N_4878);
or U5157 (N_5157,N_4765,N_4937);
and U5158 (N_5158,N_4589,N_4803);
nand U5159 (N_5159,N_4988,N_4541);
and U5160 (N_5160,N_4705,N_4677);
nor U5161 (N_5161,N_4741,N_4939);
or U5162 (N_5162,N_4824,N_4975);
nor U5163 (N_5163,N_4519,N_4645);
and U5164 (N_5164,N_4646,N_4608);
nor U5165 (N_5165,N_4865,N_4678);
and U5166 (N_5166,N_4826,N_4550);
nand U5167 (N_5167,N_4818,N_4886);
and U5168 (N_5168,N_4617,N_4790);
nor U5169 (N_5169,N_4680,N_4658);
nand U5170 (N_5170,N_4596,N_4807);
nor U5171 (N_5171,N_4894,N_4666);
or U5172 (N_5172,N_4976,N_4915);
nand U5173 (N_5173,N_4882,N_4525);
nor U5174 (N_5174,N_4659,N_4782);
nor U5175 (N_5175,N_4775,N_4528);
or U5176 (N_5176,N_4859,N_4848);
nor U5177 (N_5177,N_4507,N_4650);
nor U5178 (N_5178,N_4819,N_4916);
nor U5179 (N_5179,N_4890,N_4967);
and U5180 (N_5180,N_4727,N_4875);
and U5181 (N_5181,N_4922,N_4834);
or U5182 (N_5182,N_4569,N_4578);
or U5183 (N_5183,N_4995,N_4817);
nand U5184 (N_5184,N_4581,N_4825);
nor U5185 (N_5185,N_4828,N_4504);
nand U5186 (N_5186,N_4543,N_4754);
or U5187 (N_5187,N_4732,N_4720);
or U5188 (N_5188,N_4508,N_4563);
nor U5189 (N_5189,N_4796,N_4540);
nand U5190 (N_5190,N_4766,N_4892);
nor U5191 (N_5191,N_4574,N_4999);
xnor U5192 (N_5192,N_4558,N_4761);
and U5193 (N_5193,N_4808,N_4547);
xor U5194 (N_5194,N_4960,N_4661);
and U5195 (N_5195,N_4788,N_4598);
or U5196 (N_5196,N_4719,N_4954);
nand U5197 (N_5197,N_4860,N_4642);
nand U5198 (N_5198,N_4913,N_4891);
and U5199 (N_5199,N_4955,N_4616);
nor U5200 (N_5200,N_4527,N_4618);
nor U5201 (N_5201,N_4518,N_4839);
nand U5202 (N_5202,N_4629,N_4780);
and U5203 (N_5203,N_4760,N_4740);
nand U5204 (N_5204,N_4858,N_4697);
nor U5205 (N_5205,N_4531,N_4797);
and U5206 (N_5206,N_4655,N_4957);
and U5207 (N_5207,N_4585,N_4643);
or U5208 (N_5208,N_4924,N_4709);
nor U5209 (N_5209,N_4653,N_4668);
nor U5210 (N_5210,N_4676,N_4634);
or U5211 (N_5211,N_4656,N_4912);
nand U5212 (N_5212,N_4874,N_4615);
nand U5213 (N_5213,N_4887,N_4749);
and U5214 (N_5214,N_4557,N_4934);
nor U5215 (N_5215,N_4889,N_4500);
and U5216 (N_5216,N_4851,N_4971);
nand U5217 (N_5217,N_4515,N_4674);
or U5218 (N_5218,N_4958,N_4654);
nand U5219 (N_5219,N_4846,N_4752);
or U5220 (N_5220,N_4735,N_4972);
nand U5221 (N_5221,N_4640,N_4623);
or U5222 (N_5222,N_4584,N_4809);
or U5223 (N_5223,N_4721,N_4943);
or U5224 (N_5224,N_4974,N_4566);
or U5225 (N_5225,N_4901,N_4977);
nor U5226 (N_5226,N_4785,N_4510);
and U5227 (N_5227,N_4753,N_4632);
and U5228 (N_5228,N_4688,N_4739);
nand U5229 (N_5229,N_4811,N_4836);
or U5230 (N_5230,N_4847,N_4879);
nand U5231 (N_5231,N_4733,N_4602);
nor U5232 (N_5232,N_4606,N_4852);
nor U5233 (N_5233,N_4679,N_4576);
nand U5234 (N_5234,N_4663,N_4699);
xor U5235 (N_5235,N_4731,N_4920);
nand U5236 (N_5236,N_4791,N_4789);
and U5237 (N_5237,N_4781,N_4777);
or U5238 (N_5238,N_4535,N_4877);
and U5239 (N_5239,N_4698,N_4595);
and U5240 (N_5240,N_4718,N_4838);
xor U5241 (N_5241,N_4900,N_4909);
nand U5242 (N_5242,N_4614,N_4862);
and U5243 (N_5243,N_4549,N_4969);
and U5244 (N_5244,N_4747,N_4682);
and U5245 (N_5245,N_4651,N_4794);
nand U5246 (N_5246,N_4904,N_4929);
nor U5247 (N_5247,N_4936,N_4546);
and U5248 (N_5248,N_4831,N_4911);
nor U5249 (N_5249,N_4579,N_4644);
or U5250 (N_5250,N_4885,N_4909);
and U5251 (N_5251,N_4680,N_4577);
or U5252 (N_5252,N_4826,N_4822);
nand U5253 (N_5253,N_4827,N_4572);
and U5254 (N_5254,N_4783,N_4760);
xnor U5255 (N_5255,N_4732,N_4622);
nand U5256 (N_5256,N_4758,N_4701);
nand U5257 (N_5257,N_4722,N_4806);
and U5258 (N_5258,N_4779,N_4757);
and U5259 (N_5259,N_4925,N_4872);
nand U5260 (N_5260,N_4728,N_4962);
nor U5261 (N_5261,N_4912,N_4545);
and U5262 (N_5262,N_4926,N_4573);
nand U5263 (N_5263,N_4980,N_4627);
or U5264 (N_5264,N_4766,N_4751);
and U5265 (N_5265,N_4885,N_4705);
nor U5266 (N_5266,N_4695,N_4609);
and U5267 (N_5267,N_4645,N_4644);
and U5268 (N_5268,N_4610,N_4866);
nand U5269 (N_5269,N_4693,N_4819);
and U5270 (N_5270,N_4539,N_4799);
nand U5271 (N_5271,N_4641,N_4674);
nand U5272 (N_5272,N_4665,N_4837);
nor U5273 (N_5273,N_4900,N_4870);
or U5274 (N_5274,N_4592,N_4794);
and U5275 (N_5275,N_4726,N_4678);
xnor U5276 (N_5276,N_4646,N_4828);
and U5277 (N_5277,N_4808,N_4868);
or U5278 (N_5278,N_4515,N_4576);
or U5279 (N_5279,N_4529,N_4922);
nor U5280 (N_5280,N_4978,N_4548);
nand U5281 (N_5281,N_4850,N_4663);
nand U5282 (N_5282,N_4509,N_4767);
nand U5283 (N_5283,N_4746,N_4992);
and U5284 (N_5284,N_4682,N_4795);
or U5285 (N_5285,N_4569,N_4594);
and U5286 (N_5286,N_4846,N_4501);
and U5287 (N_5287,N_4903,N_4860);
and U5288 (N_5288,N_4508,N_4719);
or U5289 (N_5289,N_4894,N_4861);
nand U5290 (N_5290,N_4762,N_4826);
and U5291 (N_5291,N_4774,N_4561);
nand U5292 (N_5292,N_4810,N_4551);
or U5293 (N_5293,N_4596,N_4729);
or U5294 (N_5294,N_4923,N_4569);
nor U5295 (N_5295,N_4688,N_4549);
and U5296 (N_5296,N_4700,N_4515);
nand U5297 (N_5297,N_4797,N_4882);
or U5298 (N_5298,N_4661,N_4570);
nor U5299 (N_5299,N_4838,N_4710);
and U5300 (N_5300,N_4994,N_4801);
or U5301 (N_5301,N_4830,N_4855);
and U5302 (N_5302,N_4549,N_4912);
nand U5303 (N_5303,N_4764,N_4682);
or U5304 (N_5304,N_4899,N_4834);
nor U5305 (N_5305,N_4794,N_4685);
nor U5306 (N_5306,N_4764,N_4707);
and U5307 (N_5307,N_4932,N_4662);
and U5308 (N_5308,N_4813,N_4868);
xnor U5309 (N_5309,N_4556,N_4789);
and U5310 (N_5310,N_4809,N_4794);
nand U5311 (N_5311,N_4725,N_4885);
nor U5312 (N_5312,N_4718,N_4530);
xor U5313 (N_5313,N_4638,N_4789);
or U5314 (N_5314,N_4748,N_4938);
nand U5315 (N_5315,N_4945,N_4919);
nand U5316 (N_5316,N_4994,N_4667);
and U5317 (N_5317,N_4751,N_4779);
nor U5318 (N_5318,N_4629,N_4585);
nand U5319 (N_5319,N_4674,N_4730);
or U5320 (N_5320,N_4906,N_4752);
xnor U5321 (N_5321,N_4888,N_4662);
nand U5322 (N_5322,N_4874,N_4553);
nor U5323 (N_5323,N_4971,N_4543);
and U5324 (N_5324,N_4839,N_4834);
and U5325 (N_5325,N_4557,N_4723);
nand U5326 (N_5326,N_4896,N_4786);
and U5327 (N_5327,N_4813,N_4971);
nor U5328 (N_5328,N_4952,N_4617);
and U5329 (N_5329,N_4565,N_4641);
or U5330 (N_5330,N_4985,N_4884);
nor U5331 (N_5331,N_4736,N_4827);
or U5332 (N_5332,N_4797,N_4866);
nand U5333 (N_5333,N_4783,N_4649);
and U5334 (N_5334,N_4613,N_4775);
nand U5335 (N_5335,N_4568,N_4955);
and U5336 (N_5336,N_4828,N_4812);
nand U5337 (N_5337,N_4904,N_4687);
nor U5338 (N_5338,N_4917,N_4809);
nor U5339 (N_5339,N_4827,N_4883);
and U5340 (N_5340,N_4996,N_4579);
or U5341 (N_5341,N_4650,N_4596);
nor U5342 (N_5342,N_4711,N_4609);
nor U5343 (N_5343,N_4697,N_4805);
and U5344 (N_5344,N_4621,N_4763);
nor U5345 (N_5345,N_4964,N_4536);
nand U5346 (N_5346,N_4525,N_4604);
nor U5347 (N_5347,N_4613,N_4688);
nor U5348 (N_5348,N_4741,N_4931);
or U5349 (N_5349,N_4685,N_4649);
nand U5350 (N_5350,N_4725,N_4974);
and U5351 (N_5351,N_4525,N_4712);
and U5352 (N_5352,N_4965,N_4572);
nand U5353 (N_5353,N_4914,N_4579);
nor U5354 (N_5354,N_4652,N_4928);
and U5355 (N_5355,N_4919,N_4509);
nand U5356 (N_5356,N_4558,N_4511);
nor U5357 (N_5357,N_4918,N_4683);
and U5358 (N_5358,N_4801,N_4544);
nor U5359 (N_5359,N_4566,N_4970);
and U5360 (N_5360,N_4652,N_4997);
or U5361 (N_5361,N_4656,N_4771);
or U5362 (N_5362,N_4581,N_4551);
nand U5363 (N_5363,N_4788,N_4698);
and U5364 (N_5364,N_4876,N_4625);
or U5365 (N_5365,N_4556,N_4982);
or U5366 (N_5366,N_4929,N_4743);
nand U5367 (N_5367,N_4691,N_4598);
nor U5368 (N_5368,N_4661,N_4617);
nor U5369 (N_5369,N_4651,N_4821);
or U5370 (N_5370,N_4583,N_4861);
nor U5371 (N_5371,N_4850,N_4935);
or U5372 (N_5372,N_4739,N_4568);
or U5373 (N_5373,N_4572,N_4701);
or U5374 (N_5374,N_4677,N_4770);
or U5375 (N_5375,N_4515,N_4920);
nand U5376 (N_5376,N_4518,N_4975);
or U5377 (N_5377,N_4987,N_4514);
and U5378 (N_5378,N_4722,N_4904);
or U5379 (N_5379,N_4842,N_4981);
or U5380 (N_5380,N_4593,N_4675);
nor U5381 (N_5381,N_4707,N_4660);
or U5382 (N_5382,N_4866,N_4971);
or U5383 (N_5383,N_4993,N_4546);
and U5384 (N_5384,N_4539,N_4962);
nand U5385 (N_5385,N_4876,N_4930);
or U5386 (N_5386,N_4694,N_4965);
nand U5387 (N_5387,N_4856,N_4984);
nand U5388 (N_5388,N_4737,N_4782);
and U5389 (N_5389,N_4561,N_4981);
or U5390 (N_5390,N_4677,N_4869);
nor U5391 (N_5391,N_4820,N_4929);
nor U5392 (N_5392,N_4523,N_4610);
and U5393 (N_5393,N_4856,N_4610);
nor U5394 (N_5394,N_4687,N_4616);
or U5395 (N_5395,N_4705,N_4840);
nand U5396 (N_5396,N_4816,N_4975);
and U5397 (N_5397,N_4875,N_4634);
and U5398 (N_5398,N_4520,N_4757);
nor U5399 (N_5399,N_4598,N_4789);
nor U5400 (N_5400,N_4856,N_4546);
nand U5401 (N_5401,N_4732,N_4857);
and U5402 (N_5402,N_4804,N_4958);
or U5403 (N_5403,N_4504,N_4526);
and U5404 (N_5404,N_4540,N_4991);
and U5405 (N_5405,N_4700,N_4605);
nand U5406 (N_5406,N_4652,N_4770);
and U5407 (N_5407,N_4530,N_4870);
and U5408 (N_5408,N_4842,N_4812);
nor U5409 (N_5409,N_4570,N_4925);
or U5410 (N_5410,N_4903,N_4916);
xnor U5411 (N_5411,N_4963,N_4994);
nor U5412 (N_5412,N_4710,N_4531);
nand U5413 (N_5413,N_4541,N_4805);
nand U5414 (N_5414,N_4607,N_4922);
and U5415 (N_5415,N_4675,N_4689);
xnor U5416 (N_5416,N_4703,N_4625);
or U5417 (N_5417,N_4804,N_4783);
nand U5418 (N_5418,N_4844,N_4732);
nand U5419 (N_5419,N_4516,N_4522);
nand U5420 (N_5420,N_4820,N_4585);
nor U5421 (N_5421,N_4820,N_4632);
and U5422 (N_5422,N_4791,N_4768);
and U5423 (N_5423,N_4592,N_4572);
and U5424 (N_5424,N_4872,N_4792);
nor U5425 (N_5425,N_4776,N_4808);
or U5426 (N_5426,N_4664,N_4680);
or U5427 (N_5427,N_4516,N_4614);
nand U5428 (N_5428,N_4757,N_4501);
nand U5429 (N_5429,N_4542,N_4893);
and U5430 (N_5430,N_4870,N_4504);
nor U5431 (N_5431,N_4589,N_4727);
nand U5432 (N_5432,N_4705,N_4860);
or U5433 (N_5433,N_4541,N_4689);
nand U5434 (N_5434,N_4953,N_4994);
and U5435 (N_5435,N_4799,N_4591);
and U5436 (N_5436,N_4833,N_4750);
nor U5437 (N_5437,N_4826,N_4515);
nand U5438 (N_5438,N_4579,N_4731);
and U5439 (N_5439,N_4995,N_4568);
nor U5440 (N_5440,N_4554,N_4946);
and U5441 (N_5441,N_4699,N_4615);
nor U5442 (N_5442,N_4880,N_4945);
and U5443 (N_5443,N_4939,N_4936);
and U5444 (N_5444,N_4566,N_4780);
xor U5445 (N_5445,N_4617,N_4546);
nor U5446 (N_5446,N_4559,N_4591);
nand U5447 (N_5447,N_4987,N_4773);
nand U5448 (N_5448,N_4750,N_4998);
or U5449 (N_5449,N_4688,N_4606);
and U5450 (N_5450,N_4970,N_4599);
and U5451 (N_5451,N_4789,N_4591);
nand U5452 (N_5452,N_4996,N_4758);
nand U5453 (N_5453,N_4889,N_4712);
nand U5454 (N_5454,N_4701,N_4712);
nand U5455 (N_5455,N_4867,N_4696);
or U5456 (N_5456,N_4771,N_4880);
nand U5457 (N_5457,N_4791,N_4578);
and U5458 (N_5458,N_4933,N_4922);
nor U5459 (N_5459,N_4523,N_4558);
and U5460 (N_5460,N_4721,N_4929);
or U5461 (N_5461,N_4958,N_4886);
nor U5462 (N_5462,N_4778,N_4618);
and U5463 (N_5463,N_4833,N_4692);
and U5464 (N_5464,N_4763,N_4578);
xnor U5465 (N_5465,N_4696,N_4888);
nand U5466 (N_5466,N_4830,N_4975);
or U5467 (N_5467,N_4836,N_4977);
and U5468 (N_5468,N_4706,N_4553);
nor U5469 (N_5469,N_4656,N_4652);
or U5470 (N_5470,N_4723,N_4661);
nor U5471 (N_5471,N_4561,N_4733);
nor U5472 (N_5472,N_4968,N_4590);
nand U5473 (N_5473,N_4732,N_4680);
or U5474 (N_5474,N_4660,N_4811);
nand U5475 (N_5475,N_4596,N_4713);
and U5476 (N_5476,N_4878,N_4964);
and U5477 (N_5477,N_4952,N_4857);
nor U5478 (N_5478,N_4986,N_4556);
or U5479 (N_5479,N_4793,N_4541);
or U5480 (N_5480,N_4593,N_4782);
and U5481 (N_5481,N_4710,N_4658);
and U5482 (N_5482,N_4693,N_4521);
and U5483 (N_5483,N_4916,N_4533);
or U5484 (N_5484,N_4629,N_4962);
and U5485 (N_5485,N_4753,N_4942);
nand U5486 (N_5486,N_4704,N_4503);
nor U5487 (N_5487,N_4920,N_4914);
and U5488 (N_5488,N_4765,N_4518);
or U5489 (N_5489,N_4611,N_4990);
nor U5490 (N_5490,N_4727,N_4785);
or U5491 (N_5491,N_4767,N_4502);
nor U5492 (N_5492,N_4945,N_4607);
nor U5493 (N_5493,N_4761,N_4500);
nand U5494 (N_5494,N_4703,N_4917);
and U5495 (N_5495,N_4501,N_4839);
and U5496 (N_5496,N_4527,N_4703);
and U5497 (N_5497,N_4920,N_4585);
nor U5498 (N_5498,N_4748,N_4529);
and U5499 (N_5499,N_4827,N_4855);
or U5500 (N_5500,N_5335,N_5208);
and U5501 (N_5501,N_5243,N_5440);
nand U5502 (N_5502,N_5284,N_5028);
xnor U5503 (N_5503,N_5390,N_5266);
and U5504 (N_5504,N_5364,N_5141);
or U5505 (N_5505,N_5238,N_5255);
nor U5506 (N_5506,N_5279,N_5408);
or U5507 (N_5507,N_5047,N_5189);
and U5508 (N_5508,N_5110,N_5326);
and U5509 (N_5509,N_5478,N_5239);
or U5510 (N_5510,N_5039,N_5345);
or U5511 (N_5511,N_5191,N_5058);
nand U5512 (N_5512,N_5249,N_5270);
and U5513 (N_5513,N_5483,N_5392);
nand U5514 (N_5514,N_5436,N_5056);
nor U5515 (N_5515,N_5385,N_5464);
and U5516 (N_5516,N_5104,N_5035);
nand U5517 (N_5517,N_5252,N_5269);
nor U5518 (N_5518,N_5219,N_5133);
and U5519 (N_5519,N_5205,N_5146);
nor U5520 (N_5520,N_5148,N_5451);
or U5521 (N_5521,N_5014,N_5293);
or U5522 (N_5522,N_5052,N_5407);
and U5523 (N_5523,N_5168,N_5202);
nor U5524 (N_5524,N_5383,N_5418);
and U5525 (N_5525,N_5493,N_5099);
nand U5526 (N_5526,N_5494,N_5457);
and U5527 (N_5527,N_5150,N_5227);
and U5528 (N_5528,N_5458,N_5049);
nor U5529 (N_5529,N_5416,N_5441);
nor U5530 (N_5530,N_5334,N_5231);
and U5531 (N_5531,N_5190,N_5404);
nand U5532 (N_5532,N_5161,N_5072);
nor U5533 (N_5533,N_5403,N_5155);
and U5534 (N_5534,N_5077,N_5406);
or U5535 (N_5535,N_5375,N_5445);
and U5536 (N_5536,N_5057,N_5398);
nand U5537 (N_5537,N_5342,N_5267);
nor U5538 (N_5538,N_5315,N_5097);
and U5539 (N_5539,N_5420,N_5157);
nand U5540 (N_5540,N_5484,N_5263);
and U5541 (N_5541,N_5068,N_5051);
and U5542 (N_5542,N_5366,N_5106);
nand U5543 (N_5543,N_5329,N_5031);
nand U5544 (N_5544,N_5181,N_5154);
or U5545 (N_5545,N_5145,N_5129);
nand U5546 (N_5546,N_5027,N_5112);
nor U5547 (N_5547,N_5492,N_5302);
nand U5548 (N_5548,N_5369,N_5461);
nor U5549 (N_5549,N_5357,N_5071);
nor U5550 (N_5550,N_5401,N_5044);
and U5551 (N_5551,N_5429,N_5025);
nand U5552 (N_5552,N_5405,N_5169);
nand U5553 (N_5553,N_5410,N_5163);
nand U5554 (N_5554,N_5138,N_5182);
and U5555 (N_5555,N_5036,N_5176);
or U5556 (N_5556,N_5479,N_5069);
nor U5557 (N_5557,N_5391,N_5498);
and U5558 (N_5558,N_5113,N_5034);
or U5559 (N_5559,N_5365,N_5199);
nand U5560 (N_5560,N_5234,N_5328);
or U5561 (N_5561,N_5108,N_5074);
xor U5562 (N_5562,N_5477,N_5188);
and U5563 (N_5563,N_5003,N_5124);
nor U5564 (N_5564,N_5229,N_5272);
or U5565 (N_5565,N_5032,N_5339);
or U5566 (N_5566,N_5307,N_5233);
nand U5567 (N_5567,N_5175,N_5485);
or U5568 (N_5568,N_5230,N_5119);
nand U5569 (N_5569,N_5139,N_5236);
nand U5570 (N_5570,N_5367,N_5096);
or U5571 (N_5571,N_5258,N_5187);
xor U5572 (N_5572,N_5241,N_5368);
or U5573 (N_5573,N_5331,N_5394);
or U5574 (N_5574,N_5497,N_5164);
and U5575 (N_5575,N_5135,N_5281);
or U5576 (N_5576,N_5434,N_5237);
nand U5577 (N_5577,N_5082,N_5374);
and U5578 (N_5578,N_5442,N_5016);
or U5579 (N_5579,N_5256,N_5211);
nand U5580 (N_5580,N_5240,N_5377);
or U5581 (N_5581,N_5271,N_5105);
nand U5582 (N_5582,N_5118,N_5005);
nor U5583 (N_5583,N_5421,N_5314);
nor U5584 (N_5584,N_5424,N_5147);
nor U5585 (N_5585,N_5162,N_5423);
nand U5586 (N_5586,N_5446,N_5431);
nand U5587 (N_5587,N_5073,N_5257);
or U5588 (N_5588,N_5012,N_5120);
nor U5589 (N_5589,N_5221,N_5319);
nand U5590 (N_5590,N_5359,N_5309);
or U5591 (N_5591,N_5166,N_5042);
xnor U5592 (N_5592,N_5471,N_5428);
nor U5593 (N_5593,N_5303,N_5397);
nand U5594 (N_5594,N_5358,N_5278);
nor U5595 (N_5595,N_5210,N_5131);
or U5596 (N_5596,N_5304,N_5351);
and U5597 (N_5597,N_5393,N_5316);
or U5598 (N_5598,N_5389,N_5473);
nor U5599 (N_5599,N_5323,N_5443);
nand U5600 (N_5600,N_5001,N_5282);
and U5601 (N_5601,N_5276,N_5399);
or U5602 (N_5602,N_5149,N_5064);
or U5603 (N_5603,N_5246,N_5450);
nand U5604 (N_5604,N_5348,N_5223);
and U5605 (N_5605,N_5158,N_5286);
nand U5606 (N_5606,N_5180,N_5062);
or U5607 (N_5607,N_5079,N_5280);
nand U5608 (N_5608,N_5136,N_5207);
and U5609 (N_5609,N_5165,N_5144);
or U5610 (N_5610,N_5381,N_5109);
nand U5611 (N_5611,N_5087,N_5121);
or U5612 (N_5612,N_5004,N_5432);
and U5613 (N_5613,N_5006,N_5475);
and U5614 (N_5614,N_5178,N_5310);
and U5615 (N_5615,N_5444,N_5117);
nor U5616 (N_5616,N_5045,N_5026);
and U5617 (N_5617,N_5482,N_5462);
nor U5618 (N_5618,N_5115,N_5107);
nand U5619 (N_5619,N_5346,N_5201);
nor U5620 (N_5620,N_5260,N_5480);
and U5621 (N_5621,N_5371,N_5018);
or U5622 (N_5622,N_5156,N_5123);
nand U5623 (N_5623,N_5100,N_5373);
or U5624 (N_5624,N_5499,N_5320);
xor U5625 (N_5625,N_5192,N_5127);
nand U5626 (N_5626,N_5384,N_5350);
nor U5627 (N_5627,N_5296,N_5220);
and U5628 (N_5628,N_5324,N_5417);
or U5629 (N_5629,N_5037,N_5299);
and U5630 (N_5630,N_5002,N_5274);
nand U5631 (N_5631,N_5453,N_5140);
nor U5632 (N_5632,N_5142,N_5327);
and U5633 (N_5633,N_5301,N_5376);
nand U5634 (N_5634,N_5019,N_5490);
and U5635 (N_5635,N_5332,N_5321);
or U5636 (N_5636,N_5218,N_5151);
and U5637 (N_5637,N_5217,N_5292);
and U5638 (N_5638,N_5290,N_5489);
nand U5639 (N_5639,N_5206,N_5195);
nor U5640 (N_5640,N_5197,N_5455);
or U5641 (N_5641,N_5395,N_5402);
nor U5642 (N_5642,N_5491,N_5128);
and U5643 (N_5643,N_5360,N_5288);
xor U5644 (N_5644,N_5244,N_5179);
nand U5645 (N_5645,N_5022,N_5352);
nor U5646 (N_5646,N_5386,N_5215);
and U5647 (N_5647,N_5040,N_5305);
and U5648 (N_5648,N_5287,N_5065);
nor U5649 (N_5649,N_5409,N_5093);
or U5650 (N_5650,N_5103,N_5043);
xor U5651 (N_5651,N_5167,N_5264);
nand U5652 (N_5652,N_5452,N_5275);
nor U5653 (N_5653,N_5033,N_5038);
and U5654 (N_5654,N_5295,N_5224);
and U5655 (N_5655,N_5426,N_5070);
xor U5656 (N_5656,N_5170,N_5363);
nor U5657 (N_5657,N_5160,N_5092);
or U5658 (N_5658,N_5472,N_5094);
and U5659 (N_5659,N_5060,N_5122);
nand U5660 (N_5660,N_5228,N_5134);
or U5661 (N_5661,N_5474,N_5300);
nor U5662 (N_5662,N_5011,N_5198);
nor U5663 (N_5663,N_5277,N_5048);
and U5664 (N_5664,N_5046,N_5388);
and U5665 (N_5665,N_5496,N_5268);
nor U5666 (N_5666,N_5468,N_5355);
nor U5667 (N_5667,N_5213,N_5341);
nor U5668 (N_5668,N_5285,N_5333);
nand U5669 (N_5669,N_5362,N_5379);
or U5670 (N_5670,N_5439,N_5283);
and U5671 (N_5671,N_5460,N_5469);
and U5672 (N_5672,N_5289,N_5415);
nor U5673 (N_5673,N_5495,N_5447);
and U5674 (N_5674,N_5265,N_5061);
nor U5675 (N_5675,N_5171,N_5214);
nor U5676 (N_5676,N_5422,N_5343);
xor U5677 (N_5677,N_5382,N_5313);
nand U5678 (N_5678,N_5130,N_5294);
nand U5679 (N_5679,N_5467,N_5259);
or U5680 (N_5680,N_5425,N_5159);
nand U5681 (N_5681,N_5338,N_5209);
xnor U5682 (N_5682,N_5029,N_5063);
xor U5683 (N_5683,N_5194,N_5095);
nand U5684 (N_5684,N_5486,N_5463);
or U5685 (N_5685,N_5449,N_5349);
nor U5686 (N_5686,N_5261,N_5347);
or U5687 (N_5687,N_5080,N_5245);
nand U5688 (N_5688,N_5091,N_5419);
nor U5689 (N_5689,N_5330,N_5396);
or U5690 (N_5690,N_5322,N_5183);
nor U5691 (N_5691,N_5273,N_5476);
nor U5692 (N_5692,N_5050,N_5066);
or U5693 (N_5693,N_5318,N_5344);
nor U5694 (N_5694,N_5325,N_5116);
or U5695 (N_5695,N_5454,N_5200);
or U5696 (N_5696,N_5174,N_5184);
nand U5697 (N_5697,N_5111,N_5488);
and U5698 (N_5698,N_5262,N_5152);
nor U5699 (N_5699,N_5185,N_5435);
nor U5700 (N_5700,N_5084,N_5186);
and U5701 (N_5701,N_5248,N_5081);
or U5702 (N_5702,N_5448,N_5204);
nand U5703 (N_5703,N_5015,N_5470);
and U5704 (N_5704,N_5177,N_5427);
nand U5705 (N_5705,N_5437,N_5212);
nand U5706 (N_5706,N_5308,N_5253);
or U5707 (N_5707,N_5235,N_5083);
and U5708 (N_5708,N_5009,N_5317);
nand U5709 (N_5709,N_5378,N_5076);
nand U5710 (N_5710,N_5078,N_5222);
and U5711 (N_5711,N_5053,N_5137);
or U5712 (N_5712,N_5242,N_5020);
xnor U5713 (N_5713,N_5125,N_5013);
and U5714 (N_5714,N_5456,N_5126);
and U5715 (N_5715,N_5132,N_5172);
or U5716 (N_5716,N_5090,N_5387);
or U5717 (N_5717,N_5054,N_5430);
nand U5718 (N_5718,N_5143,N_5250);
nor U5719 (N_5719,N_5251,N_5459);
nand U5720 (N_5720,N_5312,N_5413);
or U5721 (N_5721,N_5088,N_5021);
and U5722 (N_5722,N_5306,N_5173);
or U5723 (N_5723,N_5196,N_5153);
or U5724 (N_5724,N_5247,N_5411);
nor U5725 (N_5725,N_5007,N_5412);
or U5726 (N_5726,N_5232,N_5370);
nand U5727 (N_5727,N_5023,N_5361);
and U5728 (N_5728,N_5008,N_5203);
nor U5729 (N_5729,N_5067,N_5059);
nor U5730 (N_5730,N_5400,N_5098);
or U5731 (N_5731,N_5010,N_5075);
or U5732 (N_5732,N_5433,N_5225);
nor U5733 (N_5733,N_5380,N_5337);
and U5734 (N_5734,N_5353,N_5226);
nand U5735 (N_5735,N_5297,N_5000);
nand U5736 (N_5736,N_5216,N_5193);
and U5737 (N_5737,N_5336,N_5372);
nor U5738 (N_5738,N_5085,N_5291);
nor U5739 (N_5739,N_5298,N_5101);
nor U5740 (N_5740,N_5089,N_5340);
nor U5741 (N_5741,N_5466,N_5354);
and U5742 (N_5742,N_5024,N_5041);
nand U5743 (N_5743,N_5114,N_5086);
nand U5744 (N_5744,N_5030,N_5102);
nand U5745 (N_5745,N_5356,N_5055);
and U5746 (N_5746,N_5311,N_5254);
nor U5747 (N_5747,N_5438,N_5414);
or U5748 (N_5748,N_5465,N_5481);
or U5749 (N_5749,N_5017,N_5487);
and U5750 (N_5750,N_5302,N_5321);
and U5751 (N_5751,N_5157,N_5288);
or U5752 (N_5752,N_5344,N_5213);
and U5753 (N_5753,N_5221,N_5302);
or U5754 (N_5754,N_5168,N_5102);
nor U5755 (N_5755,N_5407,N_5207);
nand U5756 (N_5756,N_5493,N_5156);
and U5757 (N_5757,N_5310,N_5207);
and U5758 (N_5758,N_5113,N_5426);
nand U5759 (N_5759,N_5195,N_5265);
or U5760 (N_5760,N_5076,N_5479);
or U5761 (N_5761,N_5027,N_5497);
or U5762 (N_5762,N_5016,N_5414);
nor U5763 (N_5763,N_5430,N_5428);
and U5764 (N_5764,N_5239,N_5363);
nor U5765 (N_5765,N_5110,N_5241);
nand U5766 (N_5766,N_5436,N_5034);
and U5767 (N_5767,N_5145,N_5177);
nor U5768 (N_5768,N_5068,N_5149);
and U5769 (N_5769,N_5206,N_5283);
or U5770 (N_5770,N_5169,N_5296);
or U5771 (N_5771,N_5000,N_5313);
and U5772 (N_5772,N_5401,N_5371);
nor U5773 (N_5773,N_5102,N_5055);
nand U5774 (N_5774,N_5387,N_5228);
and U5775 (N_5775,N_5046,N_5188);
nand U5776 (N_5776,N_5361,N_5231);
and U5777 (N_5777,N_5448,N_5121);
or U5778 (N_5778,N_5237,N_5005);
nand U5779 (N_5779,N_5160,N_5096);
or U5780 (N_5780,N_5142,N_5464);
or U5781 (N_5781,N_5221,N_5091);
and U5782 (N_5782,N_5213,N_5457);
and U5783 (N_5783,N_5291,N_5190);
or U5784 (N_5784,N_5039,N_5481);
and U5785 (N_5785,N_5245,N_5410);
or U5786 (N_5786,N_5326,N_5157);
and U5787 (N_5787,N_5286,N_5437);
xor U5788 (N_5788,N_5412,N_5190);
and U5789 (N_5789,N_5359,N_5160);
nand U5790 (N_5790,N_5015,N_5030);
nor U5791 (N_5791,N_5334,N_5354);
nor U5792 (N_5792,N_5098,N_5386);
or U5793 (N_5793,N_5255,N_5438);
or U5794 (N_5794,N_5249,N_5300);
and U5795 (N_5795,N_5126,N_5439);
and U5796 (N_5796,N_5035,N_5023);
or U5797 (N_5797,N_5001,N_5247);
nand U5798 (N_5798,N_5405,N_5074);
nor U5799 (N_5799,N_5293,N_5483);
nor U5800 (N_5800,N_5422,N_5293);
or U5801 (N_5801,N_5096,N_5196);
or U5802 (N_5802,N_5308,N_5319);
nor U5803 (N_5803,N_5182,N_5060);
nand U5804 (N_5804,N_5336,N_5234);
nor U5805 (N_5805,N_5429,N_5001);
and U5806 (N_5806,N_5206,N_5484);
nor U5807 (N_5807,N_5418,N_5456);
and U5808 (N_5808,N_5219,N_5093);
or U5809 (N_5809,N_5146,N_5416);
or U5810 (N_5810,N_5081,N_5311);
nor U5811 (N_5811,N_5179,N_5498);
or U5812 (N_5812,N_5331,N_5051);
and U5813 (N_5813,N_5165,N_5337);
and U5814 (N_5814,N_5470,N_5233);
and U5815 (N_5815,N_5118,N_5250);
nand U5816 (N_5816,N_5375,N_5424);
nand U5817 (N_5817,N_5213,N_5144);
xnor U5818 (N_5818,N_5319,N_5152);
nand U5819 (N_5819,N_5113,N_5464);
and U5820 (N_5820,N_5375,N_5328);
and U5821 (N_5821,N_5098,N_5139);
nand U5822 (N_5822,N_5000,N_5147);
and U5823 (N_5823,N_5177,N_5155);
or U5824 (N_5824,N_5251,N_5256);
nand U5825 (N_5825,N_5473,N_5421);
nand U5826 (N_5826,N_5407,N_5243);
or U5827 (N_5827,N_5076,N_5207);
nand U5828 (N_5828,N_5169,N_5430);
or U5829 (N_5829,N_5191,N_5337);
and U5830 (N_5830,N_5121,N_5129);
and U5831 (N_5831,N_5298,N_5120);
or U5832 (N_5832,N_5278,N_5123);
or U5833 (N_5833,N_5112,N_5279);
or U5834 (N_5834,N_5496,N_5204);
and U5835 (N_5835,N_5334,N_5262);
nor U5836 (N_5836,N_5161,N_5238);
nand U5837 (N_5837,N_5193,N_5162);
or U5838 (N_5838,N_5382,N_5197);
nand U5839 (N_5839,N_5499,N_5163);
or U5840 (N_5840,N_5041,N_5380);
nand U5841 (N_5841,N_5065,N_5261);
or U5842 (N_5842,N_5202,N_5114);
or U5843 (N_5843,N_5053,N_5038);
nand U5844 (N_5844,N_5166,N_5357);
nand U5845 (N_5845,N_5455,N_5191);
nor U5846 (N_5846,N_5460,N_5393);
and U5847 (N_5847,N_5287,N_5387);
nand U5848 (N_5848,N_5244,N_5498);
nor U5849 (N_5849,N_5245,N_5383);
nor U5850 (N_5850,N_5272,N_5318);
and U5851 (N_5851,N_5497,N_5277);
nor U5852 (N_5852,N_5352,N_5153);
nand U5853 (N_5853,N_5450,N_5404);
xor U5854 (N_5854,N_5194,N_5131);
nand U5855 (N_5855,N_5398,N_5116);
or U5856 (N_5856,N_5414,N_5161);
and U5857 (N_5857,N_5272,N_5160);
and U5858 (N_5858,N_5205,N_5153);
or U5859 (N_5859,N_5009,N_5111);
nor U5860 (N_5860,N_5118,N_5126);
or U5861 (N_5861,N_5032,N_5187);
nand U5862 (N_5862,N_5288,N_5002);
nand U5863 (N_5863,N_5323,N_5237);
or U5864 (N_5864,N_5371,N_5209);
and U5865 (N_5865,N_5056,N_5004);
nor U5866 (N_5866,N_5059,N_5316);
nand U5867 (N_5867,N_5097,N_5274);
and U5868 (N_5868,N_5164,N_5299);
nor U5869 (N_5869,N_5069,N_5233);
nand U5870 (N_5870,N_5487,N_5232);
or U5871 (N_5871,N_5114,N_5083);
or U5872 (N_5872,N_5393,N_5451);
nand U5873 (N_5873,N_5388,N_5053);
nor U5874 (N_5874,N_5302,N_5006);
nor U5875 (N_5875,N_5426,N_5165);
or U5876 (N_5876,N_5324,N_5189);
or U5877 (N_5877,N_5389,N_5128);
or U5878 (N_5878,N_5461,N_5418);
nor U5879 (N_5879,N_5301,N_5156);
or U5880 (N_5880,N_5235,N_5353);
and U5881 (N_5881,N_5163,N_5067);
and U5882 (N_5882,N_5461,N_5339);
nand U5883 (N_5883,N_5334,N_5358);
nand U5884 (N_5884,N_5376,N_5124);
and U5885 (N_5885,N_5016,N_5468);
nand U5886 (N_5886,N_5310,N_5424);
and U5887 (N_5887,N_5018,N_5362);
and U5888 (N_5888,N_5054,N_5400);
nand U5889 (N_5889,N_5210,N_5043);
or U5890 (N_5890,N_5259,N_5469);
or U5891 (N_5891,N_5455,N_5107);
nor U5892 (N_5892,N_5159,N_5461);
nand U5893 (N_5893,N_5286,N_5200);
nor U5894 (N_5894,N_5234,N_5297);
nor U5895 (N_5895,N_5480,N_5126);
or U5896 (N_5896,N_5100,N_5430);
and U5897 (N_5897,N_5462,N_5265);
nor U5898 (N_5898,N_5009,N_5253);
and U5899 (N_5899,N_5271,N_5277);
or U5900 (N_5900,N_5192,N_5108);
and U5901 (N_5901,N_5426,N_5030);
or U5902 (N_5902,N_5075,N_5287);
and U5903 (N_5903,N_5195,N_5220);
and U5904 (N_5904,N_5349,N_5164);
nor U5905 (N_5905,N_5063,N_5130);
nand U5906 (N_5906,N_5368,N_5105);
and U5907 (N_5907,N_5180,N_5332);
nand U5908 (N_5908,N_5117,N_5365);
nor U5909 (N_5909,N_5468,N_5405);
or U5910 (N_5910,N_5135,N_5177);
nand U5911 (N_5911,N_5287,N_5274);
nor U5912 (N_5912,N_5190,N_5165);
or U5913 (N_5913,N_5271,N_5159);
nor U5914 (N_5914,N_5185,N_5409);
and U5915 (N_5915,N_5137,N_5303);
nor U5916 (N_5916,N_5206,N_5348);
or U5917 (N_5917,N_5198,N_5238);
and U5918 (N_5918,N_5165,N_5113);
nand U5919 (N_5919,N_5413,N_5108);
nand U5920 (N_5920,N_5485,N_5478);
and U5921 (N_5921,N_5257,N_5173);
and U5922 (N_5922,N_5199,N_5348);
nand U5923 (N_5923,N_5492,N_5458);
or U5924 (N_5924,N_5060,N_5252);
nand U5925 (N_5925,N_5314,N_5488);
or U5926 (N_5926,N_5188,N_5117);
nand U5927 (N_5927,N_5076,N_5008);
or U5928 (N_5928,N_5216,N_5287);
and U5929 (N_5929,N_5253,N_5327);
nor U5930 (N_5930,N_5239,N_5167);
nor U5931 (N_5931,N_5221,N_5269);
or U5932 (N_5932,N_5386,N_5057);
and U5933 (N_5933,N_5224,N_5250);
nor U5934 (N_5934,N_5130,N_5367);
and U5935 (N_5935,N_5127,N_5018);
or U5936 (N_5936,N_5246,N_5249);
nand U5937 (N_5937,N_5311,N_5063);
nand U5938 (N_5938,N_5297,N_5471);
nand U5939 (N_5939,N_5213,N_5206);
or U5940 (N_5940,N_5142,N_5328);
and U5941 (N_5941,N_5207,N_5124);
nand U5942 (N_5942,N_5307,N_5464);
or U5943 (N_5943,N_5057,N_5352);
nand U5944 (N_5944,N_5217,N_5295);
nand U5945 (N_5945,N_5177,N_5088);
nor U5946 (N_5946,N_5083,N_5334);
nand U5947 (N_5947,N_5078,N_5344);
or U5948 (N_5948,N_5251,N_5257);
or U5949 (N_5949,N_5177,N_5019);
or U5950 (N_5950,N_5198,N_5137);
nor U5951 (N_5951,N_5044,N_5029);
nor U5952 (N_5952,N_5403,N_5135);
or U5953 (N_5953,N_5237,N_5329);
xor U5954 (N_5954,N_5357,N_5227);
xor U5955 (N_5955,N_5250,N_5467);
nor U5956 (N_5956,N_5477,N_5291);
nand U5957 (N_5957,N_5141,N_5476);
or U5958 (N_5958,N_5086,N_5318);
or U5959 (N_5959,N_5085,N_5407);
and U5960 (N_5960,N_5271,N_5154);
nand U5961 (N_5961,N_5280,N_5451);
or U5962 (N_5962,N_5302,N_5352);
nand U5963 (N_5963,N_5033,N_5136);
nor U5964 (N_5964,N_5329,N_5141);
and U5965 (N_5965,N_5121,N_5349);
nor U5966 (N_5966,N_5470,N_5377);
or U5967 (N_5967,N_5460,N_5115);
or U5968 (N_5968,N_5163,N_5019);
or U5969 (N_5969,N_5024,N_5033);
and U5970 (N_5970,N_5191,N_5121);
nand U5971 (N_5971,N_5321,N_5022);
xor U5972 (N_5972,N_5107,N_5392);
nand U5973 (N_5973,N_5168,N_5496);
and U5974 (N_5974,N_5483,N_5372);
xnor U5975 (N_5975,N_5221,N_5137);
and U5976 (N_5976,N_5251,N_5308);
and U5977 (N_5977,N_5144,N_5364);
nor U5978 (N_5978,N_5005,N_5383);
or U5979 (N_5979,N_5012,N_5153);
nor U5980 (N_5980,N_5368,N_5276);
and U5981 (N_5981,N_5395,N_5282);
nand U5982 (N_5982,N_5358,N_5109);
nor U5983 (N_5983,N_5382,N_5025);
or U5984 (N_5984,N_5400,N_5142);
or U5985 (N_5985,N_5230,N_5116);
or U5986 (N_5986,N_5420,N_5435);
nand U5987 (N_5987,N_5401,N_5439);
and U5988 (N_5988,N_5110,N_5385);
or U5989 (N_5989,N_5029,N_5395);
or U5990 (N_5990,N_5447,N_5150);
nor U5991 (N_5991,N_5261,N_5257);
and U5992 (N_5992,N_5024,N_5218);
or U5993 (N_5993,N_5153,N_5434);
nand U5994 (N_5994,N_5109,N_5172);
or U5995 (N_5995,N_5292,N_5012);
and U5996 (N_5996,N_5278,N_5484);
nand U5997 (N_5997,N_5085,N_5095);
nor U5998 (N_5998,N_5053,N_5422);
or U5999 (N_5999,N_5499,N_5439);
nor U6000 (N_6000,N_5777,N_5690);
and U6001 (N_6001,N_5829,N_5557);
nand U6002 (N_6002,N_5889,N_5576);
and U6003 (N_6003,N_5731,N_5669);
nand U6004 (N_6004,N_5886,N_5679);
nor U6005 (N_6005,N_5890,N_5602);
nor U6006 (N_6006,N_5951,N_5756);
nor U6007 (N_6007,N_5677,N_5661);
nor U6008 (N_6008,N_5521,N_5845);
nor U6009 (N_6009,N_5538,N_5788);
or U6010 (N_6010,N_5820,N_5981);
nor U6011 (N_6011,N_5701,N_5581);
nor U6012 (N_6012,N_5684,N_5902);
and U6013 (N_6013,N_5543,N_5587);
nand U6014 (N_6014,N_5773,N_5834);
nand U6015 (N_6015,N_5640,N_5595);
or U6016 (N_6016,N_5863,N_5974);
and U6017 (N_6017,N_5843,N_5645);
nand U6018 (N_6018,N_5720,N_5940);
or U6019 (N_6019,N_5934,N_5597);
nor U6020 (N_6020,N_5753,N_5852);
or U6021 (N_6021,N_5901,N_5651);
nand U6022 (N_6022,N_5751,N_5582);
or U6023 (N_6023,N_5765,N_5665);
and U6024 (N_6024,N_5642,N_5999);
nand U6025 (N_6025,N_5818,N_5618);
or U6026 (N_6026,N_5688,N_5947);
or U6027 (N_6027,N_5639,N_5949);
and U6028 (N_6028,N_5938,N_5807);
and U6029 (N_6029,N_5969,N_5917);
or U6030 (N_6030,N_5859,N_5752);
nand U6031 (N_6031,N_5839,N_5687);
nand U6032 (N_6032,N_5727,N_5821);
and U6033 (N_6033,N_5626,N_5911);
and U6034 (N_6034,N_5790,N_5896);
nand U6035 (N_6035,N_5736,N_5563);
nor U6036 (N_6036,N_5923,N_5776);
and U6037 (N_6037,N_5604,N_5881);
and U6038 (N_6038,N_5990,N_5786);
or U6039 (N_6039,N_5551,N_5635);
nand U6040 (N_6040,N_5875,N_5854);
or U6041 (N_6041,N_5713,N_5833);
or U6042 (N_6042,N_5771,N_5714);
or U6043 (N_6043,N_5608,N_5919);
or U6044 (N_6044,N_5691,N_5780);
and U6045 (N_6045,N_5916,N_5517);
nor U6046 (N_6046,N_5998,N_5828);
nand U6047 (N_6047,N_5957,N_5953);
or U6048 (N_6048,N_5932,N_5656);
and U6049 (N_6049,N_5747,N_5680);
nor U6050 (N_6050,N_5678,N_5900);
and U6051 (N_6051,N_5585,N_5993);
nand U6052 (N_6052,N_5866,N_5583);
nor U6053 (N_6053,N_5697,N_5700);
and U6054 (N_6054,N_5841,N_5758);
nor U6055 (N_6055,N_5897,N_5696);
or U6056 (N_6056,N_5681,N_5813);
nor U6057 (N_6057,N_5819,N_5927);
nor U6058 (N_6058,N_5518,N_5762);
or U6059 (N_6059,N_5768,N_5692);
nor U6060 (N_6060,N_5532,N_5598);
and U6061 (N_6061,N_5507,N_5805);
nand U6062 (N_6062,N_5750,N_5593);
nand U6063 (N_6063,N_5827,N_5825);
nand U6064 (N_6064,N_5908,N_5944);
nor U6065 (N_6065,N_5997,N_5530);
xor U6066 (N_6066,N_5577,N_5966);
nor U6067 (N_6067,N_5505,N_5667);
or U6068 (N_6068,N_5888,N_5516);
and U6069 (N_6069,N_5924,N_5766);
nor U6070 (N_6070,N_5670,N_5874);
nor U6071 (N_6071,N_5826,N_5726);
nor U6072 (N_6072,N_5718,N_5848);
nand U6073 (N_6073,N_5809,N_5560);
xor U6074 (N_6074,N_5745,N_5878);
nand U6075 (N_6075,N_5935,N_5509);
nand U6076 (N_6076,N_5501,N_5569);
or U6077 (N_6077,N_5784,N_5894);
or U6078 (N_6078,N_5971,N_5785);
nor U6079 (N_6079,N_5967,N_5794);
nand U6080 (N_6080,N_5553,N_5512);
nand U6081 (N_6081,N_5955,N_5710);
and U6082 (N_6082,N_5570,N_5973);
nor U6083 (N_6083,N_5636,N_5571);
and U6084 (N_6084,N_5939,N_5504);
nand U6085 (N_6085,N_5895,N_5907);
or U6086 (N_6086,N_5616,N_5673);
and U6087 (N_6087,N_5580,N_5686);
nand U6088 (N_6088,N_5808,N_5860);
nor U6089 (N_6089,N_5989,N_5711);
or U6090 (N_6090,N_5948,N_5849);
nand U6091 (N_6091,N_5926,N_5883);
or U6092 (N_6092,N_5950,N_5613);
or U6093 (N_6093,N_5767,N_5801);
nor U6094 (N_6094,N_5757,N_5921);
nand U6095 (N_6095,N_5510,N_5740);
nor U6096 (N_6096,N_5545,N_5755);
nor U6097 (N_6097,N_5905,N_5659);
or U6098 (N_6098,N_5842,N_5864);
nand U6099 (N_6099,N_5601,N_5666);
nand U6100 (N_6100,N_5943,N_5742);
nor U6101 (N_6101,N_5522,N_5527);
nor U6102 (N_6102,N_5572,N_5706);
xor U6103 (N_6103,N_5664,N_5929);
nor U6104 (N_6104,N_5632,N_5719);
and U6105 (N_6105,N_5945,N_5937);
and U6106 (N_6106,N_5946,N_5591);
nand U6107 (N_6107,N_5520,N_5975);
nand U6108 (N_6108,N_5564,N_5619);
and U6109 (N_6109,N_5609,N_5803);
nand U6110 (N_6110,N_5868,N_5856);
nand U6111 (N_6111,N_5717,N_5528);
nand U6112 (N_6112,N_5554,N_5853);
or U6113 (N_6113,N_5574,N_5987);
and U6114 (N_6114,N_5738,N_5732);
nor U6115 (N_6115,N_5796,N_5658);
or U6116 (N_6116,N_5857,N_5599);
and U6117 (N_6117,N_5832,N_5892);
or U6118 (N_6118,N_5844,N_5728);
xnor U6119 (N_6119,N_5579,N_5693);
and U6120 (N_6120,N_5565,N_5793);
and U6121 (N_6121,N_5815,N_5649);
and U6122 (N_6122,N_5566,N_5723);
nand U6123 (N_6123,N_5634,N_5631);
nand U6124 (N_6124,N_5643,N_5741);
nor U6125 (N_6125,N_5850,N_5871);
nor U6126 (N_6126,N_5672,N_5920);
or U6127 (N_6127,N_5630,N_5623);
or U6128 (N_6128,N_5622,N_5748);
nand U6129 (N_6129,N_5676,N_5712);
and U6130 (N_6130,N_5781,N_5983);
nand U6131 (N_6131,N_5739,N_5912);
or U6132 (N_6132,N_5858,N_5968);
and U6133 (N_6133,N_5986,N_5596);
nor U6134 (N_6134,N_5823,N_5698);
or U6135 (N_6135,N_5590,N_5514);
nor U6136 (N_6136,N_5822,N_5746);
nor U6137 (N_6137,N_5531,N_5737);
nand U6138 (N_6138,N_5715,N_5637);
and U6139 (N_6139,N_5734,N_5627);
and U6140 (N_6140,N_5972,N_5963);
or U6141 (N_6141,N_5559,N_5562);
nand U6142 (N_6142,N_5707,N_5539);
and U6143 (N_6143,N_5760,N_5526);
and U6144 (N_6144,N_5502,N_5996);
and U6145 (N_6145,N_5847,N_5840);
nand U6146 (N_6146,N_5699,N_5918);
nor U6147 (N_6147,N_5544,N_5876);
nand U6148 (N_6148,N_5754,N_5668);
nand U6149 (N_6149,N_5513,N_5804);
or U6150 (N_6150,N_5814,N_5958);
or U6151 (N_6151,N_5759,N_5855);
nor U6152 (N_6152,N_5952,N_5708);
and U6153 (N_6153,N_5542,N_5641);
nor U6154 (N_6154,N_5671,N_5798);
or U6155 (N_6155,N_5617,N_5561);
nor U6156 (N_6156,N_5709,N_5647);
and U6157 (N_6157,N_5533,N_5744);
nand U6158 (N_6158,N_5933,N_5870);
nor U6159 (N_6159,N_5956,N_5795);
nor U6160 (N_6160,N_5615,N_5913);
and U6161 (N_6161,N_5705,N_5685);
nand U6162 (N_6162,N_5980,N_5729);
nor U6163 (N_6163,N_5730,N_5600);
or U6164 (N_6164,N_5772,N_5869);
or U6165 (N_6165,N_5592,N_5650);
nor U6166 (N_6166,N_5578,N_5936);
or U6167 (N_6167,N_5694,N_5928);
nand U6168 (N_6168,N_5534,N_5769);
nand U6169 (N_6169,N_5519,N_5515);
and U6170 (N_6170,N_5607,N_5824);
and U6171 (N_6171,N_5702,N_5594);
or U6172 (N_6172,N_5941,N_5761);
and U6173 (N_6173,N_5584,N_5898);
or U6174 (N_6174,N_5552,N_5909);
and U6175 (N_6175,N_5644,N_5979);
nand U6176 (N_6176,N_5621,N_5537);
nand U6177 (N_6177,N_5774,N_5589);
and U6178 (N_6178,N_5962,N_5872);
nand U6179 (N_6179,N_5851,N_5978);
or U6180 (N_6180,N_5994,N_5877);
and U6181 (N_6181,N_5704,N_5861);
nor U6182 (N_6182,N_5646,N_5653);
and U6183 (N_6183,N_5547,N_5573);
xor U6184 (N_6184,N_5503,N_5887);
and U6185 (N_6185,N_5838,N_5524);
and U6186 (N_6186,N_5903,N_5846);
and U6187 (N_6187,N_5633,N_5942);
nor U6188 (N_6188,N_5612,N_5882);
nor U6189 (N_6189,N_5799,N_5893);
nor U6190 (N_6190,N_5914,N_5995);
nand U6191 (N_6191,N_5610,N_5770);
nor U6192 (N_6192,N_5764,N_5660);
or U6193 (N_6193,N_5689,N_5862);
nor U6194 (N_6194,N_5663,N_5568);
or U6195 (N_6195,N_5541,N_5558);
or U6196 (N_6196,N_5638,N_5523);
or U6197 (N_6197,N_5508,N_5906);
and U6198 (N_6198,N_5873,N_5654);
nand U6199 (N_6199,N_5586,N_5792);
or U6200 (N_6200,N_5812,N_5791);
nand U6201 (N_6201,N_5970,N_5724);
nor U6202 (N_6202,N_5606,N_5683);
nand U6203 (N_6203,N_5749,N_5817);
or U6204 (N_6204,N_5797,N_5500);
and U6205 (N_6205,N_5954,N_5783);
and U6206 (N_6206,N_5614,N_5960);
nor U6207 (N_6207,N_5703,N_5787);
or U6208 (N_6208,N_5735,N_5611);
and U6209 (N_6209,N_5992,N_5961);
nor U6210 (N_6210,N_5535,N_5984);
nand U6211 (N_6211,N_5620,N_5567);
nor U6212 (N_6212,N_5985,N_5778);
and U6213 (N_6213,N_5930,N_5743);
or U6214 (N_6214,N_5550,N_5721);
nand U6215 (N_6215,N_5775,N_5695);
and U6216 (N_6216,N_5965,N_5657);
nor U6217 (N_6217,N_5763,N_5977);
and U6218 (N_6218,N_5540,N_5899);
or U6219 (N_6219,N_5915,N_5733);
nand U6220 (N_6220,N_5603,N_5782);
nand U6221 (N_6221,N_5867,N_5555);
nor U6222 (N_6222,N_5536,N_5529);
nand U6223 (N_6223,N_5625,N_5991);
nand U6224 (N_6224,N_5811,N_5879);
nand U6225 (N_6225,N_5648,N_5605);
nor U6226 (N_6226,N_5722,N_5556);
and U6227 (N_6227,N_5588,N_5988);
nand U6228 (N_6228,N_5837,N_5810);
or U6229 (N_6229,N_5629,N_5885);
or U6230 (N_6230,N_5836,N_5674);
nand U6231 (N_6231,N_5976,N_5891);
or U6232 (N_6232,N_5662,N_5931);
and U6233 (N_6233,N_5925,N_5865);
nor U6234 (N_6234,N_5628,N_5884);
or U6235 (N_6235,N_5816,N_5682);
nor U6236 (N_6236,N_5982,N_5800);
or U6237 (N_6237,N_5506,N_5922);
and U6238 (N_6238,N_5789,N_5725);
or U6239 (N_6239,N_5525,N_5549);
nor U6240 (N_6240,N_5652,N_5716);
or U6241 (N_6241,N_5779,N_5835);
and U6242 (N_6242,N_5831,N_5675);
or U6243 (N_6243,N_5959,N_5830);
nor U6244 (N_6244,N_5964,N_5910);
or U6245 (N_6245,N_5806,N_5548);
or U6246 (N_6246,N_5575,N_5546);
and U6247 (N_6247,N_5904,N_5655);
nor U6248 (N_6248,N_5802,N_5511);
nand U6249 (N_6249,N_5880,N_5624);
nor U6250 (N_6250,N_5850,N_5770);
xor U6251 (N_6251,N_5945,N_5578);
nor U6252 (N_6252,N_5821,N_5567);
or U6253 (N_6253,N_5766,N_5803);
or U6254 (N_6254,N_5569,N_5656);
nand U6255 (N_6255,N_5906,N_5911);
nand U6256 (N_6256,N_5720,N_5674);
nor U6257 (N_6257,N_5732,N_5681);
nand U6258 (N_6258,N_5657,N_5883);
and U6259 (N_6259,N_5955,N_5841);
nor U6260 (N_6260,N_5818,N_5918);
nand U6261 (N_6261,N_5676,N_5789);
nand U6262 (N_6262,N_5962,N_5969);
nor U6263 (N_6263,N_5562,N_5675);
nand U6264 (N_6264,N_5629,N_5851);
nand U6265 (N_6265,N_5848,N_5660);
nand U6266 (N_6266,N_5797,N_5844);
or U6267 (N_6267,N_5772,N_5948);
and U6268 (N_6268,N_5874,N_5699);
or U6269 (N_6269,N_5579,N_5949);
or U6270 (N_6270,N_5583,N_5850);
nand U6271 (N_6271,N_5635,N_5707);
nor U6272 (N_6272,N_5834,N_5763);
xor U6273 (N_6273,N_5555,N_5815);
or U6274 (N_6274,N_5997,N_5924);
nor U6275 (N_6275,N_5718,N_5962);
or U6276 (N_6276,N_5646,N_5883);
and U6277 (N_6277,N_5751,N_5507);
nand U6278 (N_6278,N_5706,N_5685);
nand U6279 (N_6279,N_5755,N_5509);
nand U6280 (N_6280,N_5657,N_5885);
nor U6281 (N_6281,N_5797,N_5894);
or U6282 (N_6282,N_5505,N_5870);
and U6283 (N_6283,N_5820,N_5595);
or U6284 (N_6284,N_5502,N_5887);
xor U6285 (N_6285,N_5939,N_5789);
nor U6286 (N_6286,N_5921,N_5885);
and U6287 (N_6287,N_5933,N_5818);
nor U6288 (N_6288,N_5798,N_5597);
nor U6289 (N_6289,N_5717,N_5774);
or U6290 (N_6290,N_5652,N_5684);
and U6291 (N_6291,N_5672,N_5784);
and U6292 (N_6292,N_5779,N_5966);
nand U6293 (N_6293,N_5832,N_5899);
nor U6294 (N_6294,N_5849,N_5823);
xor U6295 (N_6295,N_5539,N_5885);
or U6296 (N_6296,N_5907,N_5505);
nand U6297 (N_6297,N_5732,N_5757);
nor U6298 (N_6298,N_5884,N_5830);
or U6299 (N_6299,N_5711,N_5745);
nor U6300 (N_6300,N_5962,N_5755);
and U6301 (N_6301,N_5890,N_5857);
and U6302 (N_6302,N_5503,N_5508);
and U6303 (N_6303,N_5617,N_5626);
nor U6304 (N_6304,N_5543,N_5885);
nand U6305 (N_6305,N_5594,N_5666);
nand U6306 (N_6306,N_5933,N_5581);
nand U6307 (N_6307,N_5735,N_5831);
or U6308 (N_6308,N_5814,N_5984);
nor U6309 (N_6309,N_5783,N_5848);
nor U6310 (N_6310,N_5511,N_5556);
nand U6311 (N_6311,N_5958,N_5831);
nor U6312 (N_6312,N_5625,N_5570);
and U6313 (N_6313,N_5793,N_5867);
or U6314 (N_6314,N_5967,N_5974);
and U6315 (N_6315,N_5593,N_5885);
nor U6316 (N_6316,N_5848,N_5599);
nand U6317 (N_6317,N_5614,N_5795);
or U6318 (N_6318,N_5690,N_5929);
or U6319 (N_6319,N_5562,N_5548);
nor U6320 (N_6320,N_5826,N_5999);
nand U6321 (N_6321,N_5733,N_5696);
or U6322 (N_6322,N_5811,N_5513);
nor U6323 (N_6323,N_5672,N_5628);
nand U6324 (N_6324,N_5880,N_5986);
and U6325 (N_6325,N_5565,N_5645);
nand U6326 (N_6326,N_5688,N_5910);
or U6327 (N_6327,N_5503,N_5639);
nor U6328 (N_6328,N_5698,N_5779);
xnor U6329 (N_6329,N_5501,N_5684);
or U6330 (N_6330,N_5879,N_5942);
and U6331 (N_6331,N_5506,N_5805);
and U6332 (N_6332,N_5794,N_5593);
or U6333 (N_6333,N_5951,N_5657);
nor U6334 (N_6334,N_5564,N_5897);
nor U6335 (N_6335,N_5840,N_5507);
nand U6336 (N_6336,N_5834,N_5967);
nand U6337 (N_6337,N_5777,N_5783);
and U6338 (N_6338,N_5679,N_5855);
or U6339 (N_6339,N_5543,N_5936);
or U6340 (N_6340,N_5551,N_5791);
nor U6341 (N_6341,N_5864,N_5798);
or U6342 (N_6342,N_5671,N_5795);
nor U6343 (N_6343,N_5708,N_5693);
nor U6344 (N_6344,N_5555,N_5964);
nand U6345 (N_6345,N_5936,N_5729);
nor U6346 (N_6346,N_5735,N_5548);
nand U6347 (N_6347,N_5958,N_5527);
nand U6348 (N_6348,N_5571,N_5574);
and U6349 (N_6349,N_5511,N_5740);
nand U6350 (N_6350,N_5648,N_5912);
and U6351 (N_6351,N_5921,N_5882);
xnor U6352 (N_6352,N_5724,N_5584);
nand U6353 (N_6353,N_5663,N_5689);
nand U6354 (N_6354,N_5854,N_5921);
and U6355 (N_6355,N_5526,N_5693);
nand U6356 (N_6356,N_5572,N_5857);
nor U6357 (N_6357,N_5655,N_5700);
nand U6358 (N_6358,N_5699,N_5948);
or U6359 (N_6359,N_5547,N_5911);
and U6360 (N_6360,N_5861,N_5848);
nand U6361 (N_6361,N_5671,N_5584);
nor U6362 (N_6362,N_5833,N_5907);
or U6363 (N_6363,N_5668,N_5884);
or U6364 (N_6364,N_5694,N_5986);
and U6365 (N_6365,N_5869,N_5864);
xor U6366 (N_6366,N_5557,N_5645);
and U6367 (N_6367,N_5905,N_5580);
nor U6368 (N_6368,N_5872,N_5638);
and U6369 (N_6369,N_5725,N_5960);
or U6370 (N_6370,N_5988,N_5625);
nand U6371 (N_6371,N_5571,N_5831);
nor U6372 (N_6372,N_5568,N_5705);
nand U6373 (N_6373,N_5788,N_5721);
and U6374 (N_6374,N_5585,N_5691);
or U6375 (N_6375,N_5664,N_5696);
nand U6376 (N_6376,N_5667,N_5587);
nor U6377 (N_6377,N_5723,N_5590);
nor U6378 (N_6378,N_5873,N_5581);
or U6379 (N_6379,N_5996,N_5924);
nor U6380 (N_6380,N_5746,N_5515);
or U6381 (N_6381,N_5701,N_5824);
or U6382 (N_6382,N_5819,N_5772);
nor U6383 (N_6383,N_5983,N_5882);
nand U6384 (N_6384,N_5581,N_5938);
nor U6385 (N_6385,N_5607,N_5868);
nand U6386 (N_6386,N_5613,N_5871);
nand U6387 (N_6387,N_5829,N_5615);
xor U6388 (N_6388,N_5505,N_5503);
or U6389 (N_6389,N_5517,N_5513);
or U6390 (N_6390,N_5666,N_5816);
or U6391 (N_6391,N_5526,N_5877);
nor U6392 (N_6392,N_5732,N_5599);
and U6393 (N_6393,N_5975,N_5922);
and U6394 (N_6394,N_5914,N_5681);
and U6395 (N_6395,N_5566,N_5701);
nand U6396 (N_6396,N_5916,N_5619);
nand U6397 (N_6397,N_5766,N_5763);
or U6398 (N_6398,N_5527,N_5596);
nor U6399 (N_6399,N_5776,N_5891);
nand U6400 (N_6400,N_5615,N_5642);
or U6401 (N_6401,N_5875,N_5988);
and U6402 (N_6402,N_5805,N_5746);
and U6403 (N_6403,N_5539,N_5867);
or U6404 (N_6404,N_5943,N_5631);
or U6405 (N_6405,N_5883,N_5725);
and U6406 (N_6406,N_5624,N_5827);
and U6407 (N_6407,N_5750,N_5537);
nand U6408 (N_6408,N_5803,N_5619);
and U6409 (N_6409,N_5853,N_5548);
or U6410 (N_6410,N_5972,N_5680);
or U6411 (N_6411,N_5589,N_5657);
nor U6412 (N_6412,N_5686,N_5954);
and U6413 (N_6413,N_5821,N_5881);
or U6414 (N_6414,N_5914,N_5831);
nand U6415 (N_6415,N_5861,N_5517);
nand U6416 (N_6416,N_5765,N_5716);
or U6417 (N_6417,N_5534,N_5868);
and U6418 (N_6418,N_5955,N_5718);
nor U6419 (N_6419,N_5672,N_5890);
nand U6420 (N_6420,N_5680,N_5627);
nand U6421 (N_6421,N_5618,N_5836);
nand U6422 (N_6422,N_5741,N_5598);
nor U6423 (N_6423,N_5922,N_5690);
nor U6424 (N_6424,N_5855,N_5842);
nor U6425 (N_6425,N_5525,N_5750);
and U6426 (N_6426,N_5525,N_5923);
and U6427 (N_6427,N_5634,N_5956);
or U6428 (N_6428,N_5974,N_5847);
and U6429 (N_6429,N_5607,N_5553);
and U6430 (N_6430,N_5792,N_5512);
or U6431 (N_6431,N_5614,N_5939);
or U6432 (N_6432,N_5870,N_5969);
nand U6433 (N_6433,N_5928,N_5763);
and U6434 (N_6434,N_5947,N_5634);
and U6435 (N_6435,N_5607,N_5522);
xnor U6436 (N_6436,N_5632,N_5740);
nor U6437 (N_6437,N_5794,N_5844);
and U6438 (N_6438,N_5543,N_5968);
nor U6439 (N_6439,N_5837,N_5671);
nor U6440 (N_6440,N_5547,N_5827);
or U6441 (N_6441,N_5700,N_5871);
xnor U6442 (N_6442,N_5967,N_5983);
nand U6443 (N_6443,N_5605,N_5663);
or U6444 (N_6444,N_5798,N_5567);
and U6445 (N_6445,N_5638,N_5586);
nor U6446 (N_6446,N_5668,N_5676);
nand U6447 (N_6447,N_5814,N_5627);
nor U6448 (N_6448,N_5916,N_5631);
nand U6449 (N_6449,N_5881,N_5786);
and U6450 (N_6450,N_5514,N_5712);
nor U6451 (N_6451,N_5580,N_5962);
nor U6452 (N_6452,N_5508,N_5718);
xor U6453 (N_6453,N_5948,N_5924);
nand U6454 (N_6454,N_5930,N_5965);
nand U6455 (N_6455,N_5744,N_5502);
xor U6456 (N_6456,N_5698,N_5731);
nor U6457 (N_6457,N_5703,N_5734);
or U6458 (N_6458,N_5857,N_5558);
and U6459 (N_6459,N_5887,N_5866);
nand U6460 (N_6460,N_5988,N_5593);
nor U6461 (N_6461,N_5686,N_5702);
nor U6462 (N_6462,N_5512,N_5624);
nand U6463 (N_6463,N_5546,N_5594);
nand U6464 (N_6464,N_5583,N_5511);
or U6465 (N_6465,N_5569,N_5867);
nand U6466 (N_6466,N_5543,N_5769);
and U6467 (N_6467,N_5885,N_5695);
or U6468 (N_6468,N_5858,N_5647);
nor U6469 (N_6469,N_5749,N_5977);
and U6470 (N_6470,N_5625,N_5774);
nor U6471 (N_6471,N_5549,N_5925);
and U6472 (N_6472,N_5995,N_5504);
and U6473 (N_6473,N_5752,N_5549);
nand U6474 (N_6474,N_5831,N_5907);
or U6475 (N_6475,N_5572,N_5945);
nor U6476 (N_6476,N_5761,N_5600);
and U6477 (N_6477,N_5962,N_5663);
or U6478 (N_6478,N_5518,N_5680);
nand U6479 (N_6479,N_5656,N_5783);
nor U6480 (N_6480,N_5986,N_5950);
nor U6481 (N_6481,N_5861,N_5639);
and U6482 (N_6482,N_5991,N_5668);
or U6483 (N_6483,N_5736,N_5661);
xnor U6484 (N_6484,N_5813,N_5895);
or U6485 (N_6485,N_5694,N_5999);
xnor U6486 (N_6486,N_5833,N_5962);
nand U6487 (N_6487,N_5823,N_5920);
nand U6488 (N_6488,N_5933,N_5724);
nor U6489 (N_6489,N_5591,N_5633);
and U6490 (N_6490,N_5654,N_5714);
nor U6491 (N_6491,N_5910,N_5915);
nor U6492 (N_6492,N_5698,N_5865);
or U6493 (N_6493,N_5953,N_5526);
nor U6494 (N_6494,N_5560,N_5807);
and U6495 (N_6495,N_5724,N_5727);
and U6496 (N_6496,N_5669,N_5971);
and U6497 (N_6497,N_5840,N_5757);
and U6498 (N_6498,N_5833,N_5634);
or U6499 (N_6499,N_5677,N_5898);
nor U6500 (N_6500,N_6355,N_6325);
nand U6501 (N_6501,N_6249,N_6434);
nor U6502 (N_6502,N_6032,N_6103);
or U6503 (N_6503,N_6343,N_6307);
or U6504 (N_6504,N_6132,N_6398);
or U6505 (N_6505,N_6273,N_6117);
and U6506 (N_6506,N_6478,N_6145);
and U6507 (N_6507,N_6148,N_6058);
and U6508 (N_6508,N_6372,N_6092);
and U6509 (N_6509,N_6040,N_6229);
nand U6510 (N_6510,N_6477,N_6067);
nor U6511 (N_6511,N_6349,N_6350);
nor U6512 (N_6512,N_6286,N_6400);
nand U6513 (N_6513,N_6115,N_6451);
nand U6514 (N_6514,N_6379,N_6134);
nor U6515 (N_6515,N_6404,N_6193);
nand U6516 (N_6516,N_6172,N_6199);
or U6517 (N_6517,N_6484,N_6001);
nor U6518 (N_6518,N_6472,N_6374);
and U6519 (N_6519,N_6321,N_6065);
or U6520 (N_6520,N_6322,N_6158);
and U6521 (N_6521,N_6353,N_6427);
or U6522 (N_6522,N_6483,N_6124);
and U6523 (N_6523,N_6051,N_6244);
nor U6524 (N_6524,N_6462,N_6498);
nor U6525 (N_6525,N_6112,N_6107);
nor U6526 (N_6526,N_6126,N_6493);
and U6527 (N_6527,N_6288,N_6463);
xor U6528 (N_6528,N_6388,N_6075);
or U6529 (N_6529,N_6086,N_6183);
nor U6530 (N_6530,N_6409,N_6176);
or U6531 (N_6531,N_6271,N_6243);
and U6532 (N_6532,N_6085,N_6200);
nor U6533 (N_6533,N_6253,N_6010);
nor U6534 (N_6534,N_6188,N_6141);
nor U6535 (N_6535,N_6245,N_6029);
and U6536 (N_6536,N_6382,N_6280);
and U6537 (N_6537,N_6308,N_6143);
or U6538 (N_6538,N_6333,N_6387);
and U6539 (N_6539,N_6386,N_6442);
nand U6540 (N_6540,N_6323,N_6088);
or U6541 (N_6541,N_6133,N_6237);
or U6542 (N_6542,N_6408,N_6282);
nand U6543 (N_6543,N_6405,N_6284);
or U6544 (N_6544,N_6482,N_6480);
and U6545 (N_6545,N_6167,N_6073);
nor U6546 (N_6546,N_6332,N_6021);
or U6547 (N_6547,N_6219,N_6044);
nand U6548 (N_6548,N_6182,N_6473);
nor U6549 (N_6549,N_6373,N_6091);
or U6550 (N_6550,N_6022,N_6429);
nor U6551 (N_6551,N_6114,N_6038);
nor U6552 (N_6552,N_6417,N_6313);
xnor U6553 (N_6553,N_6142,N_6125);
or U6554 (N_6554,N_6450,N_6383);
xnor U6555 (N_6555,N_6055,N_6069);
and U6556 (N_6556,N_6053,N_6234);
or U6557 (N_6557,N_6415,N_6389);
or U6558 (N_6558,N_6329,N_6033);
nor U6559 (N_6559,N_6302,N_6163);
and U6560 (N_6560,N_6147,N_6265);
nor U6561 (N_6561,N_6440,N_6093);
nand U6562 (N_6562,N_6187,N_6410);
and U6563 (N_6563,N_6403,N_6359);
nor U6564 (N_6564,N_6407,N_6251);
nor U6565 (N_6565,N_6102,N_6207);
nor U6566 (N_6566,N_6424,N_6334);
nand U6567 (N_6567,N_6023,N_6454);
or U6568 (N_6568,N_6306,N_6411);
nand U6569 (N_6569,N_6294,N_6241);
nand U6570 (N_6570,N_6337,N_6211);
nand U6571 (N_6571,N_6290,N_6303);
and U6572 (N_6572,N_6105,N_6214);
or U6573 (N_6573,N_6223,N_6311);
and U6574 (N_6574,N_6377,N_6293);
or U6575 (N_6575,N_6458,N_6178);
or U6576 (N_6576,N_6213,N_6423);
and U6577 (N_6577,N_6250,N_6020);
nand U6578 (N_6578,N_6314,N_6448);
nor U6579 (N_6579,N_6231,N_6270);
and U6580 (N_6580,N_6456,N_6426);
or U6581 (N_6581,N_6089,N_6104);
and U6582 (N_6582,N_6481,N_6138);
or U6583 (N_6583,N_6192,N_6452);
nand U6584 (N_6584,N_6196,N_6479);
nand U6585 (N_6585,N_6468,N_6239);
nor U6586 (N_6586,N_6340,N_6292);
nor U6587 (N_6587,N_6003,N_6057);
and U6588 (N_6588,N_6376,N_6257);
nor U6589 (N_6589,N_6018,N_6489);
nor U6590 (N_6590,N_6464,N_6371);
nor U6591 (N_6591,N_6399,N_6179);
and U6592 (N_6592,N_6165,N_6397);
or U6593 (N_6593,N_6246,N_6430);
nand U6594 (N_6594,N_6202,N_6390);
nor U6595 (N_6595,N_6146,N_6443);
nand U6596 (N_6596,N_6064,N_6221);
and U6597 (N_6597,N_6151,N_6395);
and U6598 (N_6598,N_6358,N_6025);
and U6599 (N_6599,N_6381,N_6283);
nand U6600 (N_6600,N_6320,N_6100);
or U6601 (N_6601,N_6275,N_6154);
nor U6602 (N_6602,N_6406,N_6242);
nand U6603 (N_6603,N_6084,N_6002);
and U6604 (N_6604,N_6037,N_6122);
nor U6605 (N_6605,N_6272,N_6296);
xor U6606 (N_6606,N_6432,N_6419);
and U6607 (N_6607,N_6418,N_6016);
nor U6608 (N_6608,N_6365,N_6378);
nor U6609 (N_6609,N_6486,N_6485);
nor U6610 (N_6610,N_6366,N_6225);
nor U6611 (N_6611,N_6299,N_6120);
nand U6612 (N_6612,N_6446,N_6228);
or U6613 (N_6613,N_6341,N_6248);
nor U6614 (N_6614,N_6420,N_6177);
nor U6615 (N_6615,N_6360,N_6068);
nor U6616 (N_6616,N_6080,N_6101);
or U6617 (N_6617,N_6471,N_6487);
and U6618 (N_6618,N_6045,N_6318);
nor U6619 (N_6619,N_6054,N_6444);
xor U6620 (N_6620,N_6465,N_6205);
and U6621 (N_6621,N_6152,N_6319);
and U6622 (N_6622,N_6123,N_6437);
and U6623 (N_6623,N_6317,N_6162);
nand U6624 (N_6624,N_6050,N_6180);
or U6625 (N_6625,N_6279,N_6166);
nor U6626 (N_6626,N_6356,N_6190);
or U6627 (N_6627,N_6140,N_6087);
nor U6628 (N_6628,N_6169,N_6339);
xnor U6629 (N_6629,N_6011,N_6157);
and U6630 (N_6630,N_6304,N_6361);
nand U6631 (N_6631,N_6474,N_6402);
and U6632 (N_6632,N_6173,N_6298);
or U6633 (N_6633,N_6276,N_6170);
and U6634 (N_6634,N_6401,N_6328);
and U6635 (N_6635,N_6074,N_6354);
nor U6636 (N_6636,N_6435,N_6149);
and U6637 (N_6637,N_6210,N_6467);
nand U6638 (N_6638,N_6077,N_6136);
nor U6639 (N_6639,N_6155,N_6197);
or U6640 (N_6640,N_6295,N_6135);
xor U6641 (N_6641,N_6305,N_6008);
nor U6642 (N_6642,N_6367,N_6364);
nor U6643 (N_6643,N_6394,N_6338);
nand U6644 (N_6644,N_6186,N_6208);
nand U6645 (N_6645,N_6052,N_6499);
nand U6646 (N_6646,N_6139,N_6150);
or U6647 (N_6647,N_6203,N_6488);
nand U6648 (N_6648,N_6153,N_6352);
or U6649 (N_6649,N_6227,N_6335);
or U6650 (N_6650,N_6384,N_6204);
nand U6651 (N_6651,N_6009,N_6344);
and U6652 (N_6652,N_6000,N_6233);
or U6653 (N_6653,N_6449,N_6005);
and U6654 (N_6654,N_6062,N_6070);
and U6655 (N_6655,N_6048,N_6056);
nor U6656 (N_6656,N_6396,N_6015);
nand U6657 (N_6657,N_6469,N_6495);
nand U6658 (N_6658,N_6269,N_6046);
and U6659 (N_6659,N_6063,N_6460);
nor U6660 (N_6660,N_6024,N_6413);
nand U6661 (N_6661,N_6240,N_6236);
and U6662 (N_6662,N_6110,N_6301);
nor U6663 (N_6663,N_6137,N_6098);
nor U6664 (N_6664,N_6119,N_6066);
nor U6665 (N_6665,N_6099,N_6433);
nor U6666 (N_6666,N_6346,N_6370);
or U6667 (N_6667,N_6031,N_6041);
and U6668 (N_6668,N_6496,N_6078);
nand U6669 (N_6669,N_6441,N_6181);
nand U6670 (N_6670,N_6289,N_6285);
and U6671 (N_6671,N_6194,N_6212);
nand U6672 (N_6672,N_6171,N_6019);
nand U6673 (N_6673,N_6189,N_6082);
and U6674 (N_6674,N_6012,N_6258);
and U6675 (N_6675,N_6006,N_6281);
or U6676 (N_6676,N_6422,N_6226);
and U6677 (N_6677,N_6235,N_6428);
nand U6678 (N_6678,N_6326,N_6267);
and U6679 (N_6679,N_6168,N_6416);
or U6680 (N_6680,N_6348,N_6079);
nand U6681 (N_6681,N_6209,N_6490);
or U6682 (N_6682,N_6109,N_6291);
or U6683 (N_6683,N_6030,N_6026);
nand U6684 (N_6684,N_6274,N_6217);
nor U6685 (N_6685,N_6042,N_6393);
nor U6686 (N_6686,N_6362,N_6252);
and U6687 (N_6687,N_6392,N_6342);
xor U6688 (N_6688,N_6095,N_6059);
or U6689 (N_6689,N_6461,N_6331);
nor U6690 (N_6690,N_6206,N_6191);
and U6691 (N_6691,N_6047,N_6264);
and U6692 (N_6692,N_6261,N_6369);
xor U6693 (N_6693,N_6238,N_6034);
or U6694 (N_6694,N_6425,N_6039);
nor U6695 (N_6695,N_6297,N_6347);
and U6696 (N_6696,N_6260,N_6439);
nor U6697 (N_6697,N_6447,N_6043);
nand U6698 (N_6698,N_6164,N_6049);
nor U6699 (N_6699,N_6014,N_6255);
or U6700 (N_6700,N_6259,N_6071);
or U6701 (N_6701,N_6113,N_6096);
nand U6702 (N_6702,N_6129,N_6310);
or U6703 (N_6703,N_6254,N_6262);
or U6704 (N_6704,N_6144,N_6108);
and U6705 (N_6705,N_6431,N_6061);
nand U6706 (N_6706,N_6131,N_6076);
and U6707 (N_6707,N_6017,N_6421);
nor U6708 (N_6708,N_6035,N_6412);
or U6709 (N_6709,N_6445,N_6111);
nand U6710 (N_6710,N_6007,N_6230);
nand U6711 (N_6711,N_6470,N_6224);
nor U6712 (N_6712,N_6156,N_6327);
and U6713 (N_6713,N_6330,N_6336);
nor U6714 (N_6714,N_6175,N_6436);
nor U6715 (N_6715,N_6013,N_6130);
nor U6716 (N_6716,N_6263,N_6459);
nand U6717 (N_6717,N_6414,N_6351);
nand U6718 (N_6718,N_6028,N_6497);
nor U6719 (N_6719,N_6309,N_6385);
nand U6720 (N_6720,N_6222,N_6195);
nand U6721 (N_6721,N_6453,N_6466);
or U6722 (N_6722,N_6345,N_6184);
nand U6723 (N_6723,N_6121,N_6004);
nand U6724 (N_6724,N_6036,N_6072);
and U6725 (N_6725,N_6218,N_6316);
nor U6726 (N_6726,N_6357,N_6368);
nand U6727 (N_6727,N_6216,N_6094);
nand U6728 (N_6728,N_6027,N_6277);
or U6729 (N_6729,N_6278,N_6060);
nor U6730 (N_6730,N_6118,N_6266);
or U6731 (N_6731,N_6174,N_6315);
nor U6732 (N_6732,N_6457,N_6375);
xnor U6733 (N_6733,N_6097,N_6160);
or U6734 (N_6734,N_6232,N_6380);
nor U6735 (N_6735,N_6185,N_6128);
and U6736 (N_6736,N_6159,N_6363);
nor U6737 (N_6737,N_6475,N_6247);
nand U6738 (N_6738,N_6491,N_6083);
nand U6739 (N_6739,N_6494,N_6438);
and U6740 (N_6740,N_6116,N_6201);
or U6741 (N_6741,N_6198,N_6391);
nand U6742 (N_6742,N_6127,N_6287);
and U6743 (N_6743,N_6220,N_6268);
nand U6744 (N_6744,N_6476,N_6161);
or U6745 (N_6745,N_6300,N_6256);
nor U6746 (N_6746,N_6215,N_6312);
or U6747 (N_6747,N_6090,N_6492);
nand U6748 (N_6748,N_6324,N_6455);
and U6749 (N_6749,N_6106,N_6081);
nor U6750 (N_6750,N_6060,N_6129);
nand U6751 (N_6751,N_6160,N_6196);
nand U6752 (N_6752,N_6422,N_6482);
nand U6753 (N_6753,N_6218,N_6194);
or U6754 (N_6754,N_6275,N_6102);
and U6755 (N_6755,N_6225,N_6481);
nor U6756 (N_6756,N_6166,N_6433);
and U6757 (N_6757,N_6463,N_6205);
nor U6758 (N_6758,N_6462,N_6387);
nand U6759 (N_6759,N_6368,N_6386);
and U6760 (N_6760,N_6301,N_6457);
or U6761 (N_6761,N_6032,N_6356);
and U6762 (N_6762,N_6296,N_6285);
nand U6763 (N_6763,N_6293,N_6464);
nand U6764 (N_6764,N_6008,N_6070);
or U6765 (N_6765,N_6206,N_6066);
nand U6766 (N_6766,N_6178,N_6014);
and U6767 (N_6767,N_6052,N_6482);
or U6768 (N_6768,N_6162,N_6059);
nand U6769 (N_6769,N_6174,N_6026);
nand U6770 (N_6770,N_6177,N_6195);
nand U6771 (N_6771,N_6389,N_6360);
nor U6772 (N_6772,N_6059,N_6305);
or U6773 (N_6773,N_6198,N_6341);
nor U6774 (N_6774,N_6410,N_6070);
or U6775 (N_6775,N_6226,N_6216);
nor U6776 (N_6776,N_6355,N_6082);
and U6777 (N_6777,N_6399,N_6483);
xnor U6778 (N_6778,N_6236,N_6157);
or U6779 (N_6779,N_6488,N_6484);
nand U6780 (N_6780,N_6085,N_6416);
nor U6781 (N_6781,N_6299,N_6103);
or U6782 (N_6782,N_6042,N_6365);
nor U6783 (N_6783,N_6015,N_6327);
nand U6784 (N_6784,N_6281,N_6362);
or U6785 (N_6785,N_6020,N_6148);
and U6786 (N_6786,N_6352,N_6270);
nor U6787 (N_6787,N_6097,N_6208);
and U6788 (N_6788,N_6252,N_6275);
and U6789 (N_6789,N_6463,N_6470);
nand U6790 (N_6790,N_6128,N_6425);
nor U6791 (N_6791,N_6273,N_6438);
or U6792 (N_6792,N_6290,N_6156);
or U6793 (N_6793,N_6286,N_6499);
and U6794 (N_6794,N_6285,N_6015);
or U6795 (N_6795,N_6395,N_6220);
nand U6796 (N_6796,N_6299,N_6202);
and U6797 (N_6797,N_6134,N_6148);
xor U6798 (N_6798,N_6309,N_6231);
nand U6799 (N_6799,N_6307,N_6102);
or U6800 (N_6800,N_6264,N_6371);
nor U6801 (N_6801,N_6256,N_6311);
nor U6802 (N_6802,N_6144,N_6466);
nor U6803 (N_6803,N_6311,N_6483);
nor U6804 (N_6804,N_6490,N_6154);
nor U6805 (N_6805,N_6287,N_6276);
or U6806 (N_6806,N_6386,N_6204);
nand U6807 (N_6807,N_6072,N_6435);
or U6808 (N_6808,N_6061,N_6378);
or U6809 (N_6809,N_6049,N_6275);
or U6810 (N_6810,N_6156,N_6041);
and U6811 (N_6811,N_6483,N_6244);
and U6812 (N_6812,N_6104,N_6223);
nor U6813 (N_6813,N_6028,N_6331);
and U6814 (N_6814,N_6189,N_6083);
and U6815 (N_6815,N_6210,N_6463);
nor U6816 (N_6816,N_6456,N_6083);
or U6817 (N_6817,N_6052,N_6115);
nor U6818 (N_6818,N_6057,N_6150);
nor U6819 (N_6819,N_6223,N_6012);
and U6820 (N_6820,N_6356,N_6020);
or U6821 (N_6821,N_6054,N_6374);
nand U6822 (N_6822,N_6459,N_6098);
and U6823 (N_6823,N_6180,N_6242);
nor U6824 (N_6824,N_6228,N_6339);
or U6825 (N_6825,N_6374,N_6390);
or U6826 (N_6826,N_6436,N_6219);
nand U6827 (N_6827,N_6154,N_6250);
nor U6828 (N_6828,N_6479,N_6151);
nor U6829 (N_6829,N_6481,N_6385);
xnor U6830 (N_6830,N_6484,N_6491);
nor U6831 (N_6831,N_6105,N_6250);
or U6832 (N_6832,N_6437,N_6159);
or U6833 (N_6833,N_6413,N_6078);
nand U6834 (N_6834,N_6279,N_6234);
and U6835 (N_6835,N_6372,N_6488);
nand U6836 (N_6836,N_6407,N_6172);
nand U6837 (N_6837,N_6208,N_6115);
nor U6838 (N_6838,N_6096,N_6466);
and U6839 (N_6839,N_6285,N_6014);
nand U6840 (N_6840,N_6167,N_6159);
and U6841 (N_6841,N_6420,N_6421);
and U6842 (N_6842,N_6363,N_6069);
or U6843 (N_6843,N_6499,N_6340);
and U6844 (N_6844,N_6385,N_6390);
nand U6845 (N_6845,N_6474,N_6191);
nand U6846 (N_6846,N_6479,N_6491);
or U6847 (N_6847,N_6063,N_6036);
and U6848 (N_6848,N_6013,N_6416);
nor U6849 (N_6849,N_6334,N_6275);
nor U6850 (N_6850,N_6306,N_6165);
and U6851 (N_6851,N_6128,N_6116);
nor U6852 (N_6852,N_6169,N_6215);
and U6853 (N_6853,N_6491,N_6492);
nor U6854 (N_6854,N_6038,N_6227);
or U6855 (N_6855,N_6289,N_6104);
and U6856 (N_6856,N_6414,N_6113);
nand U6857 (N_6857,N_6341,N_6441);
xor U6858 (N_6858,N_6186,N_6147);
or U6859 (N_6859,N_6372,N_6302);
nand U6860 (N_6860,N_6218,N_6155);
nand U6861 (N_6861,N_6198,N_6218);
and U6862 (N_6862,N_6367,N_6103);
or U6863 (N_6863,N_6028,N_6222);
nand U6864 (N_6864,N_6297,N_6438);
or U6865 (N_6865,N_6110,N_6386);
nor U6866 (N_6866,N_6364,N_6051);
nand U6867 (N_6867,N_6154,N_6063);
and U6868 (N_6868,N_6388,N_6480);
and U6869 (N_6869,N_6203,N_6389);
nor U6870 (N_6870,N_6244,N_6312);
nor U6871 (N_6871,N_6042,N_6050);
nand U6872 (N_6872,N_6367,N_6029);
and U6873 (N_6873,N_6290,N_6295);
or U6874 (N_6874,N_6193,N_6362);
nand U6875 (N_6875,N_6461,N_6140);
or U6876 (N_6876,N_6457,N_6493);
nand U6877 (N_6877,N_6392,N_6455);
and U6878 (N_6878,N_6184,N_6283);
nand U6879 (N_6879,N_6493,N_6003);
nand U6880 (N_6880,N_6287,N_6371);
and U6881 (N_6881,N_6020,N_6393);
or U6882 (N_6882,N_6279,N_6172);
or U6883 (N_6883,N_6294,N_6392);
and U6884 (N_6884,N_6463,N_6339);
or U6885 (N_6885,N_6455,N_6372);
or U6886 (N_6886,N_6002,N_6321);
or U6887 (N_6887,N_6226,N_6173);
nor U6888 (N_6888,N_6144,N_6075);
and U6889 (N_6889,N_6286,N_6361);
or U6890 (N_6890,N_6126,N_6245);
or U6891 (N_6891,N_6346,N_6442);
xor U6892 (N_6892,N_6480,N_6454);
nor U6893 (N_6893,N_6150,N_6189);
and U6894 (N_6894,N_6239,N_6141);
nand U6895 (N_6895,N_6277,N_6395);
nor U6896 (N_6896,N_6453,N_6403);
nor U6897 (N_6897,N_6097,N_6054);
nor U6898 (N_6898,N_6006,N_6037);
or U6899 (N_6899,N_6226,N_6071);
and U6900 (N_6900,N_6284,N_6445);
or U6901 (N_6901,N_6207,N_6378);
or U6902 (N_6902,N_6488,N_6003);
and U6903 (N_6903,N_6475,N_6432);
xnor U6904 (N_6904,N_6422,N_6250);
nor U6905 (N_6905,N_6001,N_6460);
and U6906 (N_6906,N_6129,N_6226);
nand U6907 (N_6907,N_6210,N_6325);
nand U6908 (N_6908,N_6216,N_6187);
and U6909 (N_6909,N_6400,N_6450);
and U6910 (N_6910,N_6403,N_6048);
and U6911 (N_6911,N_6216,N_6104);
nand U6912 (N_6912,N_6354,N_6301);
nand U6913 (N_6913,N_6158,N_6079);
and U6914 (N_6914,N_6227,N_6409);
and U6915 (N_6915,N_6470,N_6259);
or U6916 (N_6916,N_6448,N_6391);
or U6917 (N_6917,N_6389,N_6386);
or U6918 (N_6918,N_6462,N_6063);
nor U6919 (N_6919,N_6428,N_6213);
nand U6920 (N_6920,N_6187,N_6284);
and U6921 (N_6921,N_6162,N_6419);
nand U6922 (N_6922,N_6211,N_6085);
nand U6923 (N_6923,N_6000,N_6327);
or U6924 (N_6924,N_6004,N_6114);
and U6925 (N_6925,N_6119,N_6140);
or U6926 (N_6926,N_6269,N_6252);
or U6927 (N_6927,N_6382,N_6483);
and U6928 (N_6928,N_6230,N_6425);
or U6929 (N_6929,N_6346,N_6467);
or U6930 (N_6930,N_6429,N_6140);
nor U6931 (N_6931,N_6000,N_6010);
and U6932 (N_6932,N_6277,N_6012);
nand U6933 (N_6933,N_6331,N_6413);
or U6934 (N_6934,N_6436,N_6402);
nand U6935 (N_6935,N_6252,N_6022);
or U6936 (N_6936,N_6399,N_6087);
nand U6937 (N_6937,N_6056,N_6185);
nand U6938 (N_6938,N_6164,N_6254);
and U6939 (N_6939,N_6409,N_6370);
or U6940 (N_6940,N_6355,N_6169);
and U6941 (N_6941,N_6400,N_6204);
or U6942 (N_6942,N_6036,N_6044);
and U6943 (N_6943,N_6048,N_6025);
and U6944 (N_6944,N_6277,N_6205);
or U6945 (N_6945,N_6105,N_6364);
nor U6946 (N_6946,N_6440,N_6429);
or U6947 (N_6947,N_6167,N_6032);
nor U6948 (N_6948,N_6018,N_6428);
or U6949 (N_6949,N_6070,N_6253);
and U6950 (N_6950,N_6374,N_6497);
and U6951 (N_6951,N_6475,N_6036);
nor U6952 (N_6952,N_6439,N_6233);
and U6953 (N_6953,N_6291,N_6366);
nor U6954 (N_6954,N_6455,N_6468);
nor U6955 (N_6955,N_6160,N_6433);
nor U6956 (N_6956,N_6055,N_6212);
and U6957 (N_6957,N_6186,N_6334);
nand U6958 (N_6958,N_6000,N_6146);
or U6959 (N_6959,N_6152,N_6396);
nor U6960 (N_6960,N_6030,N_6050);
or U6961 (N_6961,N_6322,N_6467);
nand U6962 (N_6962,N_6089,N_6323);
nor U6963 (N_6963,N_6328,N_6206);
nand U6964 (N_6964,N_6015,N_6280);
nor U6965 (N_6965,N_6485,N_6349);
or U6966 (N_6966,N_6153,N_6096);
xor U6967 (N_6967,N_6018,N_6164);
and U6968 (N_6968,N_6365,N_6482);
nand U6969 (N_6969,N_6459,N_6032);
or U6970 (N_6970,N_6426,N_6317);
and U6971 (N_6971,N_6256,N_6074);
xor U6972 (N_6972,N_6292,N_6280);
and U6973 (N_6973,N_6498,N_6256);
nor U6974 (N_6974,N_6285,N_6207);
and U6975 (N_6975,N_6058,N_6389);
nand U6976 (N_6976,N_6159,N_6205);
nor U6977 (N_6977,N_6396,N_6465);
nor U6978 (N_6978,N_6359,N_6395);
nor U6979 (N_6979,N_6044,N_6419);
and U6980 (N_6980,N_6416,N_6375);
nand U6981 (N_6981,N_6006,N_6029);
or U6982 (N_6982,N_6115,N_6092);
nor U6983 (N_6983,N_6161,N_6174);
nand U6984 (N_6984,N_6083,N_6063);
nor U6985 (N_6985,N_6483,N_6045);
nand U6986 (N_6986,N_6146,N_6176);
nand U6987 (N_6987,N_6004,N_6290);
or U6988 (N_6988,N_6486,N_6353);
nand U6989 (N_6989,N_6208,N_6041);
and U6990 (N_6990,N_6041,N_6422);
nor U6991 (N_6991,N_6083,N_6413);
nand U6992 (N_6992,N_6013,N_6156);
or U6993 (N_6993,N_6128,N_6452);
or U6994 (N_6994,N_6025,N_6430);
nand U6995 (N_6995,N_6140,N_6351);
nand U6996 (N_6996,N_6088,N_6343);
nand U6997 (N_6997,N_6077,N_6153);
nor U6998 (N_6998,N_6347,N_6058);
or U6999 (N_6999,N_6349,N_6112);
and U7000 (N_7000,N_6571,N_6564);
or U7001 (N_7001,N_6990,N_6609);
nor U7002 (N_7002,N_6755,N_6854);
and U7003 (N_7003,N_6579,N_6934);
nand U7004 (N_7004,N_6667,N_6615);
and U7005 (N_7005,N_6610,N_6563);
and U7006 (N_7006,N_6668,N_6617);
or U7007 (N_7007,N_6820,N_6558);
nand U7008 (N_7008,N_6989,N_6559);
nand U7009 (N_7009,N_6605,N_6687);
nor U7010 (N_7010,N_6987,N_6601);
nor U7011 (N_7011,N_6731,N_6603);
nor U7012 (N_7012,N_6707,N_6500);
and U7013 (N_7013,N_6710,N_6676);
and U7014 (N_7014,N_6748,N_6672);
xnor U7015 (N_7015,N_6588,N_6914);
or U7016 (N_7016,N_6915,N_6646);
or U7017 (N_7017,N_6518,N_6907);
or U7018 (N_7018,N_6575,N_6850);
or U7019 (N_7019,N_6507,N_6639);
and U7020 (N_7020,N_6726,N_6597);
and U7021 (N_7021,N_6911,N_6691);
or U7022 (N_7022,N_6595,N_6832);
nand U7023 (N_7023,N_6774,N_6883);
or U7024 (N_7024,N_6930,N_6730);
nand U7025 (N_7025,N_6951,N_6947);
and U7026 (N_7026,N_6943,N_6742);
or U7027 (N_7027,N_6577,N_6538);
or U7028 (N_7028,N_6621,N_6815);
nor U7029 (N_7029,N_6512,N_6517);
and U7030 (N_7030,N_6897,N_6771);
nand U7031 (N_7031,N_6949,N_6878);
and U7032 (N_7032,N_6808,N_6953);
nand U7033 (N_7033,N_6890,N_6527);
or U7034 (N_7034,N_6873,N_6945);
nand U7035 (N_7035,N_6670,N_6806);
nor U7036 (N_7036,N_6862,N_6846);
and U7037 (N_7037,N_6524,N_6939);
nand U7038 (N_7038,N_6932,N_6838);
and U7039 (N_7039,N_6598,N_6789);
nor U7040 (N_7040,N_6999,N_6860);
nand U7041 (N_7041,N_6810,N_6938);
or U7042 (N_7042,N_6622,N_6582);
or U7043 (N_7043,N_6965,N_6940);
or U7044 (N_7044,N_6887,N_6505);
and U7045 (N_7045,N_6535,N_6809);
nor U7046 (N_7046,N_6991,N_6828);
nor U7047 (N_7047,N_6787,N_6712);
nor U7048 (N_7048,N_6711,N_6766);
nor U7049 (N_7049,N_6544,N_6585);
nand U7050 (N_7050,N_6813,N_6851);
nand U7051 (N_7051,N_6560,N_6665);
and U7052 (N_7052,N_6642,N_6977);
or U7053 (N_7053,N_6664,N_6791);
or U7054 (N_7054,N_6529,N_6592);
nor U7055 (N_7055,N_6904,N_6863);
or U7056 (N_7056,N_6916,N_6894);
or U7057 (N_7057,N_6929,N_6866);
and U7058 (N_7058,N_6636,N_6542);
nand U7059 (N_7059,N_6754,N_6761);
and U7060 (N_7060,N_6960,N_6650);
nor U7061 (N_7061,N_6533,N_6669);
or U7062 (N_7062,N_6777,N_6974);
or U7063 (N_7063,N_6578,N_6912);
nor U7064 (N_7064,N_6825,N_6853);
nor U7065 (N_7065,N_6632,N_6752);
nor U7066 (N_7066,N_6537,N_6798);
nor U7067 (N_7067,N_6674,N_6756);
nand U7068 (N_7068,N_6901,N_6782);
nor U7069 (N_7069,N_6709,N_6562);
or U7070 (N_7070,N_6841,N_6555);
or U7071 (N_7071,N_6843,N_6995);
nor U7072 (N_7072,N_6986,N_6623);
nand U7073 (N_7073,N_6652,N_6703);
and U7074 (N_7074,N_6746,N_6685);
nor U7075 (N_7075,N_6727,N_6784);
nor U7076 (N_7076,N_6768,N_6513);
and U7077 (N_7077,N_6701,N_6865);
nor U7078 (N_7078,N_6587,N_6928);
and U7079 (N_7079,N_6658,N_6614);
or U7080 (N_7080,N_6902,N_6735);
nand U7081 (N_7081,N_6565,N_6600);
and U7082 (N_7082,N_6728,N_6879);
or U7083 (N_7083,N_6681,N_6881);
and U7084 (N_7084,N_6637,N_6504);
nand U7085 (N_7085,N_6647,N_6633);
or U7086 (N_7086,N_6998,N_6526);
or U7087 (N_7087,N_6796,N_6590);
nand U7088 (N_7088,N_6516,N_6747);
and U7089 (N_7089,N_6606,N_6856);
nand U7090 (N_7090,N_6830,N_6584);
nand U7091 (N_7091,N_6839,N_6522);
nor U7092 (N_7092,N_6935,N_6797);
and U7093 (N_7093,N_6635,N_6968);
or U7094 (N_7094,N_6973,N_6908);
or U7095 (N_7095,N_6762,N_6539);
nor U7096 (N_7096,N_6591,N_6552);
and U7097 (N_7097,N_6985,N_6740);
nand U7098 (N_7098,N_6741,N_6611);
nand U7099 (N_7099,N_6607,N_6714);
nor U7100 (N_7100,N_6697,N_6675);
nand U7101 (N_7101,N_6634,N_6534);
and U7102 (N_7102,N_6984,N_6899);
nor U7103 (N_7103,N_6586,N_6790);
nand U7104 (N_7104,N_6630,N_6952);
nor U7105 (N_7105,N_6720,N_6765);
or U7106 (N_7106,N_6905,N_6624);
and U7107 (N_7107,N_6566,N_6868);
and U7108 (N_7108,N_6918,N_6925);
and U7109 (N_7109,N_6982,N_6895);
nand U7110 (N_7110,N_6981,N_6959);
nor U7111 (N_7111,N_6817,N_6657);
and U7112 (N_7112,N_6931,N_6716);
and U7113 (N_7113,N_6706,N_6785);
nand U7114 (N_7114,N_6722,N_6645);
and U7115 (N_7115,N_6975,N_6718);
and U7116 (N_7116,N_6869,N_6547);
nor U7117 (N_7117,N_6719,N_6961);
nor U7118 (N_7118,N_6779,N_6698);
nor U7119 (N_7119,N_6807,N_6957);
nor U7120 (N_7120,N_6677,N_6690);
or U7121 (N_7121,N_6996,N_6508);
nor U7122 (N_7122,N_6651,N_6704);
and U7123 (N_7123,N_6780,N_6858);
or U7124 (N_7124,N_6955,N_6909);
and U7125 (N_7125,N_6962,N_6644);
and U7126 (N_7126,N_6653,N_6772);
or U7127 (N_7127,N_6760,N_6655);
nor U7128 (N_7128,N_6778,N_6978);
nor U7129 (N_7129,N_6919,N_6723);
or U7130 (N_7130,N_6786,N_6800);
and U7131 (N_7131,N_6910,N_6845);
nand U7132 (N_7132,N_6745,N_6572);
or U7133 (N_7133,N_6525,N_6662);
or U7134 (N_7134,N_6521,N_6568);
or U7135 (N_7135,N_6979,N_6835);
nor U7136 (N_7136,N_6549,N_6725);
nand U7137 (N_7137,N_6656,N_6570);
and U7138 (N_7138,N_6971,N_6849);
and U7139 (N_7139,N_6581,N_6898);
nor U7140 (N_7140,N_6573,N_6666);
and U7141 (N_7141,N_6802,N_6738);
and U7142 (N_7142,N_6744,N_6649);
and U7143 (N_7143,N_6702,N_6805);
nor U7144 (N_7144,N_6926,N_6792);
nor U7145 (N_7145,N_6861,N_6734);
nand U7146 (N_7146,N_6576,N_6814);
and U7147 (N_7147,N_6801,N_6659);
or U7148 (N_7148,N_6503,N_6885);
xor U7149 (N_7149,N_6888,N_6988);
or U7150 (N_7150,N_6859,N_6520);
and U7151 (N_7151,N_6750,N_6942);
nor U7152 (N_7152,N_6705,N_6874);
nor U7153 (N_7153,N_6794,N_6678);
and U7154 (N_7154,N_6751,N_6688);
and U7155 (N_7155,N_6580,N_6821);
and U7156 (N_7156,N_6654,N_6506);
or U7157 (N_7157,N_6546,N_6620);
nor U7158 (N_7158,N_6837,N_6826);
nand U7159 (N_7159,N_6773,N_6956);
nand U7160 (N_7160,N_6502,N_6767);
or U7161 (N_7161,N_6557,N_6848);
nor U7162 (N_7162,N_6561,N_6950);
nor U7163 (N_7163,N_6689,N_6827);
and U7164 (N_7164,N_6671,N_6640);
nand U7165 (N_7165,N_6924,N_6550);
and U7166 (N_7166,N_6680,N_6864);
nand U7167 (N_7167,N_6855,N_6927);
or U7168 (N_7168,N_6663,N_6625);
or U7169 (N_7169,N_6872,N_6840);
and U7170 (N_7170,N_6770,N_6531);
nor U7171 (N_7171,N_6834,N_6913);
and U7172 (N_7172,N_6695,N_6892);
and U7173 (N_7173,N_6569,N_6692);
nor U7174 (N_7174,N_6842,N_6966);
or U7175 (N_7175,N_6641,N_6889);
nor U7176 (N_7176,N_6867,N_6548);
nand U7177 (N_7177,N_6759,N_6886);
nand U7178 (N_7178,N_6847,N_6583);
and U7179 (N_7179,N_6992,N_6937);
and U7180 (N_7180,N_6963,N_6660);
nand U7181 (N_7181,N_6501,N_6857);
nand U7182 (N_7182,N_6509,N_6593);
and U7183 (N_7183,N_6922,N_6661);
and U7184 (N_7184,N_6696,N_6523);
and U7185 (N_7185,N_6763,N_6733);
xor U7186 (N_7186,N_6682,N_6540);
nor U7187 (N_7187,N_6638,N_6969);
or U7188 (N_7188,N_6612,N_6749);
nand U7189 (N_7189,N_6967,N_6684);
nor U7190 (N_7190,N_6994,N_6941);
nand U7191 (N_7191,N_6515,N_6627);
and U7192 (N_7192,N_6876,N_6831);
or U7193 (N_7193,N_6877,N_6764);
nor U7194 (N_7194,N_6532,N_6954);
and U7195 (N_7195,N_6514,N_6844);
and U7196 (N_7196,N_6788,N_6753);
or U7197 (N_7197,N_6739,N_6970);
nor U7198 (N_7198,N_6713,N_6519);
nand U7199 (N_7199,N_6643,N_6729);
xor U7200 (N_7200,N_6958,N_6781);
nor U7201 (N_7201,N_6554,N_6743);
nand U7202 (N_7202,N_6948,N_6896);
nand U7203 (N_7203,N_6510,N_6804);
nand U7204 (N_7204,N_6604,N_6757);
and U7205 (N_7205,N_6946,N_6811);
nor U7206 (N_7206,N_6818,N_6545);
or U7207 (N_7207,N_6983,N_6699);
xor U7208 (N_7208,N_6708,N_6944);
nor U7209 (N_7209,N_6819,N_6921);
nand U7210 (N_7210,N_6602,N_6700);
nand U7211 (N_7211,N_6616,N_6721);
and U7212 (N_7212,N_6769,N_6776);
nand U7213 (N_7213,N_6528,N_6822);
or U7214 (N_7214,N_6833,N_6715);
or U7215 (N_7215,N_6906,N_6619);
and U7216 (N_7216,N_6875,N_6823);
nor U7217 (N_7217,N_6732,N_6511);
and U7218 (N_7218,N_6836,N_6758);
nand U7219 (N_7219,N_6972,N_6829);
or U7220 (N_7220,N_6824,N_6936);
or U7221 (N_7221,N_6795,N_6693);
or U7222 (N_7222,N_6686,N_6553);
or U7223 (N_7223,N_6629,N_6536);
nand U7224 (N_7224,N_6717,N_6631);
and U7225 (N_7225,N_6736,N_6980);
nand U7226 (N_7226,N_6997,N_6923);
or U7227 (N_7227,N_6920,N_6530);
or U7228 (N_7228,N_6993,N_6683);
nand U7229 (N_7229,N_6812,N_6903);
xnor U7230 (N_7230,N_6880,N_6673);
nand U7231 (N_7231,N_6933,N_6599);
and U7232 (N_7232,N_6917,N_6589);
nor U7233 (N_7233,N_6543,N_6882);
and U7234 (N_7234,N_6541,N_6793);
xor U7235 (N_7235,N_6799,N_6574);
and U7236 (N_7236,N_6556,N_6618);
nand U7237 (N_7237,N_6884,N_6613);
or U7238 (N_7238,N_6964,N_6871);
nor U7239 (N_7239,N_6775,N_6628);
or U7240 (N_7240,N_6648,N_6596);
nand U7241 (N_7241,N_6737,N_6852);
nor U7242 (N_7242,N_6803,N_6694);
nand U7243 (N_7243,N_6567,N_6893);
or U7244 (N_7244,N_6783,N_6594);
nand U7245 (N_7245,N_6976,N_6891);
nor U7246 (N_7246,N_6608,N_6870);
nor U7247 (N_7247,N_6679,N_6816);
and U7248 (N_7248,N_6626,N_6551);
and U7249 (N_7249,N_6724,N_6900);
or U7250 (N_7250,N_6578,N_6525);
nor U7251 (N_7251,N_6755,N_6859);
nand U7252 (N_7252,N_6973,N_6626);
or U7253 (N_7253,N_6977,N_6867);
or U7254 (N_7254,N_6521,N_6941);
xnor U7255 (N_7255,N_6523,N_6838);
nand U7256 (N_7256,N_6940,N_6703);
nand U7257 (N_7257,N_6573,N_6534);
and U7258 (N_7258,N_6546,N_6930);
nor U7259 (N_7259,N_6962,N_6508);
nor U7260 (N_7260,N_6837,N_6617);
xnor U7261 (N_7261,N_6928,N_6709);
or U7262 (N_7262,N_6615,N_6866);
nand U7263 (N_7263,N_6674,N_6997);
or U7264 (N_7264,N_6654,N_6697);
nand U7265 (N_7265,N_6711,N_6902);
nand U7266 (N_7266,N_6594,N_6839);
or U7267 (N_7267,N_6696,N_6861);
and U7268 (N_7268,N_6873,N_6741);
xor U7269 (N_7269,N_6847,N_6648);
nor U7270 (N_7270,N_6880,N_6793);
nand U7271 (N_7271,N_6516,N_6869);
nor U7272 (N_7272,N_6530,N_6592);
and U7273 (N_7273,N_6789,N_6997);
nand U7274 (N_7274,N_6568,N_6911);
nor U7275 (N_7275,N_6782,N_6851);
xor U7276 (N_7276,N_6834,N_6756);
nand U7277 (N_7277,N_6807,N_6546);
nand U7278 (N_7278,N_6648,N_6557);
and U7279 (N_7279,N_6987,N_6534);
nor U7280 (N_7280,N_6677,N_6502);
nor U7281 (N_7281,N_6844,N_6795);
or U7282 (N_7282,N_6669,N_6821);
and U7283 (N_7283,N_6691,N_6842);
and U7284 (N_7284,N_6932,N_6907);
and U7285 (N_7285,N_6863,N_6531);
nand U7286 (N_7286,N_6676,N_6905);
nand U7287 (N_7287,N_6614,N_6738);
nand U7288 (N_7288,N_6928,N_6573);
nor U7289 (N_7289,N_6859,N_6642);
nor U7290 (N_7290,N_6864,N_6500);
or U7291 (N_7291,N_6984,N_6705);
and U7292 (N_7292,N_6590,N_6826);
or U7293 (N_7293,N_6543,N_6819);
and U7294 (N_7294,N_6742,N_6712);
nand U7295 (N_7295,N_6849,N_6944);
nand U7296 (N_7296,N_6630,N_6789);
or U7297 (N_7297,N_6898,N_6981);
nor U7298 (N_7298,N_6539,N_6821);
or U7299 (N_7299,N_6714,N_6908);
or U7300 (N_7300,N_6561,N_6771);
or U7301 (N_7301,N_6972,N_6614);
nand U7302 (N_7302,N_6669,N_6841);
nor U7303 (N_7303,N_6977,N_6561);
or U7304 (N_7304,N_6912,N_6628);
and U7305 (N_7305,N_6632,N_6562);
and U7306 (N_7306,N_6699,N_6856);
nor U7307 (N_7307,N_6743,N_6884);
or U7308 (N_7308,N_6624,N_6645);
or U7309 (N_7309,N_6971,N_6685);
or U7310 (N_7310,N_6672,N_6626);
and U7311 (N_7311,N_6889,N_6721);
xor U7312 (N_7312,N_6744,N_6794);
and U7313 (N_7313,N_6640,N_6616);
or U7314 (N_7314,N_6655,N_6958);
nand U7315 (N_7315,N_6845,N_6626);
and U7316 (N_7316,N_6551,N_6778);
or U7317 (N_7317,N_6811,N_6994);
or U7318 (N_7318,N_6841,N_6553);
or U7319 (N_7319,N_6677,N_6816);
or U7320 (N_7320,N_6730,N_6775);
or U7321 (N_7321,N_6517,N_6865);
nor U7322 (N_7322,N_6984,N_6571);
and U7323 (N_7323,N_6686,N_6810);
nor U7324 (N_7324,N_6678,N_6765);
or U7325 (N_7325,N_6841,N_6739);
and U7326 (N_7326,N_6593,N_6938);
and U7327 (N_7327,N_6570,N_6580);
and U7328 (N_7328,N_6797,N_6663);
nor U7329 (N_7329,N_6611,N_6663);
nand U7330 (N_7330,N_6846,N_6818);
and U7331 (N_7331,N_6927,N_6916);
and U7332 (N_7332,N_6753,N_6743);
nor U7333 (N_7333,N_6699,N_6576);
nor U7334 (N_7334,N_6533,N_6997);
nor U7335 (N_7335,N_6945,N_6880);
nor U7336 (N_7336,N_6832,N_6579);
nor U7337 (N_7337,N_6787,N_6933);
and U7338 (N_7338,N_6871,N_6550);
nor U7339 (N_7339,N_6594,N_6502);
and U7340 (N_7340,N_6606,N_6890);
nand U7341 (N_7341,N_6936,N_6702);
nand U7342 (N_7342,N_6920,N_6932);
nand U7343 (N_7343,N_6960,N_6840);
or U7344 (N_7344,N_6826,N_6908);
nand U7345 (N_7345,N_6614,N_6999);
or U7346 (N_7346,N_6690,N_6841);
or U7347 (N_7347,N_6588,N_6693);
nand U7348 (N_7348,N_6506,N_6847);
and U7349 (N_7349,N_6571,N_6730);
nand U7350 (N_7350,N_6798,N_6752);
nand U7351 (N_7351,N_6535,N_6845);
and U7352 (N_7352,N_6574,N_6621);
or U7353 (N_7353,N_6510,N_6695);
and U7354 (N_7354,N_6971,N_6794);
nand U7355 (N_7355,N_6915,N_6692);
nand U7356 (N_7356,N_6777,N_6867);
nand U7357 (N_7357,N_6842,N_6879);
nor U7358 (N_7358,N_6843,N_6511);
nor U7359 (N_7359,N_6929,N_6740);
nand U7360 (N_7360,N_6515,N_6992);
or U7361 (N_7361,N_6853,N_6559);
and U7362 (N_7362,N_6735,N_6805);
and U7363 (N_7363,N_6770,N_6591);
and U7364 (N_7364,N_6891,N_6836);
or U7365 (N_7365,N_6895,N_6586);
nand U7366 (N_7366,N_6568,N_6556);
nor U7367 (N_7367,N_6864,N_6781);
nor U7368 (N_7368,N_6681,N_6856);
nand U7369 (N_7369,N_6856,N_6916);
nor U7370 (N_7370,N_6520,N_6878);
and U7371 (N_7371,N_6883,N_6978);
nand U7372 (N_7372,N_6853,N_6528);
and U7373 (N_7373,N_6566,N_6857);
or U7374 (N_7374,N_6537,N_6746);
and U7375 (N_7375,N_6796,N_6560);
and U7376 (N_7376,N_6832,N_6625);
and U7377 (N_7377,N_6729,N_6648);
and U7378 (N_7378,N_6816,N_6564);
and U7379 (N_7379,N_6975,N_6941);
and U7380 (N_7380,N_6850,N_6811);
or U7381 (N_7381,N_6620,N_6596);
nand U7382 (N_7382,N_6576,N_6579);
nand U7383 (N_7383,N_6557,N_6512);
or U7384 (N_7384,N_6595,N_6528);
nand U7385 (N_7385,N_6625,N_6837);
and U7386 (N_7386,N_6663,N_6689);
nand U7387 (N_7387,N_6708,N_6929);
nor U7388 (N_7388,N_6551,N_6912);
and U7389 (N_7389,N_6946,N_6692);
or U7390 (N_7390,N_6810,N_6805);
xnor U7391 (N_7391,N_6794,N_6637);
or U7392 (N_7392,N_6990,N_6805);
and U7393 (N_7393,N_6967,N_6769);
nor U7394 (N_7394,N_6631,N_6653);
nor U7395 (N_7395,N_6613,N_6677);
nor U7396 (N_7396,N_6660,N_6621);
and U7397 (N_7397,N_6519,N_6866);
or U7398 (N_7398,N_6599,N_6847);
nor U7399 (N_7399,N_6821,N_6607);
and U7400 (N_7400,N_6513,N_6997);
and U7401 (N_7401,N_6801,N_6631);
or U7402 (N_7402,N_6958,N_6721);
or U7403 (N_7403,N_6685,N_6875);
nand U7404 (N_7404,N_6654,N_6544);
nor U7405 (N_7405,N_6541,N_6995);
nand U7406 (N_7406,N_6722,N_6508);
or U7407 (N_7407,N_6608,N_6542);
and U7408 (N_7408,N_6669,N_6891);
nor U7409 (N_7409,N_6535,N_6713);
nor U7410 (N_7410,N_6525,N_6666);
nor U7411 (N_7411,N_6607,N_6536);
and U7412 (N_7412,N_6588,N_6713);
nor U7413 (N_7413,N_6664,N_6518);
nand U7414 (N_7414,N_6688,N_6944);
or U7415 (N_7415,N_6986,N_6535);
xnor U7416 (N_7416,N_6561,N_6547);
nor U7417 (N_7417,N_6671,N_6655);
and U7418 (N_7418,N_6508,N_6914);
nand U7419 (N_7419,N_6981,N_6634);
nor U7420 (N_7420,N_6548,N_6960);
nand U7421 (N_7421,N_6840,N_6539);
and U7422 (N_7422,N_6995,N_6953);
nand U7423 (N_7423,N_6649,N_6714);
nor U7424 (N_7424,N_6825,N_6863);
or U7425 (N_7425,N_6512,N_6958);
nor U7426 (N_7426,N_6891,N_6647);
and U7427 (N_7427,N_6500,N_6523);
nand U7428 (N_7428,N_6871,N_6958);
or U7429 (N_7429,N_6998,N_6700);
nor U7430 (N_7430,N_6562,N_6970);
nor U7431 (N_7431,N_6933,N_6658);
nor U7432 (N_7432,N_6855,N_6759);
or U7433 (N_7433,N_6593,N_6780);
and U7434 (N_7434,N_6618,N_6577);
nand U7435 (N_7435,N_6679,N_6672);
nand U7436 (N_7436,N_6535,N_6769);
nand U7437 (N_7437,N_6899,N_6634);
nor U7438 (N_7438,N_6825,N_6583);
and U7439 (N_7439,N_6996,N_6624);
nand U7440 (N_7440,N_6967,N_6626);
or U7441 (N_7441,N_6512,N_6666);
nor U7442 (N_7442,N_6873,N_6917);
nor U7443 (N_7443,N_6559,N_6578);
or U7444 (N_7444,N_6637,N_6508);
and U7445 (N_7445,N_6719,N_6559);
or U7446 (N_7446,N_6688,N_6625);
or U7447 (N_7447,N_6639,N_6609);
nor U7448 (N_7448,N_6642,N_6543);
and U7449 (N_7449,N_6878,N_6923);
nand U7450 (N_7450,N_6517,N_6762);
nor U7451 (N_7451,N_6589,N_6791);
nor U7452 (N_7452,N_6579,N_6782);
or U7453 (N_7453,N_6958,N_6929);
and U7454 (N_7454,N_6963,N_6668);
and U7455 (N_7455,N_6759,N_6535);
nand U7456 (N_7456,N_6757,N_6559);
nand U7457 (N_7457,N_6702,N_6983);
nand U7458 (N_7458,N_6798,N_6674);
nor U7459 (N_7459,N_6976,N_6989);
and U7460 (N_7460,N_6956,N_6693);
nand U7461 (N_7461,N_6740,N_6730);
and U7462 (N_7462,N_6572,N_6909);
or U7463 (N_7463,N_6871,N_6859);
or U7464 (N_7464,N_6722,N_6706);
xnor U7465 (N_7465,N_6896,N_6789);
or U7466 (N_7466,N_6882,N_6601);
and U7467 (N_7467,N_6793,N_6549);
nand U7468 (N_7468,N_6712,N_6854);
xnor U7469 (N_7469,N_6602,N_6657);
nor U7470 (N_7470,N_6996,N_6946);
nor U7471 (N_7471,N_6694,N_6985);
or U7472 (N_7472,N_6722,N_6768);
or U7473 (N_7473,N_6687,N_6612);
nor U7474 (N_7474,N_6644,N_6702);
nand U7475 (N_7475,N_6704,N_6693);
and U7476 (N_7476,N_6987,N_6684);
or U7477 (N_7477,N_6900,N_6828);
and U7478 (N_7478,N_6577,N_6787);
or U7479 (N_7479,N_6724,N_6782);
nor U7480 (N_7480,N_6917,N_6753);
nor U7481 (N_7481,N_6839,N_6599);
xor U7482 (N_7482,N_6573,N_6720);
and U7483 (N_7483,N_6948,N_6842);
and U7484 (N_7484,N_6939,N_6608);
nand U7485 (N_7485,N_6848,N_6734);
or U7486 (N_7486,N_6744,N_6928);
or U7487 (N_7487,N_6550,N_6735);
or U7488 (N_7488,N_6872,N_6557);
nor U7489 (N_7489,N_6504,N_6883);
xor U7490 (N_7490,N_6749,N_6989);
nor U7491 (N_7491,N_6803,N_6673);
or U7492 (N_7492,N_6557,N_6715);
nand U7493 (N_7493,N_6729,N_6798);
nor U7494 (N_7494,N_6519,N_6504);
nand U7495 (N_7495,N_6614,N_6750);
or U7496 (N_7496,N_6562,N_6602);
nand U7497 (N_7497,N_6906,N_6931);
nand U7498 (N_7498,N_6590,N_6848);
nor U7499 (N_7499,N_6913,N_6962);
and U7500 (N_7500,N_7208,N_7419);
or U7501 (N_7501,N_7036,N_7453);
or U7502 (N_7502,N_7213,N_7214);
nor U7503 (N_7503,N_7312,N_7079);
nor U7504 (N_7504,N_7329,N_7115);
and U7505 (N_7505,N_7047,N_7318);
or U7506 (N_7506,N_7444,N_7072);
nand U7507 (N_7507,N_7090,N_7068);
nor U7508 (N_7508,N_7161,N_7244);
and U7509 (N_7509,N_7305,N_7059);
or U7510 (N_7510,N_7249,N_7424);
nor U7511 (N_7511,N_7000,N_7468);
nor U7512 (N_7512,N_7186,N_7466);
nand U7513 (N_7513,N_7357,N_7374);
nand U7514 (N_7514,N_7464,N_7232);
and U7515 (N_7515,N_7053,N_7015);
and U7516 (N_7516,N_7099,N_7471);
nand U7517 (N_7517,N_7302,N_7494);
or U7518 (N_7518,N_7369,N_7029);
or U7519 (N_7519,N_7486,N_7288);
nand U7520 (N_7520,N_7070,N_7485);
and U7521 (N_7521,N_7060,N_7028);
nor U7522 (N_7522,N_7102,N_7146);
or U7523 (N_7523,N_7103,N_7283);
or U7524 (N_7524,N_7414,N_7465);
and U7525 (N_7525,N_7174,N_7258);
or U7526 (N_7526,N_7474,N_7076);
or U7527 (N_7527,N_7257,N_7215);
nand U7528 (N_7528,N_7135,N_7452);
or U7529 (N_7529,N_7091,N_7206);
or U7530 (N_7530,N_7181,N_7341);
xor U7531 (N_7531,N_7024,N_7347);
or U7532 (N_7532,N_7114,N_7477);
or U7533 (N_7533,N_7385,N_7293);
and U7534 (N_7534,N_7432,N_7198);
and U7535 (N_7535,N_7360,N_7346);
or U7536 (N_7536,N_7314,N_7254);
nor U7537 (N_7537,N_7250,N_7247);
nand U7538 (N_7538,N_7204,N_7307);
and U7539 (N_7539,N_7025,N_7016);
nor U7540 (N_7540,N_7140,N_7380);
or U7541 (N_7541,N_7132,N_7119);
or U7542 (N_7542,N_7363,N_7163);
or U7543 (N_7543,N_7252,N_7229);
or U7544 (N_7544,N_7101,N_7006);
or U7545 (N_7545,N_7106,N_7231);
nor U7546 (N_7546,N_7027,N_7441);
or U7547 (N_7547,N_7343,N_7075);
and U7548 (N_7548,N_7086,N_7460);
and U7549 (N_7549,N_7221,N_7150);
nor U7550 (N_7550,N_7165,N_7224);
nor U7551 (N_7551,N_7100,N_7001);
nand U7552 (N_7552,N_7040,N_7497);
and U7553 (N_7553,N_7118,N_7488);
and U7554 (N_7554,N_7223,N_7131);
and U7555 (N_7555,N_7473,N_7290);
or U7556 (N_7556,N_7183,N_7317);
nand U7557 (N_7557,N_7005,N_7331);
nand U7558 (N_7558,N_7242,N_7160);
xor U7559 (N_7559,N_7203,N_7484);
xor U7560 (N_7560,N_7097,N_7058);
and U7561 (N_7561,N_7342,N_7406);
and U7562 (N_7562,N_7299,N_7435);
nand U7563 (N_7563,N_7201,N_7173);
nand U7564 (N_7564,N_7442,N_7427);
nor U7565 (N_7565,N_7169,N_7194);
nand U7566 (N_7566,N_7462,N_7145);
and U7567 (N_7567,N_7216,N_7467);
nand U7568 (N_7568,N_7316,N_7308);
nor U7569 (N_7569,N_7272,N_7275);
nand U7570 (N_7570,N_7378,N_7260);
nand U7571 (N_7571,N_7255,N_7478);
nor U7572 (N_7572,N_7049,N_7123);
nand U7573 (N_7573,N_7425,N_7124);
nor U7574 (N_7574,N_7413,N_7407);
and U7575 (N_7575,N_7062,N_7356);
or U7576 (N_7576,N_7322,N_7368);
nand U7577 (N_7577,N_7311,N_7315);
nor U7578 (N_7578,N_7271,N_7041);
nor U7579 (N_7579,N_7365,N_7212);
and U7580 (N_7580,N_7210,N_7021);
nand U7581 (N_7581,N_7192,N_7039);
and U7582 (N_7582,N_7134,N_7243);
nor U7583 (N_7583,N_7143,N_7248);
or U7584 (N_7584,N_7129,N_7415);
nand U7585 (N_7585,N_7202,N_7093);
xor U7586 (N_7586,N_7426,N_7164);
or U7587 (N_7587,N_7321,N_7351);
nand U7588 (N_7588,N_7045,N_7375);
and U7589 (N_7589,N_7285,N_7189);
or U7590 (N_7590,N_7050,N_7328);
nand U7591 (N_7591,N_7463,N_7089);
or U7592 (N_7592,N_7377,N_7267);
or U7593 (N_7593,N_7239,N_7037);
and U7594 (N_7594,N_7402,N_7372);
or U7595 (N_7595,N_7176,N_7107);
nor U7596 (N_7596,N_7226,N_7480);
or U7597 (N_7597,N_7482,N_7352);
nor U7598 (N_7598,N_7423,N_7383);
and U7599 (N_7599,N_7324,N_7297);
or U7600 (N_7600,N_7392,N_7491);
nand U7601 (N_7601,N_7187,N_7227);
and U7602 (N_7602,N_7168,N_7038);
or U7603 (N_7603,N_7437,N_7273);
nand U7604 (N_7604,N_7067,N_7044);
or U7605 (N_7605,N_7069,N_7220);
and U7606 (N_7606,N_7270,N_7004);
nand U7607 (N_7607,N_7136,N_7063);
and U7608 (N_7608,N_7191,N_7085);
nand U7609 (N_7609,N_7125,N_7055);
nand U7610 (N_7610,N_7457,N_7128);
or U7611 (N_7611,N_7498,N_7219);
or U7612 (N_7612,N_7420,N_7188);
nor U7613 (N_7613,N_7370,N_7459);
and U7614 (N_7614,N_7338,N_7389);
nand U7615 (N_7615,N_7263,N_7117);
and U7616 (N_7616,N_7278,N_7417);
nor U7617 (N_7617,N_7153,N_7019);
or U7618 (N_7618,N_7083,N_7003);
nor U7619 (N_7619,N_7008,N_7111);
or U7620 (N_7620,N_7366,N_7151);
nand U7621 (N_7621,N_7388,N_7031);
or U7622 (N_7622,N_7051,N_7475);
nor U7623 (N_7623,N_7496,N_7429);
or U7624 (N_7624,N_7358,N_7443);
or U7625 (N_7625,N_7384,N_7295);
or U7626 (N_7626,N_7489,N_7193);
xor U7627 (N_7627,N_7061,N_7287);
or U7628 (N_7628,N_7133,N_7411);
or U7629 (N_7629,N_7057,N_7479);
nand U7630 (N_7630,N_7304,N_7233);
nand U7631 (N_7631,N_7200,N_7362);
or U7632 (N_7632,N_7238,N_7418);
nor U7633 (N_7633,N_7492,N_7121);
nor U7634 (N_7634,N_7098,N_7422);
xor U7635 (N_7635,N_7236,N_7148);
or U7636 (N_7636,N_7337,N_7447);
and U7637 (N_7637,N_7197,N_7178);
nand U7638 (N_7638,N_7276,N_7237);
or U7639 (N_7639,N_7167,N_7323);
nand U7640 (N_7640,N_7394,N_7159);
nand U7641 (N_7641,N_7112,N_7359);
or U7642 (N_7642,N_7172,N_7222);
and U7643 (N_7643,N_7280,N_7012);
or U7644 (N_7644,N_7274,N_7472);
and U7645 (N_7645,N_7157,N_7364);
nor U7646 (N_7646,N_7376,N_7399);
and U7647 (N_7647,N_7033,N_7234);
and U7648 (N_7648,N_7412,N_7043);
xnor U7649 (N_7649,N_7251,N_7456);
nor U7650 (N_7650,N_7026,N_7355);
or U7651 (N_7651,N_7373,N_7387);
or U7652 (N_7652,N_7109,N_7259);
xor U7653 (N_7653,N_7409,N_7179);
nand U7654 (N_7654,N_7266,N_7240);
and U7655 (N_7655,N_7269,N_7014);
and U7656 (N_7656,N_7077,N_7393);
and U7657 (N_7657,N_7281,N_7013);
and U7658 (N_7658,N_7301,N_7032);
or U7659 (N_7659,N_7074,N_7023);
nand U7660 (N_7660,N_7306,N_7339);
nor U7661 (N_7661,N_7064,N_7158);
or U7662 (N_7662,N_7400,N_7190);
and U7663 (N_7663,N_7078,N_7166);
nor U7664 (N_7664,N_7386,N_7279);
nand U7665 (N_7665,N_7154,N_7088);
and U7666 (N_7666,N_7211,N_7310);
nand U7667 (N_7667,N_7350,N_7262);
or U7668 (N_7668,N_7289,N_7007);
or U7669 (N_7669,N_7449,N_7298);
and U7670 (N_7670,N_7175,N_7199);
nand U7671 (N_7671,N_7431,N_7319);
nor U7672 (N_7672,N_7430,N_7034);
nor U7673 (N_7673,N_7408,N_7141);
nand U7674 (N_7674,N_7230,N_7397);
and U7675 (N_7675,N_7461,N_7225);
and U7676 (N_7676,N_7180,N_7499);
or U7677 (N_7677,N_7009,N_7433);
and U7678 (N_7678,N_7137,N_7440);
and U7679 (N_7679,N_7235,N_7035);
nor U7680 (N_7680,N_7171,N_7303);
or U7681 (N_7681,N_7391,N_7218);
nand U7682 (N_7682,N_7084,N_7495);
and U7683 (N_7683,N_7265,N_7048);
or U7684 (N_7684,N_7205,N_7139);
nor U7685 (N_7685,N_7030,N_7361);
nand U7686 (N_7686,N_7428,N_7052);
nor U7687 (N_7687,N_7327,N_7439);
nor U7688 (N_7688,N_7054,N_7113);
or U7689 (N_7689,N_7284,N_7487);
nand U7690 (N_7690,N_7095,N_7142);
and U7691 (N_7691,N_7066,N_7092);
or U7692 (N_7692,N_7185,N_7349);
nand U7693 (N_7693,N_7381,N_7152);
nand U7694 (N_7694,N_7082,N_7367);
xnor U7695 (N_7695,N_7002,N_7481);
nor U7696 (N_7696,N_7046,N_7320);
nor U7697 (N_7697,N_7010,N_7081);
nand U7698 (N_7698,N_7291,N_7261);
nor U7699 (N_7699,N_7104,N_7110);
nand U7700 (N_7700,N_7195,N_7020);
nor U7701 (N_7701,N_7436,N_7127);
nor U7702 (N_7702,N_7184,N_7277);
nand U7703 (N_7703,N_7445,N_7268);
and U7704 (N_7704,N_7410,N_7094);
or U7705 (N_7705,N_7348,N_7416);
or U7706 (N_7706,N_7313,N_7434);
and U7707 (N_7707,N_7379,N_7450);
or U7708 (N_7708,N_7116,N_7476);
nand U7709 (N_7709,N_7490,N_7493);
and U7710 (N_7710,N_7087,N_7353);
nand U7711 (N_7711,N_7228,N_7332);
nand U7712 (N_7712,N_7382,N_7403);
xor U7713 (N_7713,N_7294,N_7105);
or U7714 (N_7714,N_7073,N_7371);
nor U7715 (N_7715,N_7483,N_7296);
nand U7716 (N_7716,N_7469,N_7451);
and U7717 (N_7717,N_7404,N_7065);
or U7718 (N_7718,N_7182,N_7401);
nand U7719 (N_7719,N_7209,N_7162);
and U7720 (N_7720,N_7264,N_7245);
nand U7721 (N_7721,N_7335,N_7071);
and U7722 (N_7722,N_7022,N_7398);
or U7723 (N_7723,N_7246,N_7042);
or U7724 (N_7724,N_7155,N_7126);
nand U7725 (N_7725,N_7446,N_7334);
nor U7726 (N_7726,N_7130,N_7241);
nand U7727 (N_7727,N_7405,N_7018);
or U7728 (N_7728,N_7345,N_7390);
or U7729 (N_7729,N_7056,N_7196);
and U7730 (N_7730,N_7454,N_7421);
or U7731 (N_7731,N_7326,N_7156);
xnor U7732 (N_7732,N_7147,N_7122);
nand U7733 (N_7733,N_7340,N_7309);
and U7734 (N_7734,N_7282,N_7344);
and U7735 (N_7735,N_7455,N_7170);
nand U7736 (N_7736,N_7149,N_7253);
nor U7737 (N_7737,N_7325,N_7177);
or U7738 (N_7738,N_7470,N_7096);
nand U7739 (N_7739,N_7438,N_7138);
nand U7740 (N_7740,N_7300,N_7396);
nor U7741 (N_7741,N_7458,N_7080);
or U7742 (N_7742,N_7336,N_7217);
nor U7743 (N_7743,N_7011,N_7017);
nor U7744 (N_7744,N_7395,N_7448);
nor U7745 (N_7745,N_7256,N_7354);
and U7746 (N_7746,N_7330,N_7207);
and U7747 (N_7747,N_7120,N_7286);
and U7748 (N_7748,N_7292,N_7108);
and U7749 (N_7749,N_7333,N_7144);
or U7750 (N_7750,N_7445,N_7392);
nand U7751 (N_7751,N_7112,N_7013);
and U7752 (N_7752,N_7460,N_7467);
and U7753 (N_7753,N_7319,N_7382);
xor U7754 (N_7754,N_7335,N_7139);
nor U7755 (N_7755,N_7106,N_7447);
nand U7756 (N_7756,N_7398,N_7259);
or U7757 (N_7757,N_7212,N_7095);
nor U7758 (N_7758,N_7351,N_7062);
nand U7759 (N_7759,N_7457,N_7313);
nand U7760 (N_7760,N_7062,N_7189);
and U7761 (N_7761,N_7071,N_7421);
nand U7762 (N_7762,N_7343,N_7494);
xor U7763 (N_7763,N_7220,N_7273);
or U7764 (N_7764,N_7440,N_7027);
nand U7765 (N_7765,N_7188,N_7021);
xor U7766 (N_7766,N_7208,N_7487);
nor U7767 (N_7767,N_7005,N_7298);
nor U7768 (N_7768,N_7196,N_7294);
nand U7769 (N_7769,N_7330,N_7013);
nand U7770 (N_7770,N_7244,N_7444);
and U7771 (N_7771,N_7034,N_7288);
or U7772 (N_7772,N_7011,N_7275);
nand U7773 (N_7773,N_7267,N_7366);
and U7774 (N_7774,N_7111,N_7084);
and U7775 (N_7775,N_7307,N_7044);
nor U7776 (N_7776,N_7243,N_7217);
nor U7777 (N_7777,N_7428,N_7434);
nor U7778 (N_7778,N_7278,N_7020);
nand U7779 (N_7779,N_7280,N_7377);
nor U7780 (N_7780,N_7331,N_7135);
or U7781 (N_7781,N_7477,N_7198);
nand U7782 (N_7782,N_7431,N_7345);
nor U7783 (N_7783,N_7309,N_7028);
nand U7784 (N_7784,N_7406,N_7226);
nor U7785 (N_7785,N_7173,N_7381);
nand U7786 (N_7786,N_7073,N_7104);
nand U7787 (N_7787,N_7036,N_7381);
nand U7788 (N_7788,N_7239,N_7049);
and U7789 (N_7789,N_7063,N_7449);
nor U7790 (N_7790,N_7435,N_7288);
nor U7791 (N_7791,N_7188,N_7059);
or U7792 (N_7792,N_7073,N_7072);
nand U7793 (N_7793,N_7318,N_7281);
or U7794 (N_7794,N_7406,N_7265);
or U7795 (N_7795,N_7106,N_7101);
or U7796 (N_7796,N_7307,N_7242);
nand U7797 (N_7797,N_7469,N_7252);
or U7798 (N_7798,N_7475,N_7097);
or U7799 (N_7799,N_7030,N_7294);
nand U7800 (N_7800,N_7414,N_7354);
nor U7801 (N_7801,N_7489,N_7405);
nor U7802 (N_7802,N_7447,N_7231);
or U7803 (N_7803,N_7264,N_7086);
and U7804 (N_7804,N_7468,N_7201);
or U7805 (N_7805,N_7439,N_7100);
nand U7806 (N_7806,N_7046,N_7005);
nor U7807 (N_7807,N_7156,N_7395);
nand U7808 (N_7808,N_7248,N_7196);
and U7809 (N_7809,N_7109,N_7264);
nor U7810 (N_7810,N_7274,N_7350);
nor U7811 (N_7811,N_7387,N_7324);
nor U7812 (N_7812,N_7081,N_7211);
and U7813 (N_7813,N_7497,N_7384);
nor U7814 (N_7814,N_7431,N_7200);
and U7815 (N_7815,N_7224,N_7437);
nand U7816 (N_7816,N_7289,N_7440);
or U7817 (N_7817,N_7157,N_7013);
nor U7818 (N_7818,N_7002,N_7438);
nor U7819 (N_7819,N_7359,N_7135);
and U7820 (N_7820,N_7291,N_7417);
nand U7821 (N_7821,N_7263,N_7431);
nor U7822 (N_7822,N_7335,N_7487);
nand U7823 (N_7823,N_7092,N_7045);
nand U7824 (N_7824,N_7076,N_7393);
nand U7825 (N_7825,N_7166,N_7052);
or U7826 (N_7826,N_7176,N_7316);
and U7827 (N_7827,N_7262,N_7461);
nand U7828 (N_7828,N_7145,N_7235);
nor U7829 (N_7829,N_7399,N_7196);
and U7830 (N_7830,N_7220,N_7133);
xnor U7831 (N_7831,N_7241,N_7221);
nand U7832 (N_7832,N_7453,N_7216);
nand U7833 (N_7833,N_7022,N_7025);
and U7834 (N_7834,N_7157,N_7353);
nand U7835 (N_7835,N_7239,N_7083);
and U7836 (N_7836,N_7444,N_7195);
and U7837 (N_7837,N_7061,N_7242);
nor U7838 (N_7838,N_7195,N_7018);
and U7839 (N_7839,N_7311,N_7478);
nand U7840 (N_7840,N_7278,N_7398);
or U7841 (N_7841,N_7350,N_7040);
or U7842 (N_7842,N_7314,N_7411);
or U7843 (N_7843,N_7455,N_7429);
and U7844 (N_7844,N_7242,N_7198);
and U7845 (N_7845,N_7040,N_7466);
or U7846 (N_7846,N_7051,N_7250);
or U7847 (N_7847,N_7062,N_7065);
or U7848 (N_7848,N_7405,N_7400);
nand U7849 (N_7849,N_7151,N_7341);
nor U7850 (N_7850,N_7348,N_7357);
or U7851 (N_7851,N_7445,N_7311);
nor U7852 (N_7852,N_7264,N_7377);
nand U7853 (N_7853,N_7167,N_7015);
or U7854 (N_7854,N_7246,N_7439);
nand U7855 (N_7855,N_7222,N_7018);
and U7856 (N_7856,N_7362,N_7436);
nor U7857 (N_7857,N_7292,N_7332);
nand U7858 (N_7858,N_7487,N_7147);
nand U7859 (N_7859,N_7007,N_7388);
or U7860 (N_7860,N_7422,N_7255);
and U7861 (N_7861,N_7206,N_7193);
or U7862 (N_7862,N_7180,N_7448);
or U7863 (N_7863,N_7375,N_7386);
nor U7864 (N_7864,N_7397,N_7414);
nor U7865 (N_7865,N_7100,N_7095);
nor U7866 (N_7866,N_7362,N_7210);
and U7867 (N_7867,N_7495,N_7170);
nor U7868 (N_7868,N_7074,N_7236);
nor U7869 (N_7869,N_7216,N_7400);
nor U7870 (N_7870,N_7011,N_7302);
nor U7871 (N_7871,N_7269,N_7298);
or U7872 (N_7872,N_7078,N_7199);
or U7873 (N_7873,N_7130,N_7385);
nand U7874 (N_7874,N_7492,N_7496);
nor U7875 (N_7875,N_7046,N_7240);
and U7876 (N_7876,N_7352,N_7186);
and U7877 (N_7877,N_7447,N_7094);
nor U7878 (N_7878,N_7195,N_7318);
and U7879 (N_7879,N_7040,N_7312);
and U7880 (N_7880,N_7054,N_7463);
and U7881 (N_7881,N_7282,N_7317);
and U7882 (N_7882,N_7467,N_7007);
and U7883 (N_7883,N_7251,N_7478);
nand U7884 (N_7884,N_7450,N_7360);
nor U7885 (N_7885,N_7050,N_7407);
and U7886 (N_7886,N_7485,N_7406);
and U7887 (N_7887,N_7319,N_7389);
or U7888 (N_7888,N_7354,N_7484);
nor U7889 (N_7889,N_7008,N_7241);
and U7890 (N_7890,N_7136,N_7061);
nand U7891 (N_7891,N_7134,N_7244);
and U7892 (N_7892,N_7390,N_7054);
nor U7893 (N_7893,N_7167,N_7491);
and U7894 (N_7894,N_7225,N_7385);
or U7895 (N_7895,N_7154,N_7091);
nor U7896 (N_7896,N_7141,N_7204);
or U7897 (N_7897,N_7057,N_7450);
or U7898 (N_7898,N_7488,N_7413);
nor U7899 (N_7899,N_7185,N_7443);
nand U7900 (N_7900,N_7276,N_7280);
or U7901 (N_7901,N_7491,N_7039);
nand U7902 (N_7902,N_7205,N_7181);
nor U7903 (N_7903,N_7301,N_7076);
or U7904 (N_7904,N_7114,N_7080);
nand U7905 (N_7905,N_7072,N_7048);
nor U7906 (N_7906,N_7451,N_7278);
nand U7907 (N_7907,N_7097,N_7439);
nand U7908 (N_7908,N_7490,N_7355);
nor U7909 (N_7909,N_7246,N_7391);
nand U7910 (N_7910,N_7215,N_7347);
and U7911 (N_7911,N_7359,N_7058);
nor U7912 (N_7912,N_7489,N_7468);
nor U7913 (N_7913,N_7321,N_7164);
and U7914 (N_7914,N_7145,N_7054);
or U7915 (N_7915,N_7218,N_7001);
nand U7916 (N_7916,N_7236,N_7091);
or U7917 (N_7917,N_7118,N_7402);
nand U7918 (N_7918,N_7195,N_7174);
nand U7919 (N_7919,N_7448,N_7388);
or U7920 (N_7920,N_7277,N_7389);
and U7921 (N_7921,N_7480,N_7245);
nor U7922 (N_7922,N_7297,N_7385);
nor U7923 (N_7923,N_7338,N_7077);
nand U7924 (N_7924,N_7386,N_7485);
and U7925 (N_7925,N_7007,N_7352);
xnor U7926 (N_7926,N_7231,N_7128);
nand U7927 (N_7927,N_7208,N_7411);
nand U7928 (N_7928,N_7121,N_7043);
nor U7929 (N_7929,N_7095,N_7435);
or U7930 (N_7930,N_7229,N_7090);
and U7931 (N_7931,N_7462,N_7474);
or U7932 (N_7932,N_7302,N_7413);
and U7933 (N_7933,N_7019,N_7471);
nand U7934 (N_7934,N_7196,N_7442);
or U7935 (N_7935,N_7047,N_7372);
and U7936 (N_7936,N_7458,N_7344);
nand U7937 (N_7937,N_7430,N_7066);
or U7938 (N_7938,N_7452,N_7326);
nand U7939 (N_7939,N_7400,N_7434);
nor U7940 (N_7940,N_7112,N_7362);
xor U7941 (N_7941,N_7404,N_7488);
nor U7942 (N_7942,N_7045,N_7250);
nor U7943 (N_7943,N_7250,N_7071);
and U7944 (N_7944,N_7264,N_7329);
or U7945 (N_7945,N_7109,N_7460);
and U7946 (N_7946,N_7128,N_7467);
or U7947 (N_7947,N_7390,N_7451);
and U7948 (N_7948,N_7445,N_7422);
and U7949 (N_7949,N_7359,N_7054);
nand U7950 (N_7950,N_7172,N_7369);
nor U7951 (N_7951,N_7085,N_7208);
xnor U7952 (N_7952,N_7428,N_7021);
or U7953 (N_7953,N_7381,N_7241);
nand U7954 (N_7954,N_7155,N_7333);
nand U7955 (N_7955,N_7412,N_7394);
or U7956 (N_7956,N_7384,N_7280);
nand U7957 (N_7957,N_7334,N_7490);
nor U7958 (N_7958,N_7435,N_7415);
and U7959 (N_7959,N_7307,N_7486);
and U7960 (N_7960,N_7353,N_7464);
and U7961 (N_7961,N_7020,N_7307);
nand U7962 (N_7962,N_7383,N_7285);
and U7963 (N_7963,N_7271,N_7318);
nand U7964 (N_7964,N_7495,N_7229);
nor U7965 (N_7965,N_7000,N_7422);
nor U7966 (N_7966,N_7229,N_7013);
and U7967 (N_7967,N_7402,N_7075);
nand U7968 (N_7968,N_7202,N_7321);
nor U7969 (N_7969,N_7140,N_7485);
nand U7970 (N_7970,N_7146,N_7221);
or U7971 (N_7971,N_7403,N_7173);
nor U7972 (N_7972,N_7019,N_7245);
nand U7973 (N_7973,N_7217,N_7097);
and U7974 (N_7974,N_7444,N_7284);
and U7975 (N_7975,N_7162,N_7303);
nand U7976 (N_7976,N_7327,N_7294);
nor U7977 (N_7977,N_7289,N_7103);
nor U7978 (N_7978,N_7040,N_7209);
or U7979 (N_7979,N_7090,N_7483);
or U7980 (N_7980,N_7479,N_7050);
and U7981 (N_7981,N_7025,N_7041);
or U7982 (N_7982,N_7481,N_7253);
or U7983 (N_7983,N_7336,N_7100);
nor U7984 (N_7984,N_7035,N_7102);
nand U7985 (N_7985,N_7360,N_7388);
nand U7986 (N_7986,N_7404,N_7245);
nand U7987 (N_7987,N_7202,N_7392);
or U7988 (N_7988,N_7285,N_7164);
or U7989 (N_7989,N_7431,N_7308);
or U7990 (N_7990,N_7122,N_7349);
nor U7991 (N_7991,N_7163,N_7490);
nor U7992 (N_7992,N_7205,N_7271);
and U7993 (N_7993,N_7413,N_7158);
or U7994 (N_7994,N_7124,N_7065);
nand U7995 (N_7995,N_7387,N_7196);
or U7996 (N_7996,N_7065,N_7131);
nand U7997 (N_7997,N_7481,N_7383);
nor U7998 (N_7998,N_7345,N_7389);
nor U7999 (N_7999,N_7359,N_7315);
nor U8000 (N_8000,N_7692,N_7539);
xnor U8001 (N_8001,N_7927,N_7857);
xnor U8002 (N_8002,N_7941,N_7704);
nand U8003 (N_8003,N_7868,N_7797);
nor U8004 (N_8004,N_7671,N_7617);
and U8005 (N_8005,N_7816,N_7728);
nor U8006 (N_8006,N_7901,N_7731);
nor U8007 (N_8007,N_7534,N_7686);
nand U8008 (N_8008,N_7934,N_7827);
nor U8009 (N_8009,N_7645,N_7609);
nor U8010 (N_8010,N_7983,N_7500);
nand U8011 (N_8011,N_7553,N_7559);
nor U8012 (N_8012,N_7806,N_7920);
nand U8013 (N_8013,N_7574,N_7864);
nand U8014 (N_8014,N_7641,N_7684);
nor U8015 (N_8015,N_7949,N_7608);
nand U8016 (N_8016,N_7952,N_7585);
or U8017 (N_8017,N_7991,N_7603);
nand U8018 (N_8018,N_7637,N_7606);
and U8019 (N_8019,N_7524,N_7943);
nor U8020 (N_8020,N_7838,N_7963);
or U8021 (N_8021,N_7848,N_7689);
nor U8022 (N_8022,N_7897,N_7834);
and U8023 (N_8023,N_7572,N_7712);
or U8024 (N_8024,N_7571,N_7577);
and U8025 (N_8025,N_7807,N_7947);
nor U8026 (N_8026,N_7674,N_7509);
nand U8027 (N_8027,N_7588,N_7974);
nor U8028 (N_8028,N_7912,N_7542);
and U8029 (N_8029,N_7656,N_7911);
nor U8030 (N_8030,N_7958,N_7681);
xnor U8031 (N_8031,N_7525,N_7812);
and U8032 (N_8032,N_7582,N_7850);
nor U8033 (N_8033,N_7937,N_7871);
or U8034 (N_8034,N_7769,N_7531);
or U8035 (N_8035,N_7616,N_7504);
and U8036 (N_8036,N_7789,N_7878);
nand U8037 (N_8037,N_7989,N_7618);
nor U8038 (N_8038,N_7701,N_7682);
nand U8039 (N_8039,N_7634,N_7560);
or U8040 (N_8040,N_7836,N_7591);
nor U8041 (N_8041,N_7554,N_7843);
nor U8042 (N_8042,N_7988,N_7640);
and U8043 (N_8043,N_7540,N_7774);
nor U8044 (N_8044,N_7971,N_7518);
or U8045 (N_8045,N_7663,N_7996);
or U8046 (N_8046,N_7700,N_7763);
nand U8047 (N_8047,N_7905,N_7826);
nand U8048 (N_8048,N_7955,N_7581);
nor U8049 (N_8049,N_7845,N_7880);
or U8050 (N_8050,N_7739,N_7725);
nor U8051 (N_8051,N_7945,N_7652);
or U8052 (N_8052,N_7638,N_7813);
nand U8053 (N_8053,N_7702,N_7820);
and U8054 (N_8054,N_7749,N_7629);
and U8055 (N_8055,N_7928,N_7825);
and U8056 (N_8056,N_7804,N_7607);
nor U8057 (N_8057,N_7872,N_7898);
nor U8058 (N_8058,N_7758,N_7977);
and U8059 (N_8059,N_7994,N_7612);
or U8060 (N_8060,N_7532,N_7876);
nor U8061 (N_8061,N_7501,N_7851);
or U8062 (N_8062,N_7926,N_7830);
nand U8063 (N_8063,N_7649,N_7558);
or U8064 (N_8064,N_7803,N_7859);
or U8065 (N_8065,N_7969,N_7661);
or U8066 (N_8066,N_7747,N_7718);
or U8067 (N_8067,N_7547,N_7879);
nand U8068 (N_8068,N_7759,N_7740);
nor U8069 (N_8069,N_7925,N_7610);
nor U8070 (N_8070,N_7894,N_7678);
and U8071 (N_8071,N_7631,N_7968);
and U8072 (N_8072,N_7683,N_7929);
and U8073 (N_8073,N_7915,N_7824);
and U8074 (N_8074,N_7787,N_7742);
and U8075 (N_8075,N_7919,N_7995);
or U8076 (N_8076,N_7999,N_7515);
nor U8077 (N_8077,N_7869,N_7556);
and U8078 (N_8078,N_7957,N_7630);
nand U8079 (N_8079,N_7873,N_7732);
nand U8080 (N_8080,N_7528,N_7858);
or U8081 (N_8081,N_7673,N_7589);
nor U8082 (N_8082,N_7844,N_7975);
and U8083 (N_8083,N_7735,N_7853);
nand U8084 (N_8084,N_7713,N_7651);
nand U8085 (N_8085,N_7579,N_7791);
or U8086 (N_8086,N_7895,N_7510);
nand U8087 (N_8087,N_7670,N_7982);
nand U8088 (N_8088,N_7782,N_7538);
nand U8089 (N_8089,N_7951,N_7802);
nand U8090 (N_8090,N_7516,N_7889);
nand U8091 (N_8091,N_7688,N_7530);
and U8092 (N_8092,N_7935,N_7865);
or U8093 (N_8093,N_7506,N_7622);
or U8094 (N_8094,N_7772,N_7940);
nor U8095 (N_8095,N_7710,N_7766);
and U8096 (N_8096,N_7993,N_7548);
or U8097 (N_8097,N_7578,N_7765);
or U8098 (N_8098,N_7907,N_7831);
or U8099 (N_8099,N_7668,N_7561);
nand U8100 (N_8100,N_7724,N_7867);
nor U8101 (N_8101,N_7964,N_7567);
nand U8102 (N_8102,N_7533,N_7696);
nand U8103 (N_8103,N_7767,N_7970);
or U8104 (N_8104,N_7833,N_7726);
or U8105 (N_8105,N_7846,N_7636);
or U8106 (N_8106,N_7817,N_7655);
and U8107 (N_8107,N_7744,N_7727);
nor U8108 (N_8108,N_7960,N_7669);
or U8109 (N_8109,N_7521,N_7882);
nor U8110 (N_8110,N_7543,N_7931);
or U8111 (N_8111,N_7601,N_7598);
nand U8112 (N_8112,N_7913,N_7593);
and U8113 (N_8113,N_7741,N_7950);
nand U8114 (N_8114,N_7523,N_7884);
xor U8115 (N_8115,N_7730,N_7755);
nor U8116 (N_8116,N_7555,N_7959);
nor U8117 (N_8117,N_7918,N_7810);
nor U8118 (N_8118,N_7738,N_7737);
and U8119 (N_8119,N_7664,N_7657);
or U8120 (N_8120,N_7733,N_7736);
and U8121 (N_8121,N_7595,N_7821);
nand U8122 (N_8122,N_7754,N_7777);
or U8123 (N_8123,N_7784,N_7566);
nor U8124 (N_8124,N_7860,N_7604);
or U8125 (N_8125,N_7788,N_7602);
nor U8126 (N_8126,N_7776,N_7854);
nand U8127 (N_8127,N_7828,N_7746);
nor U8128 (N_8128,N_7680,N_7753);
nor U8129 (N_8129,N_7537,N_7786);
and U8130 (N_8130,N_7529,N_7679);
nor U8131 (N_8131,N_7541,N_7717);
nand U8132 (N_8132,N_7667,N_7832);
nor U8133 (N_8133,N_7847,N_7768);
nor U8134 (N_8134,N_7779,N_7502);
xnor U8135 (N_8135,N_7930,N_7508);
nand U8136 (N_8136,N_7849,N_7714);
and U8137 (N_8137,N_7852,N_7557);
nor U8138 (N_8138,N_7505,N_7773);
or U8139 (N_8139,N_7881,N_7590);
or U8140 (N_8140,N_7794,N_7583);
nand U8141 (N_8141,N_7587,N_7902);
nand U8142 (N_8142,N_7805,N_7980);
and U8143 (N_8143,N_7514,N_7984);
and U8144 (N_8144,N_7778,N_7801);
or U8145 (N_8145,N_7966,N_7695);
and U8146 (N_8146,N_7708,N_7908);
nand U8147 (N_8147,N_7676,N_7948);
nand U8148 (N_8148,N_7517,N_7811);
nand U8149 (N_8149,N_7644,N_7596);
and U8150 (N_8150,N_7623,N_7584);
or U8151 (N_8151,N_7760,N_7793);
or U8152 (N_8152,N_7808,N_7716);
nand U8153 (N_8153,N_7976,N_7917);
and U8154 (N_8154,N_7647,N_7900);
nor U8155 (N_8155,N_7750,N_7745);
nand U8156 (N_8156,N_7707,N_7814);
nand U8157 (N_8157,N_7906,N_7899);
or U8158 (N_8158,N_7795,N_7693);
nor U8159 (N_8159,N_7874,N_7762);
nand U8160 (N_8160,N_7904,N_7719);
and U8161 (N_8161,N_7697,N_7550);
nand U8162 (N_8162,N_7809,N_7563);
nor U8163 (N_8163,N_7705,N_7870);
or U8164 (N_8164,N_7594,N_7761);
nor U8165 (N_8165,N_7822,N_7823);
nor U8166 (N_8166,N_7792,N_7997);
nand U8167 (N_8167,N_7863,N_7648);
nor U8168 (N_8168,N_7672,N_7565);
nor U8169 (N_8169,N_7665,N_7544);
nor U8170 (N_8170,N_7654,N_7513);
nand U8171 (N_8171,N_7921,N_7706);
or U8172 (N_8172,N_7723,N_7756);
or U8173 (N_8173,N_7562,N_7896);
nor U8174 (N_8174,N_7620,N_7944);
nor U8175 (N_8175,N_7837,N_7576);
nor U8176 (N_8176,N_7862,N_7546);
nor U8177 (N_8177,N_7666,N_7998);
nor U8178 (N_8178,N_7936,N_7883);
or U8179 (N_8179,N_7646,N_7903);
and U8180 (N_8180,N_7967,N_7615);
and U8181 (N_8181,N_7924,N_7751);
and U8182 (N_8182,N_7597,N_7633);
nor U8183 (N_8183,N_7796,N_7614);
nor U8184 (N_8184,N_7938,N_7660);
nand U8185 (N_8185,N_7771,N_7545);
and U8186 (N_8186,N_7711,N_7829);
or U8187 (N_8187,N_7650,N_7892);
nand U8188 (N_8188,N_7839,N_7687);
and U8189 (N_8189,N_7992,N_7990);
nor U8190 (N_8190,N_7722,N_7659);
or U8191 (N_8191,N_7570,N_7987);
or U8192 (N_8192,N_7962,N_7694);
nor U8193 (N_8193,N_7621,N_7658);
nand U8194 (N_8194,N_7914,N_7549);
and U8195 (N_8195,N_7653,N_7662);
and U8196 (N_8196,N_7972,N_7757);
and U8197 (N_8197,N_7709,N_7527);
or U8198 (N_8198,N_7922,N_7798);
or U8199 (N_8199,N_7875,N_7942);
nand U8200 (N_8200,N_7627,N_7973);
or U8201 (N_8201,N_7819,N_7978);
and U8202 (N_8202,N_7799,N_7564);
and U8203 (N_8203,N_7939,N_7785);
nor U8204 (N_8204,N_7520,N_7632);
nand U8205 (N_8205,N_7923,N_7507);
and U8206 (N_8206,N_7780,N_7586);
or U8207 (N_8207,N_7592,N_7573);
or U8208 (N_8208,N_7985,N_7835);
and U8209 (N_8209,N_7552,N_7519);
or U8210 (N_8210,N_7961,N_7599);
and U8211 (N_8211,N_7690,N_7979);
nand U8212 (N_8212,N_7703,N_7512);
or U8213 (N_8213,N_7526,N_7783);
nor U8214 (N_8214,N_7536,N_7818);
nand U8215 (N_8215,N_7885,N_7770);
and U8216 (N_8216,N_7635,N_7691);
nor U8217 (N_8217,N_7861,N_7841);
or U8218 (N_8218,N_7790,N_7568);
nand U8219 (N_8219,N_7626,N_7628);
nand U8220 (N_8220,N_7916,N_7856);
or U8221 (N_8221,N_7932,N_7625);
nor U8222 (N_8222,N_7600,N_7752);
and U8223 (N_8223,N_7748,N_7954);
nand U8224 (N_8224,N_7986,N_7677);
nor U8225 (N_8225,N_7840,N_7956);
or U8226 (N_8226,N_7619,N_7953);
nor U8227 (N_8227,N_7887,N_7729);
or U8228 (N_8228,N_7580,N_7800);
and U8229 (N_8229,N_7720,N_7698);
and U8230 (N_8230,N_7877,N_7909);
and U8231 (N_8231,N_7775,N_7981);
nor U8232 (N_8232,N_7522,N_7715);
nand U8233 (N_8233,N_7743,N_7699);
xnor U8234 (N_8234,N_7685,N_7890);
nand U8235 (N_8235,N_7842,N_7721);
nor U8236 (N_8236,N_7611,N_7535);
nand U8237 (N_8237,N_7815,N_7503);
nand U8238 (N_8238,N_7605,N_7511);
and U8239 (N_8239,N_7891,N_7575);
and U8240 (N_8240,N_7910,N_7886);
or U8241 (N_8241,N_7642,N_7893);
and U8242 (N_8242,N_7675,N_7639);
and U8243 (N_8243,N_7933,N_7551);
or U8244 (N_8244,N_7764,N_7888);
and U8245 (N_8245,N_7734,N_7613);
and U8246 (N_8246,N_7781,N_7643);
and U8247 (N_8247,N_7624,N_7866);
nand U8248 (N_8248,N_7855,N_7965);
nor U8249 (N_8249,N_7946,N_7569);
nor U8250 (N_8250,N_7704,N_7993);
xnor U8251 (N_8251,N_7574,N_7631);
and U8252 (N_8252,N_7737,N_7947);
nand U8253 (N_8253,N_7584,N_7626);
nand U8254 (N_8254,N_7556,N_7714);
nand U8255 (N_8255,N_7723,N_7716);
nand U8256 (N_8256,N_7526,N_7863);
and U8257 (N_8257,N_7768,N_7656);
and U8258 (N_8258,N_7882,N_7878);
or U8259 (N_8259,N_7847,N_7592);
or U8260 (N_8260,N_7814,N_7975);
and U8261 (N_8261,N_7812,N_7733);
or U8262 (N_8262,N_7619,N_7682);
or U8263 (N_8263,N_7576,N_7634);
and U8264 (N_8264,N_7809,N_7804);
nor U8265 (N_8265,N_7728,N_7593);
nor U8266 (N_8266,N_7688,N_7851);
and U8267 (N_8267,N_7855,N_7746);
and U8268 (N_8268,N_7709,N_7940);
nand U8269 (N_8269,N_7770,N_7677);
and U8270 (N_8270,N_7720,N_7669);
nand U8271 (N_8271,N_7818,N_7929);
and U8272 (N_8272,N_7597,N_7894);
or U8273 (N_8273,N_7714,N_7544);
and U8274 (N_8274,N_7806,N_7985);
or U8275 (N_8275,N_7540,N_7863);
nor U8276 (N_8276,N_7578,N_7981);
or U8277 (N_8277,N_7527,N_7644);
nand U8278 (N_8278,N_7941,N_7836);
nand U8279 (N_8279,N_7710,N_7514);
nand U8280 (N_8280,N_7505,N_7941);
nand U8281 (N_8281,N_7738,N_7687);
or U8282 (N_8282,N_7599,N_7529);
xor U8283 (N_8283,N_7746,N_7780);
nor U8284 (N_8284,N_7658,N_7579);
or U8285 (N_8285,N_7765,N_7550);
or U8286 (N_8286,N_7912,N_7775);
and U8287 (N_8287,N_7694,N_7532);
nor U8288 (N_8288,N_7698,N_7519);
nand U8289 (N_8289,N_7882,N_7613);
nor U8290 (N_8290,N_7559,N_7644);
and U8291 (N_8291,N_7896,N_7943);
nand U8292 (N_8292,N_7719,N_7582);
and U8293 (N_8293,N_7541,N_7969);
nand U8294 (N_8294,N_7643,N_7607);
nor U8295 (N_8295,N_7526,N_7841);
nor U8296 (N_8296,N_7787,N_7781);
or U8297 (N_8297,N_7993,N_7568);
or U8298 (N_8298,N_7568,N_7782);
nor U8299 (N_8299,N_7692,N_7904);
nand U8300 (N_8300,N_7516,N_7843);
or U8301 (N_8301,N_7715,N_7935);
or U8302 (N_8302,N_7871,N_7997);
nor U8303 (N_8303,N_7782,N_7730);
or U8304 (N_8304,N_7607,N_7919);
nor U8305 (N_8305,N_7644,N_7751);
nand U8306 (N_8306,N_7545,N_7567);
nand U8307 (N_8307,N_7899,N_7969);
and U8308 (N_8308,N_7834,N_7502);
nor U8309 (N_8309,N_7675,N_7914);
and U8310 (N_8310,N_7829,N_7953);
or U8311 (N_8311,N_7578,N_7626);
and U8312 (N_8312,N_7556,N_7905);
nand U8313 (N_8313,N_7881,N_7940);
nor U8314 (N_8314,N_7673,N_7798);
or U8315 (N_8315,N_7810,N_7852);
nand U8316 (N_8316,N_7590,N_7661);
or U8317 (N_8317,N_7718,N_7710);
or U8318 (N_8318,N_7648,N_7799);
or U8319 (N_8319,N_7768,N_7636);
nor U8320 (N_8320,N_7812,N_7850);
nand U8321 (N_8321,N_7659,N_7936);
nor U8322 (N_8322,N_7842,N_7690);
nor U8323 (N_8323,N_7872,N_7684);
and U8324 (N_8324,N_7953,N_7885);
nor U8325 (N_8325,N_7984,N_7546);
nand U8326 (N_8326,N_7555,N_7786);
nor U8327 (N_8327,N_7664,N_7554);
nand U8328 (N_8328,N_7805,N_7839);
nor U8329 (N_8329,N_7562,N_7696);
and U8330 (N_8330,N_7567,N_7934);
nor U8331 (N_8331,N_7835,N_7747);
or U8332 (N_8332,N_7892,N_7518);
nand U8333 (N_8333,N_7854,N_7957);
nand U8334 (N_8334,N_7567,N_7579);
or U8335 (N_8335,N_7631,N_7620);
and U8336 (N_8336,N_7738,N_7808);
nor U8337 (N_8337,N_7693,N_7662);
or U8338 (N_8338,N_7801,N_7854);
and U8339 (N_8339,N_7949,N_7866);
nand U8340 (N_8340,N_7861,N_7582);
or U8341 (N_8341,N_7701,N_7521);
nor U8342 (N_8342,N_7854,N_7737);
nor U8343 (N_8343,N_7844,N_7705);
nor U8344 (N_8344,N_7613,N_7545);
nor U8345 (N_8345,N_7698,N_7530);
and U8346 (N_8346,N_7568,N_7588);
and U8347 (N_8347,N_7700,N_7735);
and U8348 (N_8348,N_7830,N_7820);
and U8349 (N_8349,N_7907,N_7678);
nand U8350 (N_8350,N_7875,N_7851);
and U8351 (N_8351,N_7914,N_7896);
and U8352 (N_8352,N_7513,N_7696);
and U8353 (N_8353,N_7932,N_7506);
nor U8354 (N_8354,N_7732,N_7574);
or U8355 (N_8355,N_7704,N_7632);
nor U8356 (N_8356,N_7657,N_7880);
or U8357 (N_8357,N_7898,N_7917);
nor U8358 (N_8358,N_7578,N_7653);
and U8359 (N_8359,N_7744,N_7664);
or U8360 (N_8360,N_7665,N_7717);
nand U8361 (N_8361,N_7970,N_7957);
or U8362 (N_8362,N_7634,N_7986);
nor U8363 (N_8363,N_7714,N_7887);
or U8364 (N_8364,N_7707,N_7616);
nor U8365 (N_8365,N_7905,N_7760);
and U8366 (N_8366,N_7866,N_7871);
or U8367 (N_8367,N_7833,N_7710);
and U8368 (N_8368,N_7612,N_7817);
and U8369 (N_8369,N_7525,N_7606);
nor U8370 (N_8370,N_7561,N_7746);
and U8371 (N_8371,N_7829,N_7781);
nand U8372 (N_8372,N_7541,N_7614);
nor U8373 (N_8373,N_7543,N_7991);
nor U8374 (N_8374,N_7759,N_7541);
nor U8375 (N_8375,N_7963,N_7598);
or U8376 (N_8376,N_7641,N_7842);
or U8377 (N_8377,N_7972,N_7848);
nor U8378 (N_8378,N_7691,N_7975);
or U8379 (N_8379,N_7522,N_7532);
or U8380 (N_8380,N_7543,N_7561);
nor U8381 (N_8381,N_7647,N_7705);
and U8382 (N_8382,N_7931,N_7517);
nor U8383 (N_8383,N_7695,N_7829);
nor U8384 (N_8384,N_7943,N_7641);
nor U8385 (N_8385,N_7777,N_7691);
nand U8386 (N_8386,N_7690,N_7977);
nor U8387 (N_8387,N_7556,N_7681);
or U8388 (N_8388,N_7952,N_7816);
and U8389 (N_8389,N_7693,N_7521);
and U8390 (N_8390,N_7864,N_7982);
nor U8391 (N_8391,N_7504,N_7887);
or U8392 (N_8392,N_7644,N_7593);
or U8393 (N_8393,N_7830,N_7827);
and U8394 (N_8394,N_7628,N_7985);
or U8395 (N_8395,N_7542,N_7552);
or U8396 (N_8396,N_7968,N_7741);
nor U8397 (N_8397,N_7857,N_7610);
nand U8398 (N_8398,N_7949,N_7886);
and U8399 (N_8399,N_7763,N_7570);
nor U8400 (N_8400,N_7914,N_7721);
or U8401 (N_8401,N_7716,N_7502);
nor U8402 (N_8402,N_7632,N_7719);
nand U8403 (N_8403,N_7721,N_7714);
and U8404 (N_8404,N_7798,N_7686);
or U8405 (N_8405,N_7714,N_7623);
nor U8406 (N_8406,N_7530,N_7574);
nor U8407 (N_8407,N_7519,N_7676);
nand U8408 (N_8408,N_7780,N_7718);
nor U8409 (N_8409,N_7911,N_7681);
and U8410 (N_8410,N_7591,N_7887);
or U8411 (N_8411,N_7785,N_7789);
nand U8412 (N_8412,N_7649,N_7719);
and U8413 (N_8413,N_7926,N_7749);
and U8414 (N_8414,N_7551,N_7907);
nand U8415 (N_8415,N_7722,N_7636);
or U8416 (N_8416,N_7635,N_7520);
nor U8417 (N_8417,N_7629,N_7815);
xnor U8418 (N_8418,N_7632,N_7842);
or U8419 (N_8419,N_7684,N_7823);
and U8420 (N_8420,N_7722,N_7755);
nor U8421 (N_8421,N_7939,N_7617);
and U8422 (N_8422,N_7994,N_7594);
and U8423 (N_8423,N_7984,N_7885);
nand U8424 (N_8424,N_7919,N_7678);
and U8425 (N_8425,N_7783,N_7588);
or U8426 (N_8426,N_7571,N_7678);
and U8427 (N_8427,N_7555,N_7971);
nand U8428 (N_8428,N_7629,N_7765);
and U8429 (N_8429,N_7725,N_7843);
and U8430 (N_8430,N_7598,N_7967);
and U8431 (N_8431,N_7503,N_7765);
or U8432 (N_8432,N_7783,N_7764);
nor U8433 (N_8433,N_7916,N_7951);
or U8434 (N_8434,N_7974,N_7636);
nand U8435 (N_8435,N_7718,N_7636);
or U8436 (N_8436,N_7583,N_7721);
or U8437 (N_8437,N_7643,N_7583);
nor U8438 (N_8438,N_7702,N_7607);
or U8439 (N_8439,N_7556,N_7525);
nor U8440 (N_8440,N_7896,N_7607);
and U8441 (N_8441,N_7823,N_7765);
nand U8442 (N_8442,N_7650,N_7544);
xnor U8443 (N_8443,N_7675,N_7729);
nand U8444 (N_8444,N_7838,N_7981);
nand U8445 (N_8445,N_7815,N_7640);
or U8446 (N_8446,N_7550,N_7952);
and U8447 (N_8447,N_7908,N_7680);
and U8448 (N_8448,N_7769,N_7526);
nor U8449 (N_8449,N_7896,N_7742);
or U8450 (N_8450,N_7941,N_7736);
nand U8451 (N_8451,N_7783,N_7805);
or U8452 (N_8452,N_7538,N_7796);
and U8453 (N_8453,N_7976,N_7724);
nand U8454 (N_8454,N_7838,N_7697);
nand U8455 (N_8455,N_7591,N_7739);
and U8456 (N_8456,N_7601,N_7853);
or U8457 (N_8457,N_7560,N_7783);
nand U8458 (N_8458,N_7892,N_7674);
xor U8459 (N_8459,N_7750,N_7738);
nand U8460 (N_8460,N_7731,N_7596);
and U8461 (N_8461,N_7537,N_7785);
nor U8462 (N_8462,N_7510,N_7507);
or U8463 (N_8463,N_7841,N_7715);
nor U8464 (N_8464,N_7908,N_7667);
or U8465 (N_8465,N_7842,N_7878);
nor U8466 (N_8466,N_7539,N_7608);
nor U8467 (N_8467,N_7527,N_7823);
and U8468 (N_8468,N_7865,N_7578);
or U8469 (N_8469,N_7977,N_7824);
nor U8470 (N_8470,N_7675,N_7759);
nand U8471 (N_8471,N_7803,N_7638);
nand U8472 (N_8472,N_7518,N_7950);
or U8473 (N_8473,N_7649,N_7573);
and U8474 (N_8474,N_7586,N_7771);
nand U8475 (N_8475,N_7551,N_7576);
nor U8476 (N_8476,N_7705,N_7569);
or U8477 (N_8477,N_7714,N_7734);
and U8478 (N_8478,N_7608,N_7632);
and U8479 (N_8479,N_7504,N_7632);
or U8480 (N_8480,N_7793,N_7777);
nand U8481 (N_8481,N_7882,N_7586);
or U8482 (N_8482,N_7883,N_7973);
or U8483 (N_8483,N_7619,N_7757);
nor U8484 (N_8484,N_7920,N_7876);
nor U8485 (N_8485,N_7798,N_7881);
nand U8486 (N_8486,N_7857,N_7554);
nand U8487 (N_8487,N_7615,N_7583);
and U8488 (N_8488,N_7930,N_7590);
and U8489 (N_8489,N_7680,N_7970);
nand U8490 (N_8490,N_7993,N_7887);
nand U8491 (N_8491,N_7858,N_7924);
nor U8492 (N_8492,N_7544,N_7846);
or U8493 (N_8493,N_7847,N_7529);
nand U8494 (N_8494,N_7587,N_7795);
and U8495 (N_8495,N_7765,N_7972);
or U8496 (N_8496,N_7911,N_7501);
xnor U8497 (N_8497,N_7790,N_7797);
or U8498 (N_8498,N_7842,N_7821);
and U8499 (N_8499,N_7760,N_7609);
or U8500 (N_8500,N_8431,N_8054);
and U8501 (N_8501,N_8383,N_8402);
nor U8502 (N_8502,N_8022,N_8356);
nand U8503 (N_8503,N_8321,N_8488);
nor U8504 (N_8504,N_8025,N_8474);
or U8505 (N_8505,N_8213,N_8389);
or U8506 (N_8506,N_8490,N_8262);
or U8507 (N_8507,N_8297,N_8441);
nand U8508 (N_8508,N_8238,N_8481);
nand U8509 (N_8509,N_8151,N_8030);
nor U8510 (N_8510,N_8182,N_8335);
or U8511 (N_8511,N_8121,N_8156);
or U8512 (N_8512,N_8198,N_8485);
or U8513 (N_8513,N_8167,N_8011);
nand U8514 (N_8514,N_8100,N_8143);
nor U8515 (N_8515,N_8043,N_8077);
nand U8516 (N_8516,N_8308,N_8332);
nor U8517 (N_8517,N_8222,N_8426);
or U8518 (N_8518,N_8207,N_8371);
and U8519 (N_8519,N_8096,N_8309);
nand U8520 (N_8520,N_8217,N_8320);
nor U8521 (N_8521,N_8081,N_8031);
nor U8522 (N_8522,N_8073,N_8285);
nand U8523 (N_8523,N_8174,N_8419);
nand U8524 (N_8524,N_8427,N_8210);
or U8525 (N_8525,N_8161,N_8041);
and U8526 (N_8526,N_8010,N_8264);
or U8527 (N_8527,N_8429,N_8281);
or U8528 (N_8528,N_8467,N_8492);
and U8529 (N_8529,N_8317,N_8486);
xor U8530 (N_8530,N_8430,N_8433);
nand U8531 (N_8531,N_8456,N_8042);
or U8532 (N_8532,N_8432,N_8376);
nor U8533 (N_8533,N_8483,N_8224);
and U8534 (N_8534,N_8076,N_8196);
nand U8535 (N_8535,N_8423,N_8105);
nor U8536 (N_8536,N_8005,N_8300);
and U8537 (N_8537,N_8214,N_8450);
and U8538 (N_8538,N_8436,N_8428);
nor U8539 (N_8539,N_8183,N_8004);
nor U8540 (N_8540,N_8453,N_8494);
or U8541 (N_8541,N_8475,N_8491);
nor U8542 (N_8542,N_8219,N_8395);
xnor U8543 (N_8543,N_8235,N_8299);
or U8544 (N_8544,N_8024,N_8343);
nand U8545 (N_8545,N_8415,N_8471);
nand U8546 (N_8546,N_8406,N_8128);
nand U8547 (N_8547,N_8257,N_8344);
nor U8548 (N_8548,N_8284,N_8218);
or U8549 (N_8549,N_8117,N_8392);
or U8550 (N_8550,N_8129,N_8092);
nor U8551 (N_8551,N_8083,N_8190);
nor U8552 (N_8552,N_8480,N_8381);
nand U8553 (N_8553,N_8448,N_8245);
nor U8554 (N_8554,N_8122,N_8274);
nor U8555 (N_8555,N_8477,N_8202);
nor U8556 (N_8556,N_8236,N_8063);
and U8557 (N_8557,N_8241,N_8007);
nor U8558 (N_8558,N_8303,N_8412);
xnor U8559 (N_8559,N_8061,N_8240);
or U8560 (N_8560,N_8055,N_8345);
or U8561 (N_8561,N_8177,N_8331);
nor U8562 (N_8562,N_8290,N_8439);
and U8563 (N_8563,N_8329,N_8088);
nor U8564 (N_8564,N_8497,N_8114);
nand U8565 (N_8565,N_8282,N_8249);
nand U8566 (N_8566,N_8197,N_8112);
nor U8567 (N_8567,N_8360,N_8178);
xor U8568 (N_8568,N_8242,N_8124);
xnor U8569 (N_8569,N_8060,N_8409);
nor U8570 (N_8570,N_8141,N_8184);
and U8571 (N_8571,N_8237,N_8080);
and U8572 (N_8572,N_8154,N_8017);
and U8573 (N_8573,N_8460,N_8078);
or U8574 (N_8574,N_8449,N_8407);
or U8575 (N_8575,N_8194,N_8384);
or U8576 (N_8576,N_8358,N_8230);
and U8577 (N_8577,N_8386,N_8050);
or U8578 (N_8578,N_8153,N_8323);
or U8579 (N_8579,N_8387,N_8414);
or U8580 (N_8580,N_8341,N_8188);
nor U8581 (N_8581,N_8035,N_8038);
and U8582 (N_8582,N_8180,N_8164);
nor U8583 (N_8583,N_8029,N_8234);
nand U8584 (N_8584,N_8179,N_8337);
nand U8585 (N_8585,N_8283,N_8499);
and U8586 (N_8586,N_8053,N_8220);
nand U8587 (N_8587,N_8251,N_8075);
nor U8588 (N_8588,N_8438,N_8170);
nor U8589 (N_8589,N_8295,N_8094);
and U8590 (N_8590,N_8229,N_8287);
and U8591 (N_8591,N_8446,N_8142);
or U8592 (N_8592,N_8018,N_8452);
and U8593 (N_8593,N_8254,N_8150);
nand U8594 (N_8594,N_8113,N_8110);
nand U8595 (N_8595,N_8135,N_8347);
and U8596 (N_8596,N_8211,N_8292);
nor U8597 (N_8597,N_8447,N_8165);
or U8598 (N_8598,N_8391,N_8136);
or U8599 (N_8599,N_8399,N_8339);
nor U8600 (N_8600,N_8111,N_8044);
or U8601 (N_8601,N_8090,N_8362);
nand U8602 (N_8602,N_8148,N_8400);
nand U8603 (N_8603,N_8118,N_8328);
or U8604 (N_8604,N_8307,N_8418);
xnor U8605 (N_8605,N_8003,N_8032);
and U8606 (N_8606,N_8265,N_8016);
and U8607 (N_8607,N_8163,N_8420);
nand U8608 (N_8608,N_8026,N_8280);
or U8609 (N_8609,N_8372,N_8355);
nor U8610 (N_8610,N_8166,N_8116);
nand U8611 (N_8611,N_8106,N_8319);
and U8612 (N_8612,N_8181,N_8065);
nand U8613 (N_8613,N_8146,N_8187);
or U8614 (N_8614,N_8324,N_8175);
or U8615 (N_8615,N_8001,N_8057);
nand U8616 (N_8616,N_8186,N_8019);
nor U8617 (N_8617,N_8195,N_8313);
xor U8618 (N_8618,N_8401,N_8033);
or U8619 (N_8619,N_8298,N_8070);
and U8620 (N_8620,N_8336,N_8014);
nand U8621 (N_8621,N_8302,N_8394);
nand U8622 (N_8622,N_8278,N_8243);
and U8623 (N_8623,N_8396,N_8206);
or U8624 (N_8624,N_8463,N_8346);
nand U8625 (N_8625,N_8468,N_8440);
and U8626 (N_8626,N_8231,N_8072);
or U8627 (N_8627,N_8125,N_8479);
nand U8628 (N_8628,N_8259,N_8487);
nand U8629 (N_8629,N_8435,N_8006);
nor U8630 (N_8630,N_8442,N_8086);
or U8631 (N_8631,N_8204,N_8233);
and U8632 (N_8632,N_8484,N_8250);
or U8633 (N_8633,N_8404,N_8338);
and U8634 (N_8634,N_8424,N_8119);
nand U8635 (N_8635,N_8138,N_8169);
nor U8636 (N_8636,N_8279,N_8068);
nor U8637 (N_8637,N_8350,N_8097);
nand U8638 (N_8638,N_8104,N_8466);
nand U8639 (N_8639,N_8291,N_8342);
nor U8640 (N_8640,N_8253,N_8215);
and U8641 (N_8641,N_8311,N_8272);
nor U8642 (N_8642,N_8212,N_8256);
nand U8643 (N_8643,N_8465,N_8071);
nand U8644 (N_8644,N_8459,N_8246);
nor U8645 (N_8645,N_8315,N_8208);
nor U8646 (N_8646,N_8227,N_8422);
nor U8647 (N_8647,N_8417,N_8365);
or U8648 (N_8648,N_8421,N_8062);
or U8649 (N_8649,N_8380,N_8367);
or U8650 (N_8650,N_8353,N_8286);
nand U8651 (N_8651,N_8046,N_8333);
nor U8652 (N_8652,N_8489,N_8434);
nand U8653 (N_8653,N_8147,N_8464);
and U8654 (N_8654,N_8093,N_8205);
or U8655 (N_8655,N_8325,N_8352);
nand U8656 (N_8656,N_8275,N_8445);
or U8657 (N_8657,N_8144,N_8052);
nor U8658 (N_8658,N_8493,N_8277);
or U8659 (N_8659,N_8162,N_8454);
nand U8660 (N_8660,N_8469,N_8099);
nor U8661 (N_8661,N_8101,N_8051);
nor U8662 (N_8662,N_8095,N_8348);
nand U8663 (N_8663,N_8322,N_8223);
nand U8664 (N_8664,N_8133,N_8260);
or U8665 (N_8665,N_8388,N_8273);
nor U8666 (N_8666,N_8385,N_8091);
or U8667 (N_8667,N_8357,N_8327);
nor U8668 (N_8668,N_8203,N_8269);
or U8669 (N_8669,N_8403,N_8107);
or U8670 (N_8670,N_8377,N_8416);
nor U8671 (N_8671,N_8020,N_8296);
or U8672 (N_8672,N_8066,N_8495);
and U8673 (N_8673,N_8390,N_8168);
nand U8674 (N_8674,N_8301,N_8123);
or U8675 (N_8675,N_8034,N_8437);
and U8676 (N_8676,N_8199,N_8192);
or U8677 (N_8677,N_8410,N_8375);
and U8678 (N_8678,N_8036,N_8369);
and U8679 (N_8679,N_8149,N_8027);
and U8680 (N_8680,N_8015,N_8374);
xnor U8681 (N_8681,N_8310,N_8102);
nand U8682 (N_8682,N_8457,N_8461);
or U8683 (N_8683,N_8498,N_8189);
or U8684 (N_8684,N_8069,N_8000);
xor U8685 (N_8685,N_8047,N_8126);
and U8686 (N_8686,N_8330,N_8193);
nand U8687 (N_8687,N_8289,N_8370);
and U8688 (N_8688,N_8258,N_8462);
nand U8689 (N_8689,N_8228,N_8012);
and U8690 (N_8690,N_8002,N_8364);
or U8691 (N_8691,N_8132,N_8120);
nand U8692 (N_8692,N_8109,N_8158);
or U8693 (N_8693,N_8444,N_8455);
nand U8694 (N_8694,N_8306,N_8305);
and U8695 (N_8695,N_8361,N_8045);
nor U8696 (N_8696,N_8368,N_8293);
nor U8697 (N_8697,N_8255,N_8009);
or U8698 (N_8698,N_8160,N_8127);
xnor U8699 (N_8699,N_8201,N_8354);
and U8700 (N_8700,N_8288,N_8397);
nand U8701 (N_8701,N_8252,N_8185);
and U8702 (N_8702,N_8226,N_8244);
nand U8703 (N_8703,N_8021,N_8108);
or U8704 (N_8704,N_8039,N_8458);
or U8705 (N_8705,N_8173,N_8340);
nand U8706 (N_8706,N_8366,N_8470);
nor U8707 (N_8707,N_8191,N_8451);
nand U8708 (N_8708,N_8496,N_8349);
or U8709 (N_8709,N_8130,N_8155);
nor U8710 (N_8710,N_8326,N_8137);
and U8711 (N_8711,N_8267,N_8221);
nor U8712 (N_8712,N_8359,N_8037);
nand U8713 (N_8713,N_8408,N_8028);
and U8714 (N_8714,N_8134,N_8263);
and U8715 (N_8715,N_8040,N_8152);
or U8716 (N_8716,N_8312,N_8216);
nand U8717 (N_8717,N_8363,N_8476);
or U8718 (N_8718,N_8085,N_8131);
and U8719 (N_8719,N_8172,N_8266);
nor U8720 (N_8720,N_8139,N_8098);
nand U8721 (N_8721,N_8425,N_8393);
nor U8722 (N_8722,N_8314,N_8304);
or U8723 (N_8723,N_8008,N_8157);
or U8724 (N_8724,N_8074,N_8176);
nand U8725 (N_8725,N_8171,N_8232);
and U8726 (N_8726,N_8209,N_8318);
or U8727 (N_8727,N_8140,N_8067);
or U8728 (N_8728,N_8261,N_8023);
or U8729 (N_8729,N_8013,N_8351);
or U8730 (N_8730,N_8316,N_8482);
nor U8731 (N_8731,N_8048,N_8239);
and U8732 (N_8732,N_8443,N_8268);
nand U8733 (N_8733,N_8145,N_8225);
and U8734 (N_8734,N_8084,N_8378);
nand U8735 (N_8735,N_8115,N_8270);
or U8736 (N_8736,N_8334,N_8200);
and U8737 (N_8737,N_8056,N_8472);
nand U8738 (N_8738,N_8064,N_8059);
nand U8739 (N_8739,N_8159,N_8248);
nor U8740 (N_8740,N_8049,N_8276);
nor U8741 (N_8741,N_8373,N_8271);
nand U8742 (N_8742,N_8382,N_8473);
nand U8743 (N_8743,N_8089,N_8413);
nor U8744 (N_8744,N_8082,N_8087);
and U8745 (N_8745,N_8379,N_8478);
nand U8746 (N_8746,N_8411,N_8405);
or U8747 (N_8747,N_8294,N_8079);
nor U8748 (N_8748,N_8058,N_8103);
or U8749 (N_8749,N_8398,N_8247);
and U8750 (N_8750,N_8023,N_8193);
and U8751 (N_8751,N_8440,N_8019);
nand U8752 (N_8752,N_8281,N_8183);
and U8753 (N_8753,N_8346,N_8096);
nand U8754 (N_8754,N_8278,N_8301);
and U8755 (N_8755,N_8265,N_8338);
nand U8756 (N_8756,N_8474,N_8207);
nand U8757 (N_8757,N_8320,N_8150);
nor U8758 (N_8758,N_8002,N_8290);
nor U8759 (N_8759,N_8064,N_8085);
nand U8760 (N_8760,N_8381,N_8020);
or U8761 (N_8761,N_8138,N_8335);
or U8762 (N_8762,N_8407,N_8324);
or U8763 (N_8763,N_8021,N_8358);
nor U8764 (N_8764,N_8443,N_8413);
and U8765 (N_8765,N_8071,N_8198);
or U8766 (N_8766,N_8220,N_8175);
nor U8767 (N_8767,N_8084,N_8179);
nand U8768 (N_8768,N_8261,N_8443);
nor U8769 (N_8769,N_8355,N_8238);
nand U8770 (N_8770,N_8375,N_8359);
and U8771 (N_8771,N_8045,N_8123);
and U8772 (N_8772,N_8158,N_8411);
and U8773 (N_8773,N_8134,N_8027);
nand U8774 (N_8774,N_8024,N_8106);
nor U8775 (N_8775,N_8494,N_8293);
nand U8776 (N_8776,N_8021,N_8200);
and U8777 (N_8777,N_8172,N_8383);
or U8778 (N_8778,N_8133,N_8414);
or U8779 (N_8779,N_8435,N_8431);
and U8780 (N_8780,N_8263,N_8462);
nor U8781 (N_8781,N_8292,N_8499);
or U8782 (N_8782,N_8311,N_8313);
or U8783 (N_8783,N_8239,N_8149);
and U8784 (N_8784,N_8199,N_8083);
nor U8785 (N_8785,N_8180,N_8219);
and U8786 (N_8786,N_8208,N_8375);
and U8787 (N_8787,N_8220,N_8332);
nand U8788 (N_8788,N_8428,N_8116);
nor U8789 (N_8789,N_8291,N_8195);
nand U8790 (N_8790,N_8141,N_8466);
or U8791 (N_8791,N_8052,N_8264);
nand U8792 (N_8792,N_8142,N_8134);
nor U8793 (N_8793,N_8468,N_8025);
nand U8794 (N_8794,N_8411,N_8308);
and U8795 (N_8795,N_8040,N_8301);
nor U8796 (N_8796,N_8461,N_8046);
nor U8797 (N_8797,N_8176,N_8225);
nand U8798 (N_8798,N_8092,N_8473);
xor U8799 (N_8799,N_8407,N_8194);
and U8800 (N_8800,N_8406,N_8492);
nor U8801 (N_8801,N_8161,N_8219);
nor U8802 (N_8802,N_8401,N_8169);
or U8803 (N_8803,N_8304,N_8035);
nor U8804 (N_8804,N_8170,N_8332);
xor U8805 (N_8805,N_8185,N_8005);
nand U8806 (N_8806,N_8385,N_8474);
nor U8807 (N_8807,N_8373,N_8320);
or U8808 (N_8808,N_8421,N_8289);
nand U8809 (N_8809,N_8285,N_8320);
or U8810 (N_8810,N_8398,N_8404);
nand U8811 (N_8811,N_8163,N_8402);
or U8812 (N_8812,N_8398,N_8320);
nor U8813 (N_8813,N_8103,N_8109);
or U8814 (N_8814,N_8311,N_8385);
nand U8815 (N_8815,N_8054,N_8108);
and U8816 (N_8816,N_8185,N_8024);
nand U8817 (N_8817,N_8468,N_8471);
or U8818 (N_8818,N_8047,N_8422);
and U8819 (N_8819,N_8091,N_8109);
nor U8820 (N_8820,N_8015,N_8187);
and U8821 (N_8821,N_8205,N_8228);
nor U8822 (N_8822,N_8477,N_8237);
or U8823 (N_8823,N_8207,N_8282);
nor U8824 (N_8824,N_8406,N_8151);
or U8825 (N_8825,N_8198,N_8051);
or U8826 (N_8826,N_8463,N_8327);
nand U8827 (N_8827,N_8112,N_8341);
or U8828 (N_8828,N_8361,N_8231);
nand U8829 (N_8829,N_8225,N_8257);
nor U8830 (N_8830,N_8100,N_8337);
nand U8831 (N_8831,N_8200,N_8161);
nand U8832 (N_8832,N_8401,N_8056);
nand U8833 (N_8833,N_8009,N_8417);
or U8834 (N_8834,N_8264,N_8188);
nor U8835 (N_8835,N_8372,N_8447);
nand U8836 (N_8836,N_8037,N_8207);
nand U8837 (N_8837,N_8399,N_8473);
nand U8838 (N_8838,N_8496,N_8082);
or U8839 (N_8839,N_8120,N_8261);
nand U8840 (N_8840,N_8356,N_8074);
xor U8841 (N_8841,N_8499,N_8335);
or U8842 (N_8842,N_8246,N_8014);
or U8843 (N_8843,N_8498,N_8246);
nand U8844 (N_8844,N_8136,N_8283);
or U8845 (N_8845,N_8426,N_8371);
nand U8846 (N_8846,N_8181,N_8323);
and U8847 (N_8847,N_8470,N_8469);
and U8848 (N_8848,N_8154,N_8301);
nand U8849 (N_8849,N_8115,N_8154);
nand U8850 (N_8850,N_8273,N_8208);
and U8851 (N_8851,N_8237,N_8318);
nor U8852 (N_8852,N_8096,N_8200);
nand U8853 (N_8853,N_8328,N_8396);
nand U8854 (N_8854,N_8323,N_8129);
nor U8855 (N_8855,N_8065,N_8417);
nor U8856 (N_8856,N_8269,N_8058);
nor U8857 (N_8857,N_8483,N_8282);
nand U8858 (N_8858,N_8175,N_8070);
nor U8859 (N_8859,N_8321,N_8318);
and U8860 (N_8860,N_8330,N_8303);
or U8861 (N_8861,N_8339,N_8492);
nor U8862 (N_8862,N_8227,N_8168);
nand U8863 (N_8863,N_8267,N_8236);
or U8864 (N_8864,N_8492,N_8400);
or U8865 (N_8865,N_8194,N_8348);
nand U8866 (N_8866,N_8381,N_8317);
nor U8867 (N_8867,N_8303,N_8241);
and U8868 (N_8868,N_8294,N_8431);
nand U8869 (N_8869,N_8271,N_8217);
or U8870 (N_8870,N_8035,N_8051);
nand U8871 (N_8871,N_8463,N_8401);
and U8872 (N_8872,N_8099,N_8426);
nor U8873 (N_8873,N_8144,N_8296);
or U8874 (N_8874,N_8087,N_8468);
and U8875 (N_8875,N_8469,N_8298);
and U8876 (N_8876,N_8358,N_8407);
and U8877 (N_8877,N_8293,N_8180);
nand U8878 (N_8878,N_8387,N_8084);
nor U8879 (N_8879,N_8426,N_8410);
and U8880 (N_8880,N_8092,N_8497);
and U8881 (N_8881,N_8401,N_8170);
or U8882 (N_8882,N_8461,N_8128);
or U8883 (N_8883,N_8266,N_8135);
nand U8884 (N_8884,N_8023,N_8422);
or U8885 (N_8885,N_8044,N_8330);
and U8886 (N_8886,N_8470,N_8221);
or U8887 (N_8887,N_8088,N_8445);
or U8888 (N_8888,N_8044,N_8368);
or U8889 (N_8889,N_8167,N_8438);
and U8890 (N_8890,N_8039,N_8422);
or U8891 (N_8891,N_8136,N_8074);
nand U8892 (N_8892,N_8292,N_8254);
nand U8893 (N_8893,N_8184,N_8038);
or U8894 (N_8894,N_8208,N_8418);
or U8895 (N_8895,N_8237,N_8252);
nor U8896 (N_8896,N_8086,N_8178);
nand U8897 (N_8897,N_8123,N_8255);
or U8898 (N_8898,N_8350,N_8452);
nor U8899 (N_8899,N_8020,N_8423);
and U8900 (N_8900,N_8044,N_8120);
or U8901 (N_8901,N_8334,N_8085);
nand U8902 (N_8902,N_8475,N_8355);
and U8903 (N_8903,N_8344,N_8236);
or U8904 (N_8904,N_8365,N_8499);
or U8905 (N_8905,N_8213,N_8396);
or U8906 (N_8906,N_8056,N_8493);
and U8907 (N_8907,N_8316,N_8050);
nor U8908 (N_8908,N_8296,N_8045);
nor U8909 (N_8909,N_8213,N_8231);
nand U8910 (N_8910,N_8423,N_8319);
nand U8911 (N_8911,N_8092,N_8058);
nand U8912 (N_8912,N_8361,N_8114);
and U8913 (N_8913,N_8406,N_8211);
nand U8914 (N_8914,N_8082,N_8078);
nor U8915 (N_8915,N_8258,N_8125);
and U8916 (N_8916,N_8218,N_8363);
and U8917 (N_8917,N_8466,N_8406);
xnor U8918 (N_8918,N_8276,N_8039);
nand U8919 (N_8919,N_8049,N_8114);
nand U8920 (N_8920,N_8084,N_8057);
nand U8921 (N_8921,N_8262,N_8153);
or U8922 (N_8922,N_8067,N_8253);
and U8923 (N_8923,N_8317,N_8128);
and U8924 (N_8924,N_8479,N_8480);
nand U8925 (N_8925,N_8371,N_8027);
and U8926 (N_8926,N_8272,N_8033);
xor U8927 (N_8927,N_8095,N_8343);
nand U8928 (N_8928,N_8318,N_8180);
nor U8929 (N_8929,N_8022,N_8097);
nor U8930 (N_8930,N_8110,N_8097);
or U8931 (N_8931,N_8006,N_8092);
and U8932 (N_8932,N_8170,N_8191);
nand U8933 (N_8933,N_8437,N_8041);
nand U8934 (N_8934,N_8070,N_8074);
and U8935 (N_8935,N_8123,N_8303);
or U8936 (N_8936,N_8392,N_8032);
xor U8937 (N_8937,N_8217,N_8447);
nor U8938 (N_8938,N_8267,N_8111);
and U8939 (N_8939,N_8323,N_8131);
xor U8940 (N_8940,N_8024,N_8370);
xor U8941 (N_8941,N_8319,N_8291);
and U8942 (N_8942,N_8199,N_8093);
and U8943 (N_8943,N_8147,N_8498);
and U8944 (N_8944,N_8385,N_8402);
or U8945 (N_8945,N_8345,N_8198);
nand U8946 (N_8946,N_8345,N_8439);
nand U8947 (N_8947,N_8112,N_8236);
or U8948 (N_8948,N_8039,N_8441);
nor U8949 (N_8949,N_8336,N_8445);
nand U8950 (N_8950,N_8017,N_8102);
or U8951 (N_8951,N_8148,N_8450);
and U8952 (N_8952,N_8295,N_8175);
nand U8953 (N_8953,N_8199,N_8291);
nand U8954 (N_8954,N_8370,N_8366);
or U8955 (N_8955,N_8417,N_8125);
or U8956 (N_8956,N_8102,N_8319);
and U8957 (N_8957,N_8351,N_8413);
or U8958 (N_8958,N_8080,N_8403);
nand U8959 (N_8959,N_8416,N_8164);
and U8960 (N_8960,N_8282,N_8389);
or U8961 (N_8961,N_8179,N_8340);
or U8962 (N_8962,N_8155,N_8272);
nand U8963 (N_8963,N_8129,N_8040);
nor U8964 (N_8964,N_8039,N_8350);
or U8965 (N_8965,N_8316,N_8246);
nor U8966 (N_8966,N_8199,N_8078);
nand U8967 (N_8967,N_8344,N_8272);
or U8968 (N_8968,N_8088,N_8400);
and U8969 (N_8969,N_8012,N_8054);
or U8970 (N_8970,N_8158,N_8421);
nand U8971 (N_8971,N_8142,N_8343);
and U8972 (N_8972,N_8342,N_8222);
nand U8973 (N_8973,N_8381,N_8350);
nor U8974 (N_8974,N_8427,N_8443);
or U8975 (N_8975,N_8161,N_8013);
xor U8976 (N_8976,N_8357,N_8493);
nor U8977 (N_8977,N_8175,N_8225);
and U8978 (N_8978,N_8436,N_8290);
nand U8979 (N_8979,N_8016,N_8198);
nor U8980 (N_8980,N_8072,N_8425);
or U8981 (N_8981,N_8209,N_8059);
or U8982 (N_8982,N_8397,N_8322);
or U8983 (N_8983,N_8114,N_8016);
and U8984 (N_8984,N_8141,N_8304);
or U8985 (N_8985,N_8341,N_8485);
and U8986 (N_8986,N_8167,N_8405);
nand U8987 (N_8987,N_8096,N_8243);
nand U8988 (N_8988,N_8027,N_8143);
or U8989 (N_8989,N_8025,N_8306);
and U8990 (N_8990,N_8162,N_8493);
nand U8991 (N_8991,N_8376,N_8289);
nor U8992 (N_8992,N_8256,N_8159);
nand U8993 (N_8993,N_8056,N_8234);
or U8994 (N_8994,N_8035,N_8148);
nand U8995 (N_8995,N_8408,N_8285);
nor U8996 (N_8996,N_8229,N_8017);
nand U8997 (N_8997,N_8430,N_8134);
or U8998 (N_8998,N_8260,N_8353);
nand U8999 (N_8999,N_8286,N_8374);
nor U9000 (N_9000,N_8815,N_8951);
and U9001 (N_9001,N_8853,N_8554);
and U9002 (N_9002,N_8580,N_8878);
nand U9003 (N_9003,N_8811,N_8506);
nand U9004 (N_9004,N_8718,N_8573);
and U9005 (N_9005,N_8653,N_8774);
and U9006 (N_9006,N_8784,N_8533);
and U9007 (N_9007,N_8619,N_8953);
and U9008 (N_9008,N_8913,N_8621);
nand U9009 (N_9009,N_8876,N_8512);
and U9010 (N_9010,N_8682,N_8751);
nand U9011 (N_9011,N_8906,N_8730);
nor U9012 (N_9012,N_8907,N_8966);
nand U9013 (N_9013,N_8814,N_8846);
or U9014 (N_9014,N_8891,N_8689);
and U9015 (N_9015,N_8500,N_8786);
and U9016 (N_9016,N_8692,N_8635);
or U9017 (N_9017,N_8560,N_8690);
nor U9018 (N_9018,N_8838,N_8525);
or U9019 (N_9019,N_8510,N_8993);
or U9020 (N_9020,N_8927,N_8680);
and U9021 (N_9021,N_8531,N_8867);
nand U9022 (N_9022,N_8979,N_8916);
nand U9023 (N_9023,N_8647,N_8576);
nor U9024 (N_9024,N_8607,N_8930);
nand U9025 (N_9025,N_8545,N_8890);
nor U9026 (N_9026,N_8790,N_8669);
nand U9027 (N_9027,N_8941,N_8599);
xor U9028 (N_9028,N_8721,N_8870);
or U9029 (N_9029,N_8577,N_8818);
and U9030 (N_9030,N_8755,N_8613);
nor U9031 (N_9031,N_8741,N_8695);
and U9032 (N_9032,N_8671,N_8706);
or U9033 (N_9033,N_8723,N_8996);
or U9034 (N_9034,N_8978,N_8575);
or U9035 (N_9035,N_8881,N_8962);
nand U9036 (N_9036,N_8795,N_8681);
or U9037 (N_9037,N_8789,N_8845);
nand U9038 (N_9038,N_8571,N_8758);
or U9039 (N_9039,N_8851,N_8915);
or U9040 (N_9040,N_8807,N_8538);
or U9041 (N_9041,N_8606,N_8691);
and U9042 (N_9042,N_8685,N_8844);
nor U9043 (N_9043,N_8816,N_8519);
and U9044 (N_9044,N_8670,N_8787);
or U9045 (N_9045,N_8656,N_8587);
nand U9046 (N_9046,N_8964,N_8739);
nor U9047 (N_9047,N_8973,N_8518);
nand U9048 (N_9048,N_8642,N_8763);
and U9049 (N_9049,N_8707,N_8897);
or U9050 (N_9050,N_8508,N_8711);
and U9051 (N_9051,N_8804,N_8841);
nand U9052 (N_9052,N_8639,N_8667);
nor U9053 (N_9053,N_8968,N_8877);
nor U9054 (N_9054,N_8534,N_8646);
and U9055 (N_9055,N_8694,N_8826);
or U9056 (N_9056,N_8701,N_8684);
or U9057 (N_9057,N_8820,N_8805);
and U9058 (N_9058,N_8988,N_8539);
nand U9059 (N_9059,N_8875,N_8594);
or U9060 (N_9060,N_8698,N_8530);
nor U9061 (N_9061,N_8579,N_8984);
nand U9062 (N_9062,N_8572,N_8983);
and U9063 (N_9063,N_8798,N_8872);
or U9064 (N_9064,N_8586,N_8710);
or U9065 (N_9065,N_8618,N_8597);
or U9066 (N_9066,N_8803,N_8849);
nor U9067 (N_9067,N_8590,N_8552);
nand U9068 (N_9068,N_8967,N_8769);
nand U9069 (N_9069,N_8743,N_8555);
nor U9070 (N_9070,N_8731,N_8782);
nor U9071 (N_9071,N_8716,N_8839);
and U9072 (N_9072,N_8529,N_8605);
and U9073 (N_9073,N_8779,N_8777);
and U9074 (N_9074,N_8862,N_8677);
nor U9075 (N_9075,N_8655,N_8687);
or U9076 (N_9076,N_8693,N_8501);
nand U9077 (N_9077,N_8752,N_8727);
or U9078 (N_9078,N_8547,N_8935);
nor U9079 (N_9079,N_8869,N_8880);
and U9080 (N_9080,N_8612,N_8654);
or U9081 (N_9081,N_8809,N_8658);
nor U9082 (N_9082,N_8527,N_8821);
or U9083 (N_9083,N_8850,N_8792);
nand U9084 (N_9084,N_8517,N_8660);
nand U9085 (N_9085,N_8936,N_8550);
and U9086 (N_9086,N_8883,N_8626);
nor U9087 (N_9087,N_8651,N_8666);
and U9088 (N_9088,N_8793,N_8561);
xnor U9089 (N_9089,N_8834,N_8788);
nor U9090 (N_9090,N_8932,N_8643);
nor U9091 (N_9091,N_8929,N_8649);
nand U9092 (N_9092,N_8520,N_8753);
and U9093 (N_9093,N_8631,N_8969);
xor U9094 (N_9094,N_8761,N_8750);
nor U9095 (N_9095,N_8933,N_8662);
xor U9096 (N_9096,N_8937,N_8970);
and U9097 (N_9097,N_8956,N_8884);
nand U9098 (N_9098,N_8601,N_8514);
and U9099 (N_9099,N_8773,N_8900);
nand U9100 (N_9100,N_8823,N_8744);
nor U9101 (N_9101,N_8544,N_8732);
and U9102 (N_9102,N_8712,N_8641);
or U9103 (N_9103,N_8563,N_8912);
or U9104 (N_9104,N_8738,N_8630);
nand U9105 (N_9105,N_8725,N_8972);
nor U9106 (N_9106,N_8925,N_8570);
or U9107 (N_9107,N_8987,N_8663);
nand U9108 (N_9108,N_8934,N_8894);
or U9109 (N_9109,N_8617,N_8622);
nand U9110 (N_9110,N_8515,N_8719);
nand U9111 (N_9111,N_8802,N_8644);
or U9112 (N_9112,N_8896,N_8952);
nor U9113 (N_9113,N_8958,N_8700);
or U9114 (N_9114,N_8724,N_8675);
or U9115 (N_9115,N_8858,N_8855);
nand U9116 (N_9116,N_8990,N_8756);
nor U9117 (N_9117,N_8516,N_8715);
and U9118 (N_9118,N_8836,N_8829);
nand U9119 (N_9119,N_8847,N_8864);
or U9120 (N_9120,N_8977,N_8948);
nand U9121 (N_9121,N_8523,N_8961);
nor U9122 (N_9122,N_8888,N_8674);
and U9123 (N_9123,N_8922,N_8859);
and U9124 (N_9124,N_8528,N_8615);
and U9125 (N_9125,N_8553,N_8556);
nand U9126 (N_9126,N_8778,N_8817);
and U9127 (N_9127,N_8797,N_8709);
or U9128 (N_9128,N_8865,N_8551);
and U9129 (N_9129,N_8980,N_8524);
nor U9130 (N_9130,N_8567,N_8998);
or U9131 (N_9131,N_8708,N_8583);
nand U9132 (N_9132,N_8799,N_8887);
and U9133 (N_9133,N_8856,N_8986);
nand U9134 (N_9134,N_8808,N_8509);
or U9135 (N_9135,N_8852,N_8854);
or U9136 (N_9136,N_8697,N_8648);
nand U9137 (N_9137,N_8920,N_8960);
nor U9138 (N_9138,N_8566,N_8945);
nand U9139 (N_9139,N_8813,N_8747);
or U9140 (N_9140,N_8754,N_8584);
nand U9141 (N_9141,N_8558,N_8535);
nor U9142 (N_9142,N_8623,N_8810);
and U9143 (N_9143,N_8921,N_8637);
or U9144 (N_9144,N_8905,N_8735);
xor U9145 (N_9145,N_8636,N_8976);
nor U9146 (N_9146,N_8902,N_8603);
or U9147 (N_9147,N_8511,N_8947);
nand U9148 (N_9148,N_8893,N_8503);
and U9149 (N_9149,N_8745,N_8771);
and U9150 (N_9150,N_8557,N_8661);
and U9151 (N_9151,N_8624,N_8608);
and U9152 (N_9152,N_8889,N_8837);
and U9153 (N_9153,N_8997,N_8886);
nand U9154 (N_9154,N_8652,N_8938);
nor U9155 (N_9155,N_8819,N_8737);
nand U9156 (N_9156,N_8722,N_8806);
nor U9157 (N_9157,N_8720,N_8688);
and U9158 (N_9158,N_8513,N_8568);
nor U9159 (N_9159,N_8895,N_8703);
and U9160 (N_9160,N_8672,N_8908);
and U9161 (N_9161,N_8504,N_8713);
or U9162 (N_9162,N_8940,N_8542);
nor U9163 (N_9163,N_8673,N_8505);
xnor U9164 (N_9164,N_8831,N_8892);
nand U9165 (N_9165,N_8871,N_8914);
and U9166 (N_9166,N_8678,N_8863);
and U9167 (N_9167,N_8800,N_8794);
or U9168 (N_9168,N_8965,N_8885);
nand U9169 (N_9169,N_8759,N_8634);
nand U9170 (N_9170,N_8657,N_8911);
nand U9171 (N_9171,N_8546,N_8740);
or U9172 (N_9172,N_8593,N_8600);
and U9173 (N_9173,N_8981,N_8812);
or U9174 (N_9174,N_8704,N_8860);
and U9175 (N_9175,N_8832,N_8780);
and U9176 (N_9176,N_8581,N_8633);
or U9177 (N_9177,N_8757,N_8596);
or U9178 (N_9178,N_8668,N_8982);
or U9179 (N_9179,N_8705,N_8923);
and U9180 (N_9180,N_8588,N_8950);
nand U9181 (N_9181,N_8582,N_8791);
nor U9182 (N_9182,N_8928,N_8944);
or U9183 (N_9183,N_8949,N_8591);
or U9184 (N_9184,N_8765,N_8614);
nor U9185 (N_9185,N_8733,N_8861);
nor U9186 (N_9186,N_8868,N_8548);
nand U9187 (N_9187,N_8676,N_8772);
nor U9188 (N_9188,N_8776,N_8728);
or U9189 (N_9189,N_8574,N_8917);
or U9190 (N_9190,N_8843,N_8899);
nor U9191 (N_9191,N_8931,N_8526);
and U9192 (N_9192,N_8645,N_8729);
and U9193 (N_9193,N_8989,N_8760);
or U9194 (N_9194,N_8939,N_8842);
or U9195 (N_9195,N_8702,N_8541);
and U9196 (N_9196,N_8901,N_8746);
and U9197 (N_9197,N_8562,N_8540);
and U9198 (N_9198,N_8683,N_8873);
or U9199 (N_9199,N_8627,N_8971);
nand U9200 (N_9200,N_8659,N_8549);
xnor U9201 (N_9201,N_8611,N_8768);
and U9202 (N_9202,N_8717,N_8825);
or U9203 (N_9203,N_8762,N_8954);
nand U9204 (N_9204,N_8764,N_8848);
nor U9205 (N_9205,N_8946,N_8828);
and U9206 (N_9206,N_8866,N_8537);
or U9207 (N_9207,N_8699,N_8918);
and U9208 (N_9208,N_8609,N_8942);
nand U9209 (N_9209,N_8726,N_8628);
or U9210 (N_9210,N_8679,N_8963);
or U9211 (N_9211,N_8502,N_8665);
nand U9212 (N_9212,N_8734,N_8592);
nand U9213 (N_9213,N_8898,N_8830);
and U9214 (N_9214,N_8766,N_8833);
or U9215 (N_9215,N_8992,N_8974);
xor U9216 (N_9216,N_8955,N_8991);
or U9217 (N_9217,N_8714,N_8565);
and U9218 (N_9218,N_8569,N_8903);
nand U9219 (N_9219,N_8783,N_8785);
nor U9220 (N_9220,N_8824,N_8604);
and U9221 (N_9221,N_8632,N_8589);
or U9222 (N_9222,N_8598,N_8595);
or U9223 (N_9223,N_8521,N_8736);
nand U9224 (N_9224,N_8742,N_8924);
or U9225 (N_9225,N_8625,N_8959);
nor U9226 (N_9226,N_8985,N_8620);
nand U9227 (N_9227,N_8840,N_8994);
xor U9228 (N_9228,N_8522,N_8882);
nor U9229 (N_9229,N_8957,N_8796);
nor U9230 (N_9230,N_8532,N_8781);
nand U9231 (N_9231,N_8919,N_8904);
or U9232 (N_9232,N_8536,N_8564);
and U9233 (N_9233,N_8749,N_8696);
nor U9234 (N_9234,N_8638,N_8578);
nand U9235 (N_9235,N_8559,N_8926);
nor U9236 (N_9236,N_8543,N_8835);
or U9237 (N_9237,N_8664,N_8801);
nand U9238 (N_9238,N_8909,N_8602);
xnor U9239 (N_9239,N_8827,N_8610);
and U9240 (N_9240,N_8507,N_8640);
or U9241 (N_9241,N_8629,N_8879);
and U9242 (N_9242,N_8616,N_8770);
xnor U9243 (N_9243,N_8775,N_8975);
nor U9244 (N_9244,N_8767,N_8686);
or U9245 (N_9245,N_8943,N_8910);
and U9246 (N_9246,N_8822,N_8874);
nand U9247 (N_9247,N_8748,N_8585);
nand U9248 (N_9248,N_8857,N_8995);
and U9249 (N_9249,N_8999,N_8650);
nor U9250 (N_9250,N_8811,N_8844);
or U9251 (N_9251,N_8678,N_8506);
nand U9252 (N_9252,N_8723,N_8671);
nand U9253 (N_9253,N_8751,N_8738);
nor U9254 (N_9254,N_8833,N_8611);
nor U9255 (N_9255,N_8784,N_8632);
or U9256 (N_9256,N_8696,N_8505);
or U9257 (N_9257,N_8671,N_8597);
or U9258 (N_9258,N_8761,N_8725);
or U9259 (N_9259,N_8752,N_8744);
nand U9260 (N_9260,N_8599,N_8604);
and U9261 (N_9261,N_8642,N_8942);
or U9262 (N_9262,N_8703,N_8571);
or U9263 (N_9263,N_8803,N_8994);
nor U9264 (N_9264,N_8725,N_8658);
nand U9265 (N_9265,N_8688,N_8915);
or U9266 (N_9266,N_8726,N_8555);
and U9267 (N_9267,N_8540,N_8517);
or U9268 (N_9268,N_8540,N_8830);
or U9269 (N_9269,N_8991,N_8993);
nand U9270 (N_9270,N_8751,N_8834);
nor U9271 (N_9271,N_8661,N_8935);
nand U9272 (N_9272,N_8524,N_8780);
nor U9273 (N_9273,N_8907,N_8803);
nand U9274 (N_9274,N_8812,N_8817);
nor U9275 (N_9275,N_8905,N_8876);
or U9276 (N_9276,N_8908,N_8679);
or U9277 (N_9277,N_8902,N_8519);
xnor U9278 (N_9278,N_8650,N_8867);
nand U9279 (N_9279,N_8987,N_8574);
and U9280 (N_9280,N_8657,N_8547);
nand U9281 (N_9281,N_8663,N_8938);
nand U9282 (N_9282,N_8848,N_8843);
nor U9283 (N_9283,N_8540,N_8604);
nand U9284 (N_9284,N_8778,N_8689);
nor U9285 (N_9285,N_8889,N_8635);
or U9286 (N_9286,N_8769,N_8578);
or U9287 (N_9287,N_8630,N_8594);
or U9288 (N_9288,N_8785,N_8501);
and U9289 (N_9289,N_8778,N_8756);
xnor U9290 (N_9290,N_8624,N_8777);
or U9291 (N_9291,N_8549,N_8748);
nor U9292 (N_9292,N_8837,N_8611);
nor U9293 (N_9293,N_8912,N_8723);
nand U9294 (N_9294,N_8623,N_8672);
nand U9295 (N_9295,N_8985,N_8581);
xor U9296 (N_9296,N_8687,N_8959);
nand U9297 (N_9297,N_8567,N_8861);
nand U9298 (N_9298,N_8928,N_8756);
xnor U9299 (N_9299,N_8967,N_8822);
nor U9300 (N_9300,N_8508,N_8838);
nor U9301 (N_9301,N_8559,N_8755);
nor U9302 (N_9302,N_8813,N_8701);
nor U9303 (N_9303,N_8678,N_8782);
and U9304 (N_9304,N_8594,N_8705);
nand U9305 (N_9305,N_8660,N_8583);
or U9306 (N_9306,N_8530,N_8598);
nor U9307 (N_9307,N_8978,N_8835);
nand U9308 (N_9308,N_8851,N_8725);
nor U9309 (N_9309,N_8814,N_8813);
xor U9310 (N_9310,N_8853,N_8914);
and U9311 (N_9311,N_8577,N_8533);
or U9312 (N_9312,N_8971,N_8905);
nand U9313 (N_9313,N_8939,N_8979);
nand U9314 (N_9314,N_8874,N_8901);
or U9315 (N_9315,N_8864,N_8576);
and U9316 (N_9316,N_8867,N_8989);
and U9317 (N_9317,N_8956,N_8540);
nor U9318 (N_9318,N_8900,N_8834);
nor U9319 (N_9319,N_8828,N_8656);
xnor U9320 (N_9320,N_8844,N_8718);
and U9321 (N_9321,N_8884,N_8559);
or U9322 (N_9322,N_8722,N_8628);
or U9323 (N_9323,N_8680,N_8533);
nand U9324 (N_9324,N_8982,N_8554);
nor U9325 (N_9325,N_8668,N_8930);
nand U9326 (N_9326,N_8944,N_8852);
nor U9327 (N_9327,N_8680,N_8777);
nor U9328 (N_9328,N_8729,N_8542);
or U9329 (N_9329,N_8623,N_8924);
or U9330 (N_9330,N_8739,N_8820);
and U9331 (N_9331,N_8641,N_8827);
nand U9332 (N_9332,N_8625,N_8742);
and U9333 (N_9333,N_8623,N_8973);
nand U9334 (N_9334,N_8938,N_8911);
or U9335 (N_9335,N_8914,N_8992);
or U9336 (N_9336,N_8607,N_8769);
or U9337 (N_9337,N_8862,N_8867);
and U9338 (N_9338,N_8958,N_8906);
or U9339 (N_9339,N_8711,N_8855);
or U9340 (N_9340,N_8553,N_8709);
and U9341 (N_9341,N_8602,N_8875);
or U9342 (N_9342,N_8675,N_8959);
nand U9343 (N_9343,N_8776,N_8963);
nor U9344 (N_9344,N_8573,N_8737);
xor U9345 (N_9345,N_8596,N_8788);
nor U9346 (N_9346,N_8667,N_8790);
or U9347 (N_9347,N_8904,N_8622);
nand U9348 (N_9348,N_8703,N_8614);
nor U9349 (N_9349,N_8895,N_8915);
and U9350 (N_9350,N_8867,N_8919);
nand U9351 (N_9351,N_8717,N_8939);
nor U9352 (N_9352,N_8520,N_8735);
and U9353 (N_9353,N_8618,N_8527);
nand U9354 (N_9354,N_8708,N_8504);
and U9355 (N_9355,N_8584,N_8523);
xnor U9356 (N_9356,N_8613,N_8820);
and U9357 (N_9357,N_8527,N_8712);
and U9358 (N_9358,N_8668,N_8900);
nand U9359 (N_9359,N_8589,N_8870);
and U9360 (N_9360,N_8526,N_8661);
nor U9361 (N_9361,N_8921,N_8608);
nand U9362 (N_9362,N_8710,N_8754);
or U9363 (N_9363,N_8895,N_8612);
nand U9364 (N_9364,N_8842,N_8700);
nor U9365 (N_9365,N_8617,N_8676);
or U9366 (N_9366,N_8709,N_8808);
or U9367 (N_9367,N_8820,N_8643);
and U9368 (N_9368,N_8687,N_8789);
xor U9369 (N_9369,N_8966,N_8691);
xnor U9370 (N_9370,N_8856,N_8803);
or U9371 (N_9371,N_8684,N_8582);
or U9372 (N_9372,N_8904,N_8894);
nand U9373 (N_9373,N_8654,N_8671);
or U9374 (N_9374,N_8762,N_8899);
and U9375 (N_9375,N_8789,N_8864);
and U9376 (N_9376,N_8848,N_8932);
nand U9377 (N_9377,N_8776,N_8745);
and U9378 (N_9378,N_8573,N_8760);
and U9379 (N_9379,N_8862,N_8935);
or U9380 (N_9380,N_8507,N_8957);
nor U9381 (N_9381,N_8752,N_8892);
nand U9382 (N_9382,N_8797,N_8901);
and U9383 (N_9383,N_8993,N_8669);
nand U9384 (N_9384,N_8550,N_8881);
or U9385 (N_9385,N_8856,N_8795);
nor U9386 (N_9386,N_8775,N_8529);
nand U9387 (N_9387,N_8837,N_8530);
and U9388 (N_9388,N_8675,N_8533);
nand U9389 (N_9389,N_8551,N_8986);
and U9390 (N_9390,N_8638,N_8866);
nand U9391 (N_9391,N_8709,N_8594);
or U9392 (N_9392,N_8607,N_8547);
nor U9393 (N_9393,N_8673,N_8541);
or U9394 (N_9394,N_8963,N_8869);
and U9395 (N_9395,N_8535,N_8524);
or U9396 (N_9396,N_8876,N_8907);
xor U9397 (N_9397,N_8668,N_8827);
nand U9398 (N_9398,N_8875,N_8758);
xor U9399 (N_9399,N_8885,N_8970);
nor U9400 (N_9400,N_8855,N_8597);
nand U9401 (N_9401,N_8951,N_8878);
or U9402 (N_9402,N_8955,N_8894);
nor U9403 (N_9403,N_8912,N_8610);
xnor U9404 (N_9404,N_8772,N_8755);
nand U9405 (N_9405,N_8982,N_8962);
and U9406 (N_9406,N_8856,N_8651);
or U9407 (N_9407,N_8762,N_8508);
and U9408 (N_9408,N_8723,N_8993);
or U9409 (N_9409,N_8571,N_8975);
nand U9410 (N_9410,N_8865,N_8656);
nor U9411 (N_9411,N_8603,N_8897);
or U9412 (N_9412,N_8668,N_8673);
and U9413 (N_9413,N_8832,N_8818);
and U9414 (N_9414,N_8613,N_8887);
and U9415 (N_9415,N_8823,N_8778);
or U9416 (N_9416,N_8752,N_8715);
nand U9417 (N_9417,N_8958,N_8855);
nand U9418 (N_9418,N_8684,N_8618);
or U9419 (N_9419,N_8840,N_8930);
nor U9420 (N_9420,N_8549,N_8566);
nand U9421 (N_9421,N_8744,N_8929);
nor U9422 (N_9422,N_8870,N_8525);
nor U9423 (N_9423,N_8925,N_8595);
nand U9424 (N_9424,N_8930,N_8578);
nor U9425 (N_9425,N_8777,N_8945);
or U9426 (N_9426,N_8911,N_8773);
and U9427 (N_9427,N_8625,N_8637);
nor U9428 (N_9428,N_8756,N_8972);
or U9429 (N_9429,N_8708,N_8636);
and U9430 (N_9430,N_8573,N_8539);
nand U9431 (N_9431,N_8830,N_8984);
nand U9432 (N_9432,N_8953,N_8954);
nand U9433 (N_9433,N_8822,N_8533);
or U9434 (N_9434,N_8888,N_8948);
nand U9435 (N_9435,N_8880,N_8801);
or U9436 (N_9436,N_8707,N_8761);
nand U9437 (N_9437,N_8698,N_8755);
or U9438 (N_9438,N_8928,N_8613);
and U9439 (N_9439,N_8773,N_8698);
or U9440 (N_9440,N_8684,N_8659);
and U9441 (N_9441,N_8514,N_8579);
and U9442 (N_9442,N_8976,N_8941);
and U9443 (N_9443,N_8792,N_8581);
nor U9444 (N_9444,N_8776,N_8983);
nor U9445 (N_9445,N_8570,N_8837);
or U9446 (N_9446,N_8664,N_8739);
or U9447 (N_9447,N_8589,N_8826);
nor U9448 (N_9448,N_8852,N_8962);
or U9449 (N_9449,N_8793,N_8931);
and U9450 (N_9450,N_8659,N_8510);
or U9451 (N_9451,N_8890,N_8913);
nand U9452 (N_9452,N_8674,N_8743);
nand U9453 (N_9453,N_8867,N_8810);
nand U9454 (N_9454,N_8739,N_8628);
or U9455 (N_9455,N_8912,N_8858);
nand U9456 (N_9456,N_8635,N_8708);
and U9457 (N_9457,N_8810,N_8551);
nor U9458 (N_9458,N_8836,N_8958);
nand U9459 (N_9459,N_8717,N_8722);
and U9460 (N_9460,N_8791,N_8799);
nor U9461 (N_9461,N_8577,N_8780);
nor U9462 (N_9462,N_8570,N_8718);
or U9463 (N_9463,N_8515,N_8830);
and U9464 (N_9464,N_8552,N_8712);
nor U9465 (N_9465,N_8713,N_8549);
nor U9466 (N_9466,N_8599,N_8913);
nor U9467 (N_9467,N_8768,N_8998);
or U9468 (N_9468,N_8649,N_8841);
and U9469 (N_9469,N_8733,N_8826);
or U9470 (N_9470,N_8566,N_8902);
nand U9471 (N_9471,N_8560,N_8946);
and U9472 (N_9472,N_8622,N_8738);
nor U9473 (N_9473,N_8938,N_8948);
nand U9474 (N_9474,N_8522,N_8806);
nand U9475 (N_9475,N_8942,N_8676);
nor U9476 (N_9476,N_8780,N_8766);
or U9477 (N_9477,N_8611,N_8671);
and U9478 (N_9478,N_8625,N_8888);
or U9479 (N_9479,N_8648,N_8993);
nor U9480 (N_9480,N_8623,N_8990);
or U9481 (N_9481,N_8806,N_8606);
or U9482 (N_9482,N_8711,N_8787);
nor U9483 (N_9483,N_8788,N_8512);
or U9484 (N_9484,N_8789,N_8744);
and U9485 (N_9485,N_8989,N_8591);
or U9486 (N_9486,N_8648,N_8949);
or U9487 (N_9487,N_8879,N_8752);
xor U9488 (N_9488,N_8620,N_8943);
nand U9489 (N_9489,N_8505,N_8902);
and U9490 (N_9490,N_8822,N_8582);
xnor U9491 (N_9491,N_8530,N_8792);
nand U9492 (N_9492,N_8921,N_8982);
and U9493 (N_9493,N_8546,N_8601);
nand U9494 (N_9494,N_8735,N_8997);
nand U9495 (N_9495,N_8764,N_8830);
nand U9496 (N_9496,N_8579,N_8893);
or U9497 (N_9497,N_8844,N_8964);
or U9498 (N_9498,N_8794,N_8614);
or U9499 (N_9499,N_8886,N_8607);
nor U9500 (N_9500,N_9203,N_9478);
nand U9501 (N_9501,N_9108,N_9315);
and U9502 (N_9502,N_9363,N_9089);
and U9503 (N_9503,N_9157,N_9133);
nand U9504 (N_9504,N_9248,N_9291);
nor U9505 (N_9505,N_9126,N_9498);
nand U9506 (N_9506,N_9264,N_9098);
and U9507 (N_9507,N_9343,N_9025);
nor U9508 (N_9508,N_9198,N_9464);
nor U9509 (N_9509,N_9068,N_9290);
nand U9510 (N_9510,N_9451,N_9204);
or U9511 (N_9511,N_9445,N_9336);
and U9512 (N_9512,N_9265,N_9365);
or U9513 (N_9513,N_9218,N_9328);
and U9514 (N_9514,N_9069,N_9073);
or U9515 (N_9515,N_9286,N_9135);
nand U9516 (N_9516,N_9128,N_9253);
and U9517 (N_9517,N_9407,N_9003);
nor U9518 (N_9518,N_9058,N_9035);
and U9519 (N_9519,N_9314,N_9334);
nand U9520 (N_9520,N_9102,N_9260);
nand U9521 (N_9521,N_9495,N_9105);
nor U9522 (N_9522,N_9369,N_9360);
nor U9523 (N_9523,N_9059,N_9116);
or U9524 (N_9524,N_9014,N_9245);
nor U9525 (N_9525,N_9016,N_9100);
or U9526 (N_9526,N_9139,N_9483);
or U9527 (N_9527,N_9084,N_9443);
nand U9528 (N_9528,N_9417,N_9404);
nor U9529 (N_9529,N_9351,N_9431);
nor U9530 (N_9530,N_9474,N_9392);
nand U9531 (N_9531,N_9383,N_9330);
nor U9532 (N_9532,N_9389,N_9430);
or U9533 (N_9533,N_9130,N_9352);
nor U9534 (N_9534,N_9162,N_9145);
and U9535 (N_9535,N_9302,N_9391);
nand U9536 (N_9536,N_9030,N_9226);
nor U9537 (N_9537,N_9420,N_9465);
or U9538 (N_9538,N_9358,N_9042);
and U9539 (N_9539,N_9038,N_9082);
nor U9540 (N_9540,N_9412,N_9378);
and U9541 (N_9541,N_9409,N_9236);
and U9542 (N_9542,N_9246,N_9466);
nand U9543 (N_9543,N_9463,N_9201);
or U9544 (N_9544,N_9239,N_9213);
nor U9545 (N_9545,N_9421,N_9097);
or U9546 (N_9546,N_9310,N_9040);
or U9547 (N_9547,N_9103,N_9499);
nand U9548 (N_9548,N_9010,N_9029);
nand U9549 (N_9549,N_9002,N_9374);
nand U9550 (N_9550,N_9362,N_9340);
and U9551 (N_9551,N_9078,N_9312);
nand U9552 (N_9552,N_9008,N_9087);
nand U9553 (N_9553,N_9491,N_9284);
and U9554 (N_9554,N_9159,N_9454);
and U9555 (N_9555,N_9181,N_9151);
nand U9556 (N_9556,N_9037,N_9234);
or U9557 (N_9557,N_9080,N_9196);
nand U9558 (N_9558,N_9429,N_9482);
or U9559 (N_9559,N_9229,N_9199);
and U9560 (N_9560,N_9366,N_9207);
or U9561 (N_9561,N_9044,N_9469);
xor U9562 (N_9562,N_9049,N_9023);
and U9563 (N_9563,N_9188,N_9109);
nand U9564 (N_9564,N_9018,N_9261);
and U9565 (N_9565,N_9273,N_9320);
and U9566 (N_9566,N_9259,N_9416);
nand U9567 (N_9567,N_9467,N_9479);
nor U9568 (N_9568,N_9460,N_9311);
xnor U9569 (N_9569,N_9047,N_9174);
and U9570 (N_9570,N_9275,N_9364);
or U9571 (N_9571,N_9442,N_9410);
nand U9572 (N_9572,N_9424,N_9013);
or U9573 (N_9573,N_9461,N_9077);
or U9574 (N_9574,N_9447,N_9434);
and U9575 (N_9575,N_9137,N_9227);
xnor U9576 (N_9576,N_9076,N_9490);
xnor U9577 (N_9577,N_9413,N_9161);
nand U9578 (N_9578,N_9393,N_9222);
and U9579 (N_9579,N_9233,N_9398);
nand U9580 (N_9580,N_9317,N_9147);
or U9581 (N_9581,N_9371,N_9171);
nor U9582 (N_9582,N_9271,N_9052);
nor U9583 (N_9583,N_9156,N_9172);
or U9584 (N_9584,N_9473,N_9210);
or U9585 (N_9585,N_9325,N_9493);
and U9586 (N_9586,N_9436,N_9160);
nor U9587 (N_9587,N_9326,N_9173);
or U9588 (N_9588,N_9065,N_9285);
or U9589 (N_9589,N_9004,N_9165);
nor U9590 (N_9590,N_9193,N_9197);
nand U9591 (N_9591,N_9152,N_9452);
nor U9592 (N_9592,N_9045,N_9486);
or U9593 (N_9593,N_9090,N_9191);
and U9594 (N_9594,N_9075,N_9299);
or U9595 (N_9595,N_9418,N_9309);
or U9596 (N_9596,N_9220,N_9189);
or U9597 (N_9597,N_9323,N_9146);
nor U9598 (N_9598,N_9489,N_9113);
or U9599 (N_9599,N_9319,N_9051);
nor U9600 (N_9600,N_9142,N_9341);
nand U9601 (N_9601,N_9295,N_9215);
nand U9602 (N_9602,N_9119,N_9433);
or U9603 (N_9603,N_9367,N_9294);
and U9604 (N_9604,N_9263,N_9122);
and U9605 (N_9605,N_9432,N_9110);
or U9606 (N_9606,N_9235,N_9257);
nand U9607 (N_9607,N_9106,N_9379);
nor U9608 (N_9608,N_9307,N_9107);
nor U9609 (N_9609,N_9134,N_9279);
nand U9610 (N_9610,N_9214,N_9179);
nand U9611 (N_9611,N_9141,N_9048);
and U9612 (N_9612,N_9439,N_9373);
xor U9613 (N_9613,N_9095,N_9096);
and U9614 (N_9614,N_9268,N_9459);
nand U9615 (N_9615,N_9298,N_9305);
nand U9616 (N_9616,N_9468,N_9167);
nand U9617 (N_9617,N_9306,N_9154);
nand U9618 (N_9618,N_9209,N_9335);
or U9619 (N_9619,N_9123,N_9289);
xor U9620 (N_9620,N_9249,N_9377);
nand U9621 (N_9621,N_9282,N_9480);
nor U9622 (N_9622,N_9175,N_9150);
nand U9623 (N_9623,N_9015,N_9354);
nand U9624 (N_9624,N_9450,N_9355);
or U9625 (N_9625,N_9212,N_9276);
nand U9626 (N_9626,N_9384,N_9496);
xor U9627 (N_9627,N_9301,N_9455);
nor U9628 (N_9628,N_9205,N_9375);
or U9629 (N_9629,N_9357,N_9308);
or U9630 (N_9630,N_9094,N_9485);
nor U9631 (N_9631,N_9085,N_9091);
nand U9632 (N_9632,N_9125,N_9086);
nand U9633 (N_9633,N_9056,N_9347);
nand U9634 (N_9634,N_9402,N_9032);
and U9635 (N_9635,N_9074,N_9121);
and U9636 (N_9636,N_9405,N_9148);
and U9637 (N_9637,N_9243,N_9269);
and U9638 (N_9638,N_9435,N_9192);
or U9639 (N_9639,N_9297,N_9345);
and U9640 (N_9640,N_9111,N_9267);
nand U9641 (N_9641,N_9228,N_9440);
nor U9642 (N_9642,N_9338,N_9396);
nor U9643 (N_9643,N_9067,N_9054);
nand U9644 (N_9644,N_9170,N_9427);
nor U9645 (N_9645,N_9361,N_9024);
and U9646 (N_9646,N_9129,N_9380);
nand U9647 (N_9647,N_9006,N_9072);
or U9648 (N_9648,N_9168,N_9441);
nor U9649 (N_9649,N_9288,N_9066);
nor U9650 (N_9650,N_9333,N_9019);
and U9651 (N_9651,N_9419,N_9316);
nor U9652 (N_9652,N_9254,N_9005);
nand U9653 (N_9653,N_9287,N_9132);
or U9654 (N_9654,N_9428,N_9256);
nor U9655 (N_9655,N_9444,N_9231);
or U9656 (N_9656,N_9406,N_9446);
and U9657 (N_9657,N_9438,N_9426);
or U9658 (N_9658,N_9223,N_9200);
or U9659 (N_9659,N_9020,N_9356);
nand U9660 (N_9660,N_9258,N_9055);
xnor U9661 (N_9661,N_9472,N_9448);
nand U9662 (N_9662,N_9488,N_9349);
and U9663 (N_9663,N_9124,N_9031);
or U9664 (N_9664,N_9017,N_9244);
and U9665 (N_9665,N_9386,N_9131);
nor U9666 (N_9666,N_9061,N_9158);
and U9667 (N_9667,N_9322,N_9321);
nand U9668 (N_9668,N_9092,N_9115);
or U9669 (N_9669,N_9238,N_9292);
and U9670 (N_9670,N_9456,N_9053);
nand U9671 (N_9671,N_9471,N_9190);
nand U9672 (N_9672,N_9118,N_9324);
or U9673 (N_9673,N_9346,N_9021);
and U9674 (N_9674,N_9387,N_9169);
nor U9675 (N_9675,N_9232,N_9164);
and U9676 (N_9676,N_9280,N_9225);
and U9677 (N_9677,N_9117,N_9425);
nor U9678 (N_9678,N_9270,N_9143);
nor U9679 (N_9679,N_9182,N_9381);
nor U9680 (N_9680,N_9337,N_9114);
or U9681 (N_9681,N_9043,N_9327);
and U9682 (N_9682,N_9492,N_9033);
nand U9683 (N_9683,N_9195,N_9278);
nand U9684 (N_9684,N_9394,N_9136);
nor U9685 (N_9685,N_9070,N_9453);
nand U9686 (N_9686,N_9385,N_9187);
or U9687 (N_9687,N_9081,N_9178);
or U9688 (N_9688,N_9208,N_9339);
or U9689 (N_9689,N_9240,N_9415);
or U9690 (N_9690,N_9303,N_9217);
nor U9691 (N_9691,N_9206,N_9283);
or U9692 (N_9692,N_9138,N_9060);
or U9693 (N_9693,N_9390,N_9046);
nor U9694 (N_9694,N_9332,N_9120);
nor U9695 (N_9695,N_9202,N_9057);
nand U9696 (N_9696,N_9153,N_9370);
nor U9697 (N_9697,N_9481,N_9062);
nand U9698 (N_9698,N_9350,N_9494);
and U9699 (N_9699,N_9101,N_9462);
and U9700 (N_9700,N_9408,N_9183);
or U9701 (N_9701,N_9262,N_9083);
or U9702 (N_9702,N_9422,N_9359);
nor U9703 (N_9703,N_9304,N_9423);
or U9704 (N_9704,N_9399,N_9009);
nor U9705 (N_9705,N_9104,N_9274);
and U9706 (N_9706,N_9112,N_9027);
nand U9707 (N_9707,N_9255,N_9395);
and U9708 (N_9708,N_9397,N_9140);
nor U9709 (N_9709,N_9093,N_9272);
nand U9710 (N_9710,N_9484,N_9458);
or U9711 (N_9711,N_9237,N_9149);
and U9712 (N_9712,N_9388,N_9039);
or U9713 (N_9713,N_9219,N_9007);
nand U9714 (N_9714,N_9403,N_9224);
nand U9715 (N_9715,N_9034,N_9176);
nand U9716 (N_9716,N_9368,N_9247);
or U9717 (N_9717,N_9250,N_9252);
nand U9718 (N_9718,N_9001,N_9266);
and U9719 (N_9719,N_9382,N_9437);
nor U9720 (N_9720,N_9163,N_9088);
or U9721 (N_9721,N_9318,N_9475);
nand U9722 (N_9722,N_9186,N_9230);
nand U9723 (N_9723,N_9411,N_9194);
nor U9724 (N_9724,N_9180,N_9071);
or U9725 (N_9725,N_9353,N_9127);
xor U9726 (N_9726,N_9177,N_9036);
nor U9727 (N_9727,N_9476,N_9216);
nor U9728 (N_9728,N_9022,N_9155);
nor U9729 (N_9729,N_9011,N_9041);
nor U9730 (N_9730,N_9331,N_9050);
and U9731 (N_9731,N_9144,N_9251);
nor U9732 (N_9732,N_9185,N_9342);
nor U9733 (N_9733,N_9064,N_9281);
and U9734 (N_9734,N_9221,N_9063);
nand U9735 (N_9735,N_9012,N_9344);
nor U9736 (N_9736,N_9372,N_9242);
nand U9737 (N_9737,N_9477,N_9400);
or U9738 (N_9738,N_9211,N_9470);
and U9739 (N_9739,N_9313,N_9166);
and U9740 (N_9740,N_9497,N_9487);
or U9741 (N_9741,N_9028,N_9401);
nand U9742 (N_9742,N_9329,N_9300);
nand U9743 (N_9743,N_9277,N_9414);
or U9744 (N_9744,N_9000,N_9026);
nand U9745 (N_9745,N_9296,N_9184);
and U9746 (N_9746,N_9449,N_9099);
and U9747 (N_9747,N_9293,N_9079);
xnor U9748 (N_9748,N_9348,N_9376);
or U9749 (N_9749,N_9241,N_9457);
nor U9750 (N_9750,N_9306,N_9446);
or U9751 (N_9751,N_9488,N_9246);
or U9752 (N_9752,N_9108,N_9455);
nor U9753 (N_9753,N_9424,N_9174);
nor U9754 (N_9754,N_9426,N_9459);
xnor U9755 (N_9755,N_9324,N_9404);
or U9756 (N_9756,N_9083,N_9462);
and U9757 (N_9757,N_9008,N_9423);
and U9758 (N_9758,N_9480,N_9107);
nor U9759 (N_9759,N_9410,N_9005);
and U9760 (N_9760,N_9176,N_9240);
nand U9761 (N_9761,N_9371,N_9168);
nand U9762 (N_9762,N_9292,N_9415);
nand U9763 (N_9763,N_9062,N_9089);
nor U9764 (N_9764,N_9119,N_9023);
nor U9765 (N_9765,N_9211,N_9101);
or U9766 (N_9766,N_9494,N_9303);
and U9767 (N_9767,N_9120,N_9169);
nand U9768 (N_9768,N_9099,N_9243);
and U9769 (N_9769,N_9216,N_9096);
and U9770 (N_9770,N_9311,N_9066);
nand U9771 (N_9771,N_9355,N_9283);
nand U9772 (N_9772,N_9056,N_9296);
and U9773 (N_9773,N_9434,N_9101);
or U9774 (N_9774,N_9231,N_9311);
or U9775 (N_9775,N_9128,N_9158);
nor U9776 (N_9776,N_9248,N_9256);
nand U9777 (N_9777,N_9478,N_9037);
nor U9778 (N_9778,N_9340,N_9281);
and U9779 (N_9779,N_9120,N_9168);
nand U9780 (N_9780,N_9003,N_9307);
nor U9781 (N_9781,N_9013,N_9365);
and U9782 (N_9782,N_9411,N_9193);
and U9783 (N_9783,N_9165,N_9096);
nor U9784 (N_9784,N_9007,N_9157);
xor U9785 (N_9785,N_9112,N_9010);
or U9786 (N_9786,N_9194,N_9313);
and U9787 (N_9787,N_9177,N_9317);
or U9788 (N_9788,N_9434,N_9317);
nand U9789 (N_9789,N_9201,N_9065);
nor U9790 (N_9790,N_9402,N_9006);
and U9791 (N_9791,N_9084,N_9263);
or U9792 (N_9792,N_9006,N_9351);
nand U9793 (N_9793,N_9373,N_9217);
and U9794 (N_9794,N_9019,N_9031);
and U9795 (N_9795,N_9019,N_9396);
nor U9796 (N_9796,N_9175,N_9279);
and U9797 (N_9797,N_9488,N_9347);
or U9798 (N_9798,N_9033,N_9152);
and U9799 (N_9799,N_9130,N_9243);
and U9800 (N_9800,N_9332,N_9440);
and U9801 (N_9801,N_9271,N_9100);
and U9802 (N_9802,N_9479,N_9356);
and U9803 (N_9803,N_9036,N_9481);
nand U9804 (N_9804,N_9448,N_9326);
nor U9805 (N_9805,N_9044,N_9205);
or U9806 (N_9806,N_9222,N_9424);
nand U9807 (N_9807,N_9050,N_9083);
and U9808 (N_9808,N_9274,N_9414);
nor U9809 (N_9809,N_9090,N_9247);
nand U9810 (N_9810,N_9282,N_9286);
nor U9811 (N_9811,N_9236,N_9242);
nor U9812 (N_9812,N_9276,N_9423);
nand U9813 (N_9813,N_9366,N_9260);
or U9814 (N_9814,N_9248,N_9302);
or U9815 (N_9815,N_9142,N_9109);
or U9816 (N_9816,N_9354,N_9450);
nand U9817 (N_9817,N_9315,N_9409);
nor U9818 (N_9818,N_9248,N_9052);
and U9819 (N_9819,N_9264,N_9191);
nand U9820 (N_9820,N_9066,N_9354);
or U9821 (N_9821,N_9308,N_9491);
or U9822 (N_9822,N_9315,N_9457);
and U9823 (N_9823,N_9094,N_9071);
and U9824 (N_9824,N_9403,N_9480);
nand U9825 (N_9825,N_9006,N_9366);
or U9826 (N_9826,N_9185,N_9290);
or U9827 (N_9827,N_9321,N_9252);
or U9828 (N_9828,N_9286,N_9416);
and U9829 (N_9829,N_9432,N_9477);
nor U9830 (N_9830,N_9224,N_9106);
nor U9831 (N_9831,N_9213,N_9081);
nor U9832 (N_9832,N_9486,N_9017);
or U9833 (N_9833,N_9370,N_9296);
and U9834 (N_9834,N_9456,N_9207);
and U9835 (N_9835,N_9048,N_9302);
and U9836 (N_9836,N_9006,N_9305);
and U9837 (N_9837,N_9060,N_9092);
nor U9838 (N_9838,N_9488,N_9227);
nor U9839 (N_9839,N_9002,N_9360);
and U9840 (N_9840,N_9233,N_9095);
nor U9841 (N_9841,N_9445,N_9206);
or U9842 (N_9842,N_9155,N_9107);
nor U9843 (N_9843,N_9368,N_9424);
nor U9844 (N_9844,N_9369,N_9332);
or U9845 (N_9845,N_9131,N_9019);
nor U9846 (N_9846,N_9454,N_9274);
nor U9847 (N_9847,N_9137,N_9206);
nand U9848 (N_9848,N_9015,N_9440);
nand U9849 (N_9849,N_9159,N_9008);
nor U9850 (N_9850,N_9179,N_9368);
nor U9851 (N_9851,N_9167,N_9173);
and U9852 (N_9852,N_9420,N_9008);
nand U9853 (N_9853,N_9296,N_9447);
nand U9854 (N_9854,N_9308,N_9181);
nor U9855 (N_9855,N_9294,N_9311);
and U9856 (N_9856,N_9099,N_9399);
and U9857 (N_9857,N_9097,N_9153);
nand U9858 (N_9858,N_9081,N_9191);
nand U9859 (N_9859,N_9039,N_9233);
nand U9860 (N_9860,N_9291,N_9191);
nor U9861 (N_9861,N_9426,N_9361);
nand U9862 (N_9862,N_9138,N_9443);
or U9863 (N_9863,N_9324,N_9122);
or U9864 (N_9864,N_9314,N_9013);
nor U9865 (N_9865,N_9141,N_9000);
nor U9866 (N_9866,N_9413,N_9417);
nand U9867 (N_9867,N_9242,N_9070);
nand U9868 (N_9868,N_9426,N_9454);
and U9869 (N_9869,N_9388,N_9181);
nand U9870 (N_9870,N_9142,N_9139);
xnor U9871 (N_9871,N_9425,N_9015);
nand U9872 (N_9872,N_9477,N_9031);
and U9873 (N_9873,N_9103,N_9303);
and U9874 (N_9874,N_9348,N_9054);
nand U9875 (N_9875,N_9064,N_9065);
or U9876 (N_9876,N_9045,N_9397);
nor U9877 (N_9877,N_9314,N_9484);
nand U9878 (N_9878,N_9256,N_9132);
and U9879 (N_9879,N_9431,N_9201);
and U9880 (N_9880,N_9452,N_9307);
nor U9881 (N_9881,N_9413,N_9129);
nand U9882 (N_9882,N_9401,N_9407);
and U9883 (N_9883,N_9044,N_9134);
nand U9884 (N_9884,N_9385,N_9401);
or U9885 (N_9885,N_9248,N_9231);
nor U9886 (N_9886,N_9221,N_9248);
and U9887 (N_9887,N_9079,N_9066);
and U9888 (N_9888,N_9196,N_9182);
nand U9889 (N_9889,N_9304,N_9378);
nor U9890 (N_9890,N_9177,N_9176);
or U9891 (N_9891,N_9213,N_9386);
nand U9892 (N_9892,N_9278,N_9461);
nor U9893 (N_9893,N_9126,N_9228);
nand U9894 (N_9894,N_9265,N_9171);
xor U9895 (N_9895,N_9069,N_9445);
nor U9896 (N_9896,N_9007,N_9414);
xor U9897 (N_9897,N_9328,N_9070);
or U9898 (N_9898,N_9266,N_9221);
nand U9899 (N_9899,N_9396,N_9411);
and U9900 (N_9900,N_9273,N_9130);
and U9901 (N_9901,N_9265,N_9211);
nor U9902 (N_9902,N_9011,N_9245);
nand U9903 (N_9903,N_9235,N_9460);
nor U9904 (N_9904,N_9247,N_9005);
nand U9905 (N_9905,N_9397,N_9169);
or U9906 (N_9906,N_9232,N_9456);
or U9907 (N_9907,N_9493,N_9454);
or U9908 (N_9908,N_9020,N_9360);
nor U9909 (N_9909,N_9431,N_9202);
or U9910 (N_9910,N_9262,N_9410);
or U9911 (N_9911,N_9065,N_9121);
nand U9912 (N_9912,N_9122,N_9468);
xnor U9913 (N_9913,N_9302,N_9115);
nor U9914 (N_9914,N_9483,N_9218);
and U9915 (N_9915,N_9152,N_9050);
nand U9916 (N_9916,N_9176,N_9402);
or U9917 (N_9917,N_9151,N_9266);
or U9918 (N_9918,N_9031,N_9108);
nand U9919 (N_9919,N_9272,N_9157);
or U9920 (N_9920,N_9292,N_9059);
xnor U9921 (N_9921,N_9270,N_9243);
nor U9922 (N_9922,N_9079,N_9255);
and U9923 (N_9923,N_9050,N_9088);
nor U9924 (N_9924,N_9245,N_9222);
nor U9925 (N_9925,N_9444,N_9001);
nor U9926 (N_9926,N_9038,N_9183);
and U9927 (N_9927,N_9101,N_9189);
nor U9928 (N_9928,N_9208,N_9418);
and U9929 (N_9929,N_9284,N_9431);
or U9930 (N_9930,N_9165,N_9187);
and U9931 (N_9931,N_9051,N_9088);
and U9932 (N_9932,N_9035,N_9120);
or U9933 (N_9933,N_9448,N_9363);
or U9934 (N_9934,N_9244,N_9169);
nand U9935 (N_9935,N_9188,N_9043);
xor U9936 (N_9936,N_9374,N_9352);
and U9937 (N_9937,N_9133,N_9092);
xnor U9938 (N_9938,N_9273,N_9411);
or U9939 (N_9939,N_9207,N_9278);
nor U9940 (N_9940,N_9031,N_9050);
nor U9941 (N_9941,N_9499,N_9377);
nor U9942 (N_9942,N_9430,N_9282);
or U9943 (N_9943,N_9247,N_9020);
nor U9944 (N_9944,N_9250,N_9205);
and U9945 (N_9945,N_9336,N_9027);
nor U9946 (N_9946,N_9045,N_9369);
nor U9947 (N_9947,N_9161,N_9213);
and U9948 (N_9948,N_9043,N_9273);
or U9949 (N_9949,N_9255,N_9324);
and U9950 (N_9950,N_9034,N_9238);
and U9951 (N_9951,N_9155,N_9004);
and U9952 (N_9952,N_9467,N_9294);
nor U9953 (N_9953,N_9168,N_9313);
nand U9954 (N_9954,N_9431,N_9207);
nand U9955 (N_9955,N_9283,N_9392);
or U9956 (N_9956,N_9288,N_9430);
nor U9957 (N_9957,N_9463,N_9171);
nand U9958 (N_9958,N_9050,N_9419);
nor U9959 (N_9959,N_9279,N_9264);
and U9960 (N_9960,N_9434,N_9072);
nor U9961 (N_9961,N_9000,N_9001);
xor U9962 (N_9962,N_9091,N_9164);
and U9963 (N_9963,N_9440,N_9182);
and U9964 (N_9964,N_9340,N_9405);
or U9965 (N_9965,N_9051,N_9283);
nor U9966 (N_9966,N_9017,N_9404);
nand U9967 (N_9967,N_9343,N_9183);
or U9968 (N_9968,N_9291,N_9363);
or U9969 (N_9969,N_9247,N_9029);
nor U9970 (N_9970,N_9173,N_9484);
nor U9971 (N_9971,N_9410,N_9306);
nand U9972 (N_9972,N_9383,N_9143);
nand U9973 (N_9973,N_9154,N_9225);
and U9974 (N_9974,N_9227,N_9110);
or U9975 (N_9975,N_9189,N_9171);
or U9976 (N_9976,N_9195,N_9130);
or U9977 (N_9977,N_9043,N_9040);
nor U9978 (N_9978,N_9023,N_9232);
nand U9979 (N_9979,N_9117,N_9489);
nand U9980 (N_9980,N_9424,N_9203);
nor U9981 (N_9981,N_9129,N_9356);
or U9982 (N_9982,N_9245,N_9387);
or U9983 (N_9983,N_9175,N_9314);
xnor U9984 (N_9984,N_9097,N_9493);
nor U9985 (N_9985,N_9318,N_9465);
or U9986 (N_9986,N_9009,N_9385);
or U9987 (N_9987,N_9052,N_9024);
nand U9988 (N_9988,N_9111,N_9372);
nor U9989 (N_9989,N_9356,N_9463);
nor U9990 (N_9990,N_9309,N_9099);
nor U9991 (N_9991,N_9124,N_9375);
and U9992 (N_9992,N_9402,N_9206);
and U9993 (N_9993,N_9486,N_9265);
and U9994 (N_9994,N_9022,N_9300);
and U9995 (N_9995,N_9268,N_9448);
and U9996 (N_9996,N_9360,N_9361);
and U9997 (N_9997,N_9214,N_9407);
or U9998 (N_9998,N_9471,N_9384);
nor U9999 (N_9999,N_9430,N_9022);
nand UO_0 (O_0,N_9851,N_9967);
and UO_1 (O_1,N_9711,N_9556);
and UO_2 (O_2,N_9715,N_9905);
or UO_3 (O_3,N_9525,N_9870);
nand UO_4 (O_4,N_9922,N_9679);
and UO_5 (O_5,N_9942,N_9595);
nor UO_6 (O_6,N_9583,N_9939);
nor UO_7 (O_7,N_9551,N_9815);
and UO_8 (O_8,N_9926,N_9607);
and UO_9 (O_9,N_9896,N_9878);
xnor UO_10 (O_10,N_9672,N_9512);
and UO_11 (O_11,N_9566,N_9991);
and UO_12 (O_12,N_9837,N_9532);
nor UO_13 (O_13,N_9568,N_9986);
and UO_14 (O_14,N_9919,N_9988);
nor UO_15 (O_15,N_9874,N_9659);
nand UO_16 (O_16,N_9574,N_9542);
nand UO_17 (O_17,N_9807,N_9702);
nand UO_18 (O_18,N_9884,N_9695);
nand UO_19 (O_19,N_9803,N_9906);
or UO_20 (O_20,N_9801,N_9567);
nor UO_21 (O_21,N_9880,N_9845);
or UO_22 (O_22,N_9752,N_9839);
or UO_23 (O_23,N_9721,N_9510);
nand UO_24 (O_24,N_9786,N_9971);
nor UO_25 (O_25,N_9630,N_9766);
xnor UO_26 (O_26,N_9718,N_9722);
nand UO_27 (O_27,N_9740,N_9825);
and UO_28 (O_28,N_9745,N_9917);
and UO_29 (O_29,N_9920,N_9729);
or UO_30 (O_30,N_9563,N_9758);
nand UO_31 (O_31,N_9938,N_9788);
and UO_32 (O_32,N_9844,N_9879);
nand UO_33 (O_33,N_9523,N_9555);
nor UO_34 (O_34,N_9772,N_9559);
and UO_35 (O_35,N_9966,N_9632);
or UO_36 (O_36,N_9813,N_9753);
and UO_37 (O_37,N_9611,N_9980);
nor UO_38 (O_38,N_9822,N_9950);
or UO_39 (O_39,N_9618,N_9796);
nor UO_40 (O_40,N_9639,N_9638);
and UO_41 (O_41,N_9776,N_9903);
and UO_42 (O_42,N_9626,N_9981);
nor UO_43 (O_43,N_9856,N_9731);
or UO_44 (O_44,N_9734,N_9936);
or UO_45 (O_45,N_9570,N_9828);
nor UO_46 (O_46,N_9516,N_9744);
or UO_47 (O_47,N_9562,N_9940);
and UO_48 (O_48,N_9558,N_9673);
and UO_49 (O_49,N_9661,N_9560);
nand UO_50 (O_50,N_9928,N_9543);
nor UO_51 (O_51,N_9864,N_9687);
xor UO_52 (O_52,N_9961,N_9685);
nor UO_53 (O_53,N_9746,N_9533);
and UO_54 (O_54,N_9728,N_9930);
and UO_55 (O_55,N_9932,N_9860);
nand UO_56 (O_56,N_9812,N_9688);
nor UO_57 (O_57,N_9600,N_9763);
and UO_58 (O_58,N_9750,N_9598);
or UO_59 (O_59,N_9768,N_9976);
nand UO_60 (O_60,N_9927,N_9652);
and UO_61 (O_61,N_9571,N_9973);
nand UO_62 (O_62,N_9624,N_9762);
or UO_63 (O_63,N_9765,N_9604);
nand UO_64 (O_64,N_9877,N_9992);
and UO_65 (O_65,N_9526,N_9984);
nor UO_66 (O_66,N_9968,N_9601);
nand UO_67 (O_67,N_9830,N_9777);
nor UO_68 (O_68,N_9681,N_9590);
nand UO_69 (O_69,N_9804,N_9811);
xor UO_70 (O_70,N_9535,N_9857);
nor UO_71 (O_71,N_9540,N_9941);
and UO_72 (O_72,N_9736,N_9541);
or UO_73 (O_73,N_9682,N_9960);
nand UO_74 (O_74,N_9627,N_9569);
and UO_75 (O_75,N_9519,N_9954);
nor UO_76 (O_76,N_9871,N_9893);
and UO_77 (O_77,N_9667,N_9645);
and UO_78 (O_78,N_9521,N_9594);
or UO_79 (O_79,N_9838,N_9931);
nor UO_80 (O_80,N_9584,N_9955);
or UO_81 (O_81,N_9885,N_9974);
or UO_82 (O_82,N_9572,N_9633);
and UO_83 (O_83,N_9610,N_9764);
xnor UO_84 (O_84,N_9958,N_9527);
xnor UO_85 (O_85,N_9622,N_9602);
nand UO_86 (O_86,N_9806,N_9505);
or UO_87 (O_87,N_9802,N_9642);
nor UO_88 (O_88,N_9897,N_9701);
or UO_89 (O_89,N_9552,N_9738);
or UO_90 (O_90,N_9588,N_9609);
and UO_91 (O_91,N_9910,N_9710);
nand UO_92 (O_92,N_9534,N_9599);
and UO_93 (O_93,N_9888,N_9606);
and UO_94 (O_94,N_9538,N_9635);
nand UO_95 (O_95,N_9749,N_9727);
and UO_96 (O_96,N_9504,N_9756);
nand UO_97 (O_97,N_9741,N_9883);
nor UO_98 (O_98,N_9615,N_9929);
or UO_99 (O_99,N_9677,N_9909);
nor UO_100 (O_100,N_9720,N_9904);
nand UO_101 (O_101,N_9549,N_9557);
and UO_102 (O_102,N_9712,N_9952);
or UO_103 (O_103,N_9513,N_9999);
nor UO_104 (O_104,N_9500,N_9658);
and UO_105 (O_105,N_9531,N_9996);
nand UO_106 (O_106,N_9869,N_9537);
or UO_107 (O_107,N_9735,N_9664);
nand UO_108 (O_108,N_9789,N_9503);
and UO_109 (O_109,N_9704,N_9824);
and UO_110 (O_110,N_9994,N_9656);
nor UO_111 (O_111,N_9732,N_9587);
nand UO_112 (O_112,N_9548,N_9866);
and UO_113 (O_113,N_9956,N_9683);
nand UO_114 (O_114,N_9945,N_9608);
nand UO_115 (O_115,N_9779,N_9717);
and UO_116 (O_116,N_9643,N_9675);
nor UO_117 (O_117,N_9709,N_9751);
nand UO_118 (O_118,N_9511,N_9809);
nor UO_119 (O_119,N_9816,N_9889);
or UO_120 (O_120,N_9619,N_9835);
and UO_121 (O_121,N_9647,N_9891);
or UO_122 (O_122,N_9923,N_9585);
and UO_123 (O_123,N_9631,N_9546);
and UO_124 (O_124,N_9817,N_9733);
nor UO_125 (O_125,N_9694,N_9578);
nand UO_126 (O_126,N_9553,N_9660);
and UO_127 (O_127,N_9818,N_9849);
or UO_128 (O_128,N_9530,N_9629);
nand UO_129 (O_129,N_9865,N_9653);
nor UO_130 (O_130,N_9693,N_9573);
nor UO_131 (O_131,N_9654,N_9515);
nor UO_132 (O_132,N_9621,N_9843);
nor UO_133 (O_133,N_9946,N_9550);
and UO_134 (O_134,N_9565,N_9886);
nor UO_135 (O_135,N_9640,N_9684);
and UO_136 (O_136,N_9668,N_9924);
nand UO_137 (O_137,N_9862,N_9698);
or UO_138 (O_138,N_9547,N_9714);
nand UO_139 (O_139,N_9603,N_9759);
or UO_140 (O_140,N_9616,N_9649);
nor UO_141 (O_141,N_9873,N_9648);
nor UO_142 (O_142,N_9666,N_9713);
and UO_143 (O_143,N_9620,N_9754);
nor UO_144 (O_144,N_9514,N_9554);
nand UO_145 (O_145,N_9576,N_9970);
or UO_146 (O_146,N_9771,N_9742);
and UO_147 (O_147,N_9882,N_9876);
and UO_148 (O_148,N_9861,N_9783);
or UO_149 (O_149,N_9833,N_9948);
or UO_150 (O_150,N_9794,N_9858);
nand UO_151 (O_151,N_9937,N_9502);
and UO_152 (O_152,N_9841,N_9826);
or UO_153 (O_153,N_9935,N_9774);
and UO_154 (O_154,N_9614,N_9997);
or UO_155 (O_155,N_9819,N_9591);
and UO_156 (O_156,N_9852,N_9898);
nand UO_157 (O_157,N_9953,N_9726);
nor UO_158 (O_158,N_9536,N_9760);
or UO_159 (O_159,N_9651,N_9829);
or UO_160 (O_160,N_9978,N_9918);
nand UO_161 (O_161,N_9969,N_9612);
nand UO_162 (O_162,N_9707,N_9690);
nor UO_163 (O_163,N_9730,N_9821);
and UO_164 (O_164,N_9650,N_9747);
and UO_165 (O_165,N_9799,N_9827);
nand UO_166 (O_166,N_9853,N_9655);
and UO_167 (O_167,N_9773,N_9913);
or UO_168 (O_168,N_9529,N_9674);
and UO_169 (O_169,N_9517,N_9872);
and UO_170 (O_170,N_9979,N_9831);
or UO_171 (O_171,N_9575,N_9805);
or UO_172 (O_172,N_9580,N_9739);
or UO_173 (O_173,N_9743,N_9680);
or UO_174 (O_174,N_9561,N_9868);
nor UO_175 (O_175,N_9703,N_9507);
or UO_176 (O_176,N_9990,N_9723);
nor UO_177 (O_177,N_9669,N_9637);
nor UO_178 (O_178,N_9836,N_9592);
nand UO_179 (O_179,N_9800,N_9847);
and UO_180 (O_180,N_9863,N_9911);
or UO_181 (O_181,N_9784,N_9887);
or UO_182 (O_182,N_9636,N_9613);
or UO_183 (O_183,N_9597,N_9671);
nor UO_184 (O_184,N_9808,N_9899);
or UO_185 (O_185,N_9989,N_9943);
nor UO_186 (O_186,N_9983,N_9907);
nor UO_187 (O_187,N_9686,N_9780);
and UO_188 (O_188,N_9716,N_9725);
xnor UO_189 (O_189,N_9892,N_9848);
nand UO_190 (O_190,N_9933,N_9975);
nor UO_191 (O_191,N_9957,N_9963);
xnor UO_192 (O_192,N_9798,N_9908);
nand UO_193 (O_193,N_9628,N_9834);
nand UO_194 (O_194,N_9987,N_9964);
nor UO_195 (O_195,N_9947,N_9916);
and UO_196 (O_196,N_9881,N_9501);
nand UO_197 (O_197,N_9593,N_9708);
nor UO_198 (O_198,N_9625,N_9782);
or UO_199 (O_199,N_9663,N_9965);
xnor UO_200 (O_200,N_9700,N_9901);
xnor UO_201 (O_201,N_9737,N_9770);
and UO_202 (O_202,N_9854,N_9912);
or UO_203 (O_203,N_9528,N_9579);
nand UO_204 (O_204,N_9775,N_9509);
and UO_205 (O_205,N_9691,N_9644);
nand UO_206 (O_206,N_9596,N_9670);
nor UO_207 (O_207,N_9544,N_9586);
nand UO_208 (O_208,N_9724,N_9894);
and UO_209 (O_209,N_9855,N_9859);
and UO_210 (O_210,N_9769,N_9832);
and UO_211 (O_211,N_9895,N_9900);
nand UO_212 (O_212,N_9944,N_9785);
and UO_213 (O_213,N_9890,N_9914);
nor UO_214 (O_214,N_9617,N_9761);
or UO_215 (O_215,N_9689,N_9792);
xor UO_216 (O_216,N_9995,N_9634);
or UO_217 (O_217,N_9678,N_9959);
and UO_218 (O_218,N_9706,N_9524);
nor UO_219 (O_219,N_9767,N_9696);
or UO_220 (O_220,N_9539,N_9699);
nand UO_221 (O_221,N_9820,N_9623);
and UO_222 (O_222,N_9795,N_9787);
nand UO_223 (O_223,N_9814,N_9577);
nand UO_224 (O_224,N_9646,N_9705);
and UO_225 (O_225,N_9949,N_9697);
nor UO_226 (O_226,N_9605,N_9921);
and UO_227 (O_227,N_9810,N_9793);
and UO_228 (O_228,N_9520,N_9676);
nand UO_229 (O_229,N_9840,N_9962);
nor UO_230 (O_230,N_9993,N_9951);
nand UO_231 (O_231,N_9915,N_9823);
nor UO_232 (O_232,N_9934,N_9985);
nor UO_233 (O_233,N_9972,N_9902);
nand UO_234 (O_234,N_9665,N_9564);
or UO_235 (O_235,N_9757,N_9977);
or UO_236 (O_236,N_9581,N_9518);
and UO_237 (O_237,N_9790,N_9508);
or UO_238 (O_238,N_9850,N_9582);
nand UO_239 (O_239,N_9781,N_9842);
and UO_240 (O_240,N_9692,N_9797);
and UO_241 (O_241,N_9755,N_9998);
nor UO_242 (O_242,N_9846,N_9867);
nand UO_243 (O_243,N_9778,N_9545);
and UO_244 (O_244,N_9506,N_9875);
and UO_245 (O_245,N_9791,N_9662);
or UO_246 (O_246,N_9982,N_9925);
nor UO_247 (O_247,N_9641,N_9719);
or UO_248 (O_248,N_9748,N_9522);
and UO_249 (O_249,N_9589,N_9657);
nor UO_250 (O_250,N_9885,N_9637);
or UO_251 (O_251,N_9519,N_9910);
nand UO_252 (O_252,N_9859,N_9871);
nand UO_253 (O_253,N_9830,N_9537);
nor UO_254 (O_254,N_9955,N_9848);
nand UO_255 (O_255,N_9722,N_9790);
and UO_256 (O_256,N_9604,N_9569);
or UO_257 (O_257,N_9773,N_9640);
and UO_258 (O_258,N_9697,N_9561);
or UO_259 (O_259,N_9990,N_9589);
and UO_260 (O_260,N_9939,N_9905);
nor UO_261 (O_261,N_9939,N_9669);
nor UO_262 (O_262,N_9502,N_9736);
and UO_263 (O_263,N_9957,N_9549);
nand UO_264 (O_264,N_9802,N_9710);
and UO_265 (O_265,N_9787,N_9623);
nor UO_266 (O_266,N_9725,N_9529);
nor UO_267 (O_267,N_9799,N_9683);
nor UO_268 (O_268,N_9723,N_9598);
nand UO_269 (O_269,N_9612,N_9679);
nand UO_270 (O_270,N_9883,N_9978);
and UO_271 (O_271,N_9502,N_9572);
or UO_272 (O_272,N_9859,N_9914);
nand UO_273 (O_273,N_9586,N_9516);
nand UO_274 (O_274,N_9559,N_9568);
or UO_275 (O_275,N_9953,N_9709);
or UO_276 (O_276,N_9922,N_9633);
or UO_277 (O_277,N_9745,N_9584);
and UO_278 (O_278,N_9713,N_9711);
nor UO_279 (O_279,N_9955,N_9527);
nor UO_280 (O_280,N_9882,N_9878);
and UO_281 (O_281,N_9879,N_9968);
and UO_282 (O_282,N_9974,N_9534);
and UO_283 (O_283,N_9536,N_9588);
and UO_284 (O_284,N_9780,N_9510);
nand UO_285 (O_285,N_9752,N_9754);
nand UO_286 (O_286,N_9844,N_9672);
or UO_287 (O_287,N_9820,N_9501);
and UO_288 (O_288,N_9677,N_9563);
nor UO_289 (O_289,N_9687,N_9636);
or UO_290 (O_290,N_9993,N_9610);
xnor UO_291 (O_291,N_9583,N_9618);
or UO_292 (O_292,N_9615,N_9851);
nor UO_293 (O_293,N_9966,N_9799);
nor UO_294 (O_294,N_9905,N_9526);
and UO_295 (O_295,N_9878,N_9541);
nor UO_296 (O_296,N_9929,N_9693);
nor UO_297 (O_297,N_9502,N_9957);
nor UO_298 (O_298,N_9781,N_9827);
nor UO_299 (O_299,N_9598,N_9552);
or UO_300 (O_300,N_9726,N_9912);
nand UO_301 (O_301,N_9808,N_9854);
nand UO_302 (O_302,N_9866,N_9847);
nor UO_303 (O_303,N_9914,N_9955);
nor UO_304 (O_304,N_9527,N_9588);
and UO_305 (O_305,N_9711,N_9591);
nor UO_306 (O_306,N_9588,N_9525);
or UO_307 (O_307,N_9725,N_9878);
or UO_308 (O_308,N_9874,N_9689);
and UO_309 (O_309,N_9516,N_9794);
and UO_310 (O_310,N_9678,N_9638);
and UO_311 (O_311,N_9698,N_9963);
and UO_312 (O_312,N_9966,N_9604);
nor UO_313 (O_313,N_9633,N_9867);
nand UO_314 (O_314,N_9529,N_9694);
nor UO_315 (O_315,N_9913,N_9770);
nor UO_316 (O_316,N_9543,N_9794);
nor UO_317 (O_317,N_9928,N_9778);
and UO_318 (O_318,N_9593,N_9676);
or UO_319 (O_319,N_9968,N_9970);
or UO_320 (O_320,N_9765,N_9680);
or UO_321 (O_321,N_9768,N_9781);
and UO_322 (O_322,N_9878,N_9877);
or UO_323 (O_323,N_9764,N_9524);
and UO_324 (O_324,N_9616,N_9881);
nor UO_325 (O_325,N_9620,N_9917);
nor UO_326 (O_326,N_9974,N_9567);
nand UO_327 (O_327,N_9621,N_9924);
and UO_328 (O_328,N_9580,N_9579);
nor UO_329 (O_329,N_9938,N_9746);
nand UO_330 (O_330,N_9606,N_9793);
or UO_331 (O_331,N_9714,N_9828);
and UO_332 (O_332,N_9732,N_9753);
and UO_333 (O_333,N_9773,N_9756);
nor UO_334 (O_334,N_9739,N_9503);
or UO_335 (O_335,N_9865,N_9647);
nand UO_336 (O_336,N_9834,N_9813);
nand UO_337 (O_337,N_9658,N_9893);
nand UO_338 (O_338,N_9994,N_9589);
nor UO_339 (O_339,N_9858,N_9944);
nor UO_340 (O_340,N_9689,N_9961);
or UO_341 (O_341,N_9861,N_9940);
or UO_342 (O_342,N_9803,N_9709);
nand UO_343 (O_343,N_9587,N_9749);
or UO_344 (O_344,N_9863,N_9512);
nand UO_345 (O_345,N_9701,N_9814);
nand UO_346 (O_346,N_9527,N_9665);
nand UO_347 (O_347,N_9886,N_9506);
and UO_348 (O_348,N_9615,N_9821);
nand UO_349 (O_349,N_9642,N_9787);
or UO_350 (O_350,N_9937,N_9501);
and UO_351 (O_351,N_9759,N_9989);
and UO_352 (O_352,N_9972,N_9512);
nor UO_353 (O_353,N_9546,N_9512);
nand UO_354 (O_354,N_9599,N_9846);
nor UO_355 (O_355,N_9928,N_9531);
nor UO_356 (O_356,N_9961,N_9645);
or UO_357 (O_357,N_9773,N_9959);
and UO_358 (O_358,N_9721,N_9956);
nand UO_359 (O_359,N_9748,N_9548);
nand UO_360 (O_360,N_9803,N_9507);
nor UO_361 (O_361,N_9953,N_9781);
or UO_362 (O_362,N_9984,N_9573);
or UO_363 (O_363,N_9849,N_9699);
nand UO_364 (O_364,N_9677,N_9627);
or UO_365 (O_365,N_9508,N_9578);
and UO_366 (O_366,N_9738,N_9530);
nand UO_367 (O_367,N_9875,N_9683);
xnor UO_368 (O_368,N_9602,N_9831);
nand UO_369 (O_369,N_9578,N_9844);
nand UO_370 (O_370,N_9556,N_9730);
or UO_371 (O_371,N_9658,N_9739);
or UO_372 (O_372,N_9871,N_9722);
and UO_373 (O_373,N_9990,N_9526);
nor UO_374 (O_374,N_9759,N_9524);
nor UO_375 (O_375,N_9719,N_9825);
or UO_376 (O_376,N_9863,N_9838);
and UO_377 (O_377,N_9687,N_9536);
and UO_378 (O_378,N_9760,N_9692);
or UO_379 (O_379,N_9927,N_9665);
or UO_380 (O_380,N_9651,N_9626);
nand UO_381 (O_381,N_9711,N_9982);
and UO_382 (O_382,N_9766,N_9922);
nand UO_383 (O_383,N_9561,N_9959);
or UO_384 (O_384,N_9697,N_9567);
or UO_385 (O_385,N_9976,N_9780);
nand UO_386 (O_386,N_9699,N_9635);
nor UO_387 (O_387,N_9962,N_9704);
and UO_388 (O_388,N_9984,N_9698);
and UO_389 (O_389,N_9650,N_9600);
nand UO_390 (O_390,N_9544,N_9598);
nor UO_391 (O_391,N_9813,N_9870);
nor UO_392 (O_392,N_9798,N_9755);
and UO_393 (O_393,N_9500,N_9790);
nand UO_394 (O_394,N_9544,N_9851);
nand UO_395 (O_395,N_9853,N_9923);
and UO_396 (O_396,N_9672,N_9559);
or UO_397 (O_397,N_9867,N_9515);
or UO_398 (O_398,N_9842,N_9589);
or UO_399 (O_399,N_9734,N_9940);
or UO_400 (O_400,N_9621,N_9540);
nor UO_401 (O_401,N_9858,N_9773);
nor UO_402 (O_402,N_9884,N_9988);
nand UO_403 (O_403,N_9958,N_9508);
and UO_404 (O_404,N_9784,N_9537);
or UO_405 (O_405,N_9929,N_9683);
nor UO_406 (O_406,N_9715,N_9830);
or UO_407 (O_407,N_9890,N_9860);
and UO_408 (O_408,N_9591,N_9799);
or UO_409 (O_409,N_9906,N_9752);
and UO_410 (O_410,N_9545,N_9724);
nand UO_411 (O_411,N_9907,N_9540);
or UO_412 (O_412,N_9862,N_9560);
nor UO_413 (O_413,N_9892,N_9602);
and UO_414 (O_414,N_9868,N_9903);
nor UO_415 (O_415,N_9548,N_9571);
or UO_416 (O_416,N_9506,N_9697);
or UO_417 (O_417,N_9790,N_9891);
and UO_418 (O_418,N_9819,N_9593);
or UO_419 (O_419,N_9532,N_9922);
or UO_420 (O_420,N_9867,N_9964);
and UO_421 (O_421,N_9765,N_9578);
nor UO_422 (O_422,N_9826,N_9613);
nor UO_423 (O_423,N_9685,N_9862);
and UO_424 (O_424,N_9597,N_9907);
or UO_425 (O_425,N_9711,N_9720);
nand UO_426 (O_426,N_9994,N_9747);
nor UO_427 (O_427,N_9526,N_9811);
and UO_428 (O_428,N_9909,N_9976);
or UO_429 (O_429,N_9858,N_9831);
and UO_430 (O_430,N_9939,N_9695);
or UO_431 (O_431,N_9542,N_9505);
nand UO_432 (O_432,N_9641,N_9648);
nor UO_433 (O_433,N_9824,N_9865);
nand UO_434 (O_434,N_9693,N_9555);
nand UO_435 (O_435,N_9965,N_9873);
and UO_436 (O_436,N_9514,N_9986);
and UO_437 (O_437,N_9648,N_9580);
nand UO_438 (O_438,N_9700,N_9727);
nor UO_439 (O_439,N_9639,N_9899);
nor UO_440 (O_440,N_9860,N_9540);
nand UO_441 (O_441,N_9862,N_9666);
or UO_442 (O_442,N_9718,N_9991);
and UO_443 (O_443,N_9907,N_9687);
or UO_444 (O_444,N_9743,N_9560);
or UO_445 (O_445,N_9722,N_9860);
and UO_446 (O_446,N_9669,N_9771);
or UO_447 (O_447,N_9736,N_9744);
and UO_448 (O_448,N_9666,N_9865);
and UO_449 (O_449,N_9765,N_9513);
xor UO_450 (O_450,N_9893,N_9621);
nor UO_451 (O_451,N_9927,N_9794);
nand UO_452 (O_452,N_9640,N_9766);
and UO_453 (O_453,N_9962,N_9527);
nor UO_454 (O_454,N_9593,N_9552);
and UO_455 (O_455,N_9549,N_9599);
nor UO_456 (O_456,N_9527,N_9750);
or UO_457 (O_457,N_9712,N_9503);
xor UO_458 (O_458,N_9684,N_9720);
nand UO_459 (O_459,N_9890,N_9597);
nor UO_460 (O_460,N_9860,N_9531);
nor UO_461 (O_461,N_9919,N_9974);
nor UO_462 (O_462,N_9839,N_9611);
and UO_463 (O_463,N_9903,N_9562);
or UO_464 (O_464,N_9874,N_9593);
and UO_465 (O_465,N_9852,N_9557);
nand UO_466 (O_466,N_9735,N_9960);
nor UO_467 (O_467,N_9850,N_9753);
nor UO_468 (O_468,N_9502,N_9546);
nor UO_469 (O_469,N_9903,N_9700);
nand UO_470 (O_470,N_9989,N_9622);
nand UO_471 (O_471,N_9856,N_9719);
and UO_472 (O_472,N_9925,N_9777);
or UO_473 (O_473,N_9923,N_9942);
nor UO_474 (O_474,N_9934,N_9677);
and UO_475 (O_475,N_9678,N_9518);
and UO_476 (O_476,N_9800,N_9944);
and UO_477 (O_477,N_9605,N_9604);
or UO_478 (O_478,N_9921,N_9733);
nand UO_479 (O_479,N_9692,N_9969);
and UO_480 (O_480,N_9641,N_9616);
and UO_481 (O_481,N_9695,N_9749);
nor UO_482 (O_482,N_9776,N_9840);
or UO_483 (O_483,N_9860,N_9974);
or UO_484 (O_484,N_9840,N_9766);
and UO_485 (O_485,N_9616,N_9859);
nor UO_486 (O_486,N_9663,N_9895);
or UO_487 (O_487,N_9995,N_9749);
nand UO_488 (O_488,N_9658,N_9689);
and UO_489 (O_489,N_9730,N_9775);
nor UO_490 (O_490,N_9923,N_9724);
nor UO_491 (O_491,N_9722,N_9817);
nor UO_492 (O_492,N_9805,N_9874);
xor UO_493 (O_493,N_9709,N_9617);
or UO_494 (O_494,N_9522,N_9588);
or UO_495 (O_495,N_9543,N_9648);
or UO_496 (O_496,N_9750,N_9606);
nor UO_497 (O_497,N_9592,N_9613);
and UO_498 (O_498,N_9582,N_9965);
or UO_499 (O_499,N_9742,N_9773);
and UO_500 (O_500,N_9504,N_9735);
and UO_501 (O_501,N_9511,N_9688);
nor UO_502 (O_502,N_9944,N_9617);
nand UO_503 (O_503,N_9625,N_9712);
nand UO_504 (O_504,N_9763,N_9780);
nand UO_505 (O_505,N_9928,N_9884);
nor UO_506 (O_506,N_9752,N_9772);
nand UO_507 (O_507,N_9782,N_9881);
nand UO_508 (O_508,N_9693,N_9819);
nor UO_509 (O_509,N_9965,N_9927);
or UO_510 (O_510,N_9583,N_9903);
or UO_511 (O_511,N_9936,N_9546);
nand UO_512 (O_512,N_9636,N_9852);
nor UO_513 (O_513,N_9737,N_9680);
or UO_514 (O_514,N_9953,N_9964);
nand UO_515 (O_515,N_9784,N_9993);
nand UO_516 (O_516,N_9699,N_9554);
nor UO_517 (O_517,N_9679,N_9890);
or UO_518 (O_518,N_9633,N_9628);
nor UO_519 (O_519,N_9699,N_9888);
nand UO_520 (O_520,N_9765,N_9754);
or UO_521 (O_521,N_9691,N_9598);
nor UO_522 (O_522,N_9562,N_9759);
or UO_523 (O_523,N_9687,N_9662);
nor UO_524 (O_524,N_9704,N_9621);
nor UO_525 (O_525,N_9798,N_9963);
nor UO_526 (O_526,N_9764,N_9934);
xnor UO_527 (O_527,N_9712,N_9793);
nand UO_528 (O_528,N_9622,N_9526);
and UO_529 (O_529,N_9878,N_9608);
and UO_530 (O_530,N_9777,N_9640);
or UO_531 (O_531,N_9716,N_9966);
nor UO_532 (O_532,N_9662,N_9671);
and UO_533 (O_533,N_9601,N_9520);
and UO_534 (O_534,N_9785,N_9887);
or UO_535 (O_535,N_9728,N_9965);
and UO_536 (O_536,N_9757,N_9914);
nand UO_537 (O_537,N_9670,N_9913);
nor UO_538 (O_538,N_9561,N_9549);
xor UO_539 (O_539,N_9735,N_9879);
nand UO_540 (O_540,N_9950,N_9512);
or UO_541 (O_541,N_9868,N_9652);
and UO_542 (O_542,N_9619,N_9813);
and UO_543 (O_543,N_9604,N_9686);
or UO_544 (O_544,N_9677,N_9525);
and UO_545 (O_545,N_9914,N_9569);
nand UO_546 (O_546,N_9900,N_9682);
and UO_547 (O_547,N_9953,N_9883);
nand UO_548 (O_548,N_9770,N_9725);
nand UO_549 (O_549,N_9681,N_9730);
nor UO_550 (O_550,N_9796,N_9633);
nor UO_551 (O_551,N_9618,N_9555);
nor UO_552 (O_552,N_9934,N_9769);
nand UO_553 (O_553,N_9813,N_9700);
nand UO_554 (O_554,N_9955,N_9919);
and UO_555 (O_555,N_9997,N_9563);
nand UO_556 (O_556,N_9858,N_9998);
or UO_557 (O_557,N_9976,N_9900);
and UO_558 (O_558,N_9531,N_9712);
nand UO_559 (O_559,N_9766,N_9777);
or UO_560 (O_560,N_9716,N_9767);
and UO_561 (O_561,N_9707,N_9727);
and UO_562 (O_562,N_9662,N_9803);
or UO_563 (O_563,N_9592,N_9817);
nand UO_564 (O_564,N_9722,N_9729);
nand UO_565 (O_565,N_9579,N_9797);
nand UO_566 (O_566,N_9661,N_9833);
nand UO_567 (O_567,N_9988,N_9873);
or UO_568 (O_568,N_9804,N_9547);
or UO_569 (O_569,N_9977,N_9923);
nand UO_570 (O_570,N_9554,N_9735);
and UO_571 (O_571,N_9831,N_9874);
or UO_572 (O_572,N_9509,N_9946);
and UO_573 (O_573,N_9542,N_9556);
or UO_574 (O_574,N_9889,N_9861);
or UO_575 (O_575,N_9986,N_9614);
nand UO_576 (O_576,N_9504,N_9637);
nor UO_577 (O_577,N_9784,N_9586);
or UO_578 (O_578,N_9929,N_9904);
nand UO_579 (O_579,N_9718,N_9955);
or UO_580 (O_580,N_9710,N_9536);
nand UO_581 (O_581,N_9501,N_9759);
and UO_582 (O_582,N_9980,N_9775);
nand UO_583 (O_583,N_9975,N_9551);
and UO_584 (O_584,N_9537,N_9895);
nor UO_585 (O_585,N_9799,N_9677);
or UO_586 (O_586,N_9527,N_9889);
nor UO_587 (O_587,N_9685,N_9872);
nand UO_588 (O_588,N_9857,N_9822);
or UO_589 (O_589,N_9519,N_9905);
and UO_590 (O_590,N_9563,N_9641);
nor UO_591 (O_591,N_9684,N_9859);
nand UO_592 (O_592,N_9690,N_9719);
nor UO_593 (O_593,N_9956,N_9713);
or UO_594 (O_594,N_9687,N_9771);
or UO_595 (O_595,N_9659,N_9649);
or UO_596 (O_596,N_9845,N_9815);
and UO_597 (O_597,N_9731,N_9957);
or UO_598 (O_598,N_9558,N_9928);
nand UO_599 (O_599,N_9790,N_9761);
nand UO_600 (O_600,N_9536,N_9523);
nor UO_601 (O_601,N_9838,N_9822);
or UO_602 (O_602,N_9883,N_9823);
or UO_603 (O_603,N_9680,N_9690);
and UO_604 (O_604,N_9897,N_9823);
and UO_605 (O_605,N_9811,N_9968);
or UO_606 (O_606,N_9903,N_9961);
nand UO_607 (O_607,N_9569,N_9624);
and UO_608 (O_608,N_9592,N_9771);
nor UO_609 (O_609,N_9820,N_9627);
nor UO_610 (O_610,N_9633,N_9619);
and UO_611 (O_611,N_9646,N_9857);
nand UO_612 (O_612,N_9928,N_9803);
or UO_613 (O_613,N_9681,N_9708);
and UO_614 (O_614,N_9722,N_9574);
nor UO_615 (O_615,N_9920,N_9573);
nand UO_616 (O_616,N_9827,N_9865);
nor UO_617 (O_617,N_9777,N_9619);
or UO_618 (O_618,N_9662,N_9983);
and UO_619 (O_619,N_9621,N_9902);
nor UO_620 (O_620,N_9806,N_9637);
nor UO_621 (O_621,N_9614,N_9585);
and UO_622 (O_622,N_9780,N_9769);
nand UO_623 (O_623,N_9598,N_9650);
nor UO_624 (O_624,N_9991,N_9992);
or UO_625 (O_625,N_9835,N_9987);
and UO_626 (O_626,N_9681,N_9787);
and UO_627 (O_627,N_9974,N_9546);
or UO_628 (O_628,N_9666,N_9793);
nand UO_629 (O_629,N_9691,N_9710);
nor UO_630 (O_630,N_9611,N_9924);
nor UO_631 (O_631,N_9668,N_9945);
xor UO_632 (O_632,N_9573,N_9595);
nand UO_633 (O_633,N_9793,N_9836);
nand UO_634 (O_634,N_9645,N_9716);
nand UO_635 (O_635,N_9744,N_9696);
or UO_636 (O_636,N_9733,N_9612);
nand UO_637 (O_637,N_9638,N_9880);
nand UO_638 (O_638,N_9611,N_9984);
nand UO_639 (O_639,N_9808,N_9633);
and UO_640 (O_640,N_9695,N_9969);
nor UO_641 (O_641,N_9936,N_9800);
or UO_642 (O_642,N_9513,N_9930);
nand UO_643 (O_643,N_9834,N_9771);
nor UO_644 (O_644,N_9665,N_9770);
or UO_645 (O_645,N_9658,N_9513);
nor UO_646 (O_646,N_9750,N_9685);
nor UO_647 (O_647,N_9998,N_9756);
and UO_648 (O_648,N_9756,N_9626);
and UO_649 (O_649,N_9869,N_9856);
nand UO_650 (O_650,N_9599,N_9613);
or UO_651 (O_651,N_9613,N_9997);
nand UO_652 (O_652,N_9967,N_9796);
or UO_653 (O_653,N_9755,N_9535);
nor UO_654 (O_654,N_9620,N_9577);
nor UO_655 (O_655,N_9571,N_9568);
and UO_656 (O_656,N_9664,N_9904);
and UO_657 (O_657,N_9882,N_9840);
and UO_658 (O_658,N_9710,N_9500);
nor UO_659 (O_659,N_9758,N_9928);
nor UO_660 (O_660,N_9627,N_9751);
or UO_661 (O_661,N_9956,N_9664);
or UO_662 (O_662,N_9601,N_9792);
nor UO_663 (O_663,N_9848,N_9672);
or UO_664 (O_664,N_9890,N_9720);
or UO_665 (O_665,N_9947,N_9802);
xnor UO_666 (O_666,N_9681,N_9788);
nand UO_667 (O_667,N_9515,N_9703);
and UO_668 (O_668,N_9809,N_9932);
nor UO_669 (O_669,N_9534,N_9703);
and UO_670 (O_670,N_9562,N_9661);
nand UO_671 (O_671,N_9532,N_9838);
nor UO_672 (O_672,N_9595,N_9940);
or UO_673 (O_673,N_9651,N_9826);
nand UO_674 (O_674,N_9725,N_9523);
and UO_675 (O_675,N_9970,N_9927);
and UO_676 (O_676,N_9972,N_9856);
nand UO_677 (O_677,N_9713,N_9640);
or UO_678 (O_678,N_9937,N_9880);
or UO_679 (O_679,N_9582,N_9763);
xor UO_680 (O_680,N_9655,N_9516);
nor UO_681 (O_681,N_9648,N_9862);
and UO_682 (O_682,N_9951,N_9955);
nand UO_683 (O_683,N_9731,N_9628);
nor UO_684 (O_684,N_9579,N_9551);
nor UO_685 (O_685,N_9670,N_9754);
nand UO_686 (O_686,N_9635,N_9721);
and UO_687 (O_687,N_9805,N_9560);
and UO_688 (O_688,N_9783,N_9872);
nand UO_689 (O_689,N_9589,N_9752);
and UO_690 (O_690,N_9801,N_9914);
nor UO_691 (O_691,N_9660,N_9510);
xor UO_692 (O_692,N_9867,N_9775);
and UO_693 (O_693,N_9829,N_9565);
nand UO_694 (O_694,N_9985,N_9954);
or UO_695 (O_695,N_9995,N_9729);
nor UO_696 (O_696,N_9828,N_9813);
and UO_697 (O_697,N_9680,N_9591);
or UO_698 (O_698,N_9900,N_9841);
or UO_699 (O_699,N_9860,N_9728);
nor UO_700 (O_700,N_9974,N_9696);
nand UO_701 (O_701,N_9748,N_9988);
nand UO_702 (O_702,N_9801,N_9948);
or UO_703 (O_703,N_9619,N_9524);
or UO_704 (O_704,N_9558,N_9930);
and UO_705 (O_705,N_9972,N_9984);
nor UO_706 (O_706,N_9593,N_9529);
and UO_707 (O_707,N_9771,N_9957);
and UO_708 (O_708,N_9584,N_9848);
or UO_709 (O_709,N_9534,N_9748);
or UO_710 (O_710,N_9580,N_9784);
and UO_711 (O_711,N_9748,N_9590);
nor UO_712 (O_712,N_9736,N_9740);
nand UO_713 (O_713,N_9672,N_9760);
nor UO_714 (O_714,N_9702,N_9726);
nand UO_715 (O_715,N_9846,N_9685);
nor UO_716 (O_716,N_9846,N_9903);
and UO_717 (O_717,N_9861,N_9886);
nor UO_718 (O_718,N_9641,N_9527);
or UO_719 (O_719,N_9666,N_9904);
nand UO_720 (O_720,N_9587,N_9551);
or UO_721 (O_721,N_9859,N_9505);
or UO_722 (O_722,N_9519,N_9699);
nand UO_723 (O_723,N_9913,N_9691);
or UO_724 (O_724,N_9920,N_9995);
or UO_725 (O_725,N_9655,N_9824);
nor UO_726 (O_726,N_9756,N_9876);
and UO_727 (O_727,N_9669,N_9968);
nand UO_728 (O_728,N_9538,N_9501);
and UO_729 (O_729,N_9581,N_9946);
and UO_730 (O_730,N_9920,N_9698);
or UO_731 (O_731,N_9801,N_9970);
nor UO_732 (O_732,N_9810,N_9843);
or UO_733 (O_733,N_9613,N_9967);
nor UO_734 (O_734,N_9741,N_9676);
and UO_735 (O_735,N_9606,N_9907);
nand UO_736 (O_736,N_9701,N_9645);
nor UO_737 (O_737,N_9833,N_9746);
and UO_738 (O_738,N_9789,N_9854);
and UO_739 (O_739,N_9904,N_9769);
and UO_740 (O_740,N_9500,N_9580);
or UO_741 (O_741,N_9969,N_9802);
nand UO_742 (O_742,N_9977,N_9994);
nor UO_743 (O_743,N_9868,N_9864);
or UO_744 (O_744,N_9912,N_9875);
nand UO_745 (O_745,N_9981,N_9765);
nand UO_746 (O_746,N_9735,N_9707);
and UO_747 (O_747,N_9759,N_9814);
nand UO_748 (O_748,N_9880,N_9671);
nand UO_749 (O_749,N_9809,N_9825);
nor UO_750 (O_750,N_9776,N_9581);
nor UO_751 (O_751,N_9965,N_9848);
nand UO_752 (O_752,N_9763,N_9945);
nor UO_753 (O_753,N_9657,N_9831);
and UO_754 (O_754,N_9560,N_9679);
xnor UO_755 (O_755,N_9529,N_9558);
xnor UO_756 (O_756,N_9780,N_9692);
or UO_757 (O_757,N_9901,N_9903);
or UO_758 (O_758,N_9901,N_9675);
nor UO_759 (O_759,N_9847,N_9896);
or UO_760 (O_760,N_9601,N_9669);
and UO_761 (O_761,N_9550,N_9675);
and UO_762 (O_762,N_9905,N_9756);
or UO_763 (O_763,N_9620,N_9884);
nand UO_764 (O_764,N_9846,N_9635);
or UO_765 (O_765,N_9695,N_9937);
nand UO_766 (O_766,N_9557,N_9977);
and UO_767 (O_767,N_9805,N_9754);
nand UO_768 (O_768,N_9764,N_9929);
nand UO_769 (O_769,N_9735,N_9824);
or UO_770 (O_770,N_9588,N_9799);
and UO_771 (O_771,N_9829,N_9869);
nor UO_772 (O_772,N_9918,N_9710);
and UO_773 (O_773,N_9841,N_9997);
nand UO_774 (O_774,N_9684,N_9606);
and UO_775 (O_775,N_9562,N_9900);
nor UO_776 (O_776,N_9908,N_9988);
nor UO_777 (O_777,N_9547,N_9793);
or UO_778 (O_778,N_9774,N_9563);
nor UO_779 (O_779,N_9907,N_9500);
and UO_780 (O_780,N_9627,N_9661);
nor UO_781 (O_781,N_9679,N_9914);
and UO_782 (O_782,N_9565,N_9833);
and UO_783 (O_783,N_9735,N_9691);
nor UO_784 (O_784,N_9582,N_9526);
or UO_785 (O_785,N_9792,N_9512);
or UO_786 (O_786,N_9806,N_9742);
nor UO_787 (O_787,N_9840,N_9870);
or UO_788 (O_788,N_9612,N_9616);
nand UO_789 (O_789,N_9622,N_9784);
nand UO_790 (O_790,N_9790,N_9911);
and UO_791 (O_791,N_9864,N_9674);
nand UO_792 (O_792,N_9546,N_9524);
and UO_793 (O_793,N_9700,N_9742);
nor UO_794 (O_794,N_9805,N_9574);
and UO_795 (O_795,N_9583,N_9685);
nor UO_796 (O_796,N_9778,N_9542);
or UO_797 (O_797,N_9796,N_9957);
and UO_798 (O_798,N_9907,N_9533);
and UO_799 (O_799,N_9636,N_9548);
and UO_800 (O_800,N_9728,N_9848);
nor UO_801 (O_801,N_9535,N_9664);
or UO_802 (O_802,N_9810,N_9873);
nor UO_803 (O_803,N_9673,N_9946);
nand UO_804 (O_804,N_9658,N_9660);
xor UO_805 (O_805,N_9524,N_9964);
nand UO_806 (O_806,N_9722,N_9677);
nand UO_807 (O_807,N_9542,N_9536);
or UO_808 (O_808,N_9887,N_9664);
nand UO_809 (O_809,N_9798,N_9612);
nand UO_810 (O_810,N_9542,N_9848);
and UO_811 (O_811,N_9536,N_9795);
or UO_812 (O_812,N_9978,N_9889);
nand UO_813 (O_813,N_9983,N_9539);
or UO_814 (O_814,N_9630,N_9621);
and UO_815 (O_815,N_9814,N_9593);
and UO_816 (O_816,N_9949,N_9919);
nor UO_817 (O_817,N_9708,N_9639);
nand UO_818 (O_818,N_9807,N_9785);
or UO_819 (O_819,N_9663,N_9931);
or UO_820 (O_820,N_9500,N_9612);
or UO_821 (O_821,N_9612,N_9547);
and UO_822 (O_822,N_9607,N_9735);
and UO_823 (O_823,N_9811,N_9689);
xor UO_824 (O_824,N_9689,N_9942);
nor UO_825 (O_825,N_9621,N_9510);
nand UO_826 (O_826,N_9795,N_9979);
and UO_827 (O_827,N_9567,N_9965);
or UO_828 (O_828,N_9859,N_9664);
nor UO_829 (O_829,N_9638,N_9800);
nand UO_830 (O_830,N_9583,N_9757);
nand UO_831 (O_831,N_9683,N_9624);
nand UO_832 (O_832,N_9552,N_9697);
nor UO_833 (O_833,N_9659,N_9534);
or UO_834 (O_834,N_9956,N_9847);
or UO_835 (O_835,N_9684,N_9934);
or UO_836 (O_836,N_9898,N_9951);
nand UO_837 (O_837,N_9669,N_9880);
nand UO_838 (O_838,N_9804,N_9933);
nor UO_839 (O_839,N_9713,N_9546);
and UO_840 (O_840,N_9514,N_9816);
or UO_841 (O_841,N_9509,N_9706);
or UO_842 (O_842,N_9590,N_9977);
or UO_843 (O_843,N_9688,N_9972);
or UO_844 (O_844,N_9721,N_9825);
nand UO_845 (O_845,N_9794,N_9761);
nand UO_846 (O_846,N_9822,N_9508);
and UO_847 (O_847,N_9740,N_9634);
nor UO_848 (O_848,N_9560,N_9526);
and UO_849 (O_849,N_9923,N_9633);
nand UO_850 (O_850,N_9749,N_9698);
xor UO_851 (O_851,N_9668,N_9629);
and UO_852 (O_852,N_9699,N_9943);
nor UO_853 (O_853,N_9570,N_9555);
and UO_854 (O_854,N_9819,N_9515);
nand UO_855 (O_855,N_9827,N_9872);
nor UO_856 (O_856,N_9940,N_9879);
and UO_857 (O_857,N_9782,N_9988);
nand UO_858 (O_858,N_9775,N_9580);
and UO_859 (O_859,N_9520,N_9711);
or UO_860 (O_860,N_9761,N_9557);
nor UO_861 (O_861,N_9985,N_9689);
or UO_862 (O_862,N_9743,N_9586);
or UO_863 (O_863,N_9954,N_9721);
and UO_864 (O_864,N_9601,N_9572);
or UO_865 (O_865,N_9969,N_9705);
and UO_866 (O_866,N_9738,N_9584);
nand UO_867 (O_867,N_9906,N_9934);
nand UO_868 (O_868,N_9527,N_9984);
nor UO_869 (O_869,N_9975,N_9583);
nand UO_870 (O_870,N_9783,N_9981);
and UO_871 (O_871,N_9693,N_9922);
nand UO_872 (O_872,N_9560,N_9736);
nor UO_873 (O_873,N_9757,N_9633);
nor UO_874 (O_874,N_9833,N_9883);
nor UO_875 (O_875,N_9979,N_9571);
or UO_876 (O_876,N_9949,N_9817);
and UO_877 (O_877,N_9995,N_9615);
or UO_878 (O_878,N_9961,N_9657);
or UO_879 (O_879,N_9695,N_9921);
nor UO_880 (O_880,N_9966,N_9979);
nor UO_881 (O_881,N_9789,N_9927);
or UO_882 (O_882,N_9976,N_9842);
and UO_883 (O_883,N_9997,N_9621);
and UO_884 (O_884,N_9951,N_9754);
or UO_885 (O_885,N_9618,N_9556);
or UO_886 (O_886,N_9539,N_9658);
or UO_887 (O_887,N_9895,N_9575);
nor UO_888 (O_888,N_9774,N_9933);
or UO_889 (O_889,N_9693,N_9548);
nand UO_890 (O_890,N_9565,N_9610);
or UO_891 (O_891,N_9858,N_9520);
and UO_892 (O_892,N_9639,N_9551);
nand UO_893 (O_893,N_9916,N_9677);
or UO_894 (O_894,N_9794,N_9584);
or UO_895 (O_895,N_9880,N_9737);
and UO_896 (O_896,N_9640,N_9581);
or UO_897 (O_897,N_9601,N_9736);
nor UO_898 (O_898,N_9552,N_9545);
nor UO_899 (O_899,N_9620,N_9889);
nor UO_900 (O_900,N_9537,N_9767);
or UO_901 (O_901,N_9544,N_9705);
nor UO_902 (O_902,N_9812,N_9780);
nor UO_903 (O_903,N_9919,N_9805);
nor UO_904 (O_904,N_9840,N_9769);
nor UO_905 (O_905,N_9908,N_9893);
nor UO_906 (O_906,N_9976,N_9748);
and UO_907 (O_907,N_9619,N_9530);
xor UO_908 (O_908,N_9596,N_9523);
or UO_909 (O_909,N_9660,N_9548);
or UO_910 (O_910,N_9872,N_9581);
nor UO_911 (O_911,N_9975,N_9834);
and UO_912 (O_912,N_9786,N_9857);
nand UO_913 (O_913,N_9956,N_9857);
and UO_914 (O_914,N_9692,N_9658);
xor UO_915 (O_915,N_9598,N_9524);
xnor UO_916 (O_916,N_9550,N_9747);
and UO_917 (O_917,N_9806,N_9980);
and UO_918 (O_918,N_9847,N_9778);
or UO_919 (O_919,N_9853,N_9911);
or UO_920 (O_920,N_9820,N_9981);
nor UO_921 (O_921,N_9980,N_9511);
or UO_922 (O_922,N_9639,N_9567);
or UO_923 (O_923,N_9949,N_9965);
nand UO_924 (O_924,N_9985,N_9996);
nor UO_925 (O_925,N_9519,N_9631);
nand UO_926 (O_926,N_9532,N_9935);
or UO_927 (O_927,N_9934,N_9631);
or UO_928 (O_928,N_9986,N_9973);
nand UO_929 (O_929,N_9568,N_9648);
or UO_930 (O_930,N_9620,N_9934);
and UO_931 (O_931,N_9706,N_9745);
nand UO_932 (O_932,N_9632,N_9704);
and UO_933 (O_933,N_9856,N_9589);
nand UO_934 (O_934,N_9883,N_9999);
and UO_935 (O_935,N_9793,N_9846);
or UO_936 (O_936,N_9804,N_9669);
nor UO_937 (O_937,N_9803,N_9533);
and UO_938 (O_938,N_9502,N_9515);
or UO_939 (O_939,N_9535,N_9929);
nand UO_940 (O_940,N_9584,N_9879);
or UO_941 (O_941,N_9729,N_9552);
and UO_942 (O_942,N_9775,N_9600);
nand UO_943 (O_943,N_9646,N_9764);
and UO_944 (O_944,N_9729,N_9806);
and UO_945 (O_945,N_9729,N_9743);
nor UO_946 (O_946,N_9898,N_9551);
and UO_947 (O_947,N_9642,N_9519);
and UO_948 (O_948,N_9643,N_9605);
xnor UO_949 (O_949,N_9864,N_9966);
and UO_950 (O_950,N_9890,N_9589);
or UO_951 (O_951,N_9536,N_9562);
and UO_952 (O_952,N_9669,N_9529);
nand UO_953 (O_953,N_9705,N_9862);
or UO_954 (O_954,N_9536,N_9857);
nand UO_955 (O_955,N_9503,N_9793);
or UO_956 (O_956,N_9585,N_9571);
or UO_957 (O_957,N_9522,N_9643);
nand UO_958 (O_958,N_9850,N_9687);
and UO_959 (O_959,N_9759,N_9564);
nand UO_960 (O_960,N_9917,N_9577);
nor UO_961 (O_961,N_9609,N_9686);
nor UO_962 (O_962,N_9660,N_9981);
or UO_963 (O_963,N_9767,N_9769);
nor UO_964 (O_964,N_9945,N_9790);
or UO_965 (O_965,N_9593,N_9794);
nand UO_966 (O_966,N_9693,N_9763);
nor UO_967 (O_967,N_9808,N_9626);
nand UO_968 (O_968,N_9520,N_9844);
nand UO_969 (O_969,N_9550,N_9882);
nor UO_970 (O_970,N_9751,N_9939);
and UO_971 (O_971,N_9897,N_9558);
or UO_972 (O_972,N_9639,N_9969);
nor UO_973 (O_973,N_9788,N_9602);
nor UO_974 (O_974,N_9914,N_9705);
and UO_975 (O_975,N_9644,N_9949);
nor UO_976 (O_976,N_9508,N_9804);
or UO_977 (O_977,N_9699,N_9996);
or UO_978 (O_978,N_9805,N_9808);
and UO_979 (O_979,N_9855,N_9675);
or UO_980 (O_980,N_9872,N_9754);
or UO_981 (O_981,N_9790,N_9933);
and UO_982 (O_982,N_9771,N_9694);
nor UO_983 (O_983,N_9723,N_9527);
nor UO_984 (O_984,N_9753,N_9891);
nor UO_985 (O_985,N_9556,N_9878);
nor UO_986 (O_986,N_9688,N_9755);
and UO_987 (O_987,N_9860,N_9876);
nor UO_988 (O_988,N_9995,N_9876);
or UO_989 (O_989,N_9865,N_9556);
nand UO_990 (O_990,N_9733,N_9573);
and UO_991 (O_991,N_9530,N_9798);
xor UO_992 (O_992,N_9649,N_9652);
nand UO_993 (O_993,N_9974,N_9509);
nand UO_994 (O_994,N_9563,N_9803);
or UO_995 (O_995,N_9684,N_9910);
or UO_996 (O_996,N_9664,N_9938);
and UO_997 (O_997,N_9778,N_9769);
nor UO_998 (O_998,N_9559,N_9997);
and UO_999 (O_999,N_9674,N_9603);
and UO_1000 (O_1000,N_9694,N_9729);
and UO_1001 (O_1001,N_9786,N_9774);
or UO_1002 (O_1002,N_9654,N_9546);
nand UO_1003 (O_1003,N_9945,N_9645);
and UO_1004 (O_1004,N_9635,N_9640);
and UO_1005 (O_1005,N_9634,N_9534);
or UO_1006 (O_1006,N_9569,N_9722);
or UO_1007 (O_1007,N_9724,N_9792);
or UO_1008 (O_1008,N_9835,N_9802);
nand UO_1009 (O_1009,N_9824,N_9722);
or UO_1010 (O_1010,N_9908,N_9600);
or UO_1011 (O_1011,N_9786,N_9725);
and UO_1012 (O_1012,N_9844,N_9834);
or UO_1013 (O_1013,N_9892,N_9869);
nand UO_1014 (O_1014,N_9684,N_9887);
nor UO_1015 (O_1015,N_9538,N_9571);
and UO_1016 (O_1016,N_9579,N_9721);
nor UO_1017 (O_1017,N_9709,N_9979);
nand UO_1018 (O_1018,N_9853,N_9575);
or UO_1019 (O_1019,N_9897,N_9924);
or UO_1020 (O_1020,N_9936,N_9884);
and UO_1021 (O_1021,N_9685,N_9814);
or UO_1022 (O_1022,N_9860,N_9911);
nor UO_1023 (O_1023,N_9698,N_9907);
or UO_1024 (O_1024,N_9916,N_9765);
nand UO_1025 (O_1025,N_9829,N_9966);
and UO_1026 (O_1026,N_9790,N_9639);
nand UO_1027 (O_1027,N_9533,N_9625);
nor UO_1028 (O_1028,N_9650,N_9997);
or UO_1029 (O_1029,N_9879,N_9860);
or UO_1030 (O_1030,N_9666,N_9719);
and UO_1031 (O_1031,N_9671,N_9675);
and UO_1032 (O_1032,N_9787,N_9663);
or UO_1033 (O_1033,N_9724,N_9989);
and UO_1034 (O_1034,N_9612,N_9825);
nand UO_1035 (O_1035,N_9946,N_9781);
and UO_1036 (O_1036,N_9618,N_9724);
nor UO_1037 (O_1037,N_9766,N_9792);
or UO_1038 (O_1038,N_9756,N_9755);
nor UO_1039 (O_1039,N_9832,N_9701);
nor UO_1040 (O_1040,N_9933,N_9993);
nor UO_1041 (O_1041,N_9656,N_9740);
and UO_1042 (O_1042,N_9773,N_9849);
and UO_1043 (O_1043,N_9517,N_9953);
and UO_1044 (O_1044,N_9646,N_9577);
nor UO_1045 (O_1045,N_9969,N_9835);
nor UO_1046 (O_1046,N_9990,N_9666);
or UO_1047 (O_1047,N_9812,N_9619);
nand UO_1048 (O_1048,N_9543,N_9732);
nand UO_1049 (O_1049,N_9806,N_9793);
nor UO_1050 (O_1050,N_9745,N_9785);
nor UO_1051 (O_1051,N_9758,N_9702);
or UO_1052 (O_1052,N_9910,N_9866);
and UO_1053 (O_1053,N_9719,N_9563);
nand UO_1054 (O_1054,N_9893,N_9588);
and UO_1055 (O_1055,N_9692,N_9632);
nor UO_1056 (O_1056,N_9523,N_9882);
nor UO_1057 (O_1057,N_9749,N_9740);
or UO_1058 (O_1058,N_9783,N_9871);
nor UO_1059 (O_1059,N_9943,N_9686);
nand UO_1060 (O_1060,N_9818,N_9528);
and UO_1061 (O_1061,N_9897,N_9896);
xor UO_1062 (O_1062,N_9834,N_9511);
nor UO_1063 (O_1063,N_9552,N_9851);
or UO_1064 (O_1064,N_9967,N_9739);
nand UO_1065 (O_1065,N_9699,N_9711);
xnor UO_1066 (O_1066,N_9944,N_9733);
and UO_1067 (O_1067,N_9607,N_9750);
and UO_1068 (O_1068,N_9821,N_9738);
and UO_1069 (O_1069,N_9503,N_9681);
and UO_1070 (O_1070,N_9805,N_9896);
nor UO_1071 (O_1071,N_9641,N_9969);
nor UO_1072 (O_1072,N_9997,N_9729);
and UO_1073 (O_1073,N_9829,N_9880);
nor UO_1074 (O_1074,N_9645,N_9610);
nand UO_1075 (O_1075,N_9884,N_9757);
and UO_1076 (O_1076,N_9891,N_9811);
and UO_1077 (O_1077,N_9704,N_9799);
xnor UO_1078 (O_1078,N_9874,N_9921);
or UO_1079 (O_1079,N_9735,N_9500);
xor UO_1080 (O_1080,N_9962,N_9641);
nor UO_1081 (O_1081,N_9963,N_9697);
nand UO_1082 (O_1082,N_9555,N_9660);
or UO_1083 (O_1083,N_9645,N_9831);
nand UO_1084 (O_1084,N_9971,N_9944);
or UO_1085 (O_1085,N_9939,N_9571);
or UO_1086 (O_1086,N_9586,N_9654);
and UO_1087 (O_1087,N_9503,N_9654);
or UO_1088 (O_1088,N_9590,N_9816);
and UO_1089 (O_1089,N_9690,N_9593);
nor UO_1090 (O_1090,N_9597,N_9581);
and UO_1091 (O_1091,N_9950,N_9558);
or UO_1092 (O_1092,N_9630,N_9917);
nor UO_1093 (O_1093,N_9715,N_9683);
nor UO_1094 (O_1094,N_9557,N_9505);
xor UO_1095 (O_1095,N_9887,N_9663);
nand UO_1096 (O_1096,N_9741,N_9938);
nor UO_1097 (O_1097,N_9962,N_9843);
nor UO_1098 (O_1098,N_9671,N_9913);
nand UO_1099 (O_1099,N_9599,N_9593);
nor UO_1100 (O_1100,N_9558,N_9602);
nor UO_1101 (O_1101,N_9946,N_9678);
and UO_1102 (O_1102,N_9980,N_9630);
and UO_1103 (O_1103,N_9639,N_9640);
or UO_1104 (O_1104,N_9902,N_9857);
nor UO_1105 (O_1105,N_9680,N_9965);
or UO_1106 (O_1106,N_9708,N_9888);
or UO_1107 (O_1107,N_9869,N_9538);
nand UO_1108 (O_1108,N_9537,N_9558);
nor UO_1109 (O_1109,N_9709,N_9887);
nand UO_1110 (O_1110,N_9806,N_9671);
nand UO_1111 (O_1111,N_9653,N_9574);
or UO_1112 (O_1112,N_9910,N_9819);
or UO_1113 (O_1113,N_9519,N_9674);
or UO_1114 (O_1114,N_9953,N_9685);
or UO_1115 (O_1115,N_9611,N_9512);
or UO_1116 (O_1116,N_9577,N_9945);
nand UO_1117 (O_1117,N_9854,N_9968);
nand UO_1118 (O_1118,N_9618,N_9767);
nor UO_1119 (O_1119,N_9810,N_9571);
and UO_1120 (O_1120,N_9572,N_9755);
nor UO_1121 (O_1121,N_9788,N_9643);
nand UO_1122 (O_1122,N_9956,N_9856);
and UO_1123 (O_1123,N_9802,N_9917);
and UO_1124 (O_1124,N_9557,N_9609);
nor UO_1125 (O_1125,N_9944,N_9705);
nand UO_1126 (O_1126,N_9828,N_9593);
and UO_1127 (O_1127,N_9666,N_9721);
nor UO_1128 (O_1128,N_9729,N_9619);
or UO_1129 (O_1129,N_9859,N_9658);
and UO_1130 (O_1130,N_9792,N_9698);
nand UO_1131 (O_1131,N_9836,N_9551);
nor UO_1132 (O_1132,N_9873,N_9606);
and UO_1133 (O_1133,N_9839,N_9624);
nor UO_1134 (O_1134,N_9647,N_9616);
nand UO_1135 (O_1135,N_9845,N_9542);
and UO_1136 (O_1136,N_9879,N_9648);
xnor UO_1137 (O_1137,N_9674,N_9855);
nand UO_1138 (O_1138,N_9547,N_9748);
nand UO_1139 (O_1139,N_9811,N_9714);
or UO_1140 (O_1140,N_9860,N_9611);
nor UO_1141 (O_1141,N_9770,N_9802);
or UO_1142 (O_1142,N_9818,N_9811);
or UO_1143 (O_1143,N_9933,N_9641);
and UO_1144 (O_1144,N_9911,N_9579);
or UO_1145 (O_1145,N_9707,N_9952);
nor UO_1146 (O_1146,N_9647,N_9518);
nand UO_1147 (O_1147,N_9826,N_9780);
or UO_1148 (O_1148,N_9885,N_9880);
and UO_1149 (O_1149,N_9932,N_9502);
nand UO_1150 (O_1150,N_9568,N_9973);
xor UO_1151 (O_1151,N_9998,N_9700);
nand UO_1152 (O_1152,N_9500,N_9635);
or UO_1153 (O_1153,N_9791,N_9617);
or UO_1154 (O_1154,N_9780,N_9875);
nand UO_1155 (O_1155,N_9575,N_9838);
or UO_1156 (O_1156,N_9554,N_9773);
or UO_1157 (O_1157,N_9679,N_9800);
and UO_1158 (O_1158,N_9752,N_9549);
or UO_1159 (O_1159,N_9990,N_9846);
nor UO_1160 (O_1160,N_9810,N_9591);
nand UO_1161 (O_1161,N_9858,N_9830);
nand UO_1162 (O_1162,N_9619,N_9900);
or UO_1163 (O_1163,N_9627,N_9588);
nor UO_1164 (O_1164,N_9655,N_9741);
or UO_1165 (O_1165,N_9958,N_9683);
nor UO_1166 (O_1166,N_9537,N_9967);
nand UO_1167 (O_1167,N_9809,N_9570);
nand UO_1168 (O_1168,N_9999,N_9726);
and UO_1169 (O_1169,N_9855,N_9827);
and UO_1170 (O_1170,N_9830,N_9932);
or UO_1171 (O_1171,N_9564,N_9638);
nand UO_1172 (O_1172,N_9515,N_9977);
and UO_1173 (O_1173,N_9684,N_9916);
or UO_1174 (O_1174,N_9522,N_9802);
nor UO_1175 (O_1175,N_9718,N_9665);
and UO_1176 (O_1176,N_9817,N_9518);
nand UO_1177 (O_1177,N_9571,N_9866);
or UO_1178 (O_1178,N_9884,N_9542);
or UO_1179 (O_1179,N_9925,N_9652);
or UO_1180 (O_1180,N_9785,N_9667);
or UO_1181 (O_1181,N_9554,N_9838);
nor UO_1182 (O_1182,N_9727,N_9618);
or UO_1183 (O_1183,N_9579,N_9616);
or UO_1184 (O_1184,N_9997,N_9875);
nand UO_1185 (O_1185,N_9612,N_9520);
nor UO_1186 (O_1186,N_9586,N_9613);
or UO_1187 (O_1187,N_9735,N_9765);
nor UO_1188 (O_1188,N_9620,N_9865);
xnor UO_1189 (O_1189,N_9731,N_9913);
and UO_1190 (O_1190,N_9728,N_9913);
or UO_1191 (O_1191,N_9520,N_9528);
and UO_1192 (O_1192,N_9637,N_9716);
and UO_1193 (O_1193,N_9811,N_9681);
nand UO_1194 (O_1194,N_9593,N_9700);
or UO_1195 (O_1195,N_9883,N_9509);
and UO_1196 (O_1196,N_9791,N_9635);
and UO_1197 (O_1197,N_9766,N_9538);
or UO_1198 (O_1198,N_9744,N_9503);
nor UO_1199 (O_1199,N_9913,N_9937);
nand UO_1200 (O_1200,N_9873,N_9555);
and UO_1201 (O_1201,N_9935,N_9578);
or UO_1202 (O_1202,N_9590,N_9743);
and UO_1203 (O_1203,N_9724,N_9566);
nand UO_1204 (O_1204,N_9869,N_9697);
nor UO_1205 (O_1205,N_9543,N_9663);
nand UO_1206 (O_1206,N_9526,N_9530);
nand UO_1207 (O_1207,N_9919,N_9695);
nand UO_1208 (O_1208,N_9783,N_9773);
and UO_1209 (O_1209,N_9792,N_9890);
or UO_1210 (O_1210,N_9862,N_9925);
nand UO_1211 (O_1211,N_9625,N_9860);
nor UO_1212 (O_1212,N_9884,N_9554);
or UO_1213 (O_1213,N_9535,N_9778);
or UO_1214 (O_1214,N_9557,N_9553);
and UO_1215 (O_1215,N_9744,N_9685);
or UO_1216 (O_1216,N_9963,N_9584);
nor UO_1217 (O_1217,N_9521,N_9737);
nand UO_1218 (O_1218,N_9954,N_9654);
and UO_1219 (O_1219,N_9787,N_9505);
or UO_1220 (O_1220,N_9655,N_9990);
and UO_1221 (O_1221,N_9806,N_9975);
or UO_1222 (O_1222,N_9501,N_9942);
nor UO_1223 (O_1223,N_9814,N_9879);
nand UO_1224 (O_1224,N_9952,N_9887);
nand UO_1225 (O_1225,N_9998,N_9995);
nand UO_1226 (O_1226,N_9965,N_9674);
and UO_1227 (O_1227,N_9881,N_9702);
nand UO_1228 (O_1228,N_9753,N_9979);
and UO_1229 (O_1229,N_9700,N_9750);
or UO_1230 (O_1230,N_9645,N_9783);
or UO_1231 (O_1231,N_9917,N_9739);
nand UO_1232 (O_1232,N_9927,N_9670);
or UO_1233 (O_1233,N_9883,N_9655);
nand UO_1234 (O_1234,N_9844,N_9949);
nor UO_1235 (O_1235,N_9820,N_9833);
or UO_1236 (O_1236,N_9916,N_9667);
or UO_1237 (O_1237,N_9580,N_9588);
nand UO_1238 (O_1238,N_9622,N_9983);
nand UO_1239 (O_1239,N_9734,N_9609);
or UO_1240 (O_1240,N_9740,N_9888);
nand UO_1241 (O_1241,N_9658,N_9524);
nand UO_1242 (O_1242,N_9968,N_9870);
nor UO_1243 (O_1243,N_9736,N_9860);
and UO_1244 (O_1244,N_9900,N_9794);
and UO_1245 (O_1245,N_9823,N_9596);
nand UO_1246 (O_1246,N_9879,N_9755);
and UO_1247 (O_1247,N_9716,N_9995);
or UO_1248 (O_1248,N_9975,N_9831);
nor UO_1249 (O_1249,N_9896,N_9568);
or UO_1250 (O_1250,N_9511,N_9997);
and UO_1251 (O_1251,N_9937,N_9956);
nor UO_1252 (O_1252,N_9764,N_9657);
and UO_1253 (O_1253,N_9683,N_9788);
and UO_1254 (O_1254,N_9831,N_9903);
and UO_1255 (O_1255,N_9904,N_9606);
or UO_1256 (O_1256,N_9856,N_9865);
or UO_1257 (O_1257,N_9945,N_9849);
and UO_1258 (O_1258,N_9570,N_9554);
or UO_1259 (O_1259,N_9971,N_9668);
and UO_1260 (O_1260,N_9998,N_9915);
or UO_1261 (O_1261,N_9630,N_9826);
and UO_1262 (O_1262,N_9901,N_9917);
or UO_1263 (O_1263,N_9697,N_9723);
or UO_1264 (O_1264,N_9541,N_9503);
or UO_1265 (O_1265,N_9527,N_9987);
or UO_1266 (O_1266,N_9961,N_9964);
nand UO_1267 (O_1267,N_9904,N_9677);
and UO_1268 (O_1268,N_9619,N_9527);
nand UO_1269 (O_1269,N_9663,N_9772);
nand UO_1270 (O_1270,N_9938,N_9511);
nand UO_1271 (O_1271,N_9837,N_9909);
nor UO_1272 (O_1272,N_9945,N_9705);
or UO_1273 (O_1273,N_9749,N_9646);
or UO_1274 (O_1274,N_9836,N_9669);
and UO_1275 (O_1275,N_9752,N_9982);
or UO_1276 (O_1276,N_9597,N_9896);
nor UO_1277 (O_1277,N_9831,N_9613);
or UO_1278 (O_1278,N_9792,N_9558);
nand UO_1279 (O_1279,N_9649,N_9678);
nor UO_1280 (O_1280,N_9840,N_9856);
nand UO_1281 (O_1281,N_9891,N_9823);
nand UO_1282 (O_1282,N_9866,N_9911);
nor UO_1283 (O_1283,N_9604,N_9509);
and UO_1284 (O_1284,N_9763,N_9720);
or UO_1285 (O_1285,N_9965,N_9604);
or UO_1286 (O_1286,N_9840,N_9722);
and UO_1287 (O_1287,N_9694,N_9816);
or UO_1288 (O_1288,N_9893,N_9697);
nand UO_1289 (O_1289,N_9538,N_9693);
nor UO_1290 (O_1290,N_9630,N_9539);
or UO_1291 (O_1291,N_9619,N_9714);
nor UO_1292 (O_1292,N_9896,N_9666);
nor UO_1293 (O_1293,N_9640,N_9871);
and UO_1294 (O_1294,N_9626,N_9664);
nor UO_1295 (O_1295,N_9527,N_9556);
and UO_1296 (O_1296,N_9813,N_9622);
and UO_1297 (O_1297,N_9534,N_9972);
nor UO_1298 (O_1298,N_9886,N_9853);
nor UO_1299 (O_1299,N_9660,N_9932);
nand UO_1300 (O_1300,N_9842,N_9830);
nor UO_1301 (O_1301,N_9828,N_9844);
and UO_1302 (O_1302,N_9524,N_9573);
or UO_1303 (O_1303,N_9659,N_9752);
nand UO_1304 (O_1304,N_9631,N_9562);
nand UO_1305 (O_1305,N_9547,N_9891);
xor UO_1306 (O_1306,N_9948,N_9974);
or UO_1307 (O_1307,N_9576,N_9932);
and UO_1308 (O_1308,N_9736,N_9850);
nand UO_1309 (O_1309,N_9517,N_9578);
nand UO_1310 (O_1310,N_9532,N_9669);
nor UO_1311 (O_1311,N_9783,N_9588);
nand UO_1312 (O_1312,N_9697,N_9819);
nand UO_1313 (O_1313,N_9746,N_9512);
and UO_1314 (O_1314,N_9757,N_9540);
nand UO_1315 (O_1315,N_9541,N_9509);
nand UO_1316 (O_1316,N_9546,N_9714);
or UO_1317 (O_1317,N_9986,N_9542);
or UO_1318 (O_1318,N_9900,N_9685);
nand UO_1319 (O_1319,N_9986,N_9956);
and UO_1320 (O_1320,N_9541,N_9683);
or UO_1321 (O_1321,N_9718,N_9881);
or UO_1322 (O_1322,N_9891,N_9539);
or UO_1323 (O_1323,N_9853,N_9506);
or UO_1324 (O_1324,N_9654,N_9590);
nor UO_1325 (O_1325,N_9772,N_9678);
nor UO_1326 (O_1326,N_9785,N_9767);
xor UO_1327 (O_1327,N_9873,N_9821);
nor UO_1328 (O_1328,N_9740,N_9872);
nor UO_1329 (O_1329,N_9706,N_9885);
nor UO_1330 (O_1330,N_9690,N_9914);
nand UO_1331 (O_1331,N_9803,N_9564);
nor UO_1332 (O_1332,N_9600,N_9836);
nand UO_1333 (O_1333,N_9580,N_9905);
or UO_1334 (O_1334,N_9958,N_9760);
and UO_1335 (O_1335,N_9981,N_9719);
and UO_1336 (O_1336,N_9963,N_9631);
nand UO_1337 (O_1337,N_9680,N_9570);
or UO_1338 (O_1338,N_9922,N_9946);
and UO_1339 (O_1339,N_9731,N_9510);
nor UO_1340 (O_1340,N_9795,N_9682);
nor UO_1341 (O_1341,N_9587,N_9528);
and UO_1342 (O_1342,N_9804,N_9934);
and UO_1343 (O_1343,N_9575,N_9654);
or UO_1344 (O_1344,N_9634,N_9695);
or UO_1345 (O_1345,N_9946,N_9658);
nand UO_1346 (O_1346,N_9884,N_9982);
nand UO_1347 (O_1347,N_9804,N_9862);
xor UO_1348 (O_1348,N_9806,N_9994);
nand UO_1349 (O_1349,N_9591,N_9549);
nor UO_1350 (O_1350,N_9899,N_9708);
nand UO_1351 (O_1351,N_9658,N_9883);
nand UO_1352 (O_1352,N_9864,N_9848);
nor UO_1353 (O_1353,N_9978,N_9726);
nand UO_1354 (O_1354,N_9679,N_9848);
and UO_1355 (O_1355,N_9539,N_9596);
or UO_1356 (O_1356,N_9593,N_9865);
nor UO_1357 (O_1357,N_9543,N_9902);
and UO_1358 (O_1358,N_9531,N_9697);
and UO_1359 (O_1359,N_9757,N_9509);
nand UO_1360 (O_1360,N_9697,N_9591);
nor UO_1361 (O_1361,N_9531,N_9505);
and UO_1362 (O_1362,N_9683,N_9724);
nor UO_1363 (O_1363,N_9952,N_9725);
or UO_1364 (O_1364,N_9813,N_9807);
nor UO_1365 (O_1365,N_9503,N_9906);
nor UO_1366 (O_1366,N_9883,N_9829);
nand UO_1367 (O_1367,N_9593,N_9675);
nand UO_1368 (O_1368,N_9506,N_9765);
or UO_1369 (O_1369,N_9786,N_9911);
nor UO_1370 (O_1370,N_9521,N_9508);
xor UO_1371 (O_1371,N_9785,N_9770);
and UO_1372 (O_1372,N_9670,N_9893);
nand UO_1373 (O_1373,N_9793,N_9838);
or UO_1374 (O_1374,N_9606,N_9519);
nor UO_1375 (O_1375,N_9612,N_9942);
or UO_1376 (O_1376,N_9639,N_9599);
or UO_1377 (O_1377,N_9937,N_9722);
nor UO_1378 (O_1378,N_9833,N_9986);
nand UO_1379 (O_1379,N_9765,N_9531);
or UO_1380 (O_1380,N_9703,N_9733);
or UO_1381 (O_1381,N_9976,N_9667);
nand UO_1382 (O_1382,N_9901,N_9502);
nor UO_1383 (O_1383,N_9555,N_9980);
and UO_1384 (O_1384,N_9707,N_9558);
nor UO_1385 (O_1385,N_9966,N_9744);
or UO_1386 (O_1386,N_9852,N_9515);
or UO_1387 (O_1387,N_9720,N_9973);
and UO_1388 (O_1388,N_9757,N_9862);
nand UO_1389 (O_1389,N_9957,N_9735);
and UO_1390 (O_1390,N_9623,N_9889);
and UO_1391 (O_1391,N_9854,N_9928);
nand UO_1392 (O_1392,N_9582,N_9665);
or UO_1393 (O_1393,N_9972,N_9659);
or UO_1394 (O_1394,N_9552,N_9711);
nor UO_1395 (O_1395,N_9777,N_9914);
and UO_1396 (O_1396,N_9673,N_9885);
or UO_1397 (O_1397,N_9522,N_9612);
nor UO_1398 (O_1398,N_9754,N_9585);
or UO_1399 (O_1399,N_9878,N_9889);
nor UO_1400 (O_1400,N_9601,N_9794);
or UO_1401 (O_1401,N_9839,N_9880);
or UO_1402 (O_1402,N_9920,N_9608);
xnor UO_1403 (O_1403,N_9852,N_9881);
xor UO_1404 (O_1404,N_9929,N_9789);
and UO_1405 (O_1405,N_9657,N_9587);
or UO_1406 (O_1406,N_9813,N_9910);
and UO_1407 (O_1407,N_9735,N_9668);
and UO_1408 (O_1408,N_9771,N_9686);
and UO_1409 (O_1409,N_9579,N_9929);
nor UO_1410 (O_1410,N_9703,N_9664);
nor UO_1411 (O_1411,N_9944,N_9734);
and UO_1412 (O_1412,N_9867,N_9720);
nor UO_1413 (O_1413,N_9834,N_9793);
or UO_1414 (O_1414,N_9814,N_9721);
and UO_1415 (O_1415,N_9818,N_9796);
nand UO_1416 (O_1416,N_9623,N_9958);
nor UO_1417 (O_1417,N_9515,N_9954);
nand UO_1418 (O_1418,N_9518,N_9630);
or UO_1419 (O_1419,N_9824,N_9703);
nand UO_1420 (O_1420,N_9607,N_9564);
nor UO_1421 (O_1421,N_9943,N_9950);
nor UO_1422 (O_1422,N_9994,N_9759);
nor UO_1423 (O_1423,N_9870,N_9861);
and UO_1424 (O_1424,N_9888,N_9722);
nor UO_1425 (O_1425,N_9730,N_9784);
nand UO_1426 (O_1426,N_9961,N_9815);
nor UO_1427 (O_1427,N_9848,N_9912);
nor UO_1428 (O_1428,N_9605,N_9573);
or UO_1429 (O_1429,N_9578,N_9957);
or UO_1430 (O_1430,N_9906,N_9867);
nand UO_1431 (O_1431,N_9756,N_9802);
or UO_1432 (O_1432,N_9872,N_9996);
or UO_1433 (O_1433,N_9555,N_9581);
nand UO_1434 (O_1434,N_9626,N_9569);
nor UO_1435 (O_1435,N_9900,N_9709);
and UO_1436 (O_1436,N_9932,N_9839);
nor UO_1437 (O_1437,N_9957,N_9868);
nand UO_1438 (O_1438,N_9577,N_9619);
or UO_1439 (O_1439,N_9670,N_9634);
and UO_1440 (O_1440,N_9677,N_9578);
or UO_1441 (O_1441,N_9711,N_9929);
nand UO_1442 (O_1442,N_9957,N_9844);
or UO_1443 (O_1443,N_9737,N_9643);
nand UO_1444 (O_1444,N_9753,N_9962);
nor UO_1445 (O_1445,N_9927,N_9909);
nand UO_1446 (O_1446,N_9900,N_9754);
or UO_1447 (O_1447,N_9827,N_9745);
nand UO_1448 (O_1448,N_9559,N_9765);
nor UO_1449 (O_1449,N_9674,N_9575);
or UO_1450 (O_1450,N_9798,N_9928);
nor UO_1451 (O_1451,N_9971,N_9989);
nand UO_1452 (O_1452,N_9914,N_9603);
and UO_1453 (O_1453,N_9575,N_9525);
or UO_1454 (O_1454,N_9844,N_9696);
nand UO_1455 (O_1455,N_9977,N_9538);
or UO_1456 (O_1456,N_9719,N_9919);
and UO_1457 (O_1457,N_9800,N_9717);
nor UO_1458 (O_1458,N_9940,N_9976);
nand UO_1459 (O_1459,N_9777,N_9683);
nor UO_1460 (O_1460,N_9657,N_9980);
or UO_1461 (O_1461,N_9903,N_9540);
nor UO_1462 (O_1462,N_9726,N_9738);
and UO_1463 (O_1463,N_9887,N_9603);
and UO_1464 (O_1464,N_9662,N_9635);
and UO_1465 (O_1465,N_9934,N_9500);
nand UO_1466 (O_1466,N_9753,N_9726);
xnor UO_1467 (O_1467,N_9568,N_9781);
and UO_1468 (O_1468,N_9549,N_9706);
nor UO_1469 (O_1469,N_9517,N_9778);
or UO_1470 (O_1470,N_9825,N_9733);
nand UO_1471 (O_1471,N_9884,N_9771);
nand UO_1472 (O_1472,N_9742,N_9994);
nand UO_1473 (O_1473,N_9570,N_9857);
or UO_1474 (O_1474,N_9992,N_9826);
or UO_1475 (O_1475,N_9565,N_9530);
xnor UO_1476 (O_1476,N_9701,N_9872);
and UO_1477 (O_1477,N_9620,N_9919);
nand UO_1478 (O_1478,N_9754,N_9569);
nand UO_1479 (O_1479,N_9916,N_9547);
and UO_1480 (O_1480,N_9566,N_9559);
and UO_1481 (O_1481,N_9814,N_9925);
nand UO_1482 (O_1482,N_9915,N_9676);
or UO_1483 (O_1483,N_9569,N_9967);
nor UO_1484 (O_1484,N_9917,N_9730);
or UO_1485 (O_1485,N_9768,N_9950);
and UO_1486 (O_1486,N_9698,N_9534);
and UO_1487 (O_1487,N_9763,N_9888);
xor UO_1488 (O_1488,N_9535,N_9508);
nand UO_1489 (O_1489,N_9746,N_9901);
nor UO_1490 (O_1490,N_9852,N_9811);
and UO_1491 (O_1491,N_9986,N_9926);
nor UO_1492 (O_1492,N_9520,N_9635);
and UO_1493 (O_1493,N_9671,N_9845);
nand UO_1494 (O_1494,N_9516,N_9834);
nor UO_1495 (O_1495,N_9952,N_9609);
nor UO_1496 (O_1496,N_9748,N_9666);
xor UO_1497 (O_1497,N_9902,N_9735);
or UO_1498 (O_1498,N_9630,N_9709);
nand UO_1499 (O_1499,N_9868,N_9545);
endmodule