module basic_1000_10000_1500_50_levels_5xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nor U0 (N_0,In_923,In_95);
or U1 (N_1,In_722,In_932);
nor U2 (N_2,In_793,In_543);
and U3 (N_3,In_720,In_541);
or U4 (N_4,In_324,In_569);
nor U5 (N_5,In_387,In_808);
xor U6 (N_6,In_8,In_386);
or U7 (N_7,In_179,In_482);
nor U8 (N_8,In_819,In_440);
and U9 (N_9,In_816,In_726);
nand U10 (N_10,In_606,In_438);
nor U11 (N_11,In_257,In_899);
nor U12 (N_12,In_293,In_553);
and U13 (N_13,In_564,In_517);
nand U14 (N_14,In_334,In_585);
or U15 (N_15,In_662,In_476);
nor U16 (N_16,In_786,In_971);
nand U17 (N_17,In_601,In_945);
xnor U18 (N_18,In_972,In_465);
nand U19 (N_19,In_629,In_667);
nand U20 (N_20,In_504,In_76);
xnor U21 (N_21,In_750,In_577);
or U22 (N_22,In_418,In_598);
nand U23 (N_23,In_396,In_420);
or U24 (N_24,In_907,In_593);
nor U25 (N_25,In_211,In_811);
nor U26 (N_26,In_616,In_44);
xnor U27 (N_27,In_153,In_207);
nor U28 (N_28,In_785,In_29);
nor U29 (N_29,In_7,In_350);
nor U30 (N_30,In_335,In_608);
nor U31 (N_31,In_617,In_214);
nor U32 (N_32,In_492,In_360);
nand U33 (N_33,In_777,In_770);
xnor U34 (N_34,In_643,In_554);
or U35 (N_35,In_957,In_312);
nand U36 (N_36,In_232,In_71);
nand U37 (N_37,In_748,In_807);
xor U38 (N_38,In_118,In_384);
or U39 (N_39,In_426,In_580);
nor U40 (N_40,In_547,In_149);
and U41 (N_41,In_823,In_186);
nor U42 (N_42,In_924,In_208);
or U43 (N_43,In_271,In_314);
nand U44 (N_44,In_172,In_925);
nand U45 (N_45,In_801,In_780);
nand U46 (N_46,In_927,In_781);
nor U47 (N_47,In_944,In_341);
nand U48 (N_48,In_472,In_666);
nand U49 (N_49,In_549,In_294);
or U50 (N_50,In_367,In_528);
xor U51 (N_51,In_249,In_728);
nor U52 (N_52,In_209,In_70);
or U53 (N_53,In_872,In_173);
nor U54 (N_54,In_653,In_347);
xor U55 (N_55,In_370,In_300);
and U56 (N_56,In_865,In_441);
or U57 (N_57,In_965,In_787);
and U58 (N_58,In_556,In_757);
nand U59 (N_59,In_52,In_741);
and U60 (N_60,In_458,In_536);
nand U61 (N_61,In_731,In_302);
xnor U62 (N_62,In_255,In_805);
nor U63 (N_63,In_560,In_698);
and U64 (N_64,In_520,In_127);
and U65 (N_65,In_216,In_835);
or U66 (N_66,In_248,In_115);
or U67 (N_67,In_909,In_631);
nand U68 (N_68,In_219,In_266);
and U69 (N_69,In_953,In_187);
nor U70 (N_70,In_125,In_298);
nand U71 (N_71,In_6,In_829);
or U72 (N_72,In_380,In_2);
nor U73 (N_73,In_678,In_57);
nor U74 (N_74,In_490,In_876);
nor U75 (N_75,In_142,In_524);
nand U76 (N_76,In_624,In_45);
xnor U77 (N_77,In_550,In_128);
xnor U78 (N_78,In_150,In_896);
nand U79 (N_79,In_412,In_670);
or U80 (N_80,In_607,In_814);
nand U81 (N_81,In_579,In_680);
nor U82 (N_82,In_462,In_604);
or U83 (N_83,In_61,In_26);
xor U84 (N_84,In_527,In_970);
and U85 (N_85,In_234,In_69);
and U86 (N_86,In_264,In_254);
nor U87 (N_87,In_514,In_727);
nor U88 (N_88,In_279,In_739);
or U89 (N_89,In_854,In_361);
nor U90 (N_90,In_831,In_41);
xor U91 (N_91,In_339,In_573);
and U92 (N_92,In_493,In_712);
or U93 (N_93,In_791,In_615);
and U94 (N_94,In_422,In_359);
or U95 (N_95,In_80,In_376);
and U96 (N_96,In_445,In_88);
or U97 (N_97,In_843,In_288);
and U98 (N_98,In_416,In_745);
or U99 (N_99,In_406,In_423);
and U100 (N_100,In_46,In_539);
or U101 (N_101,In_735,In_926);
or U102 (N_102,In_84,In_405);
or U103 (N_103,In_960,In_181);
or U104 (N_104,In_623,In_852);
nor U105 (N_105,In_375,In_922);
nand U106 (N_106,In_867,In_883);
xnor U107 (N_107,In_931,In_632);
and U108 (N_108,In_72,In_437);
nor U109 (N_109,In_329,In_851);
xnor U110 (N_110,In_190,In_451);
nand U111 (N_111,In_578,In_729);
xor U112 (N_112,In_900,In_352);
or U113 (N_113,In_73,In_240);
nor U114 (N_114,In_428,In_993);
xor U115 (N_115,In_51,In_351);
nor U116 (N_116,In_431,In_817);
xor U117 (N_117,In_589,In_319);
or U118 (N_118,In_552,In_677);
and U119 (N_119,In_169,In_4);
nor U120 (N_120,In_820,In_599);
xnor U121 (N_121,In_145,In_914);
nand U122 (N_122,In_12,In_143);
xnor U123 (N_123,In_200,In_855);
nand U124 (N_124,In_982,In_175);
nor U125 (N_125,In_252,In_622);
or U126 (N_126,In_471,In_345);
or U127 (N_127,In_964,In_268);
or U128 (N_128,In_975,In_101);
and U129 (N_129,In_663,In_419);
or U130 (N_130,In_290,In_691);
and U131 (N_131,In_586,In_424);
or U132 (N_132,In_20,In_133);
nor U133 (N_133,In_320,In_301);
nor U134 (N_134,In_508,In_934);
and U135 (N_135,In_998,In_296);
or U136 (N_136,In_938,In_174);
xor U137 (N_137,In_860,In_815);
nor U138 (N_138,In_291,In_762);
or U139 (N_139,In_809,In_463);
nand U140 (N_140,In_58,In_763);
and U141 (N_141,In_223,In_795);
and U142 (N_142,In_671,In_346);
or U143 (N_143,In_503,In_409);
nand U144 (N_144,In_790,In_806);
nand U145 (N_145,In_701,In_272);
and U146 (N_146,In_747,In_902);
and U147 (N_147,In_168,In_994);
nor U148 (N_148,In_789,In_263);
and U149 (N_149,In_507,In_713);
or U150 (N_150,In_141,In_603);
nand U151 (N_151,In_930,In_723);
nor U152 (N_152,In_937,In_292);
nand U153 (N_153,In_442,In_3);
and U154 (N_154,In_81,In_129);
nand U155 (N_155,In_697,In_68);
and U156 (N_156,In_102,In_571);
or U157 (N_157,In_810,In_170);
nor U158 (N_158,In_25,In_222);
and U159 (N_159,In_134,In_344);
and U160 (N_160,In_397,In_297);
or U161 (N_161,In_160,In_191);
nor U162 (N_162,In_479,In_875);
and U163 (N_163,In_199,In_878);
nor U164 (N_164,In_995,In_233);
nor U165 (N_165,In_605,In_918);
or U166 (N_166,In_919,In_980);
nand U167 (N_167,In_36,In_706);
xor U168 (N_168,In_498,In_837);
nor U169 (N_169,In_398,In_193);
nor U170 (N_170,In_391,In_824);
and U171 (N_171,In_383,In_353);
and U172 (N_172,In_453,In_655);
nor U173 (N_173,In_163,In_885);
xor U174 (N_174,In_338,In_449);
nor U175 (N_175,In_116,In_866);
nand U176 (N_176,In_262,In_530);
or U177 (N_177,In_66,In_983);
and U178 (N_178,In_682,In_826);
nor U179 (N_179,In_83,In_22);
or U180 (N_180,In_113,In_847);
nor U181 (N_181,In_640,In_773);
nor U182 (N_182,In_912,In_794);
or U183 (N_183,In_516,In_651);
nor U184 (N_184,In_105,In_182);
or U185 (N_185,In_488,In_48);
or U186 (N_186,In_390,In_323);
nor U187 (N_187,In_486,In_892);
nand U188 (N_188,In_707,In_844);
nand U189 (N_189,In_752,In_18);
nand U190 (N_190,In_326,In_743);
or U191 (N_191,In_628,In_716);
nor U192 (N_192,In_736,In_531);
and U193 (N_193,In_669,In_974);
nor U194 (N_194,In_411,In_124);
and U195 (N_195,In_771,In_196);
nand U196 (N_196,In_470,In_792);
nor U197 (N_197,In_685,In_568);
nor U198 (N_198,In_404,In_385);
and U199 (N_199,In_991,In_331);
nand U200 (N_200,In_260,N_0);
and U201 (N_201,In_967,In_859);
or U202 (N_202,In_333,N_114);
or U203 (N_203,In_270,In_475);
and U204 (N_204,In_704,In_849);
nor U205 (N_205,In_126,N_185);
or U206 (N_206,In_523,N_52);
nand U207 (N_207,N_58,In_802);
and U208 (N_208,In_389,In_921);
or U209 (N_209,In_821,In_446);
xor U210 (N_210,N_41,In_473);
and U211 (N_211,In_342,In_718);
nor U212 (N_212,In_863,In_277);
nand U213 (N_213,In_35,In_611);
nand U214 (N_214,In_308,In_581);
nor U215 (N_215,N_192,N_59);
nor U216 (N_216,In_646,In_929);
nor U217 (N_217,In_559,In_702);
nand U218 (N_218,In_621,In_348);
and U219 (N_219,In_987,N_117);
nor U220 (N_220,N_92,In_904);
or U221 (N_221,In_337,In_658);
nand U222 (N_222,In_590,N_179);
nand U223 (N_223,In_372,N_169);
nand U224 (N_224,In_861,N_61);
nand U225 (N_225,In_891,In_638);
and U226 (N_226,In_395,In_284);
nor U227 (N_227,In_138,N_109);
and U228 (N_228,N_172,In_761);
xor U229 (N_229,N_77,In_235);
nand U230 (N_230,In_695,In_19);
and U231 (N_231,In_410,In_903);
nand U232 (N_232,In_85,N_123);
nor U233 (N_233,In_267,N_14);
nor U234 (N_234,In_874,In_619);
xor U235 (N_235,In_484,In_584);
or U236 (N_236,In_176,In_120);
nand U237 (N_237,In_185,In_103);
nand U238 (N_238,In_215,N_76);
or U239 (N_239,N_103,N_176);
nor U240 (N_240,In_307,In_782);
and U241 (N_241,In_227,In_167);
nor U242 (N_242,In_220,In_474);
nand U243 (N_243,In_562,N_140);
or U244 (N_244,In_951,N_136);
nand U245 (N_245,In_49,In_299);
and U246 (N_246,In_454,In_64);
nand U247 (N_247,In_933,In_151);
nor U248 (N_248,In_947,In_496);
and U249 (N_249,In_368,In_690);
and U250 (N_250,In_123,In_97);
nand U251 (N_251,In_668,In_740);
nor U252 (N_252,In_700,In_0);
xor U253 (N_253,In_286,In_778);
nor U254 (N_254,In_911,In_526);
nor U255 (N_255,N_170,N_127);
nor U256 (N_256,In_660,N_190);
nor U257 (N_257,In_112,In_724);
nand U258 (N_258,In_461,N_183);
xnor U259 (N_259,In_156,N_95);
nand U260 (N_260,N_152,In_717);
nand U261 (N_261,N_101,N_50);
nor U262 (N_262,N_175,N_142);
and U263 (N_263,In_540,In_23);
nor U264 (N_264,N_7,In_576);
or U265 (N_265,In_274,In_106);
nand U266 (N_266,In_439,In_521);
nor U267 (N_267,N_13,In_228);
nor U268 (N_268,N_33,In_834);
xor U269 (N_269,N_65,In_575);
nor U270 (N_270,In_204,In_11);
and U271 (N_271,In_665,In_131);
nor U272 (N_272,In_489,N_73);
nor U273 (N_273,N_199,In_251);
nor U274 (N_274,N_108,In_229);
and U275 (N_275,N_111,In_765);
nand U276 (N_276,In_906,In_501);
nor U277 (N_277,N_44,In_137);
or U278 (N_278,In_961,In_65);
or U279 (N_279,N_187,In_379);
nor U280 (N_280,In_37,In_194);
nand U281 (N_281,In_758,In_317);
nor U282 (N_282,In_466,In_981);
nor U283 (N_283,In_864,In_650);
nand U284 (N_284,N_97,N_189);
or U285 (N_285,In_647,N_34);
and U286 (N_286,N_198,N_6);
and U287 (N_287,In_694,N_47);
nand U288 (N_288,In_511,N_78);
nor U289 (N_289,N_146,In_881);
and U290 (N_290,N_107,In_833);
nand U291 (N_291,In_546,In_672);
nor U292 (N_292,In_9,In_448);
nor U293 (N_293,N_66,In_230);
nand U294 (N_294,In_402,In_467);
or U295 (N_295,In_818,In_977);
nor U296 (N_296,In_845,In_281);
and U297 (N_297,In_407,In_800);
or U298 (N_298,In_572,In_525);
nand U299 (N_299,In_681,In_537);
nor U300 (N_300,In_400,In_839);
xor U301 (N_301,In_948,In_639);
xnor U302 (N_302,In_566,In_378);
nand U303 (N_303,In_17,In_804);
nand U304 (N_304,N_151,In_495);
nand U305 (N_305,In_245,N_35);
nor U306 (N_306,In_478,In_869);
or U307 (N_307,In_563,In_633);
or U308 (N_308,N_121,In_171);
or U309 (N_309,In_969,In_675);
and U310 (N_310,In_146,In_783);
or U311 (N_311,In_460,In_148);
nor U312 (N_312,N_17,In_77);
nor U313 (N_313,In_853,In_278);
or U314 (N_314,In_985,In_946);
or U315 (N_315,In_813,N_102);
xor U316 (N_316,In_180,N_133);
and U317 (N_317,In_798,In_121);
nor U318 (N_318,In_958,N_163);
nor U319 (N_319,N_31,N_148);
nand U320 (N_320,In_648,N_12);
or U321 (N_321,In_797,N_113);
and U322 (N_322,In_555,In_283);
xnor U323 (N_323,N_23,N_124);
nand U324 (N_324,In_738,N_141);
xor U325 (N_325,In_287,In_188);
and U326 (N_326,In_110,In_221);
nor U327 (N_327,In_699,In_888);
and U328 (N_328,In_303,In_827);
xor U329 (N_329,In_313,In_889);
and U330 (N_330,In_157,N_67);
nor U331 (N_331,In_886,In_74);
and U332 (N_332,N_37,In_388);
nand U333 (N_333,In_714,N_168);
or U334 (N_334,N_90,In_79);
nand U335 (N_335,In_862,In_588);
xnor U336 (N_336,In_705,In_538);
and U337 (N_337,In_905,N_54);
nor U338 (N_338,In_674,In_16);
nand U339 (N_339,In_369,In_901);
or U340 (N_340,In_432,In_354);
nand U341 (N_341,N_119,In_28);
nand U342 (N_342,In_183,In_487);
or U343 (N_343,In_96,N_63);
nor U344 (N_344,In_224,In_92);
nand U345 (N_345,In_93,N_69);
or U346 (N_346,In_98,In_627);
and U347 (N_347,In_710,N_157);
nor U348 (N_348,In_491,In_54);
nand U349 (N_349,In_14,In_494);
or U350 (N_350,In_349,In_15);
and U351 (N_351,In_371,In_202);
nand U352 (N_352,In_836,N_164);
xnor U353 (N_353,In_656,In_165);
and U354 (N_354,N_24,In_362);
xnor U355 (N_355,In_213,In_596);
and U356 (N_356,In_403,N_155);
or U357 (N_357,N_167,In_893);
nand U358 (N_358,In_630,N_70);
or U359 (N_359,N_85,N_147);
xor U360 (N_360,In_989,In_444);
or U361 (N_361,In_122,N_72);
nor U362 (N_362,N_138,In_842);
and U363 (N_363,In_365,In_62);
nor U364 (N_364,In_772,In_258);
nand U365 (N_365,In_684,In_104);
nand U366 (N_366,N_60,N_48);
or U367 (N_367,In_430,In_509);
nor U368 (N_368,In_968,In_529);
xnor U369 (N_369,In_756,In_55);
nand U370 (N_370,In_898,N_182);
xnor U371 (N_371,In_594,In_356);
nand U372 (N_372,N_188,In_415);
nor U373 (N_373,In_477,In_764);
nand U374 (N_374,In_275,In_90);
or U375 (N_375,In_197,N_162);
or U376 (N_376,In_749,In_828);
nand U377 (N_377,In_256,In_47);
nor U378 (N_378,In_321,In_237);
or U379 (N_379,In_979,In_602);
and U380 (N_380,In_34,In_357);
nand U381 (N_381,In_392,N_40);
or U382 (N_382,In_94,In_942);
xnor U383 (N_383,In_950,In_734);
and U384 (N_384,In_686,In_499);
nor U385 (N_385,In_746,In_978);
and U386 (N_386,In_205,In_305);
nand U387 (N_387,In_609,In_330);
nand U388 (N_388,N_84,N_53);
and U389 (N_389,In_830,In_506);
xnor U390 (N_390,In_943,In_519);
nand U391 (N_391,N_129,N_2);
nor U392 (N_392,In_613,N_145);
xor U393 (N_393,In_954,N_82);
or U394 (N_394,In_261,N_26);
nor U395 (N_395,In_464,N_150);
nand U396 (N_396,N_154,N_193);
xnor U397 (N_397,N_75,In_162);
and U398 (N_398,In_433,In_597);
and U399 (N_399,In_799,In_687);
nor U400 (N_400,In_328,N_393);
and U401 (N_401,N_57,In_309);
and U402 (N_402,In_210,In_542);
nand U403 (N_403,In_189,N_391);
nand U404 (N_404,In_32,N_342);
and U405 (N_405,In_114,N_372);
and U406 (N_406,In_469,In_719);
or U407 (N_407,In_119,N_9);
nand U408 (N_408,N_348,In_626);
and U409 (N_409,In_742,N_128);
nor U410 (N_410,N_325,In_897);
nand U411 (N_411,In_429,In_587);
or U412 (N_412,In_139,In_644);
nor U413 (N_413,N_22,In_38);
and U414 (N_414,In_246,In_657);
nor U415 (N_415,In_166,N_280);
or U416 (N_416,N_200,N_390);
and U417 (N_417,N_287,N_16);
or U418 (N_418,N_302,N_171);
nand U419 (N_419,N_247,In_53);
or U420 (N_420,In_873,N_281);
or U421 (N_421,N_27,N_62);
nand U422 (N_422,N_210,N_290);
or U423 (N_423,N_366,N_202);
or U424 (N_424,N_49,N_364);
nor U425 (N_425,In_203,N_327);
xnor U426 (N_426,N_367,N_100);
and U427 (N_427,In_30,In_887);
or U428 (N_428,N_355,N_347);
or U429 (N_429,N_268,N_174);
nand U430 (N_430,In_636,In_269);
or U431 (N_431,In_567,In_689);
and U432 (N_432,N_293,In_238);
and U433 (N_433,N_134,N_297);
nand U434 (N_434,N_258,In_289);
and U435 (N_435,N_385,N_265);
and U436 (N_436,In_976,In_544);
and U437 (N_437,In_625,N_292);
and U438 (N_438,In_140,In_225);
nor U439 (N_439,N_311,In_417);
nor U440 (N_440,N_106,N_51);
or U441 (N_441,N_328,N_143);
or U442 (N_442,In_195,N_389);
nor U443 (N_443,N_278,N_384);
and U444 (N_444,In_614,In_239);
or U445 (N_445,N_36,N_296);
or U446 (N_446,In_620,In_936);
xnor U447 (N_447,N_243,In_868);
xor U448 (N_448,In_10,N_110);
and U449 (N_449,In_177,N_212);
xor U450 (N_450,N_392,N_1);
xnor U451 (N_451,N_369,N_120);
nand U452 (N_452,N_153,In_822);
and U453 (N_453,N_21,N_375);
and U454 (N_454,In_692,In_192);
or U455 (N_455,In_915,N_261);
or U456 (N_456,N_87,In_534);
or U457 (N_457,In_641,N_105);
nor U458 (N_458,In_642,In_340);
nand U459 (N_459,In_393,N_228);
xor U460 (N_460,In_949,N_159);
nand U461 (N_461,In_877,In_939);
and U462 (N_462,In_618,N_232);
and U463 (N_463,N_276,In_973);
and U464 (N_464,N_266,In_768);
nand U465 (N_465,In_455,N_309);
and U466 (N_466,In_435,N_178);
xor U467 (N_467,In_708,In_242);
nor U468 (N_468,N_98,N_245);
nand U469 (N_469,N_371,N_131);
and U470 (N_470,In_468,In_217);
nand U471 (N_471,N_259,In_732);
nor U472 (N_472,In_117,In_751);
and U473 (N_473,In_941,In_992);
nand U474 (N_474,N_217,In_427);
xnor U475 (N_475,N_126,N_349);
xor U476 (N_476,In_374,N_213);
nor U477 (N_477,In_664,N_286);
nand U478 (N_478,N_71,N_180);
nor U479 (N_479,N_397,N_219);
or U480 (N_480,In_709,N_201);
nor U481 (N_481,In_583,N_195);
or U482 (N_482,In_693,In_50);
or U483 (N_483,In_755,In_295);
nor U484 (N_484,In_890,N_194);
nand U485 (N_485,In_421,N_354);
nand U486 (N_486,In_952,N_104);
nor U487 (N_487,N_320,In_108);
or U488 (N_488,N_222,N_365);
and U489 (N_489,N_186,N_387);
nand U490 (N_490,N_3,In_908);
nand U491 (N_491,In_510,In_986);
or U492 (N_492,In_282,N_386);
nor U493 (N_493,In_659,N_319);
nand U494 (N_494,N_305,N_56);
or U495 (N_495,N_359,In_154);
or U496 (N_496,N_206,In_776);
and U497 (N_497,N_32,In_443);
xor U498 (N_498,In_654,In_744);
nand U499 (N_499,N_83,N_197);
or U500 (N_500,In_990,In_250);
nor U501 (N_501,In_247,In_497);
and U502 (N_502,N_283,In_60);
nand U503 (N_503,In_363,In_730);
xnor U504 (N_504,N_244,N_362);
and U505 (N_505,In_21,N_313);
nor U506 (N_506,In_43,In_725);
nand U507 (N_507,N_318,In_610);
nand U508 (N_508,In_592,N_28);
and U509 (N_509,N_272,N_322);
and U510 (N_510,N_271,N_330);
nand U511 (N_511,N_288,N_227);
and U512 (N_512,N_135,In_155);
and U513 (N_513,In_343,In_858);
or U514 (N_514,In_522,In_280);
nand U515 (N_515,N_38,In_40);
nor U516 (N_516,In_336,In_273);
nand U517 (N_517,In_645,N_373);
or U518 (N_518,N_149,In_414);
xnor U519 (N_519,In_955,In_107);
xnor U520 (N_520,N_235,In_457);
or U521 (N_521,N_214,In_152);
nand U522 (N_522,In_450,In_355);
and U523 (N_523,In_988,In_39);
and U524 (N_524,In_381,N_312);
nand U525 (N_525,In_533,In_879);
nor U526 (N_526,In_505,In_769);
nor U527 (N_527,In_784,N_350);
nand U528 (N_528,In_963,In_637);
nor U529 (N_529,In_882,N_166);
nor U530 (N_530,N_204,N_184);
nor U531 (N_531,N_380,N_29);
nand U532 (N_532,In_158,In_318);
nor U533 (N_533,In_373,N_116);
and U534 (N_534,In_456,N_360);
nand U535 (N_535,N_308,In_136);
and U536 (N_536,N_326,In_966);
nor U537 (N_537,N_256,N_399);
nand U538 (N_538,In_452,In_100);
nor U539 (N_539,In_377,N_310);
nor U540 (N_540,N_226,N_262);
nand U541 (N_541,N_161,In_327);
and U542 (N_542,N_55,N_335);
nand U543 (N_543,N_315,N_345);
and U544 (N_544,N_91,In_754);
or U545 (N_545,In_364,In_848);
or U546 (N_546,N_99,N_115);
nand U547 (N_547,N_282,In_759);
or U548 (N_548,N_254,N_216);
and U549 (N_549,N_398,In_56);
and U550 (N_550,N_18,N_253);
nand U551 (N_551,In_306,N_274);
nand U552 (N_552,N_264,In_316);
xnor U553 (N_553,In_135,N_8);
and U554 (N_554,N_291,N_181);
xnor U555 (N_555,N_267,In_676);
xor U556 (N_556,In_600,N_361);
xor U557 (N_557,N_341,In_688);
xor U558 (N_558,In_253,In_24);
nor U559 (N_559,N_370,N_81);
or U560 (N_560,N_86,N_45);
nand U561 (N_561,N_316,In_766);
nor U562 (N_562,In_673,N_139);
or U563 (N_563,N_203,In_159);
xor U564 (N_564,In_447,N_234);
or U565 (N_565,In_894,In_259);
nand U566 (N_566,In_480,N_173);
nand U567 (N_567,In_870,In_753);
or U568 (N_568,N_196,In_696);
or U569 (N_569,N_363,N_333);
and U570 (N_570,In_999,In_164);
and U571 (N_571,N_329,In_75);
or U572 (N_572,N_351,In_27);
nand U573 (N_573,In_265,In_161);
and U574 (N_574,N_112,In_42);
nand U575 (N_575,N_277,N_257);
xor U576 (N_576,In_997,In_413);
and U577 (N_577,In_825,N_158);
or U578 (N_578,In_59,N_379);
nor U579 (N_579,In_871,In_856);
nor U580 (N_580,In_767,N_4);
or U581 (N_581,In_485,In_803);
or U582 (N_582,N_383,N_220);
nor U583 (N_583,In_737,In_178);
and U584 (N_584,In_425,In_850);
or U585 (N_585,N_337,N_376);
and U586 (N_586,In_703,In_111);
and U587 (N_587,In_832,N_314);
xor U588 (N_588,In_612,In_532);
or U589 (N_589,N_299,N_279);
or U590 (N_590,In_332,In_775);
or U591 (N_591,N_249,In_78);
nor U592 (N_592,N_74,N_269);
nand U593 (N_593,In_206,In_962);
and U594 (N_594,N_246,N_30);
or U595 (N_595,In_557,In_788);
nor U596 (N_596,In_796,N_225);
or U597 (N_597,In_570,In_201);
nand U598 (N_598,N_248,In_733);
nor U599 (N_599,In_500,N_10);
nor U600 (N_600,N_535,In_401);
nand U601 (N_601,N_496,In_880);
xor U602 (N_602,N_125,N_597);
nand U603 (N_603,In_399,N_475);
xnor U604 (N_604,N_533,In_582);
nor U605 (N_605,N_39,N_593);
xor U606 (N_606,N_301,N_374);
and U607 (N_607,N_473,N_414);
or U608 (N_608,N_357,N_523);
nand U609 (N_609,In_322,In_241);
and U610 (N_610,In_13,N_88);
nand U611 (N_611,N_300,N_455);
and U612 (N_612,N_527,N_295);
nor U613 (N_613,In_231,N_550);
nor U614 (N_614,N_426,N_252);
nand U615 (N_615,N_517,N_553);
or U616 (N_616,N_324,N_510);
nor U617 (N_617,N_427,N_431);
nand U618 (N_618,In_31,N_462);
nand U619 (N_619,N_515,N_564);
nand U620 (N_620,N_94,N_516);
or U621 (N_621,N_211,N_558);
and U622 (N_622,N_569,N_207);
nor U623 (N_623,N_263,In_649);
nor U624 (N_624,N_423,N_514);
and U625 (N_625,In_857,N_549);
xnor U626 (N_626,In_548,In_198);
nor U627 (N_627,In_984,N_260);
and U628 (N_628,N_334,N_599);
and U629 (N_629,In_147,In_226);
nand U630 (N_630,N_338,In_89);
nand U631 (N_631,N_493,N_420);
and U632 (N_632,N_501,N_500);
and U633 (N_633,In_545,N_466);
nor U634 (N_634,N_237,N_89);
or U635 (N_635,N_526,N_518);
and U636 (N_636,N_424,N_415);
nand U637 (N_637,In_276,N_445);
nand U638 (N_638,N_488,N_544);
and U639 (N_639,N_487,In_63);
xor U640 (N_640,N_578,N_574);
or U641 (N_641,N_444,N_433);
nor U642 (N_642,N_394,N_490);
or U643 (N_643,N_537,N_470);
nor U644 (N_644,N_570,In_82);
nand U645 (N_645,N_540,N_575);
or U646 (N_646,N_479,In_774);
nor U647 (N_647,N_421,N_306);
nand U648 (N_648,In_518,In_551);
or U649 (N_649,In_459,N_25);
nand U650 (N_650,N_534,N_581);
xnor U651 (N_651,N_340,N_582);
nand U652 (N_652,N_580,N_284);
nor U653 (N_653,N_11,N_562);
xor U654 (N_654,N_443,N_144);
or U655 (N_655,N_457,N_242);
and U656 (N_656,N_46,N_42);
xor U657 (N_657,In_928,N_241);
xor U658 (N_658,N_539,N_556);
xnor U659 (N_659,N_441,N_560);
or U660 (N_660,N_595,N_405);
nor U661 (N_661,N_118,N_538);
and U662 (N_662,N_449,N_303);
nand U663 (N_663,N_471,N_437);
xor U664 (N_664,In_436,In_408);
nor U665 (N_665,N_402,In_87);
nor U666 (N_666,In_304,N_452);
xnor U667 (N_667,N_43,N_579);
or U668 (N_668,N_307,In_512);
xnor U669 (N_669,In_956,N_250);
nor U670 (N_670,In_502,N_439);
and U671 (N_671,N_5,In_236);
or U672 (N_672,N_592,N_587);
xor U673 (N_673,N_417,N_548);
or U674 (N_674,N_381,N_484);
nor U675 (N_675,N_451,N_339);
and U676 (N_676,N_543,In_1);
and U677 (N_677,In_935,N_572);
nand U678 (N_678,N_396,In_917);
nand U679 (N_679,N_446,N_568);
or U680 (N_680,In_481,N_561);
nand U681 (N_681,N_450,N_525);
xor U682 (N_682,N_416,In_243);
and U683 (N_683,N_401,N_505);
or U684 (N_684,In_315,N_494);
xnor U685 (N_685,N_130,In_838);
or U686 (N_686,In_591,N_542);
or U687 (N_687,In_5,N_270);
and U688 (N_688,N_463,N_498);
and U689 (N_689,N_481,N_547);
or U690 (N_690,N_502,In_483);
or U691 (N_691,N_406,In_561);
and U692 (N_692,N_331,N_410);
and U693 (N_693,N_240,N_289);
nand U694 (N_694,N_236,N_545);
xnor U695 (N_695,N_499,N_456);
nand U696 (N_696,N_590,N_522);
nand U697 (N_697,N_573,N_96);
and U698 (N_698,N_317,In_920);
nor U699 (N_699,N_275,N_68);
nand U700 (N_700,N_555,N_156);
nor U701 (N_701,In_812,In_325);
or U702 (N_702,N_509,N_304);
nor U703 (N_703,N_215,N_532);
nand U704 (N_704,N_20,N_511);
or U705 (N_705,N_565,N_513);
nand U706 (N_706,N_589,In_109);
or U707 (N_707,In_144,In_382);
xnor U708 (N_708,N_378,N_594);
nor U709 (N_709,N_434,N_476);
and U710 (N_710,N_436,In_99);
and U711 (N_711,In_565,N_435);
and U712 (N_712,In_895,N_478);
nor U713 (N_713,N_122,N_448);
nand U714 (N_714,N_80,In_715);
nor U715 (N_715,In_574,In_683);
nor U716 (N_716,N_346,In_959);
xor U717 (N_717,N_521,In_218);
nor U718 (N_718,N_400,In_884);
nand U719 (N_719,N_388,In_846);
or U720 (N_720,N_591,N_588);
nor U721 (N_721,In_67,N_503);
and U722 (N_722,In_513,N_485);
nor U723 (N_723,N_554,In_515);
nor U724 (N_724,In_996,In_558);
or U725 (N_725,In_244,In_634);
nand U726 (N_726,N_177,N_352);
nor U727 (N_727,N_529,N_559);
or U728 (N_728,N_418,N_429);
and U729 (N_729,In_394,N_404);
nand U730 (N_730,N_407,In_212);
or U731 (N_731,In_840,In_310);
or U732 (N_732,N_413,N_409);
nand U733 (N_733,N_356,In_184);
nor U734 (N_734,N_382,N_425);
nand U735 (N_735,N_508,In_130);
or U736 (N_736,N_422,N_229);
or U737 (N_737,N_403,In_366);
and U738 (N_738,N_321,N_93);
or U739 (N_739,In_679,N_165);
nand U740 (N_740,N_438,N_551);
or U741 (N_741,N_208,N_598);
nor U742 (N_742,N_353,N_137);
xor U743 (N_743,In_434,N_395);
xor U744 (N_744,N_497,In_358);
and U745 (N_745,N_482,N_469);
or U746 (N_746,N_571,N_530);
or U747 (N_747,In_910,N_464);
nand U748 (N_748,In_661,N_221);
nor U749 (N_749,In_916,N_577);
xor U750 (N_750,N_454,N_492);
nand U751 (N_751,In_311,N_358);
and U752 (N_752,In_132,N_459);
and U753 (N_753,N_480,N_467);
and U754 (N_754,N_458,N_368);
nand U755 (N_755,In_595,In_91);
and U756 (N_756,N_432,N_524);
and U757 (N_757,N_19,N_453);
and U758 (N_758,N_412,In_33);
and U759 (N_759,N_512,N_566);
and U760 (N_760,N_251,N_546);
or U761 (N_761,In_535,N_64);
nand U762 (N_762,In_635,N_468);
and U763 (N_763,N_218,In_760);
nand U764 (N_764,N_344,N_584);
nor U765 (N_765,N_255,N_483);
or U766 (N_766,N_411,N_336);
or U767 (N_767,N_531,N_472);
nand U768 (N_768,N_536,N_583);
and U769 (N_769,N_223,In_913);
nand U770 (N_770,N_567,N_486);
or U771 (N_771,N_160,In_940);
xor U772 (N_772,N_552,N_528);
nor U773 (N_773,N_596,N_491);
and U774 (N_774,In_652,N_460);
nand U775 (N_775,N_440,N_520);
nand U776 (N_776,N_285,N_224);
nand U777 (N_777,N_541,N_79);
nand U778 (N_778,N_585,N_442);
nand U779 (N_779,N_408,N_477);
nor U780 (N_780,In_86,N_209);
nor U781 (N_781,N_332,In_711);
or U782 (N_782,N_519,N_586);
nand U783 (N_783,N_504,N_563);
nor U784 (N_784,N_576,N_233);
nor U785 (N_785,N_430,In_285);
and U786 (N_786,N_230,N_15);
nand U787 (N_787,N_298,N_239);
nand U788 (N_788,N_238,N_191);
nand U789 (N_789,N_447,In_721);
xor U790 (N_790,N_474,N_205);
nor U791 (N_791,N_343,N_428);
nand U792 (N_792,In_841,N_273);
nor U793 (N_793,N_465,N_461);
nand U794 (N_794,In_779,N_231);
and U795 (N_795,N_495,N_557);
xnor U796 (N_796,N_419,N_506);
xnor U797 (N_797,N_507,N_489);
and U798 (N_798,N_294,N_132);
nor U799 (N_799,N_377,N_323);
nor U800 (N_800,N_739,N_692);
nand U801 (N_801,N_762,N_766);
nor U802 (N_802,N_676,N_732);
or U803 (N_803,N_615,N_784);
nor U804 (N_804,N_665,N_715);
or U805 (N_805,N_771,N_672);
xor U806 (N_806,N_610,N_608);
xor U807 (N_807,N_668,N_798);
nand U808 (N_808,N_792,N_746);
nand U809 (N_809,N_708,N_768);
nor U810 (N_810,N_656,N_643);
or U811 (N_811,N_677,N_655);
and U812 (N_812,N_754,N_639);
nand U813 (N_813,N_737,N_662);
or U814 (N_814,N_783,N_764);
xnor U815 (N_815,N_620,N_795);
and U816 (N_816,N_735,N_648);
nand U817 (N_817,N_631,N_791);
nor U818 (N_818,N_763,N_779);
nand U819 (N_819,N_765,N_743);
and U820 (N_820,N_785,N_638);
nor U821 (N_821,N_790,N_748);
nor U822 (N_822,N_691,N_724);
or U823 (N_823,N_703,N_788);
nand U824 (N_824,N_759,N_720);
and U825 (N_825,N_757,N_617);
or U826 (N_826,N_714,N_742);
or U827 (N_827,N_761,N_778);
nand U828 (N_828,N_797,N_770);
or U829 (N_829,N_604,N_728);
and U830 (N_830,N_796,N_680);
xor U831 (N_831,N_725,N_736);
and U832 (N_832,N_693,N_637);
xor U833 (N_833,N_695,N_666);
and U834 (N_834,N_602,N_646);
nor U835 (N_835,N_729,N_696);
or U836 (N_836,N_682,N_740);
nor U837 (N_837,N_683,N_750);
nor U838 (N_838,N_640,N_701);
xor U839 (N_839,N_647,N_654);
or U840 (N_840,N_711,N_606);
nor U841 (N_841,N_653,N_685);
nor U842 (N_842,N_670,N_799);
and U843 (N_843,N_689,N_726);
or U844 (N_844,N_721,N_710);
and U845 (N_845,N_658,N_684);
or U846 (N_846,N_687,N_704);
nand U847 (N_847,N_694,N_649);
nor U848 (N_848,N_747,N_712);
nand U849 (N_849,N_702,N_776);
nand U850 (N_850,N_652,N_622);
or U851 (N_851,N_787,N_751);
or U852 (N_852,N_623,N_635);
nor U853 (N_853,N_699,N_744);
nor U854 (N_854,N_777,N_773);
or U855 (N_855,N_794,N_698);
nor U856 (N_856,N_719,N_674);
nor U857 (N_857,N_786,N_645);
or U858 (N_858,N_756,N_769);
nor U859 (N_859,N_612,N_772);
or U860 (N_860,N_621,N_650);
nor U861 (N_861,N_686,N_774);
and U862 (N_862,N_767,N_624);
and U863 (N_863,N_709,N_734);
or U864 (N_864,N_660,N_738);
nand U865 (N_865,N_664,N_760);
and U866 (N_866,N_630,N_629);
xnor U867 (N_867,N_789,N_793);
nand U868 (N_868,N_611,N_755);
nor U869 (N_869,N_633,N_716);
or U870 (N_870,N_758,N_781);
or U871 (N_871,N_659,N_673);
or U872 (N_872,N_613,N_727);
xor U873 (N_873,N_632,N_634);
and U874 (N_874,N_661,N_636);
or U875 (N_875,N_609,N_671);
and U876 (N_876,N_700,N_741);
nor U877 (N_877,N_679,N_625);
nor U878 (N_878,N_697,N_619);
nand U879 (N_879,N_723,N_675);
nand U880 (N_880,N_681,N_600);
nor U881 (N_881,N_780,N_753);
nor U882 (N_882,N_745,N_718);
nor U883 (N_883,N_657,N_603);
nor U884 (N_884,N_717,N_607);
and U885 (N_885,N_628,N_706);
nor U886 (N_886,N_713,N_722);
and U887 (N_887,N_618,N_626);
and U888 (N_888,N_775,N_678);
nand U889 (N_889,N_688,N_614);
and U890 (N_890,N_644,N_651);
and U891 (N_891,N_605,N_749);
and U892 (N_892,N_641,N_669);
nand U893 (N_893,N_731,N_601);
nand U894 (N_894,N_733,N_705);
and U895 (N_895,N_616,N_627);
or U896 (N_896,N_663,N_642);
xnor U897 (N_897,N_782,N_667);
or U898 (N_898,N_730,N_752);
nor U899 (N_899,N_690,N_707);
and U900 (N_900,N_630,N_626);
nor U901 (N_901,N_638,N_716);
nand U902 (N_902,N_751,N_659);
xnor U903 (N_903,N_659,N_797);
or U904 (N_904,N_744,N_621);
nand U905 (N_905,N_651,N_700);
nand U906 (N_906,N_789,N_621);
xor U907 (N_907,N_653,N_752);
nand U908 (N_908,N_631,N_605);
and U909 (N_909,N_626,N_726);
nor U910 (N_910,N_776,N_670);
or U911 (N_911,N_677,N_637);
and U912 (N_912,N_640,N_672);
nand U913 (N_913,N_677,N_659);
or U914 (N_914,N_712,N_782);
and U915 (N_915,N_741,N_733);
nor U916 (N_916,N_701,N_704);
nor U917 (N_917,N_743,N_720);
xnor U918 (N_918,N_713,N_654);
or U919 (N_919,N_689,N_760);
or U920 (N_920,N_719,N_749);
nand U921 (N_921,N_611,N_743);
or U922 (N_922,N_602,N_770);
or U923 (N_923,N_641,N_633);
or U924 (N_924,N_704,N_770);
or U925 (N_925,N_734,N_731);
nand U926 (N_926,N_657,N_785);
nor U927 (N_927,N_737,N_790);
and U928 (N_928,N_705,N_706);
nor U929 (N_929,N_789,N_672);
xor U930 (N_930,N_723,N_667);
nand U931 (N_931,N_740,N_625);
and U932 (N_932,N_742,N_691);
or U933 (N_933,N_723,N_631);
or U934 (N_934,N_637,N_777);
nand U935 (N_935,N_715,N_736);
or U936 (N_936,N_795,N_718);
and U937 (N_937,N_682,N_659);
nand U938 (N_938,N_743,N_641);
nand U939 (N_939,N_644,N_749);
or U940 (N_940,N_693,N_702);
nand U941 (N_941,N_751,N_649);
or U942 (N_942,N_683,N_758);
nand U943 (N_943,N_781,N_704);
or U944 (N_944,N_706,N_753);
and U945 (N_945,N_784,N_767);
or U946 (N_946,N_721,N_715);
nand U947 (N_947,N_706,N_723);
nor U948 (N_948,N_698,N_788);
nor U949 (N_949,N_789,N_629);
nand U950 (N_950,N_781,N_716);
or U951 (N_951,N_721,N_783);
and U952 (N_952,N_700,N_742);
nor U953 (N_953,N_622,N_636);
nand U954 (N_954,N_761,N_608);
and U955 (N_955,N_677,N_738);
nand U956 (N_956,N_750,N_618);
nor U957 (N_957,N_726,N_606);
xnor U958 (N_958,N_704,N_625);
nor U959 (N_959,N_733,N_651);
nor U960 (N_960,N_628,N_681);
nand U961 (N_961,N_711,N_799);
or U962 (N_962,N_670,N_758);
nand U963 (N_963,N_602,N_742);
or U964 (N_964,N_653,N_650);
nand U965 (N_965,N_761,N_663);
or U966 (N_966,N_675,N_705);
or U967 (N_967,N_703,N_608);
xnor U968 (N_968,N_781,N_755);
nand U969 (N_969,N_635,N_705);
nor U970 (N_970,N_782,N_756);
nand U971 (N_971,N_675,N_646);
nor U972 (N_972,N_680,N_784);
and U973 (N_973,N_768,N_605);
nand U974 (N_974,N_780,N_719);
nor U975 (N_975,N_636,N_697);
xnor U976 (N_976,N_633,N_747);
nor U977 (N_977,N_657,N_682);
nand U978 (N_978,N_664,N_722);
and U979 (N_979,N_790,N_639);
or U980 (N_980,N_662,N_630);
and U981 (N_981,N_754,N_649);
nor U982 (N_982,N_692,N_645);
nor U983 (N_983,N_713,N_753);
nand U984 (N_984,N_654,N_776);
and U985 (N_985,N_629,N_713);
nor U986 (N_986,N_746,N_730);
or U987 (N_987,N_736,N_753);
or U988 (N_988,N_605,N_704);
nand U989 (N_989,N_696,N_775);
and U990 (N_990,N_747,N_625);
or U991 (N_991,N_796,N_688);
nand U992 (N_992,N_621,N_711);
and U993 (N_993,N_778,N_631);
nor U994 (N_994,N_710,N_738);
and U995 (N_995,N_766,N_720);
xnor U996 (N_996,N_625,N_614);
or U997 (N_997,N_735,N_697);
and U998 (N_998,N_671,N_663);
nor U999 (N_999,N_738,N_685);
nor U1000 (N_1000,N_834,N_981);
nor U1001 (N_1001,N_831,N_818);
nor U1002 (N_1002,N_908,N_815);
nand U1003 (N_1003,N_878,N_976);
and U1004 (N_1004,N_935,N_968);
nand U1005 (N_1005,N_881,N_999);
and U1006 (N_1006,N_995,N_846);
and U1007 (N_1007,N_905,N_966);
or U1008 (N_1008,N_915,N_925);
and U1009 (N_1009,N_807,N_939);
xnor U1010 (N_1010,N_986,N_940);
and U1011 (N_1011,N_893,N_911);
or U1012 (N_1012,N_802,N_953);
and U1013 (N_1013,N_960,N_851);
nand U1014 (N_1014,N_829,N_882);
nand U1015 (N_1015,N_970,N_870);
and U1016 (N_1016,N_858,N_926);
xnor U1017 (N_1017,N_990,N_856);
nand U1018 (N_1018,N_890,N_848);
and U1019 (N_1019,N_934,N_988);
nand U1020 (N_1020,N_866,N_900);
or U1021 (N_1021,N_936,N_888);
and U1022 (N_1022,N_869,N_924);
nand U1023 (N_1023,N_942,N_898);
and U1024 (N_1024,N_983,N_806);
and U1025 (N_1025,N_808,N_827);
nand U1026 (N_1026,N_862,N_810);
nor U1027 (N_1027,N_956,N_883);
xor U1028 (N_1028,N_933,N_957);
or U1029 (N_1029,N_974,N_941);
or U1030 (N_1030,N_919,N_863);
or U1031 (N_1031,N_916,N_978);
xor U1032 (N_1032,N_906,N_964);
nor U1033 (N_1033,N_948,N_950);
or U1034 (N_1034,N_910,N_821);
xnor U1035 (N_1035,N_838,N_989);
or U1036 (N_1036,N_892,N_850);
or U1037 (N_1037,N_813,N_857);
nor U1038 (N_1038,N_843,N_938);
xnor U1039 (N_1039,N_822,N_947);
xnor U1040 (N_1040,N_969,N_820);
nand U1041 (N_1041,N_996,N_841);
nor U1042 (N_1042,N_994,N_823);
or U1043 (N_1043,N_971,N_868);
and U1044 (N_1044,N_932,N_979);
and U1045 (N_1045,N_958,N_965);
and U1046 (N_1046,N_904,N_800);
and U1047 (N_1047,N_842,N_853);
or U1048 (N_1048,N_861,N_975);
nor U1049 (N_1049,N_879,N_812);
nor U1050 (N_1050,N_951,N_859);
nand U1051 (N_1051,N_804,N_997);
or U1052 (N_1052,N_887,N_828);
and U1053 (N_1053,N_959,N_961);
nand U1054 (N_1054,N_907,N_944);
nand U1055 (N_1055,N_872,N_927);
or U1056 (N_1056,N_921,N_962);
nand U1057 (N_1057,N_946,N_897);
and U1058 (N_1058,N_895,N_844);
or U1059 (N_1059,N_805,N_832);
or U1060 (N_1060,N_903,N_922);
or U1061 (N_1061,N_918,N_836);
or U1062 (N_1062,N_884,N_867);
nand U1063 (N_1063,N_977,N_849);
nand U1064 (N_1064,N_991,N_937);
nor U1065 (N_1065,N_967,N_803);
nor U1066 (N_1066,N_901,N_817);
nor U1067 (N_1067,N_814,N_877);
nand U1068 (N_1068,N_839,N_913);
xor U1069 (N_1069,N_830,N_992);
nand U1070 (N_1070,N_837,N_801);
nor U1071 (N_1071,N_902,N_826);
xor U1072 (N_1072,N_825,N_917);
nor U1073 (N_1073,N_949,N_987);
xnor U1074 (N_1074,N_816,N_931);
or U1075 (N_1075,N_845,N_993);
and U1076 (N_1076,N_833,N_840);
or U1077 (N_1077,N_972,N_896);
nand U1078 (N_1078,N_847,N_955);
xnor U1079 (N_1079,N_860,N_912);
xnor U1080 (N_1080,N_928,N_899);
or U1081 (N_1081,N_909,N_929);
nand U1082 (N_1082,N_880,N_980);
and U1083 (N_1083,N_835,N_963);
and U1084 (N_1084,N_852,N_809);
and U1085 (N_1085,N_945,N_885);
nand U1086 (N_1086,N_854,N_824);
or U1087 (N_1087,N_855,N_865);
or U1088 (N_1088,N_954,N_982);
or U1089 (N_1089,N_894,N_923);
nor U1090 (N_1090,N_875,N_874);
or U1091 (N_1091,N_819,N_891);
and U1092 (N_1092,N_914,N_886);
nor U1093 (N_1093,N_984,N_930);
nand U1094 (N_1094,N_943,N_985);
xnor U1095 (N_1095,N_871,N_864);
xor U1096 (N_1096,N_973,N_876);
xnor U1097 (N_1097,N_873,N_811);
nor U1098 (N_1098,N_920,N_952);
or U1099 (N_1099,N_998,N_889);
or U1100 (N_1100,N_909,N_896);
and U1101 (N_1101,N_937,N_827);
nand U1102 (N_1102,N_936,N_915);
and U1103 (N_1103,N_844,N_954);
nand U1104 (N_1104,N_858,N_920);
or U1105 (N_1105,N_857,N_840);
xnor U1106 (N_1106,N_842,N_829);
or U1107 (N_1107,N_862,N_983);
nor U1108 (N_1108,N_943,N_915);
nor U1109 (N_1109,N_813,N_829);
nand U1110 (N_1110,N_995,N_913);
nor U1111 (N_1111,N_938,N_970);
or U1112 (N_1112,N_842,N_932);
nand U1113 (N_1113,N_952,N_858);
nor U1114 (N_1114,N_808,N_895);
nor U1115 (N_1115,N_890,N_825);
nor U1116 (N_1116,N_837,N_941);
or U1117 (N_1117,N_937,N_911);
nor U1118 (N_1118,N_861,N_823);
nand U1119 (N_1119,N_966,N_825);
nand U1120 (N_1120,N_876,N_816);
nor U1121 (N_1121,N_918,N_872);
or U1122 (N_1122,N_833,N_945);
or U1123 (N_1123,N_824,N_993);
nor U1124 (N_1124,N_991,N_878);
and U1125 (N_1125,N_810,N_894);
and U1126 (N_1126,N_909,N_931);
or U1127 (N_1127,N_910,N_961);
and U1128 (N_1128,N_802,N_874);
nand U1129 (N_1129,N_856,N_927);
or U1130 (N_1130,N_927,N_981);
xnor U1131 (N_1131,N_994,N_851);
nor U1132 (N_1132,N_980,N_814);
or U1133 (N_1133,N_871,N_974);
nand U1134 (N_1134,N_892,N_856);
nand U1135 (N_1135,N_993,N_924);
or U1136 (N_1136,N_985,N_880);
nor U1137 (N_1137,N_833,N_978);
nand U1138 (N_1138,N_949,N_806);
or U1139 (N_1139,N_997,N_846);
nand U1140 (N_1140,N_909,N_977);
or U1141 (N_1141,N_978,N_879);
or U1142 (N_1142,N_873,N_800);
nand U1143 (N_1143,N_908,N_872);
nor U1144 (N_1144,N_888,N_980);
nand U1145 (N_1145,N_949,N_940);
nor U1146 (N_1146,N_814,N_826);
or U1147 (N_1147,N_873,N_850);
nand U1148 (N_1148,N_940,N_868);
nand U1149 (N_1149,N_847,N_808);
nand U1150 (N_1150,N_824,N_948);
and U1151 (N_1151,N_801,N_889);
or U1152 (N_1152,N_932,N_936);
nand U1153 (N_1153,N_996,N_853);
nand U1154 (N_1154,N_816,N_903);
or U1155 (N_1155,N_939,N_888);
and U1156 (N_1156,N_833,N_809);
nand U1157 (N_1157,N_849,N_902);
or U1158 (N_1158,N_821,N_928);
nor U1159 (N_1159,N_978,N_856);
nand U1160 (N_1160,N_882,N_949);
and U1161 (N_1161,N_909,N_961);
xor U1162 (N_1162,N_847,N_821);
or U1163 (N_1163,N_976,N_877);
xnor U1164 (N_1164,N_811,N_917);
nand U1165 (N_1165,N_852,N_842);
nand U1166 (N_1166,N_807,N_806);
and U1167 (N_1167,N_857,N_994);
nand U1168 (N_1168,N_930,N_866);
nor U1169 (N_1169,N_804,N_842);
nor U1170 (N_1170,N_861,N_806);
nand U1171 (N_1171,N_900,N_966);
xor U1172 (N_1172,N_981,N_964);
and U1173 (N_1173,N_886,N_981);
or U1174 (N_1174,N_890,N_806);
nor U1175 (N_1175,N_937,N_934);
nand U1176 (N_1176,N_863,N_890);
or U1177 (N_1177,N_805,N_919);
and U1178 (N_1178,N_862,N_967);
nand U1179 (N_1179,N_933,N_866);
xor U1180 (N_1180,N_995,N_873);
and U1181 (N_1181,N_931,N_927);
nand U1182 (N_1182,N_847,N_909);
or U1183 (N_1183,N_952,N_841);
nor U1184 (N_1184,N_843,N_969);
and U1185 (N_1185,N_902,N_968);
nor U1186 (N_1186,N_890,N_891);
nor U1187 (N_1187,N_987,N_925);
and U1188 (N_1188,N_926,N_911);
nor U1189 (N_1189,N_997,N_861);
and U1190 (N_1190,N_998,N_985);
xor U1191 (N_1191,N_935,N_807);
and U1192 (N_1192,N_858,N_891);
nor U1193 (N_1193,N_897,N_973);
and U1194 (N_1194,N_991,N_837);
nor U1195 (N_1195,N_876,N_886);
and U1196 (N_1196,N_816,N_906);
xor U1197 (N_1197,N_881,N_852);
and U1198 (N_1198,N_949,N_989);
nand U1199 (N_1199,N_928,N_842);
or U1200 (N_1200,N_1187,N_1042);
or U1201 (N_1201,N_1127,N_1087);
and U1202 (N_1202,N_1168,N_1098);
nand U1203 (N_1203,N_1033,N_1173);
xnor U1204 (N_1204,N_1001,N_1156);
nand U1205 (N_1205,N_1015,N_1162);
nand U1206 (N_1206,N_1124,N_1140);
and U1207 (N_1207,N_1150,N_1163);
nor U1208 (N_1208,N_1021,N_1073);
nand U1209 (N_1209,N_1103,N_1059);
or U1210 (N_1210,N_1078,N_1153);
and U1211 (N_1211,N_1025,N_1097);
and U1212 (N_1212,N_1167,N_1071);
nand U1213 (N_1213,N_1100,N_1142);
nor U1214 (N_1214,N_1169,N_1111);
nand U1215 (N_1215,N_1003,N_1175);
nand U1216 (N_1216,N_1063,N_1113);
nand U1217 (N_1217,N_1010,N_1046);
and U1218 (N_1218,N_1037,N_1096);
or U1219 (N_1219,N_1084,N_1028);
or U1220 (N_1220,N_1136,N_1160);
nand U1221 (N_1221,N_1045,N_1104);
or U1222 (N_1222,N_1065,N_1008);
or U1223 (N_1223,N_1023,N_1157);
nor U1224 (N_1224,N_1102,N_1064);
nor U1225 (N_1225,N_1088,N_1129);
nand U1226 (N_1226,N_1004,N_1151);
nand U1227 (N_1227,N_1132,N_1165);
nand U1228 (N_1228,N_1043,N_1112);
nand U1229 (N_1229,N_1161,N_1182);
nand U1230 (N_1230,N_1079,N_1198);
and U1231 (N_1231,N_1119,N_1170);
or U1232 (N_1232,N_1070,N_1013);
and U1233 (N_1233,N_1032,N_1116);
and U1234 (N_1234,N_1190,N_1130);
and U1235 (N_1235,N_1176,N_1194);
nand U1236 (N_1236,N_1031,N_1081);
xor U1237 (N_1237,N_1179,N_1086);
nand U1238 (N_1238,N_1141,N_1094);
and U1239 (N_1239,N_1185,N_1137);
or U1240 (N_1240,N_1089,N_1083);
xor U1241 (N_1241,N_1044,N_1177);
nor U1242 (N_1242,N_1007,N_1125);
or U1243 (N_1243,N_1148,N_1074);
or U1244 (N_1244,N_1060,N_1047);
or U1245 (N_1245,N_1099,N_1134);
nand U1246 (N_1246,N_1155,N_1183);
nor U1247 (N_1247,N_1106,N_1020);
or U1248 (N_1248,N_1051,N_1154);
nor U1249 (N_1249,N_1159,N_1039);
nand U1250 (N_1250,N_1038,N_1006);
and U1251 (N_1251,N_1012,N_1196);
nand U1252 (N_1252,N_1055,N_1143);
or U1253 (N_1253,N_1067,N_1091);
xor U1254 (N_1254,N_1075,N_1062);
and U1255 (N_1255,N_1199,N_1195);
xnor U1256 (N_1256,N_1192,N_1061);
and U1257 (N_1257,N_1191,N_1178);
and U1258 (N_1258,N_1107,N_1002);
or U1259 (N_1259,N_1114,N_1054);
and U1260 (N_1260,N_1164,N_1068);
and U1261 (N_1261,N_1057,N_1066);
and U1262 (N_1262,N_1034,N_1174);
nand U1263 (N_1263,N_1026,N_1108);
and U1264 (N_1264,N_1128,N_1093);
nand U1265 (N_1265,N_1069,N_1058);
and U1266 (N_1266,N_1095,N_1048);
nor U1267 (N_1267,N_1105,N_1080);
nor U1268 (N_1268,N_1166,N_1120);
and U1269 (N_1269,N_1077,N_1030);
and U1270 (N_1270,N_1117,N_1109);
or U1271 (N_1271,N_1115,N_1139);
nand U1272 (N_1272,N_1040,N_1035);
or U1273 (N_1273,N_1009,N_1052);
or U1274 (N_1274,N_1122,N_1180);
nor U1275 (N_1275,N_1158,N_1029);
and U1276 (N_1276,N_1076,N_1147);
xor U1277 (N_1277,N_1022,N_1110);
or U1278 (N_1278,N_1138,N_1181);
nand U1279 (N_1279,N_1144,N_1171);
nor U1280 (N_1280,N_1050,N_1049);
nand U1281 (N_1281,N_1197,N_1131);
and U1282 (N_1282,N_1090,N_1149);
or U1283 (N_1283,N_1027,N_1172);
or U1284 (N_1284,N_1085,N_1005);
nand U1285 (N_1285,N_1123,N_1121);
or U1286 (N_1286,N_1024,N_1082);
and U1287 (N_1287,N_1017,N_1135);
and U1288 (N_1288,N_1072,N_1019);
and U1289 (N_1289,N_1053,N_1016);
or U1290 (N_1290,N_1133,N_1118);
or U1291 (N_1291,N_1189,N_1056);
nand U1292 (N_1292,N_1146,N_1014);
nor U1293 (N_1293,N_1092,N_1184);
nand U1294 (N_1294,N_1126,N_1041);
nor U1295 (N_1295,N_1152,N_1011);
nor U1296 (N_1296,N_1186,N_1193);
nand U1297 (N_1297,N_1101,N_1188);
or U1298 (N_1298,N_1036,N_1145);
or U1299 (N_1299,N_1000,N_1018);
or U1300 (N_1300,N_1168,N_1078);
nor U1301 (N_1301,N_1105,N_1152);
or U1302 (N_1302,N_1090,N_1150);
nor U1303 (N_1303,N_1040,N_1088);
nand U1304 (N_1304,N_1176,N_1005);
nand U1305 (N_1305,N_1052,N_1024);
or U1306 (N_1306,N_1114,N_1174);
nor U1307 (N_1307,N_1059,N_1166);
nand U1308 (N_1308,N_1178,N_1021);
and U1309 (N_1309,N_1074,N_1139);
or U1310 (N_1310,N_1198,N_1098);
and U1311 (N_1311,N_1003,N_1010);
nor U1312 (N_1312,N_1050,N_1144);
xor U1313 (N_1313,N_1018,N_1006);
nor U1314 (N_1314,N_1191,N_1073);
or U1315 (N_1315,N_1035,N_1100);
and U1316 (N_1316,N_1178,N_1176);
nand U1317 (N_1317,N_1004,N_1061);
nand U1318 (N_1318,N_1057,N_1106);
or U1319 (N_1319,N_1102,N_1072);
or U1320 (N_1320,N_1093,N_1034);
nor U1321 (N_1321,N_1086,N_1020);
nor U1322 (N_1322,N_1071,N_1108);
or U1323 (N_1323,N_1050,N_1181);
nor U1324 (N_1324,N_1138,N_1152);
and U1325 (N_1325,N_1197,N_1134);
or U1326 (N_1326,N_1031,N_1012);
or U1327 (N_1327,N_1055,N_1094);
nand U1328 (N_1328,N_1028,N_1116);
nor U1329 (N_1329,N_1068,N_1133);
and U1330 (N_1330,N_1013,N_1076);
nor U1331 (N_1331,N_1049,N_1036);
and U1332 (N_1332,N_1191,N_1141);
xor U1333 (N_1333,N_1181,N_1099);
nor U1334 (N_1334,N_1085,N_1105);
or U1335 (N_1335,N_1132,N_1113);
nand U1336 (N_1336,N_1050,N_1114);
and U1337 (N_1337,N_1161,N_1149);
or U1338 (N_1338,N_1125,N_1114);
nor U1339 (N_1339,N_1165,N_1121);
and U1340 (N_1340,N_1175,N_1002);
nor U1341 (N_1341,N_1043,N_1197);
nand U1342 (N_1342,N_1075,N_1004);
nor U1343 (N_1343,N_1042,N_1148);
and U1344 (N_1344,N_1061,N_1181);
and U1345 (N_1345,N_1174,N_1171);
nor U1346 (N_1346,N_1168,N_1129);
or U1347 (N_1347,N_1004,N_1190);
nand U1348 (N_1348,N_1172,N_1032);
and U1349 (N_1349,N_1016,N_1035);
or U1350 (N_1350,N_1074,N_1032);
and U1351 (N_1351,N_1049,N_1162);
and U1352 (N_1352,N_1115,N_1035);
nand U1353 (N_1353,N_1099,N_1177);
nor U1354 (N_1354,N_1153,N_1149);
nand U1355 (N_1355,N_1069,N_1139);
and U1356 (N_1356,N_1094,N_1047);
and U1357 (N_1357,N_1157,N_1052);
nand U1358 (N_1358,N_1067,N_1076);
nor U1359 (N_1359,N_1184,N_1055);
nor U1360 (N_1360,N_1004,N_1097);
nand U1361 (N_1361,N_1059,N_1087);
and U1362 (N_1362,N_1138,N_1050);
xor U1363 (N_1363,N_1074,N_1093);
nand U1364 (N_1364,N_1068,N_1191);
or U1365 (N_1365,N_1032,N_1071);
or U1366 (N_1366,N_1197,N_1196);
and U1367 (N_1367,N_1035,N_1157);
and U1368 (N_1368,N_1016,N_1112);
and U1369 (N_1369,N_1179,N_1080);
and U1370 (N_1370,N_1085,N_1034);
xor U1371 (N_1371,N_1144,N_1089);
nor U1372 (N_1372,N_1010,N_1160);
or U1373 (N_1373,N_1193,N_1058);
and U1374 (N_1374,N_1043,N_1016);
or U1375 (N_1375,N_1045,N_1173);
nor U1376 (N_1376,N_1178,N_1014);
or U1377 (N_1377,N_1079,N_1139);
or U1378 (N_1378,N_1077,N_1081);
nor U1379 (N_1379,N_1112,N_1113);
or U1380 (N_1380,N_1172,N_1115);
nand U1381 (N_1381,N_1126,N_1138);
nor U1382 (N_1382,N_1169,N_1141);
and U1383 (N_1383,N_1104,N_1041);
nand U1384 (N_1384,N_1059,N_1036);
and U1385 (N_1385,N_1127,N_1149);
or U1386 (N_1386,N_1170,N_1149);
nor U1387 (N_1387,N_1108,N_1155);
and U1388 (N_1388,N_1050,N_1175);
and U1389 (N_1389,N_1013,N_1088);
nor U1390 (N_1390,N_1090,N_1111);
or U1391 (N_1391,N_1064,N_1158);
nor U1392 (N_1392,N_1199,N_1148);
or U1393 (N_1393,N_1038,N_1145);
nand U1394 (N_1394,N_1153,N_1117);
xor U1395 (N_1395,N_1025,N_1064);
or U1396 (N_1396,N_1167,N_1124);
or U1397 (N_1397,N_1151,N_1181);
xor U1398 (N_1398,N_1132,N_1064);
nor U1399 (N_1399,N_1071,N_1139);
or U1400 (N_1400,N_1240,N_1256);
nor U1401 (N_1401,N_1284,N_1386);
nor U1402 (N_1402,N_1359,N_1371);
nand U1403 (N_1403,N_1220,N_1332);
and U1404 (N_1404,N_1327,N_1385);
and U1405 (N_1405,N_1306,N_1219);
and U1406 (N_1406,N_1211,N_1381);
nor U1407 (N_1407,N_1325,N_1206);
xnor U1408 (N_1408,N_1244,N_1213);
nand U1409 (N_1409,N_1315,N_1217);
nor U1410 (N_1410,N_1216,N_1391);
nor U1411 (N_1411,N_1369,N_1223);
and U1412 (N_1412,N_1235,N_1299);
nor U1413 (N_1413,N_1342,N_1328);
nand U1414 (N_1414,N_1203,N_1307);
xnor U1415 (N_1415,N_1287,N_1312);
and U1416 (N_1416,N_1208,N_1343);
nor U1417 (N_1417,N_1265,N_1282);
nand U1418 (N_1418,N_1224,N_1279);
nand U1419 (N_1419,N_1326,N_1276);
or U1420 (N_1420,N_1358,N_1255);
nor U1421 (N_1421,N_1237,N_1229);
nor U1422 (N_1422,N_1201,N_1399);
nand U1423 (N_1423,N_1210,N_1338);
and U1424 (N_1424,N_1238,N_1314);
or U1425 (N_1425,N_1200,N_1370);
nor U1426 (N_1426,N_1274,N_1245);
or U1427 (N_1427,N_1310,N_1364);
xor U1428 (N_1428,N_1266,N_1356);
or U1429 (N_1429,N_1335,N_1300);
nor U1430 (N_1430,N_1375,N_1372);
and U1431 (N_1431,N_1225,N_1374);
and U1432 (N_1432,N_1316,N_1227);
nor U1433 (N_1433,N_1344,N_1340);
and U1434 (N_1434,N_1383,N_1251);
nor U1435 (N_1435,N_1348,N_1246);
nand U1436 (N_1436,N_1302,N_1204);
or U1437 (N_1437,N_1352,N_1331);
or U1438 (N_1438,N_1259,N_1322);
nand U1439 (N_1439,N_1323,N_1263);
xnor U1440 (N_1440,N_1324,N_1289);
nor U1441 (N_1441,N_1269,N_1260);
nand U1442 (N_1442,N_1239,N_1257);
nor U1443 (N_1443,N_1268,N_1387);
or U1444 (N_1444,N_1295,N_1347);
nand U1445 (N_1445,N_1397,N_1281);
or U1446 (N_1446,N_1311,N_1275);
and U1447 (N_1447,N_1336,N_1360);
nand U1448 (N_1448,N_1277,N_1267);
or U1449 (N_1449,N_1258,N_1226);
nand U1450 (N_1450,N_1320,N_1373);
or U1451 (N_1451,N_1393,N_1313);
nor U1452 (N_1452,N_1233,N_1228);
nor U1453 (N_1453,N_1304,N_1218);
or U1454 (N_1454,N_1272,N_1384);
and U1455 (N_1455,N_1354,N_1388);
or U1456 (N_1456,N_1288,N_1234);
nand U1457 (N_1457,N_1247,N_1390);
nor U1458 (N_1458,N_1292,N_1243);
nor U1459 (N_1459,N_1330,N_1207);
nor U1460 (N_1460,N_1341,N_1377);
xor U1461 (N_1461,N_1270,N_1365);
and U1462 (N_1462,N_1396,N_1232);
xor U1463 (N_1463,N_1221,N_1293);
nand U1464 (N_1464,N_1273,N_1366);
nand U1465 (N_1465,N_1309,N_1361);
nor U1466 (N_1466,N_1298,N_1242);
xor U1467 (N_1467,N_1337,N_1205);
nand U1468 (N_1468,N_1253,N_1296);
nand U1469 (N_1469,N_1318,N_1264);
and U1470 (N_1470,N_1395,N_1280);
nand U1471 (N_1471,N_1346,N_1249);
nand U1472 (N_1472,N_1236,N_1286);
nor U1473 (N_1473,N_1367,N_1290);
nor U1474 (N_1474,N_1376,N_1261);
and U1475 (N_1475,N_1317,N_1212);
or U1476 (N_1476,N_1394,N_1378);
nand U1477 (N_1477,N_1355,N_1241);
nor U1478 (N_1478,N_1334,N_1252);
nand U1479 (N_1479,N_1329,N_1230);
and U1480 (N_1480,N_1214,N_1301);
nor U1481 (N_1481,N_1283,N_1303);
and U1482 (N_1482,N_1362,N_1345);
nand U1483 (N_1483,N_1285,N_1250);
nand U1484 (N_1484,N_1339,N_1380);
or U1485 (N_1485,N_1368,N_1308);
and U1486 (N_1486,N_1351,N_1215);
nand U1487 (N_1487,N_1271,N_1222);
or U1488 (N_1488,N_1254,N_1231);
and U1489 (N_1489,N_1379,N_1357);
xnor U1490 (N_1490,N_1389,N_1319);
and U1491 (N_1491,N_1333,N_1392);
or U1492 (N_1492,N_1349,N_1278);
nor U1493 (N_1493,N_1294,N_1398);
or U1494 (N_1494,N_1262,N_1209);
or U1495 (N_1495,N_1291,N_1202);
nor U1496 (N_1496,N_1248,N_1382);
nand U1497 (N_1497,N_1305,N_1363);
nor U1498 (N_1498,N_1353,N_1297);
nand U1499 (N_1499,N_1350,N_1321);
xor U1500 (N_1500,N_1355,N_1330);
or U1501 (N_1501,N_1336,N_1318);
or U1502 (N_1502,N_1218,N_1200);
nand U1503 (N_1503,N_1281,N_1226);
nor U1504 (N_1504,N_1207,N_1276);
nor U1505 (N_1505,N_1399,N_1214);
or U1506 (N_1506,N_1378,N_1201);
xor U1507 (N_1507,N_1345,N_1325);
and U1508 (N_1508,N_1330,N_1288);
and U1509 (N_1509,N_1256,N_1307);
and U1510 (N_1510,N_1295,N_1284);
and U1511 (N_1511,N_1228,N_1356);
nor U1512 (N_1512,N_1233,N_1215);
or U1513 (N_1513,N_1230,N_1248);
or U1514 (N_1514,N_1350,N_1281);
nor U1515 (N_1515,N_1326,N_1252);
nand U1516 (N_1516,N_1297,N_1372);
or U1517 (N_1517,N_1355,N_1329);
nand U1518 (N_1518,N_1297,N_1329);
nand U1519 (N_1519,N_1357,N_1261);
xnor U1520 (N_1520,N_1348,N_1289);
and U1521 (N_1521,N_1288,N_1278);
nor U1522 (N_1522,N_1348,N_1336);
nor U1523 (N_1523,N_1397,N_1358);
and U1524 (N_1524,N_1241,N_1358);
nor U1525 (N_1525,N_1314,N_1293);
or U1526 (N_1526,N_1320,N_1344);
nor U1527 (N_1527,N_1267,N_1324);
nand U1528 (N_1528,N_1315,N_1337);
nand U1529 (N_1529,N_1246,N_1248);
nor U1530 (N_1530,N_1325,N_1351);
nand U1531 (N_1531,N_1393,N_1341);
nand U1532 (N_1532,N_1377,N_1236);
or U1533 (N_1533,N_1207,N_1326);
and U1534 (N_1534,N_1375,N_1301);
or U1535 (N_1535,N_1367,N_1265);
nor U1536 (N_1536,N_1317,N_1373);
nor U1537 (N_1537,N_1336,N_1246);
nor U1538 (N_1538,N_1252,N_1317);
nand U1539 (N_1539,N_1211,N_1310);
nor U1540 (N_1540,N_1234,N_1229);
nand U1541 (N_1541,N_1309,N_1211);
and U1542 (N_1542,N_1252,N_1311);
or U1543 (N_1543,N_1325,N_1375);
nand U1544 (N_1544,N_1394,N_1317);
nor U1545 (N_1545,N_1239,N_1354);
and U1546 (N_1546,N_1382,N_1345);
nor U1547 (N_1547,N_1202,N_1390);
nand U1548 (N_1548,N_1397,N_1254);
or U1549 (N_1549,N_1364,N_1313);
or U1550 (N_1550,N_1309,N_1381);
nor U1551 (N_1551,N_1384,N_1217);
xnor U1552 (N_1552,N_1215,N_1246);
and U1553 (N_1553,N_1241,N_1224);
nand U1554 (N_1554,N_1239,N_1394);
and U1555 (N_1555,N_1349,N_1247);
nand U1556 (N_1556,N_1381,N_1258);
xnor U1557 (N_1557,N_1364,N_1263);
nor U1558 (N_1558,N_1397,N_1396);
nand U1559 (N_1559,N_1296,N_1301);
nand U1560 (N_1560,N_1308,N_1312);
and U1561 (N_1561,N_1277,N_1246);
nor U1562 (N_1562,N_1344,N_1261);
and U1563 (N_1563,N_1238,N_1301);
nand U1564 (N_1564,N_1261,N_1282);
nand U1565 (N_1565,N_1335,N_1329);
nand U1566 (N_1566,N_1326,N_1293);
or U1567 (N_1567,N_1387,N_1290);
and U1568 (N_1568,N_1270,N_1233);
or U1569 (N_1569,N_1372,N_1299);
or U1570 (N_1570,N_1386,N_1251);
and U1571 (N_1571,N_1393,N_1354);
or U1572 (N_1572,N_1223,N_1220);
nor U1573 (N_1573,N_1206,N_1240);
and U1574 (N_1574,N_1226,N_1291);
or U1575 (N_1575,N_1344,N_1268);
or U1576 (N_1576,N_1246,N_1292);
and U1577 (N_1577,N_1286,N_1358);
nor U1578 (N_1578,N_1342,N_1262);
or U1579 (N_1579,N_1386,N_1319);
nand U1580 (N_1580,N_1301,N_1258);
nand U1581 (N_1581,N_1368,N_1306);
nand U1582 (N_1582,N_1308,N_1302);
nand U1583 (N_1583,N_1215,N_1270);
or U1584 (N_1584,N_1325,N_1235);
or U1585 (N_1585,N_1261,N_1337);
nand U1586 (N_1586,N_1395,N_1350);
nand U1587 (N_1587,N_1361,N_1348);
or U1588 (N_1588,N_1220,N_1387);
nand U1589 (N_1589,N_1394,N_1219);
nand U1590 (N_1590,N_1357,N_1247);
and U1591 (N_1591,N_1312,N_1268);
xor U1592 (N_1592,N_1210,N_1244);
and U1593 (N_1593,N_1258,N_1385);
nor U1594 (N_1594,N_1344,N_1238);
nor U1595 (N_1595,N_1389,N_1224);
nand U1596 (N_1596,N_1280,N_1290);
xnor U1597 (N_1597,N_1390,N_1281);
or U1598 (N_1598,N_1332,N_1359);
xor U1599 (N_1599,N_1324,N_1319);
nand U1600 (N_1600,N_1461,N_1556);
nand U1601 (N_1601,N_1458,N_1439);
nor U1602 (N_1602,N_1516,N_1489);
nand U1603 (N_1603,N_1468,N_1583);
or U1604 (N_1604,N_1557,N_1412);
or U1605 (N_1605,N_1543,N_1418);
nand U1606 (N_1606,N_1416,N_1525);
and U1607 (N_1607,N_1490,N_1586);
nor U1608 (N_1608,N_1435,N_1579);
nand U1609 (N_1609,N_1502,N_1574);
and U1610 (N_1610,N_1441,N_1484);
nor U1611 (N_1611,N_1413,N_1582);
nor U1612 (N_1612,N_1560,N_1510);
and U1613 (N_1613,N_1514,N_1428);
nand U1614 (N_1614,N_1408,N_1425);
or U1615 (N_1615,N_1555,N_1464);
nand U1616 (N_1616,N_1528,N_1546);
or U1617 (N_1617,N_1496,N_1550);
or U1618 (N_1618,N_1478,N_1492);
nand U1619 (N_1619,N_1457,N_1553);
and U1620 (N_1620,N_1466,N_1533);
and U1621 (N_1621,N_1411,N_1534);
or U1622 (N_1622,N_1540,N_1563);
and U1623 (N_1623,N_1575,N_1436);
nor U1624 (N_1624,N_1498,N_1409);
or U1625 (N_1625,N_1432,N_1548);
or U1626 (N_1626,N_1505,N_1410);
xnor U1627 (N_1627,N_1415,N_1472);
and U1628 (N_1628,N_1508,N_1549);
xnor U1629 (N_1629,N_1482,N_1530);
or U1630 (N_1630,N_1519,N_1437);
and U1631 (N_1631,N_1451,N_1477);
or U1632 (N_1632,N_1531,N_1513);
nand U1633 (N_1633,N_1573,N_1442);
and U1634 (N_1634,N_1561,N_1568);
and U1635 (N_1635,N_1598,N_1544);
nor U1636 (N_1636,N_1558,N_1536);
nand U1637 (N_1637,N_1438,N_1571);
and U1638 (N_1638,N_1517,N_1597);
nor U1639 (N_1639,N_1471,N_1421);
nand U1640 (N_1640,N_1542,N_1520);
nor U1641 (N_1641,N_1515,N_1479);
xnor U1642 (N_1642,N_1587,N_1493);
nor U1643 (N_1643,N_1580,N_1456);
xor U1644 (N_1644,N_1446,N_1578);
and U1645 (N_1645,N_1404,N_1527);
nor U1646 (N_1646,N_1591,N_1547);
nand U1647 (N_1647,N_1552,N_1566);
xor U1648 (N_1648,N_1402,N_1440);
and U1649 (N_1649,N_1585,N_1538);
nand U1650 (N_1650,N_1599,N_1504);
or U1651 (N_1651,N_1433,N_1567);
nor U1652 (N_1652,N_1541,N_1511);
nor U1653 (N_1653,N_1532,N_1523);
or U1654 (N_1654,N_1562,N_1590);
nand U1655 (N_1655,N_1450,N_1455);
nand U1656 (N_1656,N_1524,N_1499);
nor U1657 (N_1657,N_1569,N_1431);
nand U1658 (N_1658,N_1494,N_1470);
or U1659 (N_1659,N_1426,N_1403);
nand U1660 (N_1660,N_1584,N_1491);
or U1661 (N_1661,N_1500,N_1414);
nand U1662 (N_1662,N_1526,N_1452);
nor U1663 (N_1663,N_1577,N_1529);
and U1664 (N_1664,N_1559,N_1592);
or U1665 (N_1665,N_1448,N_1488);
and U1666 (N_1666,N_1521,N_1429);
nor U1667 (N_1667,N_1475,N_1463);
nand U1668 (N_1668,N_1588,N_1424);
xor U1669 (N_1669,N_1509,N_1434);
or U1670 (N_1670,N_1443,N_1422);
and U1671 (N_1671,N_1564,N_1503);
nand U1672 (N_1672,N_1427,N_1483);
nand U1673 (N_1673,N_1487,N_1581);
nor U1674 (N_1674,N_1576,N_1565);
or U1675 (N_1675,N_1430,N_1594);
or U1676 (N_1676,N_1537,N_1518);
and U1677 (N_1677,N_1593,N_1405);
nor U1678 (N_1678,N_1485,N_1423);
xor U1679 (N_1679,N_1417,N_1449);
and U1680 (N_1680,N_1453,N_1465);
xor U1681 (N_1681,N_1460,N_1444);
and U1682 (N_1682,N_1407,N_1539);
nor U1683 (N_1683,N_1551,N_1570);
or U1684 (N_1684,N_1420,N_1486);
nand U1685 (N_1685,N_1535,N_1506);
and U1686 (N_1686,N_1400,N_1545);
nor U1687 (N_1687,N_1522,N_1469);
and U1688 (N_1688,N_1474,N_1596);
nand U1689 (N_1689,N_1462,N_1419);
and U1690 (N_1690,N_1480,N_1401);
nor U1691 (N_1691,N_1481,N_1454);
nand U1692 (N_1692,N_1497,N_1589);
and U1693 (N_1693,N_1572,N_1476);
xor U1694 (N_1694,N_1447,N_1512);
xnor U1695 (N_1695,N_1507,N_1495);
nand U1696 (N_1696,N_1467,N_1445);
and U1697 (N_1697,N_1406,N_1554);
or U1698 (N_1698,N_1473,N_1595);
or U1699 (N_1699,N_1501,N_1459);
and U1700 (N_1700,N_1428,N_1517);
and U1701 (N_1701,N_1468,N_1504);
or U1702 (N_1702,N_1473,N_1425);
or U1703 (N_1703,N_1525,N_1454);
nor U1704 (N_1704,N_1506,N_1541);
nand U1705 (N_1705,N_1551,N_1550);
nand U1706 (N_1706,N_1451,N_1426);
or U1707 (N_1707,N_1503,N_1416);
xor U1708 (N_1708,N_1503,N_1480);
and U1709 (N_1709,N_1554,N_1573);
and U1710 (N_1710,N_1449,N_1476);
nor U1711 (N_1711,N_1599,N_1417);
and U1712 (N_1712,N_1537,N_1469);
nor U1713 (N_1713,N_1459,N_1465);
or U1714 (N_1714,N_1543,N_1533);
nand U1715 (N_1715,N_1539,N_1449);
or U1716 (N_1716,N_1450,N_1472);
and U1717 (N_1717,N_1436,N_1494);
xor U1718 (N_1718,N_1447,N_1525);
xnor U1719 (N_1719,N_1493,N_1469);
and U1720 (N_1720,N_1580,N_1491);
or U1721 (N_1721,N_1418,N_1550);
and U1722 (N_1722,N_1566,N_1457);
and U1723 (N_1723,N_1472,N_1495);
and U1724 (N_1724,N_1515,N_1599);
or U1725 (N_1725,N_1404,N_1572);
xor U1726 (N_1726,N_1405,N_1509);
or U1727 (N_1727,N_1585,N_1540);
or U1728 (N_1728,N_1505,N_1572);
or U1729 (N_1729,N_1408,N_1440);
and U1730 (N_1730,N_1582,N_1562);
nand U1731 (N_1731,N_1532,N_1539);
nor U1732 (N_1732,N_1552,N_1461);
or U1733 (N_1733,N_1560,N_1442);
or U1734 (N_1734,N_1566,N_1556);
nor U1735 (N_1735,N_1484,N_1430);
nand U1736 (N_1736,N_1560,N_1456);
or U1737 (N_1737,N_1424,N_1426);
or U1738 (N_1738,N_1476,N_1422);
and U1739 (N_1739,N_1418,N_1554);
nor U1740 (N_1740,N_1573,N_1566);
or U1741 (N_1741,N_1471,N_1534);
and U1742 (N_1742,N_1457,N_1564);
or U1743 (N_1743,N_1578,N_1475);
or U1744 (N_1744,N_1507,N_1448);
nor U1745 (N_1745,N_1486,N_1413);
nand U1746 (N_1746,N_1524,N_1446);
and U1747 (N_1747,N_1499,N_1416);
xnor U1748 (N_1748,N_1408,N_1585);
and U1749 (N_1749,N_1599,N_1484);
and U1750 (N_1750,N_1456,N_1577);
nor U1751 (N_1751,N_1422,N_1423);
nand U1752 (N_1752,N_1522,N_1566);
xor U1753 (N_1753,N_1408,N_1545);
nor U1754 (N_1754,N_1540,N_1504);
and U1755 (N_1755,N_1448,N_1556);
nand U1756 (N_1756,N_1496,N_1529);
or U1757 (N_1757,N_1410,N_1422);
nand U1758 (N_1758,N_1493,N_1577);
nand U1759 (N_1759,N_1596,N_1523);
nand U1760 (N_1760,N_1449,N_1489);
nor U1761 (N_1761,N_1590,N_1595);
nand U1762 (N_1762,N_1450,N_1409);
nor U1763 (N_1763,N_1407,N_1526);
nor U1764 (N_1764,N_1448,N_1447);
nand U1765 (N_1765,N_1512,N_1584);
or U1766 (N_1766,N_1543,N_1466);
and U1767 (N_1767,N_1567,N_1531);
and U1768 (N_1768,N_1430,N_1455);
xnor U1769 (N_1769,N_1423,N_1594);
nor U1770 (N_1770,N_1559,N_1553);
and U1771 (N_1771,N_1561,N_1403);
and U1772 (N_1772,N_1577,N_1409);
and U1773 (N_1773,N_1414,N_1423);
nand U1774 (N_1774,N_1535,N_1454);
and U1775 (N_1775,N_1446,N_1570);
or U1776 (N_1776,N_1480,N_1505);
and U1777 (N_1777,N_1513,N_1538);
and U1778 (N_1778,N_1492,N_1575);
xor U1779 (N_1779,N_1560,N_1587);
and U1780 (N_1780,N_1518,N_1538);
nor U1781 (N_1781,N_1531,N_1446);
or U1782 (N_1782,N_1523,N_1401);
and U1783 (N_1783,N_1510,N_1526);
nor U1784 (N_1784,N_1516,N_1533);
nor U1785 (N_1785,N_1563,N_1527);
or U1786 (N_1786,N_1574,N_1549);
or U1787 (N_1787,N_1568,N_1519);
nand U1788 (N_1788,N_1537,N_1501);
or U1789 (N_1789,N_1475,N_1577);
nor U1790 (N_1790,N_1588,N_1423);
and U1791 (N_1791,N_1457,N_1485);
nor U1792 (N_1792,N_1528,N_1569);
and U1793 (N_1793,N_1592,N_1575);
or U1794 (N_1794,N_1584,N_1582);
and U1795 (N_1795,N_1571,N_1588);
and U1796 (N_1796,N_1529,N_1501);
nor U1797 (N_1797,N_1455,N_1413);
nand U1798 (N_1798,N_1579,N_1419);
or U1799 (N_1799,N_1436,N_1582);
and U1800 (N_1800,N_1670,N_1613);
nor U1801 (N_1801,N_1674,N_1718);
and U1802 (N_1802,N_1799,N_1754);
nand U1803 (N_1803,N_1702,N_1777);
nor U1804 (N_1804,N_1774,N_1685);
nand U1805 (N_1805,N_1601,N_1672);
xor U1806 (N_1806,N_1679,N_1719);
nor U1807 (N_1807,N_1713,N_1639);
or U1808 (N_1808,N_1642,N_1616);
or U1809 (N_1809,N_1664,N_1614);
and U1810 (N_1810,N_1689,N_1740);
xor U1811 (N_1811,N_1705,N_1603);
xor U1812 (N_1812,N_1759,N_1757);
xnor U1813 (N_1813,N_1786,N_1645);
nand U1814 (N_1814,N_1608,N_1605);
nand U1815 (N_1815,N_1658,N_1791);
nor U1816 (N_1816,N_1765,N_1681);
nand U1817 (N_1817,N_1646,N_1634);
xnor U1818 (N_1818,N_1723,N_1694);
nand U1819 (N_1819,N_1652,N_1633);
xnor U1820 (N_1820,N_1732,N_1751);
nor U1821 (N_1821,N_1738,N_1714);
nand U1822 (N_1822,N_1688,N_1660);
and U1823 (N_1823,N_1687,N_1675);
or U1824 (N_1824,N_1650,N_1797);
and U1825 (N_1825,N_1742,N_1769);
nand U1826 (N_1826,N_1612,N_1678);
xnor U1827 (N_1827,N_1607,N_1782);
xor U1828 (N_1828,N_1620,N_1625);
nor U1829 (N_1829,N_1667,N_1695);
nand U1830 (N_1830,N_1651,N_1699);
nor U1831 (N_1831,N_1771,N_1728);
nor U1832 (N_1832,N_1710,N_1731);
and U1833 (N_1833,N_1730,N_1647);
nand U1834 (N_1834,N_1789,N_1609);
and U1835 (N_1835,N_1635,N_1746);
nor U1836 (N_1836,N_1764,N_1669);
or U1837 (N_1837,N_1690,N_1680);
or U1838 (N_1838,N_1706,N_1700);
nand U1839 (N_1839,N_1767,N_1632);
nand U1840 (N_1840,N_1733,N_1693);
xor U1841 (N_1841,N_1661,N_1788);
or U1842 (N_1842,N_1737,N_1643);
or U1843 (N_1843,N_1677,N_1743);
xor U1844 (N_1844,N_1692,N_1659);
or U1845 (N_1845,N_1709,N_1766);
or U1846 (N_1846,N_1768,N_1739);
or U1847 (N_1847,N_1711,N_1747);
nor U1848 (N_1848,N_1626,N_1729);
nand U1849 (N_1849,N_1798,N_1668);
nor U1850 (N_1850,N_1644,N_1734);
nand U1851 (N_1851,N_1686,N_1655);
and U1852 (N_1852,N_1794,N_1630);
nor U1853 (N_1853,N_1785,N_1621);
nand U1854 (N_1854,N_1665,N_1629);
nor U1855 (N_1855,N_1758,N_1755);
and U1856 (N_1856,N_1727,N_1779);
nor U1857 (N_1857,N_1796,N_1671);
nand U1858 (N_1858,N_1673,N_1624);
nor U1859 (N_1859,N_1648,N_1781);
or U1860 (N_1860,N_1745,N_1795);
and U1861 (N_1861,N_1666,N_1749);
or U1862 (N_1862,N_1707,N_1683);
nand U1863 (N_1863,N_1638,N_1750);
nor U1864 (N_1864,N_1783,N_1619);
or U1865 (N_1865,N_1610,N_1762);
and U1866 (N_1866,N_1721,N_1691);
and U1867 (N_1867,N_1703,N_1604);
nor U1868 (N_1868,N_1752,N_1676);
or U1869 (N_1869,N_1627,N_1631);
and U1870 (N_1870,N_1623,N_1708);
and U1871 (N_1871,N_1663,N_1773);
xor U1872 (N_1872,N_1717,N_1726);
or U1873 (N_1873,N_1617,N_1784);
or U1874 (N_1874,N_1761,N_1760);
nand U1875 (N_1875,N_1600,N_1780);
nor U1876 (N_1876,N_1720,N_1715);
nand U1877 (N_1877,N_1772,N_1641);
and U1878 (N_1878,N_1763,N_1770);
nand U1879 (N_1879,N_1776,N_1649);
nor U1880 (N_1880,N_1640,N_1793);
or U1881 (N_1881,N_1744,N_1722);
nand U1882 (N_1882,N_1778,N_1622);
nand U1883 (N_1883,N_1735,N_1654);
and U1884 (N_1884,N_1637,N_1682);
and U1885 (N_1885,N_1790,N_1724);
and U1886 (N_1886,N_1662,N_1712);
nand U1887 (N_1887,N_1696,N_1725);
and U1888 (N_1888,N_1602,N_1704);
nor U1889 (N_1889,N_1787,N_1792);
nand U1890 (N_1890,N_1684,N_1698);
or U1891 (N_1891,N_1628,N_1741);
or U1892 (N_1892,N_1748,N_1756);
xor U1893 (N_1893,N_1615,N_1775);
xnor U1894 (N_1894,N_1701,N_1618);
or U1895 (N_1895,N_1657,N_1636);
and U1896 (N_1896,N_1656,N_1611);
nor U1897 (N_1897,N_1753,N_1697);
nor U1898 (N_1898,N_1716,N_1653);
and U1899 (N_1899,N_1736,N_1606);
or U1900 (N_1900,N_1679,N_1738);
and U1901 (N_1901,N_1762,N_1607);
nand U1902 (N_1902,N_1651,N_1687);
nand U1903 (N_1903,N_1776,N_1780);
or U1904 (N_1904,N_1735,N_1694);
or U1905 (N_1905,N_1653,N_1765);
and U1906 (N_1906,N_1765,N_1606);
nand U1907 (N_1907,N_1672,N_1751);
or U1908 (N_1908,N_1616,N_1675);
nor U1909 (N_1909,N_1697,N_1635);
nor U1910 (N_1910,N_1613,N_1699);
or U1911 (N_1911,N_1668,N_1600);
or U1912 (N_1912,N_1700,N_1631);
or U1913 (N_1913,N_1628,N_1714);
and U1914 (N_1914,N_1701,N_1733);
nor U1915 (N_1915,N_1606,N_1639);
nor U1916 (N_1916,N_1778,N_1620);
and U1917 (N_1917,N_1608,N_1752);
nor U1918 (N_1918,N_1720,N_1749);
nand U1919 (N_1919,N_1738,N_1757);
and U1920 (N_1920,N_1727,N_1654);
nor U1921 (N_1921,N_1652,N_1617);
and U1922 (N_1922,N_1708,N_1629);
nand U1923 (N_1923,N_1637,N_1606);
and U1924 (N_1924,N_1677,N_1793);
nor U1925 (N_1925,N_1658,N_1628);
nand U1926 (N_1926,N_1726,N_1718);
xor U1927 (N_1927,N_1735,N_1665);
nor U1928 (N_1928,N_1617,N_1621);
nand U1929 (N_1929,N_1653,N_1750);
and U1930 (N_1930,N_1701,N_1600);
and U1931 (N_1931,N_1662,N_1635);
nor U1932 (N_1932,N_1773,N_1757);
xnor U1933 (N_1933,N_1629,N_1747);
or U1934 (N_1934,N_1771,N_1614);
and U1935 (N_1935,N_1615,N_1694);
nor U1936 (N_1936,N_1698,N_1769);
xor U1937 (N_1937,N_1659,N_1686);
nand U1938 (N_1938,N_1706,N_1613);
nand U1939 (N_1939,N_1711,N_1684);
or U1940 (N_1940,N_1651,N_1762);
or U1941 (N_1941,N_1758,N_1660);
nand U1942 (N_1942,N_1616,N_1796);
and U1943 (N_1943,N_1763,N_1624);
nand U1944 (N_1944,N_1728,N_1733);
and U1945 (N_1945,N_1794,N_1702);
nand U1946 (N_1946,N_1652,N_1610);
nor U1947 (N_1947,N_1659,N_1633);
or U1948 (N_1948,N_1788,N_1753);
nand U1949 (N_1949,N_1631,N_1723);
and U1950 (N_1950,N_1683,N_1614);
nor U1951 (N_1951,N_1729,N_1602);
nand U1952 (N_1952,N_1607,N_1687);
or U1953 (N_1953,N_1601,N_1610);
or U1954 (N_1954,N_1740,N_1665);
and U1955 (N_1955,N_1628,N_1635);
nor U1956 (N_1956,N_1765,N_1750);
nor U1957 (N_1957,N_1786,N_1663);
nand U1958 (N_1958,N_1755,N_1625);
and U1959 (N_1959,N_1696,N_1626);
nor U1960 (N_1960,N_1754,N_1735);
nand U1961 (N_1961,N_1641,N_1634);
nand U1962 (N_1962,N_1757,N_1701);
and U1963 (N_1963,N_1645,N_1798);
and U1964 (N_1964,N_1661,N_1659);
or U1965 (N_1965,N_1616,N_1614);
and U1966 (N_1966,N_1611,N_1747);
or U1967 (N_1967,N_1650,N_1612);
or U1968 (N_1968,N_1775,N_1789);
nor U1969 (N_1969,N_1650,N_1745);
nor U1970 (N_1970,N_1633,N_1729);
and U1971 (N_1971,N_1603,N_1659);
or U1972 (N_1972,N_1691,N_1656);
and U1973 (N_1973,N_1737,N_1612);
nor U1974 (N_1974,N_1670,N_1635);
nor U1975 (N_1975,N_1744,N_1628);
or U1976 (N_1976,N_1664,N_1702);
and U1977 (N_1977,N_1608,N_1672);
and U1978 (N_1978,N_1637,N_1614);
or U1979 (N_1979,N_1670,N_1787);
xor U1980 (N_1980,N_1619,N_1710);
xor U1981 (N_1981,N_1781,N_1662);
nor U1982 (N_1982,N_1612,N_1613);
nand U1983 (N_1983,N_1752,N_1708);
or U1984 (N_1984,N_1688,N_1687);
and U1985 (N_1985,N_1679,N_1605);
nand U1986 (N_1986,N_1721,N_1780);
and U1987 (N_1987,N_1784,N_1717);
and U1988 (N_1988,N_1752,N_1631);
nor U1989 (N_1989,N_1792,N_1689);
or U1990 (N_1990,N_1706,N_1682);
and U1991 (N_1991,N_1741,N_1622);
or U1992 (N_1992,N_1758,N_1712);
nor U1993 (N_1993,N_1626,N_1676);
and U1994 (N_1994,N_1715,N_1670);
nand U1995 (N_1995,N_1742,N_1655);
and U1996 (N_1996,N_1616,N_1709);
or U1997 (N_1997,N_1640,N_1750);
or U1998 (N_1998,N_1747,N_1698);
or U1999 (N_1999,N_1703,N_1774);
and U2000 (N_2000,N_1839,N_1865);
and U2001 (N_2001,N_1949,N_1935);
nor U2002 (N_2002,N_1928,N_1892);
and U2003 (N_2003,N_1805,N_1912);
nor U2004 (N_2004,N_1983,N_1859);
nand U2005 (N_2005,N_1988,N_1994);
xor U2006 (N_2006,N_1885,N_1884);
or U2007 (N_2007,N_1960,N_1840);
or U2008 (N_2008,N_1851,N_1899);
or U2009 (N_2009,N_1973,N_1990);
nor U2010 (N_2010,N_1802,N_1804);
nand U2011 (N_2011,N_1958,N_1801);
nand U2012 (N_2012,N_1893,N_1843);
or U2013 (N_2013,N_1933,N_1909);
xor U2014 (N_2014,N_1830,N_1882);
and U2015 (N_2015,N_1929,N_1809);
and U2016 (N_2016,N_1931,N_1905);
nor U2017 (N_2017,N_1992,N_1901);
nor U2018 (N_2018,N_1820,N_1985);
nand U2019 (N_2019,N_1854,N_1846);
and U2020 (N_2020,N_1926,N_1991);
or U2021 (N_2021,N_1902,N_1955);
nor U2022 (N_2022,N_1925,N_1816);
nand U2023 (N_2023,N_1808,N_1922);
nand U2024 (N_2024,N_1944,N_1824);
nand U2025 (N_2025,N_1908,N_1996);
nor U2026 (N_2026,N_1858,N_1860);
and U2027 (N_2027,N_1976,N_1867);
xnor U2028 (N_2028,N_1880,N_1962);
nor U2029 (N_2029,N_1980,N_1900);
and U2030 (N_2030,N_1965,N_1868);
and U2031 (N_2031,N_1982,N_1815);
nor U2032 (N_2032,N_1924,N_1853);
nor U2033 (N_2033,N_1930,N_1869);
or U2034 (N_2034,N_1817,N_1827);
or U2035 (N_2035,N_1977,N_1981);
nor U2036 (N_2036,N_1857,N_1891);
and U2037 (N_2037,N_1995,N_1812);
or U2038 (N_2038,N_1806,N_1975);
or U2039 (N_2039,N_1946,N_1932);
xor U2040 (N_2040,N_1837,N_1948);
nor U2041 (N_2041,N_1898,N_1941);
or U2042 (N_2042,N_1813,N_1997);
nor U2043 (N_2043,N_1819,N_1870);
or U2044 (N_2044,N_1845,N_1942);
nor U2045 (N_2045,N_1896,N_1842);
nor U2046 (N_2046,N_1957,N_1886);
and U2047 (N_2047,N_1823,N_1807);
or U2048 (N_2048,N_1852,N_1921);
nand U2049 (N_2049,N_1906,N_1974);
nand U2050 (N_2050,N_1923,N_1826);
nor U2051 (N_2051,N_1879,N_1895);
and U2052 (N_2052,N_1876,N_1822);
and U2053 (N_2053,N_1864,N_1866);
xor U2054 (N_2054,N_1940,N_1943);
xor U2055 (N_2055,N_1874,N_1938);
nor U2056 (N_2056,N_1832,N_1849);
and U2057 (N_2057,N_1881,N_1951);
or U2058 (N_2058,N_1966,N_1835);
nand U2059 (N_2059,N_1978,N_1836);
nor U2060 (N_2060,N_1916,N_1862);
xnor U2061 (N_2061,N_1829,N_1918);
nand U2062 (N_2062,N_1877,N_1959);
and U2063 (N_2063,N_1844,N_1831);
or U2064 (N_2064,N_1999,N_1917);
and U2065 (N_2065,N_1936,N_1847);
or U2066 (N_2066,N_1800,N_1937);
and U2067 (N_2067,N_1889,N_1961);
nor U2068 (N_2068,N_1971,N_1903);
nor U2069 (N_2069,N_1972,N_1863);
xor U2070 (N_2070,N_1915,N_1927);
or U2071 (N_2071,N_1911,N_1848);
or U2072 (N_2072,N_1811,N_1968);
nor U2073 (N_2073,N_1970,N_1821);
or U2074 (N_2074,N_1894,N_1952);
or U2075 (N_2075,N_1803,N_1913);
and U2076 (N_2076,N_1883,N_1838);
and U2077 (N_2077,N_1956,N_1963);
nand U2078 (N_2078,N_1871,N_1834);
nor U2079 (N_2079,N_1998,N_1910);
and U2080 (N_2080,N_1861,N_1856);
or U2081 (N_2081,N_1914,N_1833);
nand U2082 (N_2082,N_1986,N_1873);
xor U2083 (N_2083,N_1945,N_1810);
or U2084 (N_2084,N_1950,N_1904);
nor U2085 (N_2085,N_1964,N_1969);
nand U2086 (N_2086,N_1993,N_1939);
or U2087 (N_2087,N_1828,N_1825);
and U2088 (N_2088,N_1855,N_1814);
nor U2089 (N_2089,N_1875,N_1907);
nor U2090 (N_2090,N_1841,N_1872);
nor U2091 (N_2091,N_1818,N_1989);
or U2092 (N_2092,N_1947,N_1967);
nand U2093 (N_2093,N_1920,N_1953);
nor U2094 (N_2094,N_1888,N_1979);
and U2095 (N_2095,N_1934,N_1919);
or U2096 (N_2096,N_1984,N_1897);
nand U2097 (N_2097,N_1890,N_1850);
nor U2098 (N_2098,N_1954,N_1987);
nand U2099 (N_2099,N_1887,N_1878);
nor U2100 (N_2100,N_1906,N_1957);
and U2101 (N_2101,N_1841,N_1914);
and U2102 (N_2102,N_1827,N_1824);
nand U2103 (N_2103,N_1899,N_1914);
or U2104 (N_2104,N_1887,N_1971);
nand U2105 (N_2105,N_1901,N_1971);
nand U2106 (N_2106,N_1992,N_1924);
or U2107 (N_2107,N_1887,N_1911);
nand U2108 (N_2108,N_1939,N_1866);
nand U2109 (N_2109,N_1993,N_1852);
and U2110 (N_2110,N_1991,N_1929);
nand U2111 (N_2111,N_1969,N_1873);
or U2112 (N_2112,N_1992,N_1951);
nand U2113 (N_2113,N_1897,N_1942);
or U2114 (N_2114,N_1836,N_1919);
and U2115 (N_2115,N_1962,N_1909);
nor U2116 (N_2116,N_1847,N_1824);
nor U2117 (N_2117,N_1920,N_1985);
or U2118 (N_2118,N_1993,N_1844);
or U2119 (N_2119,N_1923,N_1924);
and U2120 (N_2120,N_1804,N_1896);
xnor U2121 (N_2121,N_1803,N_1935);
nand U2122 (N_2122,N_1842,N_1837);
and U2123 (N_2123,N_1836,N_1812);
or U2124 (N_2124,N_1820,N_1922);
or U2125 (N_2125,N_1925,N_1878);
or U2126 (N_2126,N_1971,N_1881);
nor U2127 (N_2127,N_1995,N_1996);
and U2128 (N_2128,N_1948,N_1830);
nor U2129 (N_2129,N_1803,N_1821);
nor U2130 (N_2130,N_1839,N_1807);
nor U2131 (N_2131,N_1855,N_1913);
nor U2132 (N_2132,N_1947,N_1843);
or U2133 (N_2133,N_1920,N_1871);
xnor U2134 (N_2134,N_1854,N_1912);
nand U2135 (N_2135,N_1974,N_1938);
nand U2136 (N_2136,N_1975,N_1831);
or U2137 (N_2137,N_1885,N_1933);
or U2138 (N_2138,N_1998,N_1958);
and U2139 (N_2139,N_1983,N_1847);
xor U2140 (N_2140,N_1911,N_1908);
nor U2141 (N_2141,N_1942,N_1903);
nand U2142 (N_2142,N_1844,N_1987);
nand U2143 (N_2143,N_1917,N_1901);
nand U2144 (N_2144,N_1812,N_1927);
nor U2145 (N_2145,N_1855,N_1988);
xor U2146 (N_2146,N_1914,N_1985);
and U2147 (N_2147,N_1940,N_1869);
nor U2148 (N_2148,N_1844,N_1967);
and U2149 (N_2149,N_1803,N_1863);
xnor U2150 (N_2150,N_1876,N_1963);
nor U2151 (N_2151,N_1933,N_1977);
nor U2152 (N_2152,N_1977,N_1901);
nor U2153 (N_2153,N_1984,N_1982);
xnor U2154 (N_2154,N_1856,N_1843);
and U2155 (N_2155,N_1996,N_1861);
or U2156 (N_2156,N_1976,N_1975);
nand U2157 (N_2157,N_1982,N_1957);
or U2158 (N_2158,N_1927,N_1941);
xor U2159 (N_2159,N_1849,N_1950);
nand U2160 (N_2160,N_1946,N_1986);
or U2161 (N_2161,N_1976,N_1979);
or U2162 (N_2162,N_1848,N_1956);
xnor U2163 (N_2163,N_1862,N_1911);
or U2164 (N_2164,N_1824,N_1818);
xor U2165 (N_2165,N_1847,N_1950);
nand U2166 (N_2166,N_1993,N_1900);
or U2167 (N_2167,N_1920,N_1947);
xnor U2168 (N_2168,N_1819,N_1973);
nand U2169 (N_2169,N_1927,N_1824);
nand U2170 (N_2170,N_1966,N_1913);
and U2171 (N_2171,N_1858,N_1800);
nor U2172 (N_2172,N_1960,N_1899);
and U2173 (N_2173,N_1830,N_1810);
xor U2174 (N_2174,N_1971,N_1908);
and U2175 (N_2175,N_1969,N_1958);
nor U2176 (N_2176,N_1832,N_1846);
and U2177 (N_2177,N_1852,N_1873);
and U2178 (N_2178,N_1897,N_1873);
nand U2179 (N_2179,N_1904,N_1929);
nor U2180 (N_2180,N_1862,N_1934);
nand U2181 (N_2181,N_1963,N_1878);
or U2182 (N_2182,N_1937,N_1824);
nor U2183 (N_2183,N_1917,N_1930);
nor U2184 (N_2184,N_1978,N_1850);
nand U2185 (N_2185,N_1866,N_1867);
or U2186 (N_2186,N_1968,N_1851);
or U2187 (N_2187,N_1887,N_1854);
and U2188 (N_2188,N_1951,N_1890);
nor U2189 (N_2189,N_1904,N_1919);
or U2190 (N_2190,N_1881,N_1985);
nand U2191 (N_2191,N_1827,N_1908);
or U2192 (N_2192,N_1955,N_1839);
nand U2193 (N_2193,N_1821,N_1861);
or U2194 (N_2194,N_1877,N_1956);
nor U2195 (N_2195,N_1868,N_1905);
nor U2196 (N_2196,N_1847,N_1949);
nor U2197 (N_2197,N_1985,N_1931);
xor U2198 (N_2198,N_1821,N_1938);
or U2199 (N_2199,N_1923,N_1908);
xor U2200 (N_2200,N_2071,N_2090);
nand U2201 (N_2201,N_2152,N_2045);
nor U2202 (N_2202,N_2157,N_2008);
nand U2203 (N_2203,N_2098,N_2002);
nand U2204 (N_2204,N_2001,N_2130);
nand U2205 (N_2205,N_2027,N_2083);
nor U2206 (N_2206,N_2145,N_2096);
or U2207 (N_2207,N_2012,N_2177);
nor U2208 (N_2208,N_2113,N_2031);
and U2209 (N_2209,N_2161,N_2184);
xor U2210 (N_2210,N_2040,N_2126);
xor U2211 (N_2211,N_2064,N_2170);
and U2212 (N_2212,N_2060,N_2165);
or U2213 (N_2213,N_2057,N_2086);
and U2214 (N_2214,N_2179,N_2114);
nor U2215 (N_2215,N_2029,N_2169);
and U2216 (N_2216,N_2021,N_2017);
nand U2217 (N_2217,N_2076,N_2058);
or U2218 (N_2218,N_2042,N_2055);
xnor U2219 (N_2219,N_2156,N_2120);
or U2220 (N_2220,N_2051,N_2011);
and U2221 (N_2221,N_2041,N_2009);
and U2222 (N_2222,N_2033,N_2054);
and U2223 (N_2223,N_2081,N_2121);
nor U2224 (N_2224,N_2149,N_2155);
or U2225 (N_2225,N_2070,N_2192);
or U2226 (N_2226,N_2139,N_2061);
and U2227 (N_2227,N_2151,N_2185);
nand U2228 (N_2228,N_2117,N_2122);
and U2229 (N_2229,N_2099,N_2043);
nor U2230 (N_2230,N_2075,N_2072);
and U2231 (N_2231,N_2162,N_2014);
nor U2232 (N_2232,N_2087,N_2148);
nor U2233 (N_2233,N_2078,N_2074);
nand U2234 (N_2234,N_2197,N_2143);
or U2235 (N_2235,N_2102,N_2023);
and U2236 (N_2236,N_2183,N_2007);
nor U2237 (N_2237,N_2127,N_2104);
nand U2238 (N_2238,N_2025,N_2188);
or U2239 (N_2239,N_2091,N_2168);
or U2240 (N_2240,N_2080,N_2039);
nand U2241 (N_2241,N_2085,N_2089);
or U2242 (N_2242,N_2174,N_2140);
nor U2243 (N_2243,N_2034,N_2144);
nor U2244 (N_2244,N_2022,N_2196);
xnor U2245 (N_2245,N_2134,N_2059);
nor U2246 (N_2246,N_2178,N_2065);
and U2247 (N_2247,N_2180,N_2082);
and U2248 (N_2248,N_2154,N_2044);
nor U2249 (N_2249,N_2147,N_2181);
or U2250 (N_2250,N_2146,N_2171);
or U2251 (N_2251,N_2173,N_2131);
nor U2252 (N_2252,N_2133,N_2084);
xor U2253 (N_2253,N_2110,N_2123);
xor U2254 (N_2254,N_2115,N_2172);
xnor U2255 (N_2255,N_2164,N_2079);
or U2256 (N_2256,N_2019,N_2046);
or U2257 (N_2257,N_2138,N_2119);
and U2258 (N_2258,N_2010,N_2056);
nand U2259 (N_2259,N_2105,N_2160);
or U2260 (N_2260,N_2063,N_2048);
and U2261 (N_2261,N_2015,N_2000);
and U2262 (N_2262,N_2189,N_2038);
or U2263 (N_2263,N_2136,N_2153);
and U2264 (N_2264,N_2124,N_2112);
or U2265 (N_2265,N_2109,N_2069);
nor U2266 (N_2266,N_2167,N_2150);
nor U2267 (N_2267,N_2032,N_2005);
and U2268 (N_2268,N_2187,N_2097);
or U2269 (N_2269,N_2067,N_2006);
xnor U2270 (N_2270,N_2036,N_2088);
nand U2271 (N_2271,N_2182,N_2186);
nor U2272 (N_2272,N_2135,N_2024);
nor U2273 (N_2273,N_2068,N_2106);
nor U2274 (N_2274,N_2132,N_2095);
nor U2275 (N_2275,N_2018,N_2016);
nor U2276 (N_2276,N_2093,N_2013);
or U2277 (N_2277,N_2107,N_2194);
nor U2278 (N_2278,N_2129,N_2195);
and U2279 (N_2279,N_2163,N_2050);
or U2280 (N_2280,N_2190,N_2193);
nor U2281 (N_2281,N_2142,N_2049);
xor U2282 (N_2282,N_2092,N_2035);
nor U2283 (N_2283,N_2159,N_2116);
nand U2284 (N_2284,N_2020,N_2028);
or U2285 (N_2285,N_2026,N_2004);
nor U2286 (N_2286,N_2191,N_2101);
nor U2287 (N_2287,N_2108,N_2166);
or U2288 (N_2288,N_2125,N_2158);
or U2289 (N_2289,N_2103,N_2141);
nand U2290 (N_2290,N_2066,N_2100);
and U2291 (N_2291,N_2062,N_2003);
and U2292 (N_2292,N_2128,N_2137);
nor U2293 (N_2293,N_2199,N_2094);
xor U2294 (N_2294,N_2111,N_2198);
or U2295 (N_2295,N_2077,N_2052);
and U2296 (N_2296,N_2037,N_2073);
nand U2297 (N_2297,N_2047,N_2176);
or U2298 (N_2298,N_2030,N_2053);
nand U2299 (N_2299,N_2118,N_2175);
nor U2300 (N_2300,N_2036,N_2057);
and U2301 (N_2301,N_2117,N_2050);
nand U2302 (N_2302,N_2121,N_2124);
or U2303 (N_2303,N_2126,N_2110);
and U2304 (N_2304,N_2049,N_2043);
or U2305 (N_2305,N_2164,N_2015);
nor U2306 (N_2306,N_2132,N_2092);
nand U2307 (N_2307,N_2018,N_2188);
or U2308 (N_2308,N_2021,N_2164);
nand U2309 (N_2309,N_2157,N_2068);
and U2310 (N_2310,N_2173,N_2140);
nor U2311 (N_2311,N_2007,N_2010);
and U2312 (N_2312,N_2152,N_2103);
nand U2313 (N_2313,N_2168,N_2159);
nor U2314 (N_2314,N_2085,N_2159);
or U2315 (N_2315,N_2166,N_2152);
nand U2316 (N_2316,N_2064,N_2138);
nor U2317 (N_2317,N_2031,N_2171);
or U2318 (N_2318,N_2122,N_2151);
or U2319 (N_2319,N_2012,N_2048);
nand U2320 (N_2320,N_2060,N_2014);
nor U2321 (N_2321,N_2125,N_2115);
nor U2322 (N_2322,N_2149,N_2031);
and U2323 (N_2323,N_2139,N_2191);
or U2324 (N_2324,N_2027,N_2142);
or U2325 (N_2325,N_2091,N_2199);
nor U2326 (N_2326,N_2008,N_2072);
nor U2327 (N_2327,N_2182,N_2058);
and U2328 (N_2328,N_2136,N_2054);
nor U2329 (N_2329,N_2136,N_2100);
and U2330 (N_2330,N_2059,N_2103);
nor U2331 (N_2331,N_2115,N_2035);
or U2332 (N_2332,N_2042,N_2156);
or U2333 (N_2333,N_2012,N_2103);
and U2334 (N_2334,N_2144,N_2140);
and U2335 (N_2335,N_2020,N_2014);
nor U2336 (N_2336,N_2133,N_2101);
and U2337 (N_2337,N_2054,N_2083);
xnor U2338 (N_2338,N_2079,N_2050);
and U2339 (N_2339,N_2031,N_2073);
nand U2340 (N_2340,N_2060,N_2124);
or U2341 (N_2341,N_2075,N_2050);
nor U2342 (N_2342,N_2032,N_2130);
or U2343 (N_2343,N_2118,N_2071);
or U2344 (N_2344,N_2104,N_2090);
nand U2345 (N_2345,N_2101,N_2131);
nor U2346 (N_2346,N_2085,N_2074);
nor U2347 (N_2347,N_2111,N_2117);
nand U2348 (N_2348,N_2145,N_2077);
or U2349 (N_2349,N_2049,N_2022);
nor U2350 (N_2350,N_2108,N_2078);
or U2351 (N_2351,N_2051,N_2109);
nor U2352 (N_2352,N_2101,N_2008);
or U2353 (N_2353,N_2045,N_2165);
nand U2354 (N_2354,N_2198,N_2010);
nand U2355 (N_2355,N_2028,N_2191);
nor U2356 (N_2356,N_2029,N_2073);
and U2357 (N_2357,N_2165,N_2177);
xnor U2358 (N_2358,N_2071,N_2078);
or U2359 (N_2359,N_2077,N_2086);
or U2360 (N_2360,N_2199,N_2092);
nor U2361 (N_2361,N_2085,N_2030);
nor U2362 (N_2362,N_2165,N_2061);
and U2363 (N_2363,N_2181,N_2021);
nor U2364 (N_2364,N_2026,N_2089);
nand U2365 (N_2365,N_2096,N_2085);
nor U2366 (N_2366,N_2037,N_2179);
xor U2367 (N_2367,N_2003,N_2193);
or U2368 (N_2368,N_2099,N_2056);
nor U2369 (N_2369,N_2042,N_2197);
xnor U2370 (N_2370,N_2074,N_2070);
or U2371 (N_2371,N_2005,N_2081);
nand U2372 (N_2372,N_2178,N_2164);
nor U2373 (N_2373,N_2038,N_2000);
nor U2374 (N_2374,N_2184,N_2010);
nor U2375 (N_2375,N_2125,N_2088);
nand U2376 (N_2376,N_2178,N_2078);
or U2377 (N_2377,N_2053,N_2046);
nor U2378 (N_2378,N_2058,N_2174);
or U2379 (N_2379,N_2044,N_2028);
and U2380 (N_2380,N_2095,N_2027);
and U2381 (N_2381,N_2066,N_2036);
or U2382 (N_2382,N_2083,N_2098);
nand U2383 (N_2383,N_2007,N_2162);
nand U2384 (N_2384,N_2126,N_2097);
and U2385 (N_2385,N_2198,N_2023);
and U2386 (N_2386,N_2034,N_2176);
and U2387 (N_2387,N_2102,N_2192);
or U2388 (N_2388,N_2064,N_2129);
nor U2389 (N_2389,N_2075,N_2154);
nand U2390 (N_2390,N_2052,N_2059);
nor U2391 (N_2391,N_2012,N_2097);
nor U2392 (N_2392,N_2022,N_2170);
xor U2393 (N_2393,N_2180,N_2167);
or U2394 (N_2394,N_2181,N_2083);
nor U2395 (N_2395,N_2184,N_2028);
nand U2396 (N_2396,N_2045,N_2162);
or U2397 (N_2397,N_2025,N_2111);
nand U2398 (N_2398,N_2052,N_2064);
and U2399 (N_2399,N_2183,N_2068);
or U2400 (N_2400,N_2285,N_2265);
or U2401 (N_2401,N_2250,N_2232);
nor U2402 (N_2402,N_2256,N_2210);
and U2403 (N_2403,N_2387,N_2398);
and U2404 (N_2404,N_2235,N_2388);
and U2405 (N_2405,N_2399,N_2268);
or U2406 (N_2406,N_2204,N_2286);
nand U2407 (N_2407,N_2230,N_2355);
xor U2408 (N_2408,N_2336,N_2375);
nand U2409 (N_2409,N_2344,N_2251);
or U2410 (N_2410,N_2284,N_2229);
nor U2411 (N_2411,N_2254,N_2221);
or U2412 (N_2412,N_2312,N_2240);
or U2413 (N_2413,N_2304,N_2224);
or U2414 (N_2414,N_2393,N_2217);
and U2415 (N_2415,N_2260,N_2363);
and U2416 (N_2416,N_2228,N_2395);
or U2417 (N_2417,N_2338,N_2319);
and U2418 (N_2418,N_2207,N_2327);
nor U2419 (N_2419,N_2323,N_2266);
xnor U2420 (N_2420,N_2314,N_2278);
nand U2421 (N_2421,N_2270,N_2328);
nor U2422 (N_2422,N_2282,N_2376);
and U2423 (N_2423,N_2258,N_2290);
nand U2424 (N_2424,N_2295,N_2369);
and U2425 (N_2425,N_2356,N_2335);
and U2426 (N_2426,N_2380,N_2236);
nor U2427 (N_2427,N_2315,N_2242);
and U2428 (N_2428,N_2340,N_2259);
xnor U2429 (N_2429,N_2365,N_2257);
and U2430 (N_2430,N_2261,N_2331);
or U2431 (N_2431,N_2384,N_2337);
nand U2432 (N_2432,N_2223,N_2354);
or U2433 (N_2433,N_2359,N_2280);
and U2434 (N_2434,N_2306,N_2377);
and U2435 (N_2435,N_2205,N_2279);
and U2436 (N_2436,N_2373,N_2238);
and U2437 (N_2437,N_2202,N_2302);
and U2438 (N_2438,N_2206,N_2283);
nand U2439 (N_2439,N_2396,N_2329);
nand U2440 (N_2440,N_2288,N_2353);
or U2441 (N_2441,N_2383,N_2267);
or U2442 (N_2442,N_2333,N_2370);
and U2443 (N_2443,N_2291,N_2303);
and U2444 (N_2444,N_2299,N_2392);
nand U2445 (N_2445,N_2200,N_2276);
or U2446 (N_2446,N_2253,N_2211);
or U2447 (N_2447,N_2362,N_2381);
nor U2448 (N_2448,N_2357,N_2339);
nor U2449 (N_2449,N_2297,N_2225);
nor U2450 (N_2450,N_2281,N_2247);
nand U2451 (N_2451,N_2390,N_2364);
nand U2452 (N_2452,N_2325,N_2255);
or U2453 (N_2453,N_2321,N_2358);
nand U2454 (N_2454,N_2378,N_2341);
and U2455 (N_2455,N_2372,N_2248);
nor U2456 (N_2456,N_2347,N_2252);
or U2457 (N_2457,N_2209,N_2226);
nand U2458 (N_2458,N_2293,N_2249);
nand U2459 (N_2459,N_2368,N_2222);
nor U2460 (N_2460,N_2241,N_2243);
nand U2461 (N_2461,N_2305,N_2214);
and U2462 (N_2462,N_2220,N_2346);
nand U2463 (N_2463,N_2345,N_2233);
or U2464 (N_2464,N_2201,N_2317);
nor U2465 (N_2465,N_2367,N_2272);
and U2466 (N_2466,N_2330,N_2213);
nand U2467 (N_2467,N_2374,N_2234);
or U2468 (N_2468,N_2382,N_2394);
xnor U2469 (N_2469,N_2227,N_2385);
nand U2470 (N_2470,N_2246,N_2318);
nand U2471 (N_2471,N_2301,N_2203);
or U2472 (N_2472,N_2273,N_2311);
nor U2473 (N_2473,N_2352,N_2215);
nor U2474 (N_2474,N_2219,N_2231);
nor U2475 (N_2475,N_2264,N_2334);
nor U2476 (N_2476,N_2391,N_2262);
or U2477 (N_2477,N_2316,N_2208);
nor U2478 (N_2478,N_2397,N_2277);
and U2479 (N_2479,N_2351,N_2307);
nor U2480 (N_2480,N_2366,N_2275);
nor U2481 (N_2481,N_2343,N_2386);
nand U2482 (N_2482,N_2292,N_2300);
nand U2483 (N_2483,N_2371,N_2310);
nor U2484 (N_2484,N_2269,N_2298);
nor U2485 (N_2485,N_2294,N_2324);
or U2486 (N_2486,N_2313,N_2245);
nor U2487 (N_2487,N_2350,N_2212);
nand U2488 (N_2488,N_2320,N_2287);
nor U2489 (N_2489,N_2263,N_2289);
or U2490 (N_2490,N_2216,N_2389);
and U2491 (N_2491,N_2361,N_2349);
and U2492 (N_2492,N_2296,N_2332);
and U2493 (N_2493,N_2322,N_2218);
nor U2494 (N_2494,N_2237,N_2244);
or U2495 (N_2495,N_2342,N_2326);
nand U2496 (N_2496,N_2271,N_2379);
or U2497 (N_2497,N_2360,N_2309);
nor U2498 (N_2498,N_2348,N_2308);
nand U2499 (N_2499,N_2239,N_2274);
nor U2500 (N_2500,N_2304,N_2247);
nand U2501 (N_2501,N_2319,N_2257);
or U2502 (N_2502,N_2388,N_2237);
xor U2503 (N_2503,N_2317,N_2343);
or U2504 (N_2504,N_2376,N_2349);
and U2505 (N_2505,N_2280,N_2333);
and U2506 (N_2506,N_2270,N_2238);
xor U2507 (N_2507,N_2359,N_2242);
or U2508 (N_2508,N_2338,N_2240);
nor U2509 (N_2509,N_2274,N_2291);
nand U2510 (N_2510,N_2348,N_2287);
and U2511 (N_2511,N_2260,N_2312);
and U2512 (N_2512,N_2286,N_2243);
nand U2513 (N_2513,N_2286,N_2255);
nand U2514 (N_2514,N_2310,N_2341);
or U2515 (N_2515,N_2345,N_2330);
and U2516 (N_2516,N_2353,N_2396);
xor U2517 (N_2517,N_2230,N_2343);
xnor U2518 (N_2518,N_2311,N_2349);
nor U2519 (N_2519,N_2321,N_2244);
or U2520 (N_2520,N_2385,N_2346);
or U2521 (N_2521,N_2276,N_2235);
nor U2522 (N_2522,N_2390,N_2328);
xor U2523 (N_2523,N_2362,N_2231);
xnor U2524 (N_2524,N_2390,N_2365);
or U2525 (N_2525,N_2209,N_2333);
or U2526 (N_2526,N_2383,N_2343);
nand U2527 (N_2527,N_2367,N_2251);
or U2528 (N_2528,N_2248,N_2395);
nand U2529 (N_2529,N_2251,N_2278);
xnor U2530 (N_2530,N_2307,N_2340);
nor U2531 (N_2531,N_2386,N_2342);
and U2532 (N_2532,N_2299,N_2317);
nor U2533 (N_2533,N_2213,N_2293);
nand U2534 (N_2534,N_2249,N_2286);
and U2535 (N_2535,N_2382,N_2305);
and U2536 (N_2536,N_2235,N_2236);
and U2537 (N_2537,N_2210,N_2292);
nand U2538 (N_2538,N_2341,N_2292);
and U2539 (N_2539,N_2320,N_2266);
or U2540 (N_2540,N_2382,N_2377);
or U2541 (N_2541,N_2304,N_2394);
xor U2542 (N_2542,N_2287,N_2235);
nand U2543 (N_2543,N_2315,N_2234);
or U2544 (N_2544,N_2281,N_2370);
or U2545 (N_2545,N_2268,N_2222);
nand U2546 (N_2546,N_2227,N_2316);
nand U2547 (N_2547,N_2281,N_2359);
and U2548 (N_2548,N_2252,N_2205);
nor U2549 (N_2549,N_2394,N_2389);
and U2550 (N_2550,N_2247,N_2287);
nand U2551 (N_2551,N_2313,N_2217);
or U2552 (N_2552,N_2208,N_2379);
nand U2553 (N_2553,N_2321,N_2240);
or U2554 (N_2554,N_2247,N_2251);
nor U2555 (N_2555,N_2366,N_2278);
or U2556 (N_2556,N_2321,N_2202);
nand U2557 (N_2557,N_2252,N_2335);
or U2558 (N_2558,N_2223,N_2226);
or U2559 (N_2559,N_2320,N_2348);
or U2560 (N_2560,N_2322,N_2389);
nor U2561 (N_2561,N_2208,N_2310);
and U2562 (N_2562,N_2263,N_2377);
nor U2563 (N_2563,N_2335,N_2201);
or U2564 (N_2564,N_2318,N_2310);
nor U2565 (N_2565,N_2283,N_2339);
or U2566 (N_2566,N_2265,N_2287);
and U2567 (N_2567,N_2339,N_2282);
and U2568 (N_2568,N_2395,N_2214);
and U2569 (N_2569,N_2208,N_2295);
nor U2570 (N_2570,N_2395,N_2385);
or U2571 (N_2571,N_2395,N_2383);
nand U2572 (N_2572,N_2281,N_2238);
nor U2573 (N_2573,N_2353,N_2319);
or U2574 (N_2574,N_2240,N_2290);
and U2575 (N_2575,N_2326,N_2265);
nor U2576 (N_2576,N_2385,N_2337);
and U2577 (N_2577,N_2245,N_2215);
or U2578 (N_2578,N_2223,N_2328);
nor U2579 (N_2579,N_2226,N_2212);
or U2580 (N_2580,N_2393,N_2273);
xor U2581 (N_2581,N_2287,N_2296);
nand U2582 (N_2582,N_2293,N_2386);
xnor U2583 (N_2583,N_2316,N_2399);
nand U2584 (N_2584,N_2306,N_2253);
or U2585 (N_2585,N_2383,N_2261);
and U2586 (N_2586,N_2227,N_2231);
and U2587 (N_2587,N_2324,N_2377);
and U2588 (N_2588,N_2396,N_2315);
and U2589 (N_2589,N_2326,N_2290);
and U2590 (N_2590,N_2215,N_2341);
and U2591 (N_2591,N_2264,N_2398);
nor U2592 (N_2592,N_2335,N_2270);
nand U2593 (N_2593,N_2201,N_2256);
nor U2594 (N_2594,N_2302,N_2286);
nand U2595 (N_2595,N_2317,N_2248);
nand U2596 (N_2596,N_2268,N_2330);
and U2597 (N_2597,N_2247,N_2313);
nand U2598 (N_2598,N_2239,N_2343);
nor U2599 (N_2599,N_2315,N_2227);
or U2600 (N_2600,N_2497,N_2511);
nand U2601 (N_2601,N_2491,N_2485);
and U2602 (N_2602,N_2577,N_2468);
and U2603 (N_2603,N_2537,N_2483);
or U2604 (N_2604,N_2569,N_2550);
and U2605 (N_2605,N_2540,N_2448);
xnor U2606 (N_2606,N_2482,N_2498);
and U2607 (N_2607,N_2514,N_2501);
or U2608 (N_2608,N_2596,N_2594);
nand U2609 (N_2609,N_2430,N_2533);
nor U2610 (N_2610,N_2456,N_2564);
xnor U2611 (N_2611,N_2422,N_2409);
xnor U2612 (N_2612,N_2476,N_2519);
nand U2613 (N_2613,N_2435,N_2432);
or U2614 (N_2614,N_2542,N_2500);
nand U2615 (N_2615,N_2428,N_2547);
or U2616 (N_2616,N_2493,N_2412);
or U2617 (N_2617,N_2565,N_2507);
nor U2618 (N_2618,N_2478,N_2591);
and U2619 (N_2619,N_2571,N_2423);
and U2620 (N_2620,N_2457,N_2568);
and U2621 (N_2621,N_2494,N_2400);
nor U2622 (N_2622,N_2469,N_2410);
or U2623 (N_2623,N_2563,N_2459);
and U2624 (N_2624,N_2477,N_2473);
nand U2625 (N_2625,N_2411,N_2525);
and U2626 (N_2626,N_2439,N_2438);
nor U2627 (N_2627,N_2492,N_2546);
and U2628 (N_2628,N_2419,N_2503);
or U2629 (N_2629,N_2513,N_2556);
nor U2630 (N_2630,N_2539,N_2445);
and U2631 (N_2631,N_2415,N_2587);
or U2632 (N_2632,N_2455,N_2532);
and U2633 (N_2633,N_2450,N_2560);
or U2634 (N_2634,N_2486,N_2461);
nor U2635 (N_2635,N_2592,N_2427);
nand U2636 (N_2636,N_2578,N_2463);
and U2637 (N_2637,N_2590,N_2488);
or U2638 (N_2638,N_2502,N_2558);
and U2639 (N_2639,N_2580,N_2443);
and U2640 (N_2640,N_2495,N_2462);
and U2641 (N_2641,N_2572,N_2480);
and U2642 (N_2642,N_2505,N_2508);
nor U2643 (N_2643,N_2417,N_2567);
nand U2644 (N_2644,N_2496,N_2487);
or U2645 (N_2645,N_2526,N_2418);
nor U2646 (N_2646,N_2466,N_2531);
nor U2647 (N_2647,N_2433,N_2545);
or U2648 (N_2648,N_2573,N_2512);
nand U2649 (N_2649,N_2566,N_2529);
nand U2650 (N_2650,N_2404,N_2579);
and U2651 (N_2651,N_2406,N_2522);
xor U2652 (N_2652,N_2451,N_2402);
nor U2653 (N_2653,N_2452,N_2447);
or U2654 (N_2654,N_2499,N_2481);
xnor U2655 (N_2655,N_2429,N_2538);
and U2656 (N_2656,N_2490,N_2517);
nand U2657 (N_2657,N_2509,N_2598);
and U2658 (N_2658,N_2504,N_2585);
xnor U2659 (N_2659,N_2437,N_2553);
and U2660 (N_2660,N_2471,N_2414);
and U2661 (N_2661,N_2520,N_2464);
nand U2662 (N_2662,N_2593,N_2555);
xnor U2663 (N_2663,N_2442,N_2407);
and U2664 (N_2664,N_2489,N_2574);
or U2665 (N_2665,N_2543,N_2589);
nor U2666 (N_2666,N_2458,N_2576);
nand U2667 (N_2667,N_2544,N_2405);
nor U2668 (N_2668,N_2584,N_2583);
nor U2669 (N_2669,N_2408,N_2424);
xnor U2670 (N_2670,N_2431,N_2582);
or U2671 (N_2671,N_2421,N_2510);
nor U2672 (N_2672,N_2425,N_2528);
nand U2673 (N_2673,N_2474,N_2470);
or U2674 (N_2674,N_2588,N_2548);
xnor U2675 (N_2675,N_2484,N_2552);
xor U2676 (N_2676,N_2527,N_2413);
nand U2677 (N_2677,N_2541,N_2465);
nor U2678 (N_2678,N_2472,N_2475);
nand U2679 (N_2679,N_2416,N_2524);
nor U2680 (N_2680,N_2454,N_2549);
nand U2681 (N_2681,N_2434,N_2403);
and U2682 (N_2682,N_2449,N_2599);
nor U2683 (N_2683,N_2516,N_2559);
nor U2684 (N_2684,N_2446,N_2595);
nand U2685 (N_2685,N_2530,N_2515);
nor U2686 (N_2686,N_2401,N_2440);
nor U2687 (N_2687,N_2441,N_2460);
xnor U2688 (N_2688,N_2436,N_2444);
or U2689 (N_2689,N_2575,N_2535);
and U2690 (N_2690,N_2479,N_2551);
and U2691 (N_2691,N_2557,N_2581);
nand U2692 (N_2692,N_2518,N_2506);
or U2693 (N_2693,N_2467,N_2586);
and U2694 (N_2694,N_2561,N_2521);
and U2695 (N_2695,N_2536,N_2534);
nand U2696 (N_2696,N_2554,N_2570);
or U2697 (N_2697,N_2597,N_2426);
nand U2698 (N_2698,N_2453,N_2420);
nor U2699 (N_2699,N_2523,N_2562);
nand U2700 (N_2700,N_2409,N_2581);
nand U2701 (N_2701,N_2440,N_2437);
nor U2702 (N_2702,N_2407,N_2457);
or U2703 (N_2703,N_2588,N_2590);
nor U2704 (N_2704,N_2490,N_2433);
or U2705 (N_2705,N_2416,N_2496);
and U2706 (N_2706,N_2569,N_2407);
and U2707 (N_2707,N_2413,N_2439);
and U2708 (N_2708,N_2462,N_2589);
or U2709 (N_2709,N_2439,N_2543);
nor U2710 (N_2710,N_2519,N_2549);
nand U2711 (N_2711,N_2497,N_2546);
nand U2712 (N_2712,N_2582,N_2473);
and U2713 (N_2713,N_2402,N_2422);
nand U2714 (N_2714,N_2421,N_2423);
or U2715 (N_2715,N_2562,N_2513);
nor U2716 (N_2716,N_2573,N_2503);
nand U2717 (N_2717,N_2480,N_2482);
and U2718 (N_2718,N_2411,N_2495);
nor U2719 (N_2719,N_2592,N_2416);
or U2720 (N_2720,N_2437,N_2456);
nand U2721 (N_2721,N_2470,N_2544);
or U2722 (N_2722,N_2577,N_2477);
or U2723 (N_2723,N_2570,N_2484);
nor U2724 (N_2724,N_2481,N_2464);
or U2725 (N_2725,N_2521,N_2484);
and U2726 (N_2726,N_2494,N_2590);
or U2727 (N_2727,N_2506,N_2404);
or U2728 (N_2728,N_2493,N_2478);
nand U2729 (N_2729,N_2594,N_2515);
nand U2730 (N_2730,N_2593,N_2474);
nor U2731 (N_2731,N_2415,N_2437);
and U2732 (N_2732,N_2591,N_2541);
nor U2733 (N_2733,N_2451,N_2404);
or U2734 (N_2734,N_2427,N_2599);
or U2735 (N_2735,N_2584,N_2423);
nor U2736 (N_2736,N_2443,N_2512);
nor U2737 (N_2737,N_2459,N_2477);
or U2738 (N_2738,N_2467,N_2536);
nor U2739 (N_2739,N_2494,N_2505);
nand U2740 (N_2740,N_2416,N_2539);
nor U2741 (N_2741,N_2595,N_2461);
xnor U2742 (N_2742,N_2482,N_2523);
nor U2743 (N_2743,N_2543,N_2524);
nor U2744 (N_2744,N_2518,N_2509);
nand U2745 (N_2745,N_2478,N_2480);
nand U2746 (N_2746,N_2500,N_2530);
nor U2747 (N_2747,N_2428,N_2484);
xnor U2748 (N_2748,N_2514,N_2530);
nor U2749 (N_2749,N_2476,N_2554);
nand U2750 (N_2750,N_2581,N_2510);
nor U2751 (N_2751,N_2464,N_2548);
or U2752 (N_2752,N_2509,N_2466);
and U2753 (N_2753,N_2443,N_2597);
or U2754 (N_2754,N_2517,N_2559);
nor U2755 (N_2755,N_2487,N_2541);
and U2756 (N_2756,N_2486,N_2562);
or U2757 (N_2757,N_2586,N_2422);
nor U2758 (N_2758,N_2564,N_2470);
nand U2759 (N_2759,N_2424,N_2452);
xnor U2760 (N_2760,N_2593,N_2539);
and U2761 (N_2761,N_2561,N_2574);
and U2762 (N_2762,N_2433,N_2437);
nand U2763 (N_2763,N_2410,N_2412);
nand U2764 (N_2764,N_2590,N_2564);
nor U2765 (N_2765,N_2503,N_2597);
and U2766 (N_2766,N_2448,N_2405);
and U2767 (N_2767,N_2533,N_2545);
or U2768 (N_2768,N_2428,N_2470);
nor U2769 (N_2769,N_2589,N_2424);
and U2770 (N_2770,N_2596,N_2499);
nand U2771 (N_2771,N_2435,N_2497);
nand U2772 (N_2772,N_2593,N_2499);
nand U2773 (N_2773,N_2484,N_2456);
nand U2774 (N_2774,N_2577,N_2418);
or U2775 (N_2775,N_2579,N_2492);
nand U2776 (N_2776,N_2467,N_2415);
or U2777 (N_2777,N_2574,N_2460);
nand U2778 (N_2778,N_2428,N_2425);
xor U2779 (N_2779,N_2544,N_2513);
and U2780 (N_2780,N_2406,N_2441);
nor U2781 (N_2781,N_2455,N_2420);
or U2782 (N_2782,N_2530,N_2424);
or U2783 (N_2783,N_2406,N_2567);
xnor U2784 (N_2784,N_2449,N_2424);
or U2785 (N_2785,N_2443,N_2538);
xnor U2786 (N_2786,N_2535,N_2568);
nor U2787 (N_2787,N_2469,N_2408);
xnor U2788 (N_2788,N_2565,N_2504);
and U2789 (N_2789,N_2578,N_2429);
nand U2790 (N_2790,N_2422,N_2427);
nor U2791 (N_2791,N_2489,N_2422);
or U2792 (N_2792,N_2596,N_2538);
nor U2793 (N_2793,N_2489,N_2459);
nor U2794 (N_2794,N_2539,N_2492);
nor U2795 (N_2795,N_2421,N_2430);
and U2796 (N_2796,N_2468,N_2490);
or U2797 (N_2797,N_2444,N_2549);
nand U2798 (N_2798,N_2530,N_2471);
nand U2799 (N_2799,N_2437,N_2509);
and U2800 (N_2800,N_2662,N_2795);
nor U2801 (N_2801,N_2734,N_2780);
nor U2802 (N_2802,N_2764,N_2718);
xnor U2803 (N_2803,N_2770,N_2774);
xnor U2804 (N_2804,N_2763,N_2619);
xor U2805 (N_2805,N_2723,N_2679);
nor U2806 (N_2806,N_2768,N_2700);
and U2807 (N_2807,N_2776,N_2706);
nor U2808 (N_2808,N_2750,N_2670);
xnor U2809 (N_2809,N_2740,N_2671);
or U2810 (N_2810,N_2663,N_2625);
or U2811 (N_2811,N_2736,N_2738);
nor U2812 (N_2812,N_2789,N_2784);
and U2813 (N_2813,N_2730,N_2712);
nand U2814 (N_2814,N_2707,N_2720);
nand U2815 (N_2815,N_2646,N_2741);
and U2816 (N_2816,N_2635,N_2749);
nor U2817 (N_2817,N_2782,N_2705);
or U2818 (N_2818,N_2628,N_2636);
nor U2819 (N_2819,N_2796,N_2673);
nand U2820 (N_2820,N_2649,N_2745);
or U2821 (N_2821,N_2665,N_2719);
nor U2822 (N_2822,N_2632,N_2684);
nor U2823 (N_2823,N_2703,N_2772);
nor U2824 (N_2824,N_2653,N_2659);
nand U2825 (N_2825,N_2666,N_2760);
or U2826 (N_2826,N_2658,N_2611);
nor U2827 (N_2827,N_2794,N_2739);
nor U2828 (N_2828,N_2689,N_2716);
and U2829 (N_2829,N_2695,N_2629);
nand U2830 (N_2830,N_2651,N_2733);
nand U2831 (N_2831,N_2773,N_2685);
and U2832 (N_2832,N_2688,N_2744);
or U2833 (N_2833,N_2645,N_2687);
and U2834 (N_2834,N_2603,N_2761);
nand U2835 (N_2835,N_2779,N_2609);
xor U2836 (N_2836,N_2708,N_2728);
and U2837 (N_2837,N_2714,N_2721);
xor U2838 (N_2838,N_2711,N_2631);
and U2839 (N_2839,N_2607,N_2614);
nor U2840 (N_2840,N_2704,N_2648);
nor U2841 (N_2841,N_2752,N_2790);
nand U2842 (N_2842,N_2642,N_2786);
or U2843 (N_2843,N_2735,N_2647);
and U2844 (N_2844,N_2604,N_2726);
or U2845 (N_2845,N_2674,N_2605);
nand U2846 (N_2846,N_2690,N_2668);
or U2847 (N_2847,N_2743,N_2681);
nand U2848 (N_2848,N_2664,N_2634);
xor U2849 (N_2849,N_2667,N_2701);
nor U2850 (N_2850,N_2637,N_2722);
or U2851 (N_2851,N_2675,N_2618);
xor U2852 (N_2852,N_2610,N_2765);
xnor U2853 (N_2853,N_2657,N_2612);
or U2854 (N_2854,N_2638,N_2613);
nand U2855 (N_2855,N_2630,N_2686);
and U2856 (N_2856,N_2669,N_2787);
and U2857 (N_2857,N_2747,N_2702);
nor U2858 (N_2858,N_2680,N_2798);
and U2859 (N_2859,N_2742,N_2724);
or U2860 (N_2860,N_2650,N_2792);
nand U2861 (N_2861,N_2771,N_2732);
or U2862 (N_2862,N_2754,N_2633);
nor U2863 (N_2863,N_2672,N_2793);
nand U2864 (N_2864,N_2602,N_2682);
nand U2865 (N_2865,N_2621,N_2640);
or U2866 (N_2866,N_2626,N_2709);
nand U2867 (N_2867,N_2710,N_2783);
or U2868 (N_2868,N_2755,N_2600);
nor U2869 (N_2869,N_2620,N_2693);
nor U2870 (N_2870,N_2616,N_2775);
nor U2871 (N_2871,N_2698,N_2762);
nand U2872 (N_2872,N_2757,N_2655);
or U2873 (N_2873,N_2641,N_2753);
xor U2874 (N_2874,N_2746,N_2785);
nand U2875 (N_2875,N_2643,N_2727);
and U2876 (N_2876,N_2627,N_2644);
or U2877 (N_2877,N_2729,N_2756);
nor U2878 (N_2878,N_2766,N_2715);
nand U2879 (N_2879,N_2737,N_2725);
nor U2880 (N_2880,N_2694,N_2606);
nand U2881 (N_2881,N_2781,N_2797);
or U2882 (N_2882,N_2692,N_2791);
nand U2883 (N_2883,N_2623,N_2691);
nand U2884 (N_2884,N_2608,N_2624);
xnor U2885 (N_2885,N_2717,N_2713);
and U2886 (N_2886,N_2759,N_2799);
or U2887 (N_2887,N_2617,N_2788);
or U2888 (N_2888,N_2601,N_2777);
and U2889 (N_2889,N_2661,N_2731);
nand U2890 (N_2890,N_2769,N_2748);
or U2891 (N_2891,N_2751,N_2699);
or U2892 (N_2892,N_2697,N_2677);
or U2893 (N_2893,N_2639,N_2678);
and U2894 (N_2894,N_2622,N_2696);
nand U2895 (N_2895,N_2615,N_2778);
nor U2896 (N_2896,N_2767,N_2676);
or U2897 (N_2897,N_2654,N_2660);
nand U2898 (N_2898,N_2758,N_2652);
nand U2899 (N_2899,N_2656,N_2683);
xor U2900 (N_2900,N_2672,N_2609);
and U2901 (N_2901,N_2711,N_2621);
xnor U2902 (N_2902,N_2760,N_2744);
nor U2903 (N_2903,N_2626,N_2700);
or U2904 (N_2904,N_2620,N_2617);
nand U2905 (N_2905,N_2628,N_2646);
and U2906 (N_2906,N_2670,N_2614);
or U2907 (N_2907,N_2624,N_2720);
xnor U2908 (N_2908,N_2653,N_2649);
or U2909 (N_2909,N_2606,N_2714);
and U2910 (N_2910,N_2664,N_2655);
nand U2911 (N_2911,N_2709,N_2722);
or U2912 (N_2912,N_2602,N_2612);
xor U2913 (N_2913,N_2682,N_2768);
and U2914 (N_2914,N_2798,N_2694);
and U2915 (N_2915,N_2781,N_2710);
nand U2916 (N_2916,N_2623,N_2705);
nor U2917 (N_2917,N_2669,N_2788);
xor U2918 (N_2918,N_2671,N_2684);
nand U2919 (N_2919,N_2687,N_2774);
or U2920 (N_2920,N_2704,N_2757);
nand U2921 (N_2921,N_2678,N_2785);
nor U2922 (N_2922,N_2727,N_2773);
and U2923 (N_2923,N_2632,N_2674);
and U2924 (N_2924,N_2707,N_2751);
nor U2925 (N_2925,N_2797,N_2746);
nor U2926 (N_2926,N_2766,N_2746);
or U2927 (N_2927,N_2718,N_2747);
nor U2928 (N_2928,N_2684,N_2613);
xor U2929 (N_2929,N_2602,N_2760);
or U2930 (N_2930,N_2760,N_2634);
or U2931 (N_2931,N_2674,N_2683);
nand U2932 (N_2932,N_2618,N_2652);
nor U2933 (N_2933,N_2797,N_2639);
nor U2934 (N_2934,N_2752,N_2649);
nand U2935 (N_2935,N_2717,N_2638);
nand U2936 (N_2936,N_2632,N_2623);
and U2937 (N_2937,N_2672,N_2687);
or U2938 (N_2938,N_2720,N_2611);
nor U2939 (N_2939,N_2779,N_2626);
nand U2940 (N_2940,N_2776,N_2763);
or U2941 (N_2941,N_2666,N_2606);
nor U2942 (N_2942,N_2746,N_2640);
nor U2943 (N_2943,N_2669,N_2713);
or U2944 (N_2944,N_2760,N_2756);
and U2945 (N_2945,N_2725,N_2775);
nor U2946 (N_2946,N_2753,N_2741);
nor U2947 (N_2947,N_2753,N_2798);
nand U2948 (N_2948,N_2626,N_2762);
nand U2949 (N_2949,N_2626,N_2620);
and U2950 (N_2950,N_2648,N_2768);
nor U2951 (N_2951,N_2709,N_2607);
or U2952 (N_2952,N_2726,N_2736);
nor U2953 (N_2953,N_2693,N_2713);
or U2954 (N_2954,N_2747,N_2776);
nand U2955 (N_2955,N_2742,N_2797);
or U2956 (N_2956,N_2750,N_2634);
and U2957 (N_2957,N_2605,N_2677);
nand U2958 (N_2958,N_2783,N_2630);
or U2959 (N_2959,N_2660,N_2748);
and U2960 (N_2960,N_2625,N_2708);
nand U2961 (N_2961,N_2734,N_2669);
nor U2962 (N_2962,N_2750,N_2793);
nor U2963 (N_2963,N_2718,N_2615);
or U2964 (N_2964,N_2690,N_2691);
nor U2965 (N_2965,N_2760,N_2699);
nand U2966 (N_2966,N_2707,N_2736);
nor U2967 (N_2967,N_2745,N_2708);
xnor U2968 (N_2968,N_2681,N_2703);
nand U2969 (N_2969,N_2694,N_2635);
and U2970 (N_2970,N_2614,N_2745);
and U2971 (N_2971,N_2668,N_2737);
nand U2972 (N_2972,N_2676,N_2758);
nor U2973 (N_2973,N_2711,N_2756);
and U2974 (N_2974,N_2717,N_2610);
nor U2975 (N_2975,N_2618,N_2771);
nor U2976 (N_2976,N_2784,N_2705);
nor U2977 (N_2977,N_2614,N_2715);
and U2978 (N_2978,N_2660,N_2799);
or U2979 (N_2979,N_2689,N_2744);
and U2980 (N_2980,N_2731,N_2663);
nor U2981 (N_2981,N_2705,N_2664);
and U2982 (N_2982,N_2637,N_2648);
nor U2983 (N_2983,N_2719,N_2768);
nor U2984 (N_2984,N_2783,N_2627);
xor U2985 (N_2985,N_2704,N_2612);
and U2986 (N_2986,N_2662,N_2733);
xor U2987 (N_2987,N_2717,N_2670);
and U2988 (N_2988,N_2785,N_2734);
nor U2989 (N_2989,N_2788,N_2779);
and U2990 (N_2990,N_2669,N_2785);
and U2991 (N_2991,N_2611,N_2790);
or U2992 (N_2992,N_2754,N_2650);
nor U2993 (N_2993,N_2639,N_2738);
and U2994 (N_2994,N_2734,N_2640);
or U2995 (N_2995,N_2683,N_2757);
and U2996 (N_2996,N_2772,N_2625);
nand U2997 (N_2997,N_2799,N_2720);
nor U2998 (N_2998,N_2646,N_2642);
nand U2999 (N_2999,N_2678,N_2645);
and U3000 (N_3000,N_2964,N_2910);
or U3001 (N_3001,N_2870,N_2831);
or U3002 (N_3002,N_2935,N_2872);
or U3003 (N_3003,N_2985,N_2943);
and U3004 (N_3004,N_2928,N_2864);
or U3005 (N_3005,N_2900,N_2820);
and U3006 (N_3006,N_2933,N_2884);
and U3007 (N_3007,N_2833,N_2902);
or U3008 (N_3008,N_2832,N_2856);
and U3009 (N_3009,N_2874,N_2887);
or U3010 (N_3010,N_2978,N_2813);
nand U3011 (N_3011,N_2814,N_2807);
nor U3012 (N_3012,N_2913,N_2901);
xnor U3013 (N_3013,N_2802,N_2827);
nor U3014 (N_3014,N_2921,N_2843);
and U3015 (N_3015,N_2898,N_2944);
nand U3016 (N_3016,N_2818,N_2883);
xnor U3017 (N_3017,N_2896,N_2936);
nor U3018 (N_3018,N_2917,N_2909);
nand U3019 (N_3019,N_2982,N_2924);
nor U3020 (N_3020,N_2894,N_2811);
xnor U3021 (N_3021,N_2834,N_2871);
nand U3022 (N_3022,N_2946,N_2812);
nor U3023 (N_3023,N_2972,N_2919);
or U3024 (N_3024,N_2889,N_2920);
nor U3025 (N_3025,N_2800,N_2912);
and U3026 (N_3026,N_2992,N_2925);
or U3027 (N_3027,N_2848,N_2923);
and U3028 (N_3028,N_2860,N_2930);
nand U3029 (N_3029,N_2955,N_2824);
or U3030 (N_3030,N_2809,N_2828);
nand U3031 (N_3031,N_2801,N_2959);
or U3032 (N_3032,N_2806,N_2966);
nand U3033 (N_3033,N_2922,N_2888);
or U3034 (N_3034,N_2890,N_2817);
nor U3035 (N_3035,N_2951,N_2918);
or U3036 (N_3036,N_2869,N_2904);
and U3037 (N_3037,N_2983,N_2839);
and U3038 (N_3038,N_2968,N_2855);
and U3039 (N_3039,N_2999,N_2875);
nor U3040 (N_3040,N_2974,N_2970);
nand U3041 (N_3041,N_2932,N_2850);
nand U3042 (N_3042,N_2892,N_2859);
or U3043 (N_3043,N_2808,N_2975);
and U3044 (N_3044,N_2963,N_2987);
or U3045 (N_3045,N_2937,N_2979);
or U3046 (N_3046,N_2914,N_2857);
xor U3047 (N_3047,N_2816,N_2981);
or U3048 (N_3048,N_2853,N_2819);
xor U3049 (N_3049,N_2891,N_2996);
nand U3050 (N_3050,N_2838,N_2886);
nand U3051 (N_3051,N_2907,N_2929);
xnor U3052 (N_3052,N_2845,N_2822);
nand U3053 (N_3053,N_2976,N_2858);
nor U3054 (N_3054,N_2849,N_2852);
and U3055 (N_3055,N_2967,N_2885);
or U3056 (N_3056,N_2837,N_2803);
nor U3057 (N_3057,N_2962,N_2863);
nand U3058 (N_3058,N_2995,N_2815);
xnor U3059 (N_3059,N_2997,N_2844);
or U3060 (N_3060,N_2942,N_2941);
and U3061 (N_3061,N_2908,N_2973);
nand U3062 (N_3062,N_2956,N_2957);
xor U3063 (N_3063,N_2940,N_2906);
and U3064 (N_3064,N_2897,N_2911);
nand U3065 (N_3065,N_2876,N_2846);
nor U3066 (N_3066,N_2950,N_2841);
nor U3067 (N_3067,N_2882,N_2879);
or U3068 (N_3068,N_2988,N_2998);
or U3069 (N_3069,N_2927,N_2905);
nand U3070 (N_3070,N_2993,N_2939);
or U3071 (N_3071,N_2862,N_2977);
nor U3072 (N_3072,N_2804,N_2934);
and U3073 (N_3073,N_2868,N_2825);
and U3074 (N_3074,N_2893,N_2805);
nor U3075 (N_3075,N_2984,N_2835);
nand U3076 (N_3076,N_2826,N_2949);
nor U3077 (N_3077,N_2865,N_2990);
nand U3078 (N_3078,N_2873,N_2961);
and U3079 (N_3079,N_2854,N_2960);
and U3080 (N_3080,N_2810,N_2836);
nor U3081 (N_3081,N_2878,N_2842);
and U3082 (N_3082,N_2880,N_2899);
nor U3083 (N_3083,N_2948,N_2823);
nor U3084 (N_3084,N_2965,N_2958);
and U3085 (N_3085,N_2952,N_2969);
xnor U3086 (N_3086,N_2840,N_2986);
nand U3087 (N_3087,N_2954,N_2980);
nor U3088 (N_3088,N_2947,N_2877);
and U3089 (N_3089,N_2821,N_2945);
nor U3090 (N_3090,N_2847,N_2866);
nand U3091 (N_3091,N_2991,N_2903);
or U3092 (N_3092,N_2926,N_2989);
and U3093 (N_3093,N_2953,N_2938);
and U3094 (N_3094,N_2915,N_2994);
nand U3095 (N_3095,N_2851,N_2971);
or U3096 (N_3096,N_2931,N_2829);
xnor U3097 (N_3097,N_2881,N_2830);
and U3098 (N_3098,N_2861,N_2916);
and U3099 (N_3099,N_2895,N_2867);
nand U3100 (N_3100,N_2952,N_2844);
or U3101 (N_3101,N_2846,N_2834);
xor U3102 (N_3102,N_2995,N_2989);
or U3103 (N_3103,N_2825,N_2929);
or U3104 (N_3104,N_2905,N_2959);
or U3105 (N_3105,N_2997,N_2912);
nor U3106 (N_3106,N_2860,N_2802);
or U3107 (N_3107,N_2856,N_2926);
nor U3108 (N_3108,N_2866,N_2815);
nor U3109 (N_3109,N_2871,N_2821);
nand U3110 (N_3110,N_2957,N_2909);
or U3111 (N_3111,N_2857,N_2808);
and U3112 (N_3112,N_2946,N_2853);
or U3113 (N_3113,N_2858,N_2841);
xnor U3114 (N_3114,N_2818,N_2933);
or U3115 (N_3115,N_2937,N_2831);
or U3116 (N_3116,N_2951,N_2978);
nor U3117 (N_3117,N_2910,N_2869);
and U3118 (N_3118,N_2861,N_2842);
nor U3119 (N_3119,N_2901,N_2938);
and U3120 (N_3120,N_2954,N_2938);
and U3121 (N_3121,N_2947,N_2975);
and U3122 (N_3122,N_2853,N_2846);
or U3123 (N_3123,N_2864,N_2902);
xor U3124 (N_3124,N_2928,N_2950);
nand U3125 (N_3125,N_2942,N_2939);
and U3126 (N_3126,N_2929,N_2977);
xnor U3127 (N_3127,N_2838,N_2896);
nor U3128 (N_3128,N_2827,N_2989);
nor U3129 (N_3129,N_2862,N_2922);
nor U3130 (N_3130,N_2837,N_2938);
and U3131 (N_3131,N_2975,N_2809);
nand U3132 (N_3132,N_2858,N_2868);
nor U3133 (N_3133,N_2905,N_2944);
nor U3134 (N_3134,N_2900,N_2897);
xor U3135 (N_3135,N_2936,N_2962);
nor U3136 (N_3136,N_2864,N_2878);
nand U3137 (N_3137,N_2936,N_2865);
nor U3138 (N_3138,N_2926,N_2964);
and U3139 (N_3139,N_2964,N_2990);
nor U3140 (N_3140,N_2863,N_2922);
nand U3141 (N_3141,N_2872,N_2930);
and U3142 (N_3142,N_2938,N_2865);
and U3143 (N_3143,N_2980,N_2978);
and U3144 (N_3144,N_2879,N_2885);
or U3145 (N_3145,N_2878,N_2973);
xnor U3146 (N_3146,N_2881,N_2989);
or U3147 (N_3147,N_2973,N_2923);
or U3148 (N_3148,N_2915,N_2883);
or U3149 (N_3149,N_2830,N_2919);
or U3150 (N_3150,N_2937,N_2982);
or U3151 (N_3151,N_2840,N_2837);
xnor U3152 (N_3152,N_2867,N_2955);
xor U3153 (N_3153,N_2968,N_2884);
or U3154 (N_3154,N_2915,N_2932);
nor U3155 (N_3155,N_2826,N_2824);
or U3156 (N_3156,N_2886,N_2929);
nor U3157 (N_3157,N_2955,N_2890);
nand U3158 (N_3158,N_2999,N_2842);
nor U3159 (N_3159,N_2843,N_2855);
and U3160 (N_3160,N_2953,N_2991);
or U3161 (N_3161,N_2991,N_2845);
nor U3162 (N_3162,N_2965,N_2811);
nor U3163 (N_3163,N_2877,N_2900);
and U3164 (N_3164,N_2978,N_2846);
nand U3165 (N_3165,N_2945,N_2909);
nand U3166 (N_3166,N_2833,N_2960);
and U3167 (N_3167,N_2817,N_2865);
nor U3168 (N_3168,N_2907,N_2973);
nand U3169 (N_3169,N_2964,N_2941);
nor U3170 (N_3170,N_2838,N_2812);
nand U3171 (N_3171,N_2817,N_2870);
and U3172 (N_3172,N_2843,N_2840);
xor U3173 (N_3173,N_2958,N_2862);
nand U3174 (N_3174,N_2801,N_2806);
nor U3175 (N_3175,N_2995,N_2878);
nand U3176 (N_3176,N_2812,N_2912);
or U3177 (N_3177,N_2889,N_2888);
or U3178 (N_3178,N_2967,N_2983);
and U3179 (N_3179,N_2925,N_2818);
nand U3180 (N_3180,N_2887,N_2968);
nor U3181 (N_3181,N_2971,N_2964);
or U3182 (N_3182,N_2864,N_2806);
or U3183 (N_3183,N_2811,N_2958);
nand U3184 (N_3184,N_2929,N_2949);
or U3185 (N_3185,N_2922,N_2986);
nand U3186 (N_3186,N_2958,N_2810);
nor U3187 (N_3187,N_2999,N_2869);
and U3188 (N_3188,N_2971,N_2993);
xor U3189 (N_3189,N_2967,N_2970);
and U3190 (N_3190,N_2924,N_2809);
nor U3191 (N_3191,N_2929,N_2931);
or U3192 (N_3192,N_2844,N_2931);
xor U3193 (N_3193,N_2871,N_2829);
nor U3194 (N_3194,N_2954,N_2959);
or U3195 (N_3195,N_2955,N_2938);
nor U3196 (N_3196,N_2862,N_2845);
or U3197 (N_3197,N_2988,N_2848);
nand U3198 (N_3198,N_2886,N_2979);
nand U3199 (N_3199,N_2922,N_2874);
and U3200 (N_3200,N_3056,N_3104);
nor U3201 (N_3201,N_3123,N_3121);
and U3202 (N_3202,N_3054,N_3167);
or U3203 (N_3203,N_3144,N_3185);
and U3204 (N_3204,N_3136,N_3083);
and U3205 (N_3205,N_3173,N_3078);
nor U3206 (N_3206,N_3036,N_3149);
or U3207 (N_3207,N_3087,N_3178);
and U3208 (N_3208,N_3009,N_3132);
or U3209 (N_3209,N_3041,N_3175);
nor U3210 (N_3210,N_3014,N_3088);
and U3211 (N_3211,N_3131,N_3118);
or U3212 (N_3212,N_3119,N_3115);
and U3213 (N_3213,N_3195,N_3057);
and U3214 (N_3214,N_3172,N_3011);
or U3215 (N_3215,N_3184,N_3092);
and U3216 (N_3216,N_3034,N_3042);
and U3217 (N_3217,N_3147,N_3063);
or U3218 (N_3218,N_3027,N_3122);
nor U3219 (N_3219,N_3045,N_3183);
and U3220 (N_3220,N_3151,N_3148);
or U3221 (N_3221,N_3055,N_3081);
and U3222 (N_3222,N_3107,N_3006);
xor U3223 (N_3223,N_3152,N_3128);
nand U3224 (N_3224,N_3052,N_3058);
nand U3225 (N_3225,N_3007,N_3032);
nor U3226 (N_3226,N_3040,N_3164);
nor U3227 (N_3227,N_3150,N_3133);
and U3228 (N_3228,N_3134,N_3158);
xor U3229 (N_3229,N_3146,N_3061);
and U3230 (N_3230,N_3156,N_3116);
nor U3231 (N_3231,N_3125,N_3129);
nor U3232 (N_3232,N_3103,N_3157);
or U3233 (N_3233,N_3168,N_3143);
or U3234 (N_3234,N_3112,N_3190);
or U3235 (N_3235,N_3002,N_3169);
nor U3236 (N_3236,N_3111,N_3139);
or U3237 (N_3237,N_3074,N_3145);
and U3238 (N_3238,N_3171,N_3000);
nand U3239 (N_3239,N_3059,N_3199);
or U3240 (N_3240,N_3015,N_3044);
nor U3241 (N_3241,N_3181,N_3065);
and U3242 (N_3242,N_3155,N_3165);
nand U3243 (N_3243,N_3094,N_3091);
nand U3244 (N_3244,N_3194,N_3035);
nand U3245 (N_3245,N_3174,N_3018);
nor U3246 (N_3246,N_3033,N_3100);
or U3247 (N_3247,N_3076,N_3024);
nand U3248 (N_3248,N_3079,N_3093);
nor U3249 (N_3249,N_3159,N_3005);
nand U3250 (N_3250,N_3126,N_3085);
nand U3251 (N_3251,N_3140,N_3026);
nor U3252 (N_3252,N_3071,N_3016);
nand U3253 (N_3253,N_3180,N_3182);
nor U3254 (N_3254,N_3021,N_3137);
nor U3255 (N_3255,N_3001,N_3120);
nor U3256 (N_3256,N_3077,N_3017);
xor U3257 (N_3257,N_3177,N_3070);
and U3258 (N_3258,N_3113,N_3028);
and U3259 (N_3259,N_3046,N_3072);
nand U3260 (N_3260,N_3019,N_3010);
nand U3261 (N_3261,N_3130,N_3060);
nand U3262 (N_3262,N_3187,N_3067);
nand U3263 (N_3263,N_3099,N_3142);
nand U3264 (N_3264,N_3038,N_3127);
nor U3265 (N_3265,N_3191,N_3189);
nand U3266 (N_3266,N_3110,N_3080);
nor U3267 (N_3267,N_3023,N_3012);
nand U3268 (N_3268,N_3029,N_3008);
and U3269 (N_3269,N_3114,N_3188);
nor U3270 (N_3270,N_3163,N_3098);
or U3271 (N_3271,N_3153,N_3004);
nand U3272 (N_3272,N_3161,N_3197);
nand U3273 (N_3273,N_3117,N_3095);
or U3274 (N_3274,N_3086,N_3073);
and U3275 (N_3275,N_3141,N_3020);
or U3276 (N_3276,N_3047,N_3037);
nand U3277 (N_3277,N_3043,N_3138);
or U3278 (N_3278,N_3075,N_3108);
and U3279 (N_3279,N_3179,N_3160);
and U3280 (N_3280,N_3124,N_3089);
or U3281 (N_3281,N_3053,N_3048);
nand U3282 (N_3282,N_3170,N_3062);
and U3283 (N_3283,N_3186,N_3051);
or U3284 (N_3284,N_3049,N_3102);
nand U3285 (N_3285,N_3166,N_3025);
and U3286 (N_3286,N_3003,N_3106);
nor U3287 (N_3287,N_3198,N_3030);
nand U3288 (N_3288,N_3154,N_3135);
xor U3289 (N_3289,N_3039,N_3176);
nand U3290 (N_3290,N_3090,N_3196);
and U3291 (N_3291,N_3066,N_3082);
nand U3292 (N_3292,N_3109,N_3069);
and U3293 (N_3293,N_3050,N_3097);
nor U3294 (N_3294,N_3105,N_3162);
nor U3295 (N_3295,N_3064,N_3096);
nand U3296 (N_3296,N_3193,N_3022);
xor U3297 (N_3297,N_3013,N_3101);
or U3298 (N_3298,N_3068,N_3031);
and U3299 (N_3299,N_3084,N_3192);
nand U3300 (N_3300,N_3098,N_3006);
or U3301 (N_3301,N_3079,N_3145);
xnor U3302 (N_3302,N_3045,N_3199);
nor U3303 (N_3303,N_3181,N_3075);
nor U3304 (N_3304,N_3154,N_3067);
or U3305 (N_3305,N_3176,N_3130);
nand U3306 (N_3306,N_3107,N_3153);
xnor U3307 (N_3307,N_3019,N_3143);
and U3308 (N_3308,N_3079,N_3187);
and U3309 (N_3309,N_3184,N_3089);
nand U3310 (N_3310,N_3060,N_3076);
or U3311 (N_3311,N_3119,N_3030);
nor U3312 (N_3312,N_3025,N_3124);
and U3313 (N_3313,N_3115,N_3053);
or U3314 (N_3314,N_3008,N_3039);
or U3315 (N_3315,N_3082,N_3142);
nand U3316 (N_3316,N_3020,N_3156);
nand U3317 (N_3317,N_3127,N_3050);
nor U3318 (N_3318,N_3144,N_3081);
and U3319 (N_3319,N_3028,N_3064);
nor U3320 (N_3320,N_3061,N_3005);
or U3321 (N_3321,N_3012,N_3053);
nor U3322 (N_3322,N_3172,N_3087);
and U3323 (N_3323,N_3104,N_3154);
nor U3324 (N_3324,N_3070,N_3105);
and U3325 (N_3325,N_3090,N_3050);
xnor U3326 (N_3326,N_3009,N_3030);
nand U3327 (N_3327,N_3197,N_3131);
or U3328 (N_3328,N_3133,N_3154);
or U3329 (N_3329,N_3150,N_3176);
nor U3330 (N_3330,N_3146,N_3155);
nor U3331 (N_3331,N_3033,N_3133);
nor U3332 (N_3332,N_3104,N_3127);
or U3333 (N_3333,N_3019,N_3187);
nor U3334 (N_3334,N_3097,N_3183);
nand U3335 (N_3335,N_3009,N_3096);
or U3336 (N_3336,N_3172,N_3196);
and U3337 (N_3337,N_3025,N_3072);
or U3338 (N_3338,N_3099,N_3115);
nor U3339 (N_3339,N_3055,N_3097);
xor U3340 (N_3340,N_3152,N_3182);
or U3341 (N_3341,N_3004,N_3019);
nor U3342 (N_3342,N_3151,N_3014);
or U3343 (N_3343,N_3118,N_3198);
nor U3344 (N_3344,N_3068,N_3021);
xnor U3345 (N_3345,N_3131,N_3033);
nand U3346 (N_3346,N_3020,N_3029);
or U3347 (N_3347,N_3100,N_3110);
nor U3348 (N_3348,N_3126,N_3014);
or U3349 (N_3349,N_3155,N_3086);
xnor U3350 (N_3350,N_3184,N_3052);
nor U3351 (N_3351,N_3052,N_3063);
nand U3352 (N_3352,N_3189,N_3180);
nor U3353 (N_3353,N_3027,N_3102);
and U3354 (N_3354,N_3085,N_3154);
and U3355 (N_3355,N_3145,N_3054);
nor U3356 (N_3356,N_3160,N_3155);
or U3357 (N_3357,N_3187,N_3005);
or U3358 (N_3358,N_3170,N_3012);
nor U3359 (N_3359,N_3087,N_3095);
nor U3360 (N_3360,N_3145,N_3051);
or U3361 (N_3361,N_3001,N_3081);
nand U3362 (N_3362,N_3164,N_3123);
nor U3363 (N_3363,N_3120,N_3116);
nand U3364 (N_3364,N_3172,N_3134);
nor U3365 (N_3365,N_3097,N_3193);
nor U3366 (N_3366,N_3061,N_3041);
or U3367 (N_3367,N_3161,N_3003);
xnor U3368 (N_3368,N_3040,N_3060);
xnor U3369 (N_3369,N_3076,N_3192);
nand U3370 (N_3370,N_3122,N_3006);
nand U3371 (N_3371,N_3145,N_3089);
and U3372 (N_3372,N_3153,N_3119);
and U3373 (N_3373,N_3191,N_3152);
nor U3374 (N_3374,N_3010,N_3182);
xor U3375 (N_3375,N_3146,N_3181);
xor U3376 (N_3376,N_3118,N_3061);
nand U3377 (N_3377,N_3079,N_3056);
xor U3378 (N_3378,N_3023,N_3110);
nand U3379 (N_3379,N_3038,N_3034);
or U3380 (N_3380,N_3024,N_3060);
nand U3381 (N_3381,N_3158,N_3088);
nand U3382 (N_3382,N_3134,N_3042);
and U3383 (N_3383,N_3147,N_3188);
or U3384 (N_3384,N_3170,N_3114);
nor U3385 (N_3385,N_3047,N_3192);
nor U3386 (N_3386,N_3190,N_3138);
or U3387 (N_3387,N_3036,N_3037);
or U3388 (N_3388,N_3157,N_3193);
or U3389 (N_3389,N_3069,N_3197);
nor U3390 (N_3390,N_3135,N_3191);
nor U3391 (N_3391,N_3095,N_3162);
or U3392 (N_3392,N_3195,N_3160);
or U3393 (N_3393,N_3153,N_3089);
nand U3394 (N_3394,N_3028,N_3196);
xnor U3395 (N_3395,N_3180,N_3173);
and U3396 (N_3396,N_3136,N_3182);
nand U3397 (N_3397,N_3133,N_3071);
nor U3398 (N_3398,N_3193,N_3152);
xnor U3399 (N_3399,N_3151,N_3152);
and U3400 (N_3400,N_3293,N_3224);
nand U3401 (N_3401,N_3313,N_3264);
and U3402 (N_3402,N_3228,N_3253);
nand U3403 (N_3403,N_3237,N_3341);
nand U3404 (N_3404,N_3235,N_3304);
nor U3405 (N_3405,N_3379,N_3392);
and U3406 (N_3406,N_3236,N_3306);
nand U3407 (N_3407,N_3377,N_3305);
xor U3408 (N_3408,N_3338,N_3321);
or U3409 (N_3409,N_3381,N_3345);
nor U3410 (N_3410,N_3245,N_3204);
xor U3411 (N_3411,N_3335,N_3353);
nor U3412 (N_3412,N_3337,N_3243);
nor U3413 (N_3413,N_3382,N_3233);
nand U3414 (N_3414,N_3297,N_3387);
nor U3415 (N_3415,N_3217,N_3358);
or U3416 (N_3416,N_3346,N_3391);
or U3417 (N_3417,N_3368,N_3316);
and U3418 (N_3418,N_3267,N_3234);
or U3419 (N_3419,N_3229,N_3397);
nor U3420 (N_3420,N_3311,N_3324);
and U3421 (N_3421,N_3290,N_3209);
and U3422 (N_3422,N_3373,N_3295);
nand U3423 (N_3423,N_3256,N_3200);
or U3424 (N_3424,N_3289,N_3269);
nand U3425 (N_3425,N_3221,N_3385);
nor U3426 (N_3426,N_3328,N_3202);
or U3427 (N_3427,N_3208,N_3238);
or U3428 (N_3428,N_3275,N_3308);
and U3429 (N_3429,N_3326,N_3260);
and U3430 (N_3430,N_3303,N_3248);
or U3431 (N_3431,N_3265,N_3323);
nand U3432 (N_3432,N_3329,N_3365);
nand U3433 (N_3433,N_3319,N_3336);
nand U3434 (N_3434,N_3299,N_3342);
xnor U3435 (N_3435,N_3332,N_3206);
xnor U3436 (N_3436,N_3291,N_3261);
nand U3437 (N_3437,N_3268,N_3259);
nand U3438 (N_3438,N_3343,N_3239);
or U3439 (N_3439,N_3327,N_3278);
nor U3440 (N_3440,N_3203,N_3384);
and U3441 (N_3441,N_3352,N_3383);
or U3442 (N_3442,N_3367,N_3252);
or U3443 (N_3443,N_3350,N_3359);
nand U3444 (N_3444,N_3271,N_3244);
or U3445 (N_3445,N_3357,N_3263);
and U3446 (N_3446,N_3280,N_3262);
nand U3447 (N_3447,N_3276,N_3210);
nand U3448 (N_3448,N_3213,N_3356);
and U3449 (N_3449,N_3273,N_3310);
nor U3450 (N_3450,N_3364,N_3201);
xnor U3451 (N_3451,N_3322,N_3362);
nand U3452 (N_3452,N_3251,N_3366);
nor U3453 (N_3453,N_3300,N_3301);
nor U3454 (N_3454,N_3219,N_3334);
nand U3455 (N_3455,N_3386,N_3287);
nand U3456 (N_3456,N_3399,N_3277);
and U3457 (N_3457,N_3348,N_3355);
nor U3458 (N_3458,N_3207,N_3257);
nor U3459 (N_3459,N_3211,N_3225);
or U3460 (N_3460,N_3226,N_3330);
or U3461 (N_3461,N_3376,N_3214);
nand U3462 (N_3462,N_3390,N_3250);
nor U3463 (N_3463,N_3254,N_3349);
nor U3464 (N_3464,N_3394,N_3242);
xor U3465 (N_3465,N_3375,N_3309);
nand U3466 (N_3466,N_3246,N_3205);
or U3467 (N_3467,N_3361,N_3292);
nand U3468 (N_3468,N_3314,N_3320);
or U3469 (N_3469,N_3231,N_3241);
nor U3470 (N_3470,N_3395,N_3249);
nor U3471 (N_3471,N_3393,N_3296);
and U3472 (N_3472,N_3247,N_3288);
nor U3473 (N_3473,N_3222,N_3216);
and U3474 (N_3474,N_3398,N_3218);
and U3475 (N_3475,N_3378,N_3220);
xor U3476 (N_3476,N_3351,N_3270);
or U3477 (N_3477,N_3258,N_3347);
and U3478 (N_3478,N_3372,N_3279);
or U3479 (N_3479,N_3339,N_3315);
and U3480 (N_3480,N_3369,N_3215);
or U3481 (N_3481,N_3232,N_3388);
or U3482 (N_3482,N_3344,N_3281);
nor U3483 (N_3483,N_3396,N_3354);
nand U3484 (N_3484,N_3227,N_3331);
or U3485 (N_3485,N_3370,N_3389);
nand U3486 (N_3486,N_3282,N_3286);
xnor U3487 (N_3487,N_3318,N_3285);
and U3488 (N_3488,N_3371,N_3298);
and U3489 (N_3489,N_3340,N_3283);
or U3490 (N_3490,N_3360,N_3302);
nand U3491 (N_3491,N_3240,N_3307);
or U3492 (N_3492,N_3363,N_3272);
and U3493 (N_3493,N_3333,N_3223);
or U3494 (N_3494,N_3325,N_3312);
nor U3495 (N_3495,N_3374,N_3230);
nor U3496 (N_3496,N_3317,N_3255);
xnor U3497 (N_3497,N_3274,N_3294);
xor U3498 (N_3498,N_3380,N_3266);
and U3499 (N_3499,N_3212,N_3284);
nand U3500 (N_3500,N_3216,N_3294);
xnor U3501 (N_3501,N_3324,N_3385);
and U3502 (N_3502,N_3324,N_3261);
or U3503 (N_3503,N_3378,N_3250);
and U3504 (N_3504,N_3277,N_3383);
or U3505 (N_3505,N_3283,N_3225);
or U3506 (N_3506,N_3379,N_3384);
nand U3507 (N_3507,N_3310,N_3201);
or U3508 (N_3508,N_3349,N_3356);
nand U3509 (N_3509,N_3272,N_3304);
nor U3510 (N_3510,N_3362,N_3264);
and U3511 (N_3511,N_3217,N_3361);
and U3512 (N_3512,N_3275,N_3316);
or U3513 (N_3513,N_3357,N_3318);
and U3514 (N_3514,N_3221,N_3344);
and U3515 (N_3515,N_3375,N_3336);
or U3516 (N_3516,N_3342,N_3308);
nand U3517 (N_3517,N_3381,N_3291);
or U3518 (N_3518,N_3253,N_3369);
and U3519 (N_3519,N_3272,N_3319);
nand U3520 (N_3520,N_3234,N_3319);
nor U3521 (N_3521,N_3224,N_3258);
and U3522 (N_3522,N_3244,N_3260);
nand U3523 (N_3523,N_3257,N_3274);
or U3524 (N_3524,N_3232,N_3332);
nor U3525 (N_3525,N_3305,N_3222);
xor U3526 (N_3526,N_3231,N_3359);
nand U3527 (N_3527,N_3318,N_3223);
nor U3528 (N_3528,N_3269,N_3366);
nand U3529 (N_3529,N_3259,N_3261);
nor U3530 (N_3530,N_3350,N_3313);
nor U3531 (N_3531,N_3239,N_3263);
xnor U3532 (N_3532,N_3287,N_3345);
or U3533 (N_3533,N_3351,N_3298);
or U3534 (N_3534,N_3361,N_3327);
nand U3535 (N_3535,N_3274,N_3270);
nand U3536 (N_3536,N_3383,N_3249);
nand U3537 (N_3537,N_3274,N_3373);
or U3538 (N_3538,N_3216,N_3305);
and U3539 (N_3539,N_3319,N_3337);
nor U3540 (N_3540,N_3329,N_3305);
and U3541 (N_3541,N_3219,N_3229);
and U3542 (N_3542,N_3202,N_3218);
nor U3543 (N_3543,N_3286,N_3233);
nor U3544 (N_3544,N_3275,N_3277);
nor U3545 (N_3545,N_3290,N_3250);
and U3546 (N_3546,N_3255,N_3269);
and U3547 (N_3547,N_3316,N_3347);
or U3548 (N_3548,N_3322,N_3209);
nor U3549 (N_3549,N_3373,N_3244);
and U3550 (N_3550,N_3396,N_3264);
or U3551 (N_3551,N_3253,N_3205);
and U3552 (N_3552,N_3303,N_3255);
nor U3553 (N_3553,N_3265,N_3322);
and U3554 (N_3554,N_3310,N_3386);
nand U3555 (N_3555,N_3332,N_3360);
and U3556 (N_3556,N_3246,N_3234);
nand U3557 (N_3557,N_3386,N_3384);
or U3558 (N_3558,N_3250,N_3215);
nand U3559 (N_3559,N_3229,N_3341);
nor U3560 (N_3560,N_3318,N_3238);
nand U3561 (N_3561,N_3320,N_3278);
or U3562 (N_3562,N_3226,N_3310);
and U3563 (N_3563,N_3359,N_3265);
and U3564 (N_3564,N_3249,N_3354);
and U3565 (N_3565,N_3394,N_3384);
or U3566 (N_3566,N_3395,N_3337);
nor U3567 (N_3567,N_3264,N_3310);
xnor U3568 (N_3568,N_3285,N_3342);
nor U3569 (N_3569,N_3292,N_3274);
or U3570 (N_3570,N_3387,N_3305);
nand U3571 (N_3571,N_3206,N_3272);
xnor U3572 (N_3572,N_3206,N_3281);
nand U3573 (N_3573,N_3392,N_3232);
nand U3574 (N_3574,N_3238,N_3269);
nand U3575 (N_3575,N_3246,N_3317);
nand U3576 (N_3576,N_3253,N_3270);
and U3577 (N_3577,N_3293,N_3353);
and U3578 (N_3578,N_3322,N_3351);
or U3579 (N_3579,N_3265,N_3341);
or U3580 (N_3580,N_3217,N_3326);
xor U3581 (N_3581,N_3213,N_3364);
and U3582 (N_3582,N_3327,N_3285);
and U3583 (N_3583,N_3209,N_3280);
xnor U3584 (N_3584,N_3202,N_3301);
nor U3585 (N_3585,N_3364,N_3285);
nor U3586 (N_3586,N_3290,N_3262);
and U3587 (N_3587,N_3346,N_3381);
nand U3588 (N_3588,N_3285,N_3333);
and U3589 (N_3589,N_3389,N_3262);
nand U3590 (N_3590,N_3372,N_3226);
nor U3591 (N_3591,N_3200,N_3355);
nor U3592 (N_3592,N_3254,N_3369);
nor U3593 (N_3593,N_3268,N_3265);
or U3594 (N_3594,N_3316,N_3287);
or U3595 (N_3595,N_3282,N_3366);
nor U3596 (N_3596,N_3233,N_3279);
or U3597 (N_3597,N_3242,N_3361);
or U3598 (N_3598,N_3389,N_3336);
nand U3599 (N_3599,N_3291,N_3225);
nor U3600 (N_3600,N_3449,N_3520);
nand U3601 (N_3601,N_3490,N_3472);
nor U3602 (N_3602,N_3536,N_3456);
and U3603 (N_3603,N_3405,N_3547);
xnor U3604 (N_3604,N_3510,N_3544);
nor U3605 (N_3605,N_3407,N_3467);
nor U3606 (N_3606,N_3403,N_3554);
xnor U3607 (N_3607,N_3441,N_3401);
and U3608 (N_3608,N_3521,N_3466);
or U3609 (N_3609,N_3528,N_3560);
or U3610 (N_3610,N_3457,N_3585);
and U3611 (N_3611,N_3553,N_3552);
nand U3612 (N_3612,N_3513,N_3481);
and U3613 (N_3613,N_3514,N_3451);
and U3614 (N_3614,N_3429,N_3478);
and U3615 (N_3615,N_3592,N_3549);
nor U3616 (N_3616,N_3580,N_3425);
or U3617 (N_3617,N_3501,N_3526);
or U3618 (N_3618,N_3414,N_3483);
or U3619 (N_3619,N_3465,N_3492);
or U3620 (N_3620,N_3445,N_3452);
nor U3621 (N_3621,N_3540,N_3402);
xnor U3622 (N_3622,N_3464,N_3594);
nor U3623 (N_3623,N_3555,N_3448);
or U3624 (N_3624,N_3506,N_3569);
nor U3625 (N_3625,N_3487,N_3596);
or U3626 (N_3626,N_3455,N_3420);
and U3627 (N_3627,N_3509,N_3539);
nor U3628 (N_3628,N_3550,N_3563);
xnor U3629 (N_3629,N_3489,N_3484);
nor U3630 (N_3630,N_3515,N_3419);
nor U3631 (N_3631,N_3568,N_3559);
nand U3632 (N_3632,N_3443,N_3562);
and U3633 (N_3633,N_3575,N_3413);
nand U3634 (N_3634,N_3565,N_3459);
nand U3635 (N_3635,N_3453,N_3422);
nor U3636 (N_3636,N_3440,N_3546);
and U3637 (N_3637,N_3548,N_3479);
nor U3638 (N_3638,N_3411,N_3423);
or U3639 (N_3639,N_3523,N_3577);
or U3640 (N_3640,N_3486,N_3545);
and U3641 (N_3641,N_3482,N_3438);
or U3642 (N_3642,N_3507,N_3535);
and U3643 (N_3643,N_3511,N_3593);
nand U3644 (N_3644,N_3541,N_3542);
nor U3645 (N_3645,N_3462,N_3532);
nand U3646 (N_3646,N_3587,N_3500);
xor U3647 (N_3647,N_3418,N_3400);
xnor U3648 (N_3648,N_3436,N_3431);
and U3649 (N_3649,N_3469,N_3473);
nor U3650 (N_3650,N_3497,N_3442);
or U3651 (N_3651,N_3446,N_3493);
or U3652 (N_3652,N_3576,N_3579);
and U3653 (N_3653,N_3599,N_3517);
nor U3654 (N_3654,N_3586,N_3537);
nor U3655 (N_3655,N_3427,N_3551);
and U3656 (N_3656,N_3426,N_3558);
nand U3657 (N_3657,N_3505,N_3404);
nand U3658 (N_3658,N_3430,N_3499);
nor U3659 (N_3659,N_3435,N_3581);
nor U3660 (N_3660,N_3471,N_3480);
and U3661 (N_3661,N_3529,N_3424);
nor U3662 (N_3662,N_3582,N_3556);
nand U3663 (N_3663,N_3460,N_3573);
nand U3664 (N_3664,N_3561,N_3463);
nand U3665 (N_3665,N_3564,N_3406);
nor U3666 (N_3666,N_3595,N_3571);
xnor U3667 (N_3667,N_3584,N_3530);
nor U3668 (N_3668,N_3572,N_3428);
or U3669 (N_3669,N_3538,N_3591);
or U3670 (N_3670,N_3409,N_3503);
and U3671 (N_3671,N_3412,N_3525);
nand U3672 (N_3672,N_3447,N_3557);
nor U3673 (N_3673,N_3476,N_3488);
xnor U3674 (N_3674,N_3508,N_3516);
nand U3675 (N_3675,N_3524,N_3421);
or U3676 (N_3676,N_3434,N_3439);
nor U3677 (N_3677,N_3410,N_3498);
nand U3678 (N_3678,N_3504,N_3531);
nand U3679 (N_3679,N_3574,N_3512);
and U3680 (N_3680,N_3458,N_3533);
nand U3681 (N_3681,N_3534,N_3475);
and U3682 (N_3682,N_3474,N_3589);
nand U3683 (N_3683,N_3543,N_3588);
and U3684 (N_3684,N_3450,N_3408);
nand U3685 (N_3685,N_3416,N_3432);
xnor U3686 (N_3686,N_3590,N_3502);
and U3687 (N_3687,N_3417,N_3527);
or U3688 (N_3688,N_3598,N_3454);
or U3689 (N_3689,N_3477,N_3444);
nand U3690 (N_3690,N_3566,N_3578);
or U3691 (N_3691,N_3461,N_3583);
nor U3692 (N_3692,N_3437,N_3597);
or U3693 (N_3693,N_3495,N_3570);
and U3694 (N_3694,N_3494,N_3567);
nand U3695 (N_3695,N_3433,N_3491);
and U3696 (N_3696,N_3496,N_3485);
and U3697 (N_3697,N_3518,N_3519);
nor U3698 (N_3698,N_3522,N_3468);
and U3699 (N_3699,N_3415,N_3470);
nand U3700 (N_3700,N_3464,N_3513);
and U3701 (N_3701,N_3438,N_3569);
nand U3702 (N_3702,N_3590,N_3471);
or U3703 (N_3703,N_3449,N_3497);
and U3704 (N_3704,N_3449,N_3561);
and U3705 (N_3705,N_3516,N_3587);
nor U3706 (N_3706,N_3437,N_3414);
nand U3707 (N_3707,N_3454,N_3507);
and U3708 (N_3708,N_3519,N_3487);
nand U3709 (N_3709,N_3455,N_3513);
or U3710 (N_3710,N_3472,N_3502);
nor U3711 (N_3711,N_3574,N_3499);
nand U3712 (N_3712,N_3438,N_3504);
nand U3713 (N_3713,N_3566,N_3576);
nor U3714 (N_3714,N_3423,N_3504);
and U3715 (N_3715,N_3510,N_3496);
nor U3716 (N_3716,N_3460,N_3542);
xor U3717 (N_3717,N_3598,N_3441);
nand U3718 (N_3718,N_3534,N_3566);
xnor U3719 (N_3719,N_3519,N_3576);
or U3720 (N_3720,N_3504,N_3427);
and U3721 (N_3721,N_3508,N_3502);
and U3722 (N_3722,N_3483,N_3590);
nand U3723 (N_3723,N_3475,N_3523);
or U3724 (N_3724,N_3475,N_3431);
and U3725 (N_3725,N_3441,N_3479);
nor U3726 (N_3726,N_3559,N_3449);
and U3727 (N_3727,N_3428,N_3599);
or U3728 (N_3728,N_3455,N_3533);
xnor U3729 (N_3729,N_3501,N_3491);
nand U3730 (N_3730,N_3550,N_3521);
nor U3731 (N_3731,N_3479,N_3598);
nand U3732 (N_3732,N_3448,N_3533);
xor U3733 (N_3733,N_3586,N_3461);
and U3734 (N_3734,N_3581,N_3524);
and U3735 (N_3735,N_3452,N_3415);
nand U3736 (N_3736,N_3577,N_3495);
nor U3737 (N_3737,N_3483,N_3559);
nor U3738 (N_3738,N_3445,N_3570);
nand U3739 (N_3739,N_3517,N_3466);
and U3740 (N_3740,N_3475,N_3501);
nand U3741 (N_3741,N_3562,N_3478);
nor U3742 (N_3742,N_3557,N_3430);
nand U3743 (N_3743,N_3426,N_3583);
nand U3744 (N_3744,N_3508,N_3549);
nand U3745 (N_3745,N_3598,N_3461);
and U3746 (N_3746,N_3582,N_3479);
xor U3747 (N_3747,N_3518,N_3500);
or U3748 (N_3748,N_3514,N_3469);
xnor U3749 (N_3749,N_3505,N_3552);
nor U3750 (N_3750,N_3409,N_3567);
nor U3751 (N_3751,N_3544,N_3431);
or U3752 (N_3752,N_3445,N_3597);
and U3753 (N_3753,N_3566,N_3563);
or U3754 (N_3754,N_3522,N_3577);
nor U3755 (N_3755,N_3483,N_3528);
nor U3756 (N_3756,N_3462,N_3488);
nand U3757 (N_3757,N_3445,N_3596);
nor U3758 (N_3758,N_3569,N_3486);
and U3759 (N_3759,N_3406,N_3524);
or U3760 (N_3760,N_3402,N_3475);
and U3761 (N_3761,N_3553,N_3486);
and U3762 (N_3762,N_3414,N_3515);
and U3763 (N_3763,N_3592,N_3479);
xor U3764 (N_3764,N_3564,N_3448);
nand U3765 (N_3765,N_3515,N_3528);
or U3766 (N_3766,N_3555,N_3443);
or U3767 (N_3767,N_3465,N_3497);
or U3768 (N_3768,N_3565,N_3519);
xor U3769 (N_3769,N_3487,N_3403);
and U3770 (N_3770,N_3499,N_3591);
or U3771 (N_3771,N_3498,N_3528);
nand U3772 (N_3772,N_3537,N_3559);
nor U3773 (N_3773,N_3553,N_3408);
or U3774 (N_3774,N_3593,N_3523);
or U3775 (N_3775,N_3403,N_3479);
and U3776 (N_3776,N_3400,N_3506);
nor U3777 (N_3777,N_3544,N_3550);
nor U3778 (N_3778,N_3519,N_3472);
nand U3779 (N_3779,N_3589,N_3500);
and U3780 (N_3780,N_3491,N_3515);
xnor U3781 (N_3781,N_3567,N_3432);
or U3782 (N_3782,N_3401,N_3429);
nand U3783 (N_3783,N_3491,N_3570);
xnor U3784 (N_3784,N_3530,N_3458);
nor U3785 (N_3785,N_3432,N_3468);
or U3786 (N_3786,N_3441,N_3550);
nand U3787 (N_3787,N_3473,N_3509);
xnor U3788 (N_3788,N_3548,N_3435);
or U3789 (N_3789,N_3517,N_3400);
nor U3790 (N_3790,N_3519,N_3507);
or U3791 (N_3791,N_3448,N_3515);
nand U3792 (N_3792,N_3594,N_3593);
or U3793 (N_3793,N_3424,N_3494);
nand U3794 (N_3794,N_3471,N_3522);
nor U3795 (N_3795,N_3433,N_3487);
or U3796 (N_3796,N_3431,N_3470);
or U3797 (N_3797,N_3445,N_3493);
and U3798 (N_3798,N_3470,N_3587);
nor U3799 (N_3799,N_3438,N_3412);
nor U3800 (N_3800,N_3633,N_3726);
nor U3801 (N_3801,N_3746,N_3761);
or U3802 (N_3802,N_3614,N_3650);
and U3803 (N_3803,N_3669,N_3735);
or U3804 (N_3804,N_3792,N_3798);
nand U3805 (N_3805,N_3613,N_3694);
nor U3806 (N_3806,N_3736,N_3672);
or U3807 (N_3807,N_3796,N_3605);
nand U3808 (N_3808,N_3739,N_3656);
nor U3809 (N_3809,N_3767,N_3634);
nand U3810 (N_3810,N_3774,N_3671);
and U3811 (N_3811,N_3619,N_3632);
nor U3812 (N_3812,N_3775,N_3799);
nand U3813 (N_3813,N_3670,N_3743);
nor U3814 (N_3814,N_3688,N_3703);
and U3815 (N_3815,N_3678,N_3795);
xnor U3816 (N_3816,N_3651,N_3716);
nor U3817 (N_3817,N_3686,N_3684);
or U3818 (N_3818,N_3717,N_3727);
nor U3819 (N_3819,N_3609,N_3759);
xor U3820 (N_3820,N_3610,N_3606);
and U3821 (N_3821,N_3756,N_3662);
nand U3822 (N_3822,N_3787,N_3778);
and U3823 (N_3823,N_3734,N_3620);
xnor U3824 (N_3824,N_3693,N_3718);
or U3825 (N_3825,N_3719,N_3770);
nor U3826 (N_3826,N_3689,N_3637);
nor U3827 (N_3827,N_3772,N_3742);
nand U3828 (N_3828,N_3607,N_3748);
nor U3829 (N_3829,N_3685,N_3704);
nor U3830 (N_3830,N_3602,N_3653);
nor U3831 (N_3831,N_3749,N_3608);
nor U3832 (N_3832,N_3700,N_3640);
nor U3833 (N_3833,N_3753,N_3728);
or U3834 (N_3834,N_3715,N_3732);
and U3835 (N_3835,N_3622,N_3713);
xor U3836 (N_3836,N_3663,N_3616);
nand U3837 (N_3837,N_3745,N_3635);
and U3838 (N_3838,N_3647,N_3665);
nor U3839 (N_3839,N_3623,N_3738);
nor U3840 (N_3840,N_3661,N_3625);
xor U3841 (N_3841,N_3757,N_3786);
xor U3842 (N_3842,N_3744,N_3681);
nand U3843 (N_3843,N_3766,N_3692);
xnor U3844 (N_3844,N_3711,N_3763);
or U3845 (N_3845,N_3636,N_3747);
nor U3846 (N_3846,N_3658,N_3789);
or U3847 (N_3847,N_3723,N_3624);
nor U3848 (N_3848,N_3649,N_3784);
nor U3849 (N_3849,N_3621,N_3724);
and U3850 (N_3850,N_3706,N_3722);
nand U3851 (N_3851,N_3675,N_3628);
or U3852 (N_3852,N_3652,N_3641);
nand U3853 (N_3853,N_3687,N_3783);
or U3854 (N_3854,N_3617,N_3643);
and U3855 (N_3855,N_3603,N_3779);
nor U3856 (N_3856,N_3730,N_3768);
nand U3857 (N_3857,N_3655,N_3710);
or U3858 (N_3858,N_3639,N_3701);
or U3859 (N_3859,N_3659,N_3611);
xor U3860 (N_3860,N_3705,N_3638);
and U3861 (N_3861,N_3752,N_3791);
or U3862 (N_3862,N_3714,N_3721);
nor U3863 (N_3863,N_3776,N_3790);
and U3864 (N_3864,N_3771,N_3618);
or U3865 (N_3865,N_3612,N_3773);
nand U3866 (N_3866,N_3777,N_3702);
nor U3867 (N_3867,N_3630,N_3712);
nor U3868 (N_3868,N_3696,N_3780);
or U3869 (N_3869,N_3601,N_3691);
or U3870 (N_3870,N_3660,N_3679);
nand U3871 (N_3871,N_3676,N_3758);
and U3872 (N_3872,N_3737,N_3668);
and U3873 (N_3873,N_3631,N_3731);
and U3874 (N_3874,N_3645,N_3754);
nand U3875 (N_3875,N_3648,N_3785);
nor U3876 (N_3876,N_3769,N_3781);
or U3877 (N_3877,N_3708,N_3765);
nor U3878 (N_3878,N_3680,N_3733);
or U3879 (N_3879,N_3697,N_3707);
nand U3880 (N_3880,N_3674,N_3627);
nand U3881 (N_3881,N_3750,N_3690);
nor U3882 (N_3882,N_3600,N_3755);
and U3883 (N_3883,N_3673,N_3654);
or U3884 (N_3884,N_3644,N_3729);
nor U3885 (N_3885,N_3698,N_3677);
nor U3886 (N_3886,N_3788,N_3760);
nor U3887 (N_3887,N_3740,N_3629);
or U3888 (N_3888,N_3626,N_3646);
or U3889 (N_3889,N_3709,N_3666);
or U3890 (N_3890,N_3615,N_3725);
and U3891 (N_3891,N_3782,N_3683);
nand U3892 (N_3892,N_3764,N_3762);
nor U3893 (N_3893,N_3794,N_3657);
and U3894 (N_3894,N_3695,N_3741);
nand U3895 (N_3895,N_3642,N_3797);
or U3896 (N_3896,N_3682,N_3793);
nand U3897 (N_3897,N_3664,N_3720);
or U3898 (N_3898,N_3751,N_3667);
nand U3899 (N_3899,N_3699,N_3604);
nand U3900 (N_3900,N_3600,N_3664);
and U3901 (N_3901,N_3711,N_3761);
or U3902 (N_3902,N_3651,N_3788);
and U3903 (N_3903,N_3673,N_3789);
and U3904 (N_3904,N_3613,N_3644);
and U3905 (N_3905,N_3764,N_3748);
nand U3906 (N_3906,N_3675,N_3772);
and U3907 (N_3907,N_3645,N_3727);
and U3908 (N_3908,N_3704,N_3664);
nand U3909 (N_3909,N_3782,N_3611);
nand U3910 (N_3910,N_3606,N_3799);
nand U3911 (N_3911,N_3734,N_3668);
nand U3912 (N_3912,N_3670,N_3607);
nand U3913 (N_3913,N_3657,N_3719);
or U3914 (N_3914,N_3640,N_3781);
or U3915 (N_3915,N_3605,N_3772);
xor U3916 (N_3916,N_3696,N_3685);
nor U3917 (N_3917,N_3760,N_3664);
xor U3918 (N_3918,N_3674,N_3719);
nor U3919 (N_3919,N_3634,N_3684);
nor U3920 (N_3920,N_3658,N_3722);
and U3921 (N_3921,N_3713,N_3625);
and U3922 (N_3922,N_3775,N_3793);
or U3923 (N_3923,N_3786,N_3783);
nor U3924 (N_3924,N_3778,N_3614);
and U3925 (N_3925,N_3781,N_3622);
and U3926 (N_3926,N_3757,N_3670);
or U3927 (N_3927,N_3701,N_3798);
nand U3928 (N_3928,N_3751,N_3716);
or U3929 (N_3929,N_3700,N_3652);
xnor U3930 (N_3930,N_3705,N_3676);
nand U3931 (N_3931,N_3738,N_3784);
nor U3932 (N_3932,N_3690,N_3602);
or U3933 (N_3933,N_3630,N_3768);
nand U3934 (N_3934,N_3782,N_3610);
xor U3935 (N_3935,N_3763,N_3629);
or U3936 (N_3936,N_3794,N_3761);
nor U3937 (N_3937,N_3780,N_3785);
nor U3938 (N_3938,N_3605,N_3725);
xor U3939 (N_3939,N_3612,N_3765);
nor U3940 (N_3940,N_3726,N_3777);
xnor U3941 (N_3941,N_3762,N_3733);
nand U3942 (N_3942,N_3682,N_3738);
nor U3943 (N_3943,N_3787,N_3738);
nand U3944 (N_3944,N_3707,N_3796);
or U3945 (N_3945,N_3636,N_3735);
nor U3946 (N_3946,N_3610,N_3604);
xor U3947 (N_3947,N_3655,N_3714);
xor U3948 (N_3948,N_3773,N_3750);
nand U3949 (N_3949,N_3792,N_3690);
and U3950 (N_3950,N_3742,N_3691);
or U3951 (N_3951,N_3617,N_3782);
nand U3952 (N_3952,N_3679,N_3699);
or U3953 (N_3953,N_3648,N_3797);
nand U3954 (N_3954,N_3756,N_3728);
or U3955 (N_3955,N_3637,N_3601);
nor U3956 (N_3956,N_3654,N_3779);
nand U3957 (N_3957,N_3669,N_3725);
or U3958 (N_3958,N_3726,N_3767);
or U3959 (N_3959,N_3640,N_3651);
nand U3960 (N_3960,N_3681,N_3682);
and U3961 (N_3961,N_3629,N_3789);
xnor U3962 (N_3962,N_3685,N_3791);
and U3963 (N_3963,N_3657,N_3795);
or U3964 (N_3964,N_3708,N_3739);
or U3965 (N_3965,N_3674,N_3790);
and U3966 (N_3966,N_3687,N_3777);
or U3967 (N_3967,N_3699,N_3771);
nor U3968 (N_3968,N_3654,N_3713);
nand U3969 (N_3969,N_3769,N_3621);
nand U3970 (N_3970,N_3784,N_3691);
nand U3971 (N_3971,N_3610,N_3673);
or U3972 (N_3972,N_3785,N_3657);
and U3973 (N_3973,N_3696,N_3716);
nor U3974 (N_3974,N_3677,N_3676);
nor U3975 (N_3975,N_3714,N_3779);
or U3976 (N_3976,N_3629,N_3750);
and U3977 (N_3977,N_3667,N_3690);
and U3978 (N_3978,N_3603,N_3674);
or U3979 (N_3979,N_3670,N_3763);
nor U3980 (N_3980,N_3736,N_3673);
xnor U3981 (N_3981,N_3714,N_3634);
nand U3982 (N_3982,N_3608,N_3793);
nand U3983 (N_3983,N_3700,N_3714);
and U3984 (N_3984,N_3724,N_3792);
nand U3985 (N_3985,N_3707,N_3686);
and U3986 (N_3986,N_3721,N_3631);
or U3987 (N_3987,N_3663,N_3740);
or U3988 (N_3988,N_3603,N_3654);
or U3989 (N_3989,N_3652,N_3658);
xnor U3990 (N_3990,N_3778,N_3774);
or U3991 (N_3991,N_3688,N_3634);
nor U3992 (N_3992,N_3668,N_3797);
xnor U3993 (N_3993,N_3696,N_3793);
and U3994 (N_3994,N_3643,N_3792);
nor U3995 (N_3995,N_3655,N_3660);
xor U3996 (N_3996,N_3789,N_3638);
nand U3997 (N_3997,N_3603,N_3634);
or U3998 (N_3998,N_3647,N_3629);
and U3999 (N_3999,N_3712,N_3677);
or U4000 (N_4000,N_3880,N_3910);
nor U4001 (N_4001,N_3891,N_3862);
nor U4002 (N_4002,N_3875,N_3907);
and U4003 (N_4003,N_3872,N_3983);
xor U4004 (N_4004,N_3896,N_3846);
and U4005 (N_4005,N_3980,N_3964);
nand U4006 (N_4006,N_3956,N_3932);
and U4007 (N_4007,N_3851,N_3975);
nor U4008 (N_4008,N_3929,N_3874);
and U4009 (N_4009,N_3840,N_3925);
and U4010 (N_4010,N_3911,N_3835);
or U4011 (N_4011,N_3999,N_3953);
and U4012 (N_4012,N_3865,N_3923);
nor U4013 (N_4013,N_3989,N_3958);
or U4014 (N_4014,N_3921,N_3856);
nand U4015 (N_4015,N_3823,N_3952);
xor U4016 (N_4016,N_3943,N_3849);
or U4017 (N_4017,N_3945,N_3931);
nor U4018 (N_4018,N_3982,N_3930);
nor U4019 (N_4019,N_3969,N_3900);
and U4020 (N_4020,N_3876,N_3811);
or U4021 (N_4021,N_3818,N_3967);
nor U4022 (N_4022,N_3904,N_3801);
and U4023 (N_4023,N_3947,N_3939);
or U4024 (N_4024,N_3981,N_3887);
nor U4025 (N_4025,N_3955,N_3869);
or U4026 (N_4026,N_3993,N_3976);
nor U4027 (N_4027,N_3936,N_3909);
or U4028 (N_4028,N_3838,N_3917);
nand U4029 (N_4029,N_3831,N_3841);
or U4030 (N_4030,N_3889,N_3863);
nand U4031 (N_4031,N_3919,N_3817);
nand U4032 (N_4032,N_3915,N_3899);
xor U4033 (N_4033,N_3822,N_3805);
and U4034 (N_4034,N_3806,N_3903);
nor U4035 (N_4035,N_3918,N_3987);
or U4036 (N_4036,N_3814,N_3803);
nand U4037 (N_4037,N_3885,N_3833);
and U4038 (N_4038,N_3912,N_3837);
nand U4039 (N_4039,N_3933,N_3834);
nand U4040 (N_4040,N_3908,N_3859);
and U4041 (N_4041,N_3860,N_3997);
nand U4042 (N_4042,N_3988,N_3973);
or U4043 (N_4043,N_3944,N_3960);
or U4044 (N_4044,N_3984,N_3820);
and U4045 (N_4045,N_3836,N_3819);
nor U4046 (N_4046,N_3961,N_3882);
and U4047 (N_4047,N_3959,N_3968);
nor U4048 (N_4048,N_3992,N_3853);
xor U4049 (N_4049,N_3893,N_3985);
nor U4050 (N_4050,N_3934,N_3867);
and U4051 (N_4051,N_3996,N_3901);
and U4052 (N_4052,N_3935,N_3857);
nand U4053 (N_4053,N_3883,N_3942);
nor U4054 (N_4054,N_3884,N_3886);
nor U4055 (N_4055,N_3965,N_3812);
nand U4056 (N_4056,N_3847,N_3892);
or U4057 (N_4057,N_3950,N_3844);
and U4058 (N_4058,N_3848,N_3825);
xor U4059 (N_4059,N_3991,N_3854);
or U4060 (N_4060,N_3873,N_3895);
nand U4061 (N_4061,N_3938,N_3824);
or U4062 (N_4062,N_3970,N_3877);
nand U4063 (N_4063,N_3902,N_3878);
nand U4064 (N_4064,N_3871,N_3894);
and U4065 (N_4065,N_3816,N_3977);
and U4066 (N_4066,N_3890,N_3828);
xor U4067 (N_4067,N_3839,N_3926);
and U4068 (N_4068,N_3821,N_3978);
or U4069 (N_4069,N_3868,N_3920);
and U4070 (N_4070,N_3864,N_3905);
nor U4071 (N_4071,N_3994,N_3951);
nand U4072 (N_4072,N_3855,N_3830);
and U4073 (N_4073,N_3852,N_3827);
or U4074 (N_4074,N_3928,N_3800);
nor U4075 (N_4075,N_3810,N_3962);
or U4076 (N_4076,N_3957,N_3924);
nor U4077 (N_4077,N_3861,N_3858);
or U4078 (N_4078,N_3898,N_3842);
and U4079 (N_4079,N_3815,N_3897);
and U4080 (N_4080,N_3946,N_3916);
nor U4081 (N_4081,N_3937,N_3971);
nand U4082 (N_4082,N_3832,N_3979);
or U4083 (N_4083,N_3949,N_3972);
and U4084 (N_4084,N_3813,N_3986);
and U4085 (N_4085,N_3843,N_3906);
and U4086 (N_4086,N_3826,N_3829);
nand U4087 (N_4087,N_3922,N_3954);
or U4088 (N_4088,N_3913,N_3914);
and U4089 (N_4089,N_3808,N_3940);
and U4090 (N_4090,N_3941,N_3995);
xor U4091 (N_4091,N_3966,N_3866);
and U4092 (N_4092,N_3809,N_3948);
nor U4093 (N_4093,N_3807,N_3879);
xor U4094 (N_4094,N_3927,N_3888);
nor U4095 (N_4095,N_3850,N_3998);
and U4096 (N_4096,N_3802,N_3870);
nand U4097 (N_4097,N_3963,N_3881);
or U4098 (N_4098,N_3804,N_3990);
or U4099 (N_4099,N_3845,N_3974);
xnor U4100 (N_4100,N_3821,N_3896);
nor U4101 (N_4101,N_3915,N_3912);
nor U4102 (N_4102,N_3818,N_3905);
or U4103 (N_4103,N_3958,N_3860);
nor U4104 (N_4104,N_3895,N_3960);
or U4105 (N_4105,N_3955,N_3969);
nand U4106 (N_4106,N_3881,N_3879);
nor U4107 (N_4107,N_3928,N_3809);
nand U4108 (N_4108,N_3957,N_3840);
nor U4109 (N_4109,N_3977,N_3829);
nor U4110 (N_4110,N_3836,N_3924);
nor U4111 (N_4111,N_3990,N_3812);
or U4112 (N_4112,N_3961,N_3837);
nor U4113 (N_4113,N_3849,N_3983);
and U4114 (N_4114,N_3821,N_3909);
and U4115 (N_4115,N_3920,N_3841);
xnor U4116 (N_4116,N_3866,N_3862);
nand U4117 (N_4117,N_3808,N_3916);
xor U4118 (N_4118,N_3977,N_3811);
nor U4119 (N_4119,N_3888,N_3983);
nand U4120 (N_4120,N_3824,N_3975);
and U4121 (N_4121,N_3823,N_3855);
nor U4122 (N_4122,N_3811,N_3853);
and U4123 (N_4123,N_3947,N_3809);
nor U4124 (N_4124,N_3887,N_3825);
nand U4125 (N_4125,N_3917,N_3808);
xnor U4126 (N_4126,N_3887,N_3828);
and U4127 (N_4127,N_3913,N_3880);
or U4128 (N_4128,N_3864,N_3993);
or U4129 (N_4129,N_3946,N_3925);
or U4130 (N_4130,N_3875,N_3813);
nor U4131 (N_4131,N_3968,N_3863);
nand U4132 (N_4132,N_3905,N_3953);
nor U4133 (N_4133,N_3897,N_3836);
nand U4134 (N_4134,N_3989,N_3977);
or U4135 (N_4135,N_3918,N_3819);
xnor U4136 (N_4136,N_3940,N_3965);
xnor U4137 (N_4137,N_3821,N_3982);
and U4138 (N_4138,N_3840,N_3853);
and U4139 (N_4139,N_3910,N_3802);
nor U4140 (N_4140,N_3966,N_3988);
nor U4141 (N_4141,N_3924,N_3939);
and U4142 (N_4142,N_3990,N_3951);
and U4143 (N_4143,N_3817,N_3999);
or U4144 (N_4144,N_3863,N_3858);
or U4145 (N_4145,N_3913,N_3984);
or U4146 (N_4146,N_3804,N_3803);
nand U4147 (N_4147,N_3865,N_3998);
nand U4148 (N_4148,N_3955,N_3925);
or U4149 (N_4149,N_3938,N_3904);
nand U4150 (N_4150,N_3823,N_3848);
nor U4151 (N_4151,N_3896,N_3872);
or U4152 (N_4152,N_3925,N_3932);
xnor U4153 (N_4153,N_3849,N_3878);
and U4154 (N_4154,N_3802,N_3919);
or U4155 (N_4155,N_3929,N_3863);
nor U4156 (N_4156,N_3883,N_3873);
and U4157 (N_4157,N_3860,N_3847);
and U4158 (N_4158,N_3915,N_3820);
or U4159 (N_4159,N_3921,N_3976);
and U4160 (N_4160,N_3952,N_3972);
or U4161 (N_4161,N_3954,N_3999);
or U4162 (N_4162,N_3894,N_3936);
nor U4163 (N_4163,N_3845,N_3927);
or U4164 (N_4164,N_3894,N_3925);
and U4165 (N_4165,N_3823,N_3917);
or U4166 (N_4166,N_3803,N_3826);
or U4167 (N_4167,N_3839,N_3865);
or U4168 (N_4168,N_3940,N_3913);
nor U4169 (N_4169,N_3920,N_3875);
nand U4170 (N_4170,N_3842,N_3970);
nand U4171 (N_4171,N_3901,N_3962);
or U4172 (N_4172,N_3824,N_3834);
and U4173 (N_4173,N_3844,N_3826);
nand U4174 (N_4174,N_3939,N_3858);
nor U4175 (N_4175,N_3889,N_3981);
or U4176 (N_4176,N_3871,N_3891);
or U4177 (N_4177,N_3960,N_3977);
xnor U4178 (N_4178,N_3827,N_3952);
and U4179 (N_4179,N_3887,N_3920);
nor U4180 (N_4180,N_3919,N_3848);
nand U4181 (N_4181,N_3901,N_3828);
or U4182 (N_4182,N_3997,N_3871);
nor U4183 (N_4183,N_3972,N_3956);
nor U4184 (N_4184,N_3858,N_3970);
and U4185 (N_4185,N_3889,N_3932);
nand U4186 (N_4186,N_3893,N_3823);
and U4187 (N_4187,N_3814,N_3977);
or U4188 (N_4188,N_3887,N_3936);
and U4189 (N_4189,N_3845,N_3893);
nor U4190 (N_4190,N_3861,N_3888);
nand U4191 (N_4191,N_3999,N_3803);
nand U4192 (N_4192,N_3963,N_3880);
nand U4193 (N_4193,N_3993,N_3895);
xor U4194 (N_4194,N_3816,N_3880);
or U4195 (N_4195,N_3929,N_3956);
xnor U4196 (N_4196,N_3962,N_3804);
and U4197 (N_4197,N_3856,N_3968);
nor U4198 (N_4198,N_3931,N_3865);
xor U4199 (N_4199,N_3957,N_3987);
and U4200 (N_4200,N_4103,N_4027);
nor U4201 (N_4201,N_4179,N_4108);
or U4202 (N_4202,N_4125,N_4147);
and U4203 (N_4203,N_4061,N_4175);
and U4204 (N_4204,N_4038,N_4170);
xnor U4205 (N_4205,N_4030,N_4031);
and U4206 (N_4206,N_4084,N_4075);
and U4207 (N_4207,N_4153,N_4109);
nor U4208 (N_4208,N_4141,N_4080);
or U4209 (N_4209,N_4195,N_4012);
and U4210 (N_4210,N_4000,N_4057);
nand U4211 (N_4211,N_4191,N_4156);
nand U4212 (N_4212,N_4100,N_4065);
nor U4213 (N_4213,N_4095,N_4094);
nand U4214 (N_4214,N_4181,N_4197);
xnor U4215 (N_4215,N_4097,N_4149);
and U4216 (N_4216,N_4107,N_4187);
xor U4217 (N_4217,N_4056,N_4172);
xor U4218 (N_4218,N_4135,N_4101);
or U4219 (N_4219,N_4035,N_4188);
nor U4220 (N_4220,N_4037,N_4159);
nand U4221 (N_4221,N_4019,N_4169);
or U4222 (N_4222,N_4011,N_4150);
nand U4223 (N_4223,N_4130,N_4196);
nand U4224 (N_4224,N_4180,N_4118);
and U4225 (N_4225,N_4124,N_4016);
or U4226 (N_4226,N_4059,N_4032);
or U4227 (N_4227,N_4166,N_4161);
nand U4228 (N_4228,N_4115,N_4071);
or U4229 (N_4229,N_4171,N_4067);
and U4230 (N_4230,N_4190,N_4041);
xor U4231 (N_4231,N_4162,N_4111);
nand U4232 (N_4232,N_4102,N_4069);
nand U4233 (N_4233,N_4114,N_4020);
or U4234 (N_4234,N_4048,N_4145);
and U4235 (N_4235,N_4157,N_4110);
and U4236 (N_4236,N_4033,N_4009);
nand U4237 (N_4237,N_4066,N_4042);
nor U4238 (N_4238,N_4052,N_4015);
xnor U4239 (N_4239,N_4178,N_4122);
or U4240 (N_4240,N_4079,N_4025);
nor U4241 (N_4241,N_4136,N_4092);
or U4242 (N_4242,N_4006,N_4082);
or U4243 (N_4243,N_4013,N_4008);
nor U4244 (N_4244,N_4173,N_4024);
or U4245 (N_4245,N_4113,N_4116);
nand U4246 (N_4246,N_4077,N_4007);
xor U4247 (N_4247,N_4026,N_4072);
or U4248 (N_4248,N_4098,N_4089);
and U4249 (N_4249,N_4164,N_4039);
or U4250 (N_4250,N_4078,N_4189);
or U4251 (N_4251,N_4152,N_4112);
or U4252 (N_4252,N_4001,N_4049);
nand U4253 (N_4253,N_4064,N_4158);
nor U4254 (N_4254,N_4083,N_4093);
nand U4255 (N_4255,N_4134,N_4129);
nor U4256 (N_4256,N_4148,N_4023);
or U4257 (N_4257,N_4045,N_4054);
nor U4258 (N_4258,N_4050,N_4002);
and U4259 (N_4259,N_4140,N_4105);
nor U4260 (N_4260,N_4167,N_4021);
nand U4261 (N_4261,N_4051,N_4198);
and U4262 (N_4262,N_4154,N_4018);
nor U4263 (N_4263,N_4183,N_4151);
nand U4264 (N_4264,N_4184,N_4090);
or U4265 (N_4265,N_4146,N_4028);
nand U4266 (N_4266,N_4099,N_4174);
and U4267 (N_4267,N_4127,N_4117);
or U4268 (N_4268,N_4055,N_4034);
nor U4269 (N_4269,N_4163,N_4058);
and U4270 (N_4270,N_4029,N_4063);
and U4271 (N_4271,N_4182,N_4168);
or U4272 (N_4272,N_4068,N_4086);
or U4273 (N_4273,N_4123,N_4005);
nor U4274 (N_4274,N_4047,N_4081);
or U4275 (N_4275,N_4036,N_4132);
nand U4276 (N_4276,N_4138,N_4194);
or U4277 (N_4277,N_4185,N_4014);
nor U4278 (N_4278,N_4096,N_4088);
nor U4279 (N_4279,N_4160,N_4104);
nor U4280 (N_4280,N_4142,N_4017);
or U4281 (N_4281,N_4165,N_4133);
nor U4282 (N_4282,N_4073,N_4053);
and U4283 (N_4283,N_4139,N_4074);
nand U4284 (N_4284,N_4062,N_4199);
and U4285 (N_4285,N_4120,N_4177);
nor U4286 (N_4286,N_4010,N_4126);
and U4287 (N_4287,N_4192,N_4176);
nor U4288 (N_4288,N_4040,N_4003);
and U4289 (N_4289,N_4060,N_4004);
nand U4290 (N_4290,N_4070,N_4091);
nand U4291 (N_4291,N_4046,N_4144);
and U4292 (N_4292,N_4076,N_4106);
nand U4293 (N_4293,N_4131,N_4022);
nor U4294 (N_4294,N_4121,N_4155);
nor U4295 (N_4295,N_4119,N_4193);
and U4296 (N_4296,N_4085,N_4143);
or U4297 (N_4297,N_4087,N_4137);
or U4298 (N_4298,N_4043,N_4128);
nand U4299 (N_4299,N_4186,N_4044);
and U4300 (N_4300,N_4028,N_4069);
nand U4301 (N_4301,N_4036,N_4022);
or U4302 (N_4302,N_4110,N_4136);
nand U4303 (N_4303,N_4022,N_4123);
xor U4304 (N_4304,N_4167,N_4081);
or U4305 (N_4305,N_4076,N_4014);
xor U4306 (N_4306,N_4091,N_4178);
nand U4307 (N_4307,N_4169,N_4059);
or U4308 (N_4308,N_4019,N_4181);
nor U4309 (N_4309,N_4177,N_4040);
nand U4310 (N_4310,N_4127,N_4028);
nor U4311 (N_4311,N_4068,N_4031);
nor U4312 (N_4312,N_4090,N_4018);
xor U4313 (N_4313,N_4050,N_4052);
nand U4314 (N_4314,N_4186,N_4019);
xor U4315 (N_4315,N_4076,N_4180);
and U4316 (N_4316,N_4126,N_4156);
nor U4317 (N_4317,N_4076,N_4191);
xnor U4318 (N_4318,N_4176,N_4004);
nor U4319 (N_4319,N_4155,N_4173);
nand U4320 (N_4320,N_4183,N_4090);
nand U4321 (N_4321,N_4104,N_4153);
or U4322 (N_4322,N_4064,N_4151);
xor U4323 (N_4323,N_4124,N_4103);
or U4324 (N_4324,N_4111,N_4180);
and U4325 (N_4325,N_4110,N_4093);
or U4326 (N_4326,N_4178,N_4194);
and U4327 (N_4327,N_4051,N_4000);
and U4328 (N_4328,N_4128,N_4191);
nor U4329 (N_4329,N_4167,N_4068);
or U4330 (N_4330,N_4145,N_4126);
nor U4331 (N_4331,N_4094,N_4147);
nand U4332 (N_4332,N_4080,N_4042);
or U4333 (N_4333,N_4090,N_4177);
or U4334 (N_4334,N_4012,N_4025);
xor U4335 (N_4335,N_4013,N_4172);
or U4336 (N_4336,N_4049,N_4185);
or U4337 (N_4337,N_4068,N_4005);
and U4338 (N_4338,N_4110,N_4064);
xor U4339 (N_4339,N_4117,N_4091);
nand U4340 (N_4340,N_4068,N_4114);
nand U4341 (N_4341,N_4127,N_4090);
xnor U4342 (N_4342,N_4152,N_4133);
and U4343 (N_4343,N_4090,N_4182);
and U4344 (N_4344,N_4042,N_4135);
nor U4345 (N_4345,N_4172,N_4196);
nor U4346 (N_4346,N_4188,N_4093);
nor U4347 (N_4347,N_4194,N_4085);
or U4348 (N_4348,N_4092,N_4190);
nand U4349 (N_4349,N_4036,N_4074);
or U4350 (N_4350,N_4195,N_4113);
and U4351 (N_4351,N_4140,N_4092);
and U4352 (N_4352,N_4124,N_4155);
and U4353 (N_4353,N_4072,N_4036);
nand U4354 (N_4354,N_4068,N_4017);
and U4355 (N_4355,N_4021,N_4097);
nand U4356 (N_4356,N_4075,N_4016);
nor U4357 (N_4357,N_4116,N_4093);
and U4358 (N_4358,N_4031,N_4003);
and U4359 (N_4359,N_4021,N_4096);
nand U4360 (N_4360,N_4043,N_4065);
nor U4361 (N_4361,N_4190,N_4168);
and U4362 (N_4362,N_4070,N_4053);
nand U4363 (N_4363,N_4018,N_4188);
xnor U4364 (N_4364,N_4018,N_4097);
xnor U4365 (N_4365,N_4088,N_4090);
or U4366 (N_4366,N_4143,N_4179);
nor U4367 (N_4367,N_4025,N_4054);
and U4368 (N_4368,N_4062,N_4156);
or U4369 (N_4369,N_4156,N_4077);
or U4370 (N_4370,N_4030,N_4139);
and U4371 (N_4371,N_4072,N_4139);
or U4372 (N_4372,N_4175,N_4090);
or U4373 (N_4373,N_4156,N_4066);
nand U4374 (N_4374,N_4032,N_4085);
or U4375 (N_4375,N_4050,N_4164);
or U4376 (N_4376,N_4090,N_4058);
nor U4377 (N_4377,N_4165,N_4172);
nand U4378 (N_4378,N_4059,N_4136);
nand U4379 (N_4379,N_4152,N_4121);
xor U4380 (N_4380,N_4094,N_4030);
nand U4381 (N_4381,N_4172,N_4048);
or U4382 (N_4382,N_4044,N_4029);
and U4383 (N_4383,N_4040,N_4055);
and U4384 (N_4384,N_4043,N_4195);
and U4385 (N_4385,N_4003,N_4101);
and U4386 (N_4386,N_4187,N_4186);
nand U4387 (N_4387,N_4021,N_4020);
xor U4388 (N_4388,N_4117,N_4050);
or U4389 (N_4389,N_4195,N_4178);
or U4390 (N_4390,N_4139,N_4199);
xnor U4391 (N_4391,N_4171,N_4132);
nor U4392 (N_4392,N_4158,N_4060);
xnor U4393 (N_4393,N_4053,N_4058);
and U4394 (N_4394,N_4029,N_4187);
nand U4395 (N_4395,N_4161,N_4034);
nand U4396 (N_4396,N_4054,N_4140);
nor U4397 (N_4397,N_4088,N_4100);
nand U4398 (N_4398,N_4142,N_4128);
xor U4399 (N_4399,N_4004,N_4030);
nand U4400 (N_4400,N_4344,N_4255);
nor U4401 (N_4401,N_4244,N_4295);
and U4402 (N_4402,N_4383,N_4284);
nor U4403 (N_4403,N_4227,N_4260);
nand U4404 (N_4404,N_4274,N_4325);
or U4405 (N_4405,N_4297,N_4275);
nor U4406 (N_4406,N_4204,N_4206);
nor U4407 (N_4407,N_4219,N_4312);
and U4408 (N_4408,N_4245,N_4369);
and U4409 (N_4409,N_4340,N_4336);
nor U4410 (N_4410,N_4286,N_4287);
and U4411 (N_4411,N_4241,N_4350);
nand U4412 (N_4412,N_4310,N_4223);
nand U4413 (N_4413,N_4311,N_4381);
or U4414 (N_4414,N_4365,N_4377);
nand U4415 (N_4415,N_4272,N_4248);
or U4416 (N_4416,N_4228,N_4237);
or U4417 (N_4417,N_4218,N_4391);
xor U4418 (N_4418,N_4349,N_4232);
or U4419 (N_4419,N_4315,N_4304);
nand U4420 (N_4420,N_4352,N_4230);
nor U4421 (N_4421,N_4302,N_4386);
nand U4422 (N_4422,N_4210,N_4225);
xnor U4423 (N_4423,N_4351,N_4392);
nor U4424 (N_4424,N_4397,N_4374);
nand U4425 (N_4425,N_4326,N_4235);
and U4426 (N_4426,N_4247,N_4305);
or U4427 (N_4427,N_4281,N_4201);
and U4428 (N_4428,N_4298,N_4373);
nor U4429 (N_4429,N_4262,N_4273);
nor U4430 (N_4430,N_4294,N_4306);
nor U4431 (N_4431,N_4327,N_4268);
nand U4432 (N_4432,N_4379,N_4334);
and U4433 (N_4433,N_4348,N_4282);
or U4434 (N_4434,N_4243,N_4320);
and U4435 (N_4435,N_4323,N_4253);
nor U4436 (N_4436,N_4222,N_4390);
or U4437 (N_4437,N_4211,N_4238);
xor U4438 (N_4438,N_4343,N_4389);
or U4439 (N_4439,N_4317,N_4293);
nor U4440 (N_4440,N_4355,N_4321);
nand U4441 (N_4441,N_4396,N_4314);
nor U4442 (N_4442,N_4398,N_4341);
and U4443 (N_4443,N_4220,N_4263);
nor U4444 (N_4444,N_4299,N_4213);
nand U4445 (N_4445,N_4217,N_4347);
xnor U4446 (N_4446,N_4361,N_4301);
or U4447 (N_4447,N_4288,N_4333);
nand U4448 (N_4448,N_4215,N_4319);
nand U4449 (N_4449,N_4208,N_4256);
nand U4450 (N_4450,N_4261,N_4360);
and U4451 (N_4451,N_4242,N_4252);
and U4452 (N_4452,N_4205,N_4357);
nor U4453 (N_4453,N_4209,N_4318);
nor U4454 (N_4454,N_4308,N_4269);
or U4455 (N_4455,N_4279,N_4385);
nand U4456 (N_4456,N_4290,N_4307);
and U4457 (N_4457,N_4337,N_4278);
or U4458 (N_4458,N_4224,N_4353);
and U4459 (N_4459,N_4324,N_4370);
or U4460 (N_4460,N_4291,N_4200);
nand U4461 (N_4461,N_4221,N_4380);
or U4462 (N_4462,N_4345,N_4229);
or U4463 (N_4463,N_4339,N_4246);
and U4464 (N_4464,N_4388,N_4330);
or U4465 (N_4465,N_4399,N_4371);
and U4466 (N_4466,N_4378,N_4250);
nand U4467 (N_4467,N_4332,N_4322);
or U4468 (N_4468,N_4292,N_4234);
nor U4469 (N_4469,N_4366,N_4328);
and U4470 (N_4470,N_4236,N_4249);
or U4471 (N_4471,N_4214,N_4316);
nand U4472 (N_4472,N_4368,N_4203);
xor U4473 (N_4473,N_4394,N_4384);
nor U4474 (N_4474,N_4202,N_4254);
nor U4475 (N_4475,N_4367,N_4372);
or U4476 (N_4476,N_4329,N_4331);
xor U4477 (N_4477,N_4354,N_4362);
or U4478 (N_4478,N_4303,N_4342);
or U4479 (N_4479,N_4338,N_4296);
nand U4480 (N_4480,N_4257,N_4393);
nor U4481 (N_4481,N_4212,N_4364);
nor U4482 (N_4482,N_4226,N_4266);
nand U4483 (N_4483,N_4356,N_4358);
and U4484 (N_4484,N_4376,N_4277);
and U4485 (N_4485,N_4280,N_4233);
and U4486 (N_4486,N_4264,N_4346);
nand U4487 (N_4487,N_4335,N_4231);
nand U4488 (N_4488,N_4265,N_4216);
or U4489 (N_4489,N_4207,N_4309);
and U4490 (N_4490,N_4276,N_4289);
nand U4491 (N_4491,N_4240,N_4283);
xnor U4492 (N_4492,N_4387,N_4363);
or U4493 (N_4493,N_4258,N_4251);
xnor U4494 (N_4494,N_4239,N_4285);
xnor U4495 (N_4495,N_4259,N_4271);
or U4496 (N_4496,N_4267,N_4382);
nor U4497 (N_4497,N_4375,N_4313);
or U4498 (N_4498,N_4395,N_4359);
or U4499 (N_4499,N_4270,N_4300);
and U4500 (N_4500,N_4383,N_4385);
xnor U4501 (N_4501,N_4379,N_4211);
and U4502 (N_4502,N_4303,N_4244);
and U4503 (N_4503,N_4323,N_4335);
xnor U4504 (N_4504,N_4248,N_4378);
and U4505 (N_4505,N_4239,N_4312);
nand U4506 (N_4506,N_4344,N_4329);
nor U4507 (N_4507,N_4379,N_4311);
nor U4508 (N_4508,N_4373,N_4270);
nand U4509 (N_4509,N_4220,N_4242);
xnor U4510 (N_4510,N_4262,N_4347);
and U4511 (N_4511,N_4320,N_4230);
or U4512 (N_4512,N_4393,N_4377);
or U4513 (N_4513,N_4256,N_4331);
xnor U4514 (N_4514,N_4284,N_4297);
or U4515 (N_4515,N_4379,N_4326);
or U4516 (N_4516,N_4318,N_4284);
nand U4517 (N_4517,N_4343,N_4230);
and U4518 (N_4518,N_4361,N_4212);
or U4519 (N_4519,N_4376,N_4354);
nor U4520 (N_4520,N_4351,N_4317);
nor U4521 (N_4521,N_4300,N_4353);
nand U4522 (N_4522,N_4255,N_4289);
or U4523 (N_4523,N_4393,N_4235);
and U4524 (N_4524,N_4343,N_4290);
nand U4525 (N_4525,N_4294,N_4389);
nand U4526 (N_4526,N_4382,N_4343);
nor U4527 (N_4527,N_4250,N_4388);
and U4528 (N_4528,N_4311,N_4272);
or U4529 (N_4529,N_4272,N_4211);
xnor U4530 (N_4530,N_4252,N_4200);
nor U4531 (N_4531,N_4353,N_4379);
and U4532 (N_4532,N_4371,N_4392);
or U4533 (N_4533,N_4248,N_4233);
xnor U4534 (N_4534,N_4240,N_4343);
nand U4535 (N_4535,N_4321,N_4356);
or U4536 (N_4536,N_4318,N_4203);
xor U4537 (N_4537,N_4207,N_4386);
and U4538 (N_4538,N_4235,N_4289);
and U4539 (N_4539,N_4213,N_4288);
or U4540 (N_4540,N_4290,N_4366);
nor U4541 (N_4541,N_4205,N_4275);
and U4542 (N_4542,N_4373,N_4219);
nor U4543 (N_4543,N_4380,N_4379);
nand U4544 (N_4544,N_4277,N_4259);
nand U4545 (N_4545,N_4368,N_4285);
nand U4546 (N_4546,N_4392,N_4223);
xnor U4547 (N_4547,N_4390,N_4282);
nor U4548 (N_4548,N_4397,N_4301);
nand U4549 (N_4549,N_4278,N_4219);
nand U4550 (N_4550,N_4346,N_4332);
nand U4551 (N_4551,N_4345,N_4298);
and U4552 (N_4552,N_4353,N_4314);
xor U4553 (N_4553,N_4238,N_4385);
or U4554 (N_4554,N_4233,N_4311);
nand U4555 (N_4555,N_4343,N_4260);
xor U4556 (N_4556,N_4213,N_4352);
nand U4557 (N_4557,N_4368,N_4259);
nand U4558 (N_4558,N_4308,N_4282);
and U4559 (N_4559,N_4341,N_4265);
and U4560 (N_4560,N_4267,N_4353);
xnor U4561 (N_4561,N_4323,N_4281);
nor U4562 (N_4562,N_4229,N_4318);
and U4563 (N_4563,N_4293,N_4330);
xnor U4564 (N_4564,N_4352,N_4322);
nand U4565 (N_4565,N_4375,N_4246);
or U4566 (N_4566,N_4314,N_4317);
nand U4567 (N_4567,N_4345,N_4225);
and U4568 (N_4568,N_4361,N_4233);
nor U4569 (N_4569,N_4335,N_4371);
xor U4570 (N_4570,N_4226,N_4358);
and U4571 (N_4571,N_4350,N_4201);
nand U4572 (N_4572,N_4232,N_4282);
nor U4573 (N_4573,N_4268,N_4226);
nor U4574 (N_4574,N_4297,N_4238);
nand U4575 (N_4575,N_4227,N_4334);
nand U4576 (N_4576,N_4219,N_4227);
nand U4577 (N_4577,N_4322,N_4335);
or U4578 (N_4578,N_4287,N_4200);
nand U4579 (N_4579,N_4355,N_4335);
or U4580 (N_4580,N_4214,N_4374);
nor U4581 (N_4581,N_4282,N_4269);
or U4582 (N_4582,N_4207,N_4336);
nand U4583 (N_4583,N_4285,N_4321);
xor U4584 (N_4584,N_4248,N_4310);
or U4585 (N_4585,N_4250,N_4316);
or U4586 (N_4586,N_4331,N_4273);
nand U4587 (N_4587,N_4379,N_4264);
nor U4588 (N_4588,N_4354,N_4217);
and U4589 (N_4589,N_4356,N_4339);
and U4590 (N_4590,N_4325,N_4337);
or U4591 (N_4591,N_4350,N_4254);
or U4592 (N_4592,N_4294,N_4234);
and U4593 (N_4593,N_4234,N_4227);
nor U4594 (N_4594,N_4227,N_4348);
nor U4595 (N_4595,N_4329,N_4251);
and U4596 (N_4596,N_4241,N_4279);
nand U4597 (N_4597,N_4342,N_4374);
or U4598 (N_4598,N_4275,N_4329);
nor U4599 (N_4599,N_4369,N_4368);
xnor U4600 (N_4600,N_4457,N_4504);
nand U4601 (N_4601,N_4443,N_4524);
or U4602 (N_4602,N_4541,N_4573);
xnor U4603 (N_4603,N_4444,N_4461);
or U4604 (N_4604,N_4431,N_4459);
nor U4605 (N_4605,N_4403,N_4533);
xnor U4606 (N_4606,N_4463,N_4590);
nand U4607 (N_4607,N_4558,N_4577);
and U4608 (N_4608,N_4572,N_4428);
nand U4609 (N_4609,N_4451,N_4465);
nor U4610 (N_4610,N_4432,N_4409);
or U4611 (N_4611,N_4442,N_4481);
or U4612 (N_4612,N_4596,N_4496);
or U4613 (N_4613,N_4405,N_4427);
nand U4614 (N_4614,N_4540,N_4489);
and U4615 (N_4615,N_4513,N_4440);
nand U4616 (N_4616,N_4532,N_4416);
or U4617 (N_4617,N_4503,N_4450);
and U4618 (N_4618,N_4401,N_4469);
nor U4619 (N_4619,N_4482,N_4458);
or U4620 (N_4620,N_4424,N_4520);
or U4621 (N_4621,N_4527,N_4507);
nor U4622 (N_4622,N_4599,N_4486);
and U4623 (N_4623,N_4546,N_4545);
nand U4624 (N_4624,N_4437,N_4502);
or U4625 (N_4625,N_4478,N_4490);
or U4626 (N_4626,N_4452,N_4438);
or U4627 (N_4627,N_4582,N_4586);
and U4628 (N_4628,N_4563,N_4480);
or U4629 (N_4629,N_4449,N_4400);
nand U4630 (N_4630,N_4580,N_4439);
nand U4631 (N_4631,N_4499,N_4514);
and U4632 (N_4632,N_4448,N_4454);
and U4633 (N_4633,N_4517,N_4571);
nand U4634 (N_4634,N_4538,N_4484);
nor U4635 (N_4635,N_4512,N_4595);
nand U4636 (N_4636,N_4570,N_4589);
nand U4637 (N_4637,N_4548,N_4472);
nand U4638 (N_4638,N_4565,N_4414);
nor U4639 (N_4639,N_4544,N_4417);
and U4640 (N_4640,N_4526,N_4568);
and U4641 (N_4641,N_4597,N_4415);
nor U4642 (N_4642,N_4521,N_4581);
nand U4643 (N_4643,N_4483,N_4466);
or U4644 (N_4644,N_4473,N_4456);
nor U4645 (N_4645,N_4475,N_4598);
nor U4646 (N_4646,N_4435,N_4426);
nand U4647 (N_4647,N_4476,N_4536);
and U4648 (N_4648,N_4460,N_4560);
nand U4649 (N_4649,N_4575,N_4569);
and U4650 (N_4650,N_4594,N_4567);
nor U4651 (N_4651,N_4584,N_4433);
or U4652 (N_4652,N_4539,N_4430);
nand U4653 (N_4653,N_4578,N_4407);
or U4654 (N_4654,N_4420,N_4550);
or U4655 (N_4655,N_4593,N_4501);
nand U4656 (N_4656,N_4508,N_4566);
nor U4657 (N_4657,N_4564,N_4553);
nor U4658 (N_4658,N_4525,N_4406);
and U4659 (N_4659,N_4434,N_4576);
or U4660 (N_4660,N_4562,N_4492);
and U4661 (N_4661,N_4474,N_4516);
and U4662 (N_4662,N_4422,N_4529);
and U4663 (N_4663,N_4429,N_4537);
or U4664 (N_4664,N_4445,N_4531);
or U4665 (N_4665,N_4518,N_4488);
nand U4666 (N_4666,N_4411,N_4418);
or U4667 (N_4667,N_4535,N_4561);
or U4668 (N_4668,N_4446,N_4425);
nor U4669 (N_4669,N_4477,N_4485);
or U4670 (N_4670,N_4505,N_4498);
or U4671 (N_4671,N_4467,N_4423);
nor U4672 (N_4672,N_4464,N_4519);
or U4673 (N_4673,N_4579,N_4412);
and U4674 (N_4674,N_4413,N_4402);
and U4675 (N_4675,N_4410,N_4551);
nor U4676 (N_4676,N_4543,N_4455);
nor U4677 (N_4677,N_4497,N_4471);
or U4678 (N_4678,N_4556,N_4549);
or U4679 (N_4679,N_4419,N_4441);
or U4680 (N_4680,N_4495,N_4404);
nand U4681 (N_4681,N_4534,N_4592);
nor U4682 (N_4682,N_4528,N_4557);
nand U4683 (N_4683,N_4506,N_4530);
and U4684 (N_4684,N_4554,N_4447);
nor U4685 (N_4685,N_4587,N_4591);
nor U4686 (N_4686,N_4523,N_4555);
nand U4687 (N_4687,N_4583,N_4552);
nor U4688 (N_4688,N_4510,N_4585);
and U4689 (N_4689,N_4494,N_4493);
and U4690 (N_4690,N_4559,N_4574);
and U4691 (N_4691,N_4547,N_4479);
or U4692 (N_4692,N_4509,N_4453);
and U4693 (N_4693,N_4470,N_4542);
nand U4694 (N_4694,N_4491,N_4408);
nor U4695 (N_4695,N_4511,N_4462);
nand U4696 (N_4696,N_4522,N_4487);
nand U4697 (N_4697,N_4468,N_4421);
nand U4698 (N_4698,N_4500,N_4588);
xnor U4699 (N_4699,N_4436,N_4515);
nor U4700 (N_4700,N_4576,N_4544);
nand U4701 (N_4701,N_4517,N_4404);
and U4702 (N_4702,N_4449,N_4458);
nor U4703 (N_4703,N_4554,N_4459);
xnor U4704 (N_4704,N_4409,N_4473);
and U4705 (N_4705,N_4475,N_4448);
and U4706 (N_4706,N_4418,N_4443);
or U4707 (N_4707,N_4515,N_4407);
nor U4708 (N_4708,N_4498,N_4510);
nor U4709 (N_4709,N_4410,N_4434);
and U4710 (N_4710,N_4437,N_4558);
and U4711 (N_4711,N_4556,N_4528);
or U4712 (N_4712,N_4458,N_4440);
nand U4713 (N_4713,N_4433,N_4535);
nor U4714 (N_4714,N_4558,N_4485);
nand U4715 (N_4715,N_4569,N_4561);
or U4716 (N_4716,N_4454,N_4561);
xor U4717 (N_4717,N_4425,N_4535);
nand U4718 (N_4718,N_4401,N_4438);
nand U4719 (N_4719,N_4448,N_4509);
or U4720 (N_4720,N_4542,N_4458);
nand U4721 (N_4721,N_4441,N_4456);
nand U4722 (N_4722,N_4520,N_4501);
or U4723 (N_4723,N_4599,N_4407);
nor U4724 (N_4724,N_4403,N_4564);
xor U4725 (N_4725,N_4424,N_4409);
nand U4726 (N_4726,N_4441,N_4559);
or U4727 (N_4727,N_4532,N_4588);
and U4728 (N_4728,N_4446,N_4555);
nand U4729 (N_4729,N_4510,N_4469);
and U4730 (N_4730,N_4424,N_4437);
or U4731 (N_4731,N_4594,N_4482);
or U4732 (N_4732,N_4476,N_4597);
or U4733 (N_4733,N_4437,N_4512);
nor U4734 (N_4734,N_4524,N_4481);
or U4735 (N_4735,N_4559,N_4434);
nor U4736 (N_4736,N_4519,N_4448);
and U4737 (N_4737,N_4476,N_4492);
nand U4738 (N_4738,N_4569,N_4596);
and U4739 (N_4739,N_4489,N_4599);
nor U4740 (N_4740,N_4450,N_4546);
nor U4741 (N_4741,N_4571,N_4405);
nand U4742 (N_4742,N_4427,N_4506);
xnor U4743 (N_4743,N_4418,N_4438);
nand U4744 (N_4744,N_4478,N_4423);
or U4745 (N_4745,N_4595,N_4559);
and U4746 (N_4746,N_4512,N_4557);
nor U4747 (N_4747,N_4411,N_4417);
or U4748 (N_4748,N_4544,N_4475);
or U4749 (N_4749,N_4427,N_4500);
nor U4750 (N_4750,N_4575,N_4531);
nand U4751 (N_4751,N_4582,N_4412);
nor U4752 (N_4752,N_4473,N_4526);
nand U4753 (N_4753,N_4591,N_4409);
nor U4754 (N_4754,N_4485,N_4434);
and U4755 (N_4755,N_4460,N_4583);
nand U4756 (N_4756,N_4413,N_4407);
or U4757 (N_4757,N_4581,N_4445);
and U4758 (N_4758,N_4539,N_4412);
or U4759 (N_4759,N_4535,N_4565);
or U4760 (N_4760,N_4552,N_4500);
xor U4761 (N_4761,N_4515,N_4443);
and U4762 (N_4762,N_4584,N_4437);
and U4763 (N_4763,N_4542,N_4430);
nor U4764 (N_4764,N_4587,N_4446);
nor U4765 (N_4765,N_4533,N_4423);
and U4766 (N_4766,N_4452,N_4596);
or U4767 (N_4767,N_4432,N_4470);
nor U4768 (N_4768,N_4509,N_4450);
nor U4769 (N_4769,N_4419,N_4434);
and U4770 (N_4770,N_4499,N_4488);
and U4771 (N_4771,N_4526,N_4405);
and U4772 (N_4772,N_4449,N_4594);
nor U4773 (N_4773,N_4427,N_4448);
or U4774 (N_4774,N_4592,N_4597);
nor U4775 (N_4775,N_4498,N_4453);
and U4776 (N_4776,N_4443,N_4444);
or U4777 (N_4777,N_4432,N_4591);
and U4778 (N_4778,N_4409,N_4406);
nor U4779 (N_4779,N_4588,N_4558);
nor U4780 (N_4780,N_4574,N_4468);
and U4781 (N_4781,N_4534,N_4573);
nand U4782 (N_4782,N_4436,N_4594);
xnor U4783 (N_4783,N_4572,N_4449);
xnor U4784 (N_4784,N_4423,N_4449);
and U4785 (N_4785,N_4404,N_4568);
and U4786 (N_4786,N_4469,N_4543);
nand U4787 (N_4787,N_4504,N_4409);
and U4788 (N_4788,N_4588,N_4466);
nor U4789 (N_4789,N_4486,N_4592);
nand U4790 (N_4790,N_4412,N_4416);
and U4791 (N_4791,N_4539,N_4477);
xnor U4792 (N_4792,N_4479,N_4487);
nor U4793 (N_4793,N_4498,N_4590);
nand U4794 (N_4794,N_4527,N_4439);
and U4795 (N_4795,N_4543,N_4548);
or U4796 (N_4796,N_4489,N_4454);
nand U4797 (N_4797,N_4440,N_4454);
nand U4798 (N_4798,N_4556,N_4553);
nand U4799 (N_4799,N_4506,N_4595);
nor U4800 (N_4800,N_4775,N_4646);
and U4801 (N_4801,N_4656,N_4625);
nor U4802 (N_4802,N_4796,N_4769);
nand U4803 (N_4803,N_4603,N_4719);
nor U4804 (N_4804,N_4676,N_4721);
nand U4805 (N_4805,N_4633,N_4681);
nand U4806 (N_4806,N_4629,N_4668);
or U4807 (N_4807,N_4732,N_4774);
nor U4808 (N_4808,N_4683,N_4688);
nor U4809 (N_4809,N_4628,N_4636);
nand U4810 (N_4810,N_4694,N_4632);
nor U4811 (N_4811,N_4674,N_4794);
nor U4812 (N_4812,N_4720,N_4704);
nor U4813 (N_4813,N_4652,N_4756);
nor U4814 (N_4814,N_4711,N_4621);
nand U4815 (N_4815,N_4785,N_4710);
and U4816 (N_4816,N_4789,N_4650);
or U4817 (N_4817,N_4618,N_4699);
or U4818 (N_4818,N_4703,N_4738);
nand U4819 (N_4819,N_4783,N_4600);
and U4820 (N_4820,N_4761,N_4651);
or U4821 (N_4821,N_4616,N_4714);
nor U4822 (N_4822,N_4638,N_4729);
nor U4823 (N_4823,N_4716,N_4731);
nor U4824 (N_4824,N_4645,N_4673);
nand U4825 (N_4825,N_4626,N_4709);
nand U4826 (N_4826,N_4772,N_4725);
and U4827 (N_4827,N_4665,N_4671);
nand U4828 (N_4828,N_4701,N_4670);
and U4829 (N_4829,N_4798,N_4792);
nor U4830 (N_4830,N_4733,N_4678);
or U4831 (N_4831,N_4797,N_4755);
or U4832 (N_4832,N_4782,N_4640);
nor U4833 (N_4833,N_4610,N_4682);
or U4834 (N_4834,N_4687,N_4727);
nor U4835 (N_4835,N_4757,N_4690);
or U4836 (N_4836,N_4728,N_4614);
nor U4837 (N_4837,N_4759,N_4740);
and U4838 (N_4838,N_4648,N_4644);
nand U4839 (N_4839,N_4639,N_4748);
or U4840 (N_4840,N_4620,N_4679);
nor U4841 (N_4841,N_4619,N_4770);
nand U4842 (N_4842,N_4764,N_4696);
nand U4843 (N_4843,N_4601,N_4784);
xnor U4844 (N_4844,N_4744,N_4691);
nor U4845 (N_4845,N_4698,N_4641);
nand U4846 (N_4846,N_4649,N_4780);
or U4847 (N_4847,N_4717,N_4654);
nand U4848 (N_4848,N_4659,N_4745);
and U4849 (N_4849,N_4675,N_4669);
or U4850 (N_4850,N_4612,N_4667);
or U4851 (N_4851,N_4773,N_4602);
xor U4852 (N_4852,N_4655,N_4760);
and U4853 (N_4853,N_4767,N_4634);
nand U4854 (N_4854,N_4677,N_4741);
and U4855 (N_4855,N_4781,N_4666);
nor U4856 (N_4856,N_4707,N_4622);
and U4857 (N_4857,N_4635,N_4611);
nand U4858 (N_4858,N_4700,N_4723);
nand U4859 (N_4859,N_4607,N_4623);
nor U4860 (N_4860,N_4786,N_4697);
nand U4861 (N_4861,N_4609,N_4795);
xnor U4862 (N_4862,N_4705,N_4712);
or U4863 (N_4863,N_4793,N_4630);
or U4864 (N_4864,N_4742,N_4647);
nor U4865 (N_4865,N_4658,N_4758);
xnor U4866 (N_4866,N_4657,N_4715);
or U4867 (N_4867,N_4664,N_4799);
or U4868 (N_4868,N_4737,N_4627);
xnor U4869 (N_4869,N_4777,N_4750);
nor U4870 (N_4870,N_4771,N_4663);
nor U4871 (N_4871,N_4672,N_4615);
and U4872 (N_4872,N_4779,N_4722);
nor U4873 (N_4873,N_4662,N_4692);
nor U4874 (N_4874,N_4787,N_4718);
nor U4875 (N_4875,N_4753,N_4752);
and U4876 (N_4876,N_4790,N_4685);
or U4877 (N_4877,N_4739,N_4735);
nand U4878 (N_4878,N_4788,N_4680);
and U4879 (N_4879,N_4693,N_4746);
nand U4880 (N_4880,N_4736,N_4762);
nand U4881 (N_4881,N_4624,N_4751);
or U4882 (N_4882,N_4747,N_4754);
nand U4883 (N_4883,N_4734,N_4708);
nor U4884 (N_4884,N_4684,N_4695);
xnor U4885 (N_4885,N_4749,N_4766);
xnor U4886 (N_4886,N_4776,N_4608);
and U4887 (N_4887,N_4778,N_4653);
nor U4888 (N_4888,N_4637,N_4613);
nand U4889 (N_4889,N_4660,N_4791);
nand U4890 (N_4890,N_4730,N_4702);
nor U4891 (N_4891,N_4689,N_4768);
nand U4892 (N_4892,N_4606,N_4604);
and U4893 (N_4893,N_4661,N_4706);
nand U4894 (N_4894,N_4724,N_4765);
nand U4895 (N_4895,N_4631,N_4726);
nor U4896 (N_4896,N_4743,N_4617);
and U4897 (N_4897,N_4605,N_4643);
and U4898 (N_4898,N_4713,N_4763);
or U4899 (N_4899,N_4642,N_4686);
or U4900 (N_4900,N_4768,N_4692);
nor U4901 (N_4901,N_4658,N_4636);
nand U4902 (N_4902,N_4627,N_4751);
and U4903 (N_4903,N_4693,N_4689);
nand U4904 (N_4904,N_4689,N_4730);
nor U4905 (N_4905,N_4671,N_4645);
and U4906 (N_4906,N_4740,N_4755);
and U4907 (N_4907,N_4741,N_4638);
nand U4908 (N_4908,N_4708,N_4755);
nor U4909 (N_4909,N_4756,N_4767);
nor U4910 (N_4910,N_4623,N_4771);
nor U4911 (N_4911,N_4653,N_4775);
or U4912 (N_4912,N_4740,N_4745);
and U4913 (N_4913,N_4796,N_4628);
xnor U4914 (N_4914,N_4615,N_4636);
nor U4915 (N_4915,N_4784,N_4788);
nor U4916 (N_4916,N_4796,N_4746);
or U4917 (N_4917,N_4684,N_4673);
and U4918 (N_4918,N_4691,N_4791);
nor U4919 (N_4919,N_4709,N_4780);
and U4920 (N_4920,N_4645,N_4688);
nor U4921 (N_4921,N_4645,N_4664);
xnor U4922 (N_4922,N_4697,N_4793);
or U4923 (N_4923,N_4642,N_4755);
nand U4924 (N_4924,N_4787,N_4606);
nand U4925 (N_4925,N_4717,N_4789);
nand U4926 (N_4926,N_4657,N_4633);
nand U4927 (N_4927,N_4734,N_4739);
and U4928 (N_4928,N_4619,N_4640);
and U4929 (N_4929,N_4662,N_4614);
or U4930 (N_4930,N_4720,N_4609);
xor U4931 (N_4931,N_4752,N_4623);
and U4932 (N_4932,N_4773,N_4740);
nor U4933 (N_4933,N_4708,N_4645);
nand U4934 (N_4934,N_4648,N_4658);
or U4935 (N_4935,N_4649,N_4631);
or U4936 (N_4936,N_4623,N_4754);
or U4937 (N_4937,N_4693,N_4695);
nand U4938 (N_4938,N_4698,N_4694);
xnor U4939 (N_4939,N_4741,N_4622);
xor U4940 (N_4940,N_4775,N_4776);
and U4941 (N_4941,N_4758,N_4702);
and U4942 (N_4942,N_4735,N_4605);
and U4943 (N_4943,N_4615,N_4789);
nand U4944 (N_4944,N_4626,N_4764);
nand U4945 (N_4945,N_4679,N_4610);
and U4946 (N_4946,N_4741,N_4791);
nand U4947 (N_4947,N_4653,N_4691);
nor U4948 (N_4948,N_4645,N_4750);
nand U4949 (N_4949,N_4764,N_4608);
and U4950 (N_4950,N_4640,N_4731);
nand U4951 (N_4951,N_4772,N_4768);
and U4952 (N_4952,N_4613,N_4646);
nor U4953 (N_4953,N_4728,N_4754);
and U4954 (N_4954,N_4754,N_4634);
or U4955 (N_4955,N_4743,N_4741);
nor U4956 (N_4956,N_4660,N_4614);
and U4957 (N_4957,N_4780,N_4745);
and U4958 (N_4958,N_4787,N_4635);
and U4959 (N_4959,N_4725,N_4717);
and U4960 (N_4960,N_4665,N_4681);
or U4961 (N_4961,N_4643,N_4707);
nor U4962 (N_4962,N_4745,N_4638);
nand U4963 (N_4963,N_4741,N_4600);
nand U4964 (N_4964,N_4656,N_4655);
xor U4965 (N_4965,N_4752,N_4777);
xnor U4966 (N_4966,N_4699,N_4774);
nand U4967 (N_4967,N_4683,N_4763);
or U4968 (N_4968,N_4626,N_4608);
nor U4969 (N_4969,N_4790,N_4731);
nor U4970 (N_4970,N_4665,N_4784);
xor U4971 (N_4971,N_4756,N_4783);
and U4972 (N_4972,N_4629,N_4655);
xnor U4973 (N_4973,N_4712,N_4620);
nor U4974 (N_4974,N_4679,N_4703);
nor U4975 (N_4975,N_4735,N_4673);
nor U4976 (N_4976,N_4620,N_4686);
or U4977 (N_4977,N_4727,N_4604);
nor U4978 (N_4978,N_4624,N_4775);
nor U4979 (N_4979,N_4694,N_4710);
nor U4980 (N_4980,N_4752,N_4712);
and U4981 (N_4981,N_4694,N_4739);
nor U4982 (N_4982,N_4658,N_4727);
nand U4983 (N_4983,N_4782,N_4692);
or U4984 (N_4984,N_4625,N_4658);
and U4985 (N_4985,N_4721,N_4640);
or U4986 (N_4986,N_4659,N_4737);
nor U4987 (N_4987,N_4699,N_4629);
or U4988 (N_4988,N_4742,N_4609);
nand U4989 (N_4989,N_4753,N_4725);
and U4990 (N_4990,N_4778,N_4708);
nand U4991 (N_4991,N_4623,N_4618);
and U4992 (N_4992,N_4694,N_4633);
nor U4993 (N_4993,N_4763,N_4735);
or U4994 (N_4994,N_4766,N_4720);
nor U4995 (N_4995,N_4776,N_4664);
nand U4996 (N_4996,N_4609,N_4743);
xor U4997 (N_4997,N_4691,N_4606);
and U4998 (N_4998,N_4720,N_4761);
nand U4999 (N_4999,N_4766,N_4689);
nand U5000 (N_5000,N_4819,N_4980);
or U5001 (N_5001,N_4909,N_4908);
and U5002 (N_5002,N_4846,N_4964);
and U5003 (N_5003,N_4917,N_4905);
xor U5004 (N_5004,N_4997,N_4887);
or U5005 (N_5005,N_4985,N_4962);
nand U5006 (N_5006,N_4914,N_4898);
or U5007 (N_5007,N_4952,N_4933);
or U5008 (N_5008,N_4948,N_4988);
nor U5009 (N_5009,N_4994,N_4950);
or U5010 (N_5010,N_4832,N_4989);
xor U5011 (N_5011,N_4886,N_4899);
nor U5012 (N_5012,N_4836,N_4961);
nor U5013 (N_5013,N_4927,N_4968);
or U5014 (N_5014,N_4834,N_4839);
nand U5015 (N_5015,N_4926,N_4871);
and U5016 (N_5016,N_4910,N_4995);
nor U5017 (N_5017,N_4855,N_4872);
xor U5018 (N_5018,N_4823,N_4960);
nor U5019 (N_5019,N_4802,N_4957);
or U5020 (N_5020,N_4857,N_4975);
or U5021 (N_5021,N_4935,N_4977);
or U5022 (N_5022,N_4825,N_4953);
and U5023 (N_5023,N_4884,N_4804);
or U5024 (N_5024,N_4851,N_4915);
nand U5025 (N_5025,N_4841,N_4937);
and U5026 (N_5026,N_4902,N_4840);
nor U5027 (N_5027,N_4852,N_4998);
nand U5028 (N_5028,N_4850,N_4882);
and U5029 (N_5029,N_4976,N_4959);
and U5030 (N_5030,N_4885,N_4981);
nor U5031 (N_5031,N_4907,N_4932);
and U5032 (N_5032,N_4939,N_4889);
nand U5033 (N_5033,N_4845,N_4904);
or U5034 (N_5034,N_4966,N_4826);
and U5035 (N_5035,N_4983,N_4955);
and U5036 (N_5036,N_4859,N_4807);
xor U5037 (N_5037,N_4811,N_4869);
or U5038 (N_5038,N_4925,N_4970);
and U5039 (N_5039,N_4987,N_4991);
nor U5040 (N_5040,N_4891,N_4813);
or U5041 (N_5041,N_4992,N_4901);
and U5042 (N_5042,N_4814,N_4809);
nor U5043 (N_5043,N_4912,N_4883);
nand U5044 (N_5044,N_4996,N_4803);
nor U5045 (N_5045,N_4956,N_4878);
nor U5046 (N_5046,N_4880,N_4843);
nand U5047 (N_5047,N_4861,N_4801);
and U5048 (N_5048,N_4892,N_4879);
or U5049 (N_5049,N_4913,N_4875);
and U5050 (N_5050,N_4903,N_4900);
nand U5051 (N_5051,N_4916,N_4863);
or U5052 (N_5052,N_4958,N_4800);
xor U5053 (N_5053,N_4810,N_4924);
and U5054 (N_5054,N_4931,N_4829);
or U5055 (N_5055,N_4947,N_4963);
nand U5056 (N_5056,N_4854,N_4816);
nand U5057 (N_5057,N_4929,N_4835);
nand U5058 (N_5058,N_4822,N_4848);
nor U5059 (N_5059,N_4860,N_4856);
xnor U5060 (N_5060,N_4847,N_4999);
nor U5061 (N_5061,N_4941,N_4918);
and U5062 (N_5062,N_4921,N_4844);
nor U5063 (N_5063,N_4853,N_4969);
nor U5064 (N_5064,N_4971,N_4945);
xnor U5065 (N_5065,N_4833,N_4895);
nor U5066 (N_5066,N_4866,N_4812);
and U5067 (N_5067,N_4808,N_4943);
xnor U5068 (N_5068,N_4894,N_4837);
or U5069 (N_5069,N_4893,N_4862);
or U5070 (N_5070,N_4890,N_4936);
nand U5071 (N_5071,N_4940,N_4865);
or U5072 (N_5072,N_4965,N_4928);
or U5073 (N_5073,N_4946,N_4831);
and U5074 (N_5074,N_4842,N_4984);
or U5075 (N_5075,N_4906,N_4858);
and U5076 (N_5076,N_4828,N_4818);
or U5077 (N_5077,N_4838,N_4954);
nor U5078 (N_5078,N_4942,N_4874);
or U5079 (N_5079,N_4923,N_4806);
or U5080 (N_5080,N_4888,N_4972);
xnor U5081 (N_5081,N_4911,N_4870);
nand U5082 (N_5082,N_4876,N_4993);
nor U5083 (N_5083,N_4821,N_4944);
and U5084 (N_5084,N_4881,N_4978);
nand U5085 (N_5085,N_4979,N_4986);
and U5086 (N_5086,N_4949,N_4951);
nand U5087 (N_5087,N_4930,N_4805);
nand U5088 (N_5088,N_4849,N_4934);
nor U5089 (N_5089,N_4896,N_4830);
and U5090 (N_5090,N_4920,N_4967);
xor U5091 (N_5091,N_4877,N_4867);
nand U5092 (N_5092,N_4873,N_4824);
or U5093 (N_5093,N_4974,N_4938);
nand U5094 (N_5094,N_4820,N_4922);
nand U5095 (N_5095,N_4897,N_4868);
xnor U5096 (N_5096,N_4919,N_4815);
and U5097 (N_5097,N_4864,N_4990);
and U5098 (N_5098,N_4982,N_4817);
or U5099 (N_5099,N_4973,N_4827);
nor U5100 (N_5100,N_4802,N_4907);
nor U5101 (N_5101,N_4839,N_4852);
nand U5102 (N_5102,N_4938,N_4885);
nand U5103 (N_5103,N_4835,N_4897);
and U5104 (N_5104,N_4818,N_4883);
or U5105 (N_5105,N_4941,N_4924);
and U5106 (N_5106,N_4846,N_4824);
nor U5107 (N_5107,N_4835,N_4914);
nand U5108 (N_5108,N_4908,N_4989);
and U5109 (N_5109,N_4871,N_4916);
and U5110 (N_5110,N_4921,N_4878);
nand U5111 (N_5111,N_4817,N_4954);
nor U5112 (N_5112,N_4900,N_4969);
xnor U5113 (N_5113,N_4830,N_4822);
nand U5114 (N_5114,N_4851,N_4914);
or U5115 (N_5115,N_4824,N_4950);
or U5116 (N_5116,N_4974,N_4887);
nor U5117 (N_5117,N_4809,N_4920);
nor U5118 (N_5118,N_4944,N_4903);
nor U5119 (N_5119,N_4900,N_4909);
nand U5120 (N_5120,N_4980,N_4806);
nor U5121 (N_5121,N_4861,N_4988);
and U5122 (N_5122,N_4962,N_4990);
and U5123 (N_5123,N_4852,N_4833);
nand U5124 (N_5124,N_4942,N_4928);
nor U5125 (N_5125,N_4894,N_4817);
nand U5126 (N_5126,N_4820,N_4983);
and U5127 (N_5127,N_4816,N_4835);
nand U5128 (N_5128,N_4964,N_4957);
xnor U5129 (N_5129,N_4991,N_4989);
and U5130 (N_5130,N_4935,N_4850);
nor U5131 (N_5131,N_4845,N_4825);
xor U5132 (N_5132,N_4968,N_4950);
nor U5133 (N_5133,N_4809,N_4834);
and U5134 (N_5134,N_4997,N_4940);
nor U5135 (N_5135,N_4923,N_4817);
and U5136 (N_5136,N_4938,N_4936);
and U5137 (N_5137,N_4902,N_4877);
nor U5138 (N_5138,N_4961,N_4984);
xnor U5139 (N_5139,N_4942,N_4840);
nand U5140 (N_5140,N_4898,N_4888);
or U5141 (N_5141,N_4952,N_4804);
or U5142 (N_5142,N_4988,N_4884);
and U5143 (N_5143,N_4987,N_4957);
nor U5144 (N_5144,N_4889,N_4881);
or U5145 (N_5145,N_4888,N_4821);
nor U5146 (N_5146,N_4961,N_4987);
nor U5147 (N_5147,N_4924,N_4866);
nor U5148 (N_5148,N_4968,N_4813);
and U5149 (N_5149,N_4910,N_4874);
or U5150 (N_5150,N_4962,N_4941);
nand U5151 (N_5151,N_4817,N_4951);
nand U5152 (N_5152,N_4856,N_4991);
nor U5153 (N_5153,N_4858,N_4938);
and U5154 (N_5154,N_4996,N_4986);
and U5155 (N_5155,N_4841,N_4910);
nor U5156 (N_5156,N_4948,N_4834);
xor U5157 (N_5157,N_4815,N_4964);
or U5158 (N_5158,N_4864,N_4981);
nand U5159 (N_5159,N_4967,N_4851);
and U5160 (N_5160,N_4944,N_4967);
and U5161 (N_5161,N_4850,N_4886);
and U5162 (N_5162,N_4916,N_4885);
and U5163 (N_5163,N_4897,N_4896);
nand U5164 (N_5164,N_4978,N_4970);
nand U5165 (N_5165,N_4965,N_4903);
or U5166 (N_5166,N_4908,N_4821);
and U5167 (N_5167,N_4837,N_4876);
nor U5168 (N_5168,N_4940,N_4993);
or U5169 (N_5169,N_4894,N_4908);
nand U5170 (N_5170,N_4977,N_4872);
or U5171 (N_5171,N_4866,N_4842);
nor U5172 (N_5172,N_4867,N_4940);
nand U5173 (N_5173,N_4985,N_4958);
nand U5174 (N_5174,N_4838,N_4858);
nand U5175 (N_5175,N_4958,N_4878);
nand U5176 (N_5176,N_4810,N_4973);
nor U5177 (N_5177,N_4929,N_4910);
nand U5178 (N_5178,N_4908,N_4907);
nor U5179 (N_5179,N_4881,N_4819);
nor U5180 (N_5180,N_4851,N_4951);
nand U5181 (N_5181,N_4995,N_4895);
xnor U5182 (N_5182,N_4806,N_4905);
and U5183 (N_5183,N_4910,N_4898);
and U5184 (N_5184,N_4825,N_4977);
nor U5185 (N_5185,N_4924,N_4846);
or U5186 (N_5186,N_4949,N_4880);
and U5187 (N_5187,N_4962,N_4824);
nor U5188 (N_5188,N_4994,N_4872);
and U5189 (N_5189,N_4842,N_4805);
and U5190 (N_5190,N_4983,N_4999);
or U5191 (N_5191,N_4963,N_4908);
nor U5192 (N_5192,N_4828,N_4817);
nand U5193 (N_5193,N_4820,N_4842);
nand U5194 (N_5194,N_4976,N_4905);
nand U5195 (N_5195,N_4965,N_4950);
and U5196 (N_5196,N_4856,N_4931);
nand U5197 (N_5197,N_4979,N_4878);
and U5198 (N_5198,N_4966,N_4927);
or U5199 (N_5199,N_4812,N_4985);
nand U5200 (N_5200,N_5158,N_5079);
nand U5201 (N_5201,N_5071,N_5074);
nand U5202 (N_5202,N_5017,N_5015);
or U5203 (N_5203,N_5160,N_5039);
or U5204 (N_5204,N_5075,N_5181);
or U5205 (N_5205,N_5185,N_5061);
and U5206 (N_5206,N_5032,N_5146);
or U5207 (N_5207,N_5053,N_5166);
or U5208 (N_5208,N_5093,N_5036);
and U5209 (N_5209,N_5000,N_5101);
or U5210 (N_5210,N_5151,N_5111);
nand U5211 (N_5211,N_5072,N_5004);
or U5212 (N_5212,N_5112,N_5139);
nor U5213 (N_5213,N_5148,N_5047);
xnor U5214 (N_5214,N_5197,N_5001);
nor U5215 (N_5215,N_5083,N_5069);
and U5216 (N_5216,N_5184,N_5175);
nor U5217 (N_5217,N_5159,N_5052);
xnor U5218 (N_5218,N_5059,N_5022);
nor U5219 (N_5219,N_5009,N_5028);
nor U5220 (N_5220,N_5149,N_5014);
nor U5221 (N_5221,N_5085,N_5051);
nand U5222 (N_5222,N_5187,N_5066);
or U5223 (N_5223,N_5141,N_5023);
and U5224 (N_5224,N_5043,N_5049);
nand U5225 (N_5225,N_5068,N_5048);
or U5226 (N_5226,N_5137,N_5124);
nor U5227 (N_5227,N_5100,N_5161);
nor U5228 (N_5228,N_5103,N_5174);
nor U5229 (N_5229,N_5044,N_5163);
and U5230 (N_5230,N_5190,N_5132);
or U5231 (N_5231,N_5038,N_5167);
nor U5232 (N_5232,N_5042,N_5171);
and U5233 (N_5233,N_5145,N_5087);
nand U5234 (N_5234,N_5193,N_5196);
nand U5235 (N_5235,N_5129,N_5063);
nand U5236 (N_5236,N_5011,N_5198);
or U5237 (N_5237,N_5055,N_5126);
and U5238 (N_5238,N_5091,N_5156);
and U5239 (N_5239,N_5188,N_5192);
nand U5240 (N_5240,N_5114,N_5153);
and U5241 (N_5241,N_5154,N_5115);
nor U5242 (N_5242,N_5064,N_5155);
and U5243 (N_5243,N_5019,N_5084);
nand U5244 (N_5244,N_5172,N_5130);
or U5245 (N_5245,N_5096,N_5033);
and U5246 (N_5246,N_5116,N_5040);
or U5247 (N_5247,N_5121,N_5058);
or U5248 (N_5248,N_5106,N_5109);
xor U5249 (N_5249,N_5199,N_5041);
and U5250 (N_5250,N_5170,N_5177);
and U5251 (N_5251,N_5088,N_5095);
nand U5252 (N_5252,N_5090,N_5108);
nor U5253 (N_5253,N_5162,N_5179);
xnor U5254 (N_5254,N_5113,N_5086);
nor U5255 (N_5255,N_5018,N_5152);
nand U5256 (N_5256,N_5120,N_5133);
and U5257 (N_5257,N_5056,N_5094);
xnor U5258 (N_5258,N_5135,N_5008);
nand U5259 (N_5259,N_5080,N_5082);
nor U5260 (N_5260,N_5076,N_5123);
or U5261 (N_5261,N_5147,N_5165);
or U5262 (N_5262,N_5183,N_5186);
nand U5263 (N_5263,N_5157,N_5099);
nor U5264 (N_5264,N_5143,N_5136);
xor U5265 (N_5265,N_5013,N_5125);
nor U5266 (N_5266,N_5150,N_5025);
nand U5267 (N_5267,N_5104,N_5142);
or U5268 (N_5268,N_5168,N_5078);
and U5269 (N_5269,N_5119,N_5169);
nor U5270 (N_5270,N_5012,N_5131);
or U5271 (N_5271,N_5105,N_5073);
and U5272 (N_5272,N_5081,N_5070);
nor U5273 (N_5273,N_5098,N_5128);
and U5274 (N_5274,N_5046,N_5002);
nor U5275 (N_5275,N_5178,N_5127);
or U5276 (N_5276,N_5020,N_5117);
nand U5277 (N_5277,N_5173,N_5024);
and U5278 (N_5278,N_5191,N_5180);
nor U5279 (N_5279,N_5050,N_5035);
nor U5280 (N_5280,N_5176,N_5060);
and U5281 (N_5281,N_5065,N_5097);
nor U5282 (N_5282,N_5189,N_5031);
nor U5283 (N_5283,N_5110,N_5107);
nand U5284 (N_5284,N_5138,N_5037);
or U5285 (N_5285,N_5164,N_5030);
nand U5286 (N_5286,N_5034,N_5054);
xnor U5287 (N_5287,N_5144,N_5194);
nor U5288 (N_5288,N_5182,N_5006);
nor U5289 (N_5289,N_5005,N_5122);
nand U5290 (N_5290,N_5016,N_5062);
or U5291 (N_5291,N_5118,N_5007);
and U5292 (N_5292,N_5045,N_5089);
and U5293 (N_5293,N_5067,N_5134);
and U5294 (N_5294,N_5010,N_5092);
nor U5295 (N_5295,N_5027,N_5003);
and U5296 (N_5296,N_5140,N_5102);
nor U5297 (N_5297,N_5195,N_5057);
nor U5298 (N_5298,N_5077,N_5021);
xnor U5299 (N_5299,N_5029,N_5026);
nor U5300 (N_5300,N_5026,N_5100);
nand U5301 (N_5301,N_5162,N_5083);
nor U5302 (N_5302,N_5071,N_5143);
nand U5303 (N_5303,N_5035,N_5024);
and U5304 (N_5304,N_5013,N_5051);
and U5305 (N_5305,N_5164,N_5097);
and U5306 (N_5306,N_5006,N_5164);
nor U5307 (N_5307,N_5179,N_5175);
nor U5308 (N_5308,N_5147,N_5011);
or U5309 (N_5309,N_5009,N_5145);
and U5310 (N_5310,N_5186,N_5173);
nor U5311 (N_5311,N_5017,N_5042);
nor U5312 (N_5312,N_5005,N_5091);
xor U5313 (N_5313,N_5182,N_5107);
and U5314 (N_5314,N_5136,N_5048);
and U5315 (N_5315,N_5165,N_5117);
nor U5316 (N_5316,N_5164,N_5142);
xnor U5317 (N_5317,N_5076,N_5053);
or U5318 (N_5318,N_5186,N_5160);
nor U5319 (N_5319,N_5050,N_5107);
nor U5320 (N_5320,N_5027,N_5133);
or U5321 (N_5321,N_5188,N_5134);
nor U5322 (N_5322,N_5106,N_5032);
and U5323 (N_5323,N_5170,N_5027);
nor U5324 (N_5324,N_5096,N_5169);
or U5325 (N_5325,N_5072,N_5162);
nand U5326 (N_5326,N_5199,N_5149);
and U5327 (N_5327,N_5007,N_5081);
xnor U5328 (N_5328,N_5167,N_5149);
or U5329 (N_5329,N_5142,N_5056);
nor U5330 (N_5330,N_5045,N_5135);
nand U5331 (N_5331,N_5006,N_5118);
and U5332 (N_5332,N_5068,N_5124);
nor U5333 (N_5333,N_5052,N_5165);
and U5334 (N_5334,N_5170,N_5115);
nand U5335 (N_5335,N_5168,N_5180);
or U5336 (N_5336,N_5189,N_5072);
nand U5337 (N_5337,N_5178,N_5038);
xnor U5338 (N_5338,N_5024,N_5027);
and U5339 (N_5339,N_5184,N_5102);
xor U5340 (N_5340,N_5188,N_5178);
nor U5341 (N_5341,N_5071,N_5193);
or U5342 (N_5342,N_5131,N_5154);
or U5343 (N_5343,N_5011,N_5001);
xnor U5344 (N_5344,N_5001,N_5120);
and U5345 (N_5345,N_5173,N_5156);
xor U5346 (N_5346,N_5064,N_5020);
and U5347 (N_5347,N_5065,N_5176);
xor U5348 (N_5348,N_5089,N_5149);
nand U5349 (N_5349,N_5017,N_5071);
nand U5350 (N_5350,N_5145,N_5031);
or U5351 (N_5351,N_5114,N_5146);
nand U5352 (N_5352,N_5020,N_5055);
nor U5353 (N_5353,N_5025,N_5154);
nor U5354 (N_5354,N_5184,N_5026);
and U5355 (N_5355,N_5025,N_5195);
nor U5356 (N_5356,N_5179,N_5183);
and U5357 (N_5357,N_5069,N_5008);
nor U5358 (N_5358,N_5171,N_5033);
nor U5359 (N_5359,N_5190,N_5108);
nor U5360 (N_5360,N_5130,N_5071);
xor U5361 (N_5361,N_5147,N_5158);
xor U5362 (N_5362,N_5192,N_5059);
and U5363 (N_5363,N_5078,N_5101);
or U5364 (N_5364,N_5008,N_5146);
xor U5365 (N_5365,N_5124,N_5199);
xor U5366 (N_5366,N_5140,N_5073);
nor U5367 (N_5367,N_5035,N_5017);
or U5368 (N_5368,N_5136,N_5104);
nand U5369 (N_5369,N_5098,N_5035);
and U5370 (N_5370,N_5126,N_5043);
nor U5371 (N_5371,N_5166,N_5035);
nor U5372 (N_5372,N_5173,N_5039);
or U5373 (N_5373,N_5017,N_5062);
nor U5374 (N_5374,N_5166,N_5023);
xnor U5375 (N_5375,N_5155,N_5098);
nand U5376 (N_5376,N_5121,N_5174);
or U5377 (N_5377,N_5175,N_5024);
or U5378 (N_5378,N_5041,N_5024);
nor U5379 (N_5379,N_5019,N_5046);
nand U5380 (N_5380,N_5080,N_5183);
or U5381 (N_5381,N_5068,N_5153);
and U5382 (N_5382,N_5117,N_5060);
and U5383 (N_5383,N_5073,N_5161);
or U5384 (N_5384,N_5181,N_5139);
and U5385 (N_5385,N_5188,N_5056);
nand U5386 (N_5386,N_5019,N_5159);
nand U5387 (N_5387,N_5128,N_5018);
nand U5388 (N_5388,N_5018,N_5019);
nor U5389 (N_5389,N_5182,N_5137);
nor U5390 (N_5390,N_5011,N_5018);
xor U5391 (N_5391,N_5117,N_5124);
or U5392 (N_5392,N_5190,N_5162);
nand U5393 (N_5393,N_5031,N_5190);
and U5394 (N_5394,N_5140,N_5187);
nand U5395 (N_5395,N_5047,N_5188);
xnor U5396 (N_5396,N_5088,N_5050);
or U5397 (N_5397,N_5189,N_5140);
nand U5398 (N_5398,N_5071,N_5147);
nor U5399 (N_5399,N_5035,N_5163);
and U5400 (N_5400,N_5329,N_5395);
nand U5401 (N_5401,N_5388,N_5332);
and U5402 (N_5402,N_5373,N_5214);
nor U5403 (N_5403,N_5305,N_5291);
or U5404 (N_5404,N_5317,N_5235);
or U5405 (N_5405,N_5245,N_5311);
or U5406 (N_5406,N_5335,N_5264);
nor U5407 (N_5407,N_5371,N_5211);
nand U5408 (N_5408,N_5308,N_5269);
nand U5409 (N_5409,N_5230,N_5328);
or U5410 (N_5410,N_5320,N_5368);
nor U5411 (N_5411,N_5326,N_5327);
or U5412 (N_5412,N_5359,N_5324);
and U5413 (N_5413,N_5398,N_5210);
xor U5414 (N_5414,N_5208,N_5321);
and U5415 (N_5415,N_5325,N_5280);
nor U5416 (N_5416,N_5382,N_5363);
nor U5417 (N_5417,N_5267,N_5310);
nor U5418 (N_5418,N_5225,N_5380);
and U5419 (N_5419,N_5216,N_5336);
xor U5420 (N_5420,N_5242,N_5222);
or U5421 (N_5421,N_5374,N_5203);
nor U5422 (N_5422,N_5362,N_5276);
and U5423 (N_5423,N_5299,N_5255);
nand U5424 (N_5424,N_5238,N_5272);
xnor U5425 (N_5425,N_5357,N_5387);
nand U5426 (N_5426,N_5370,N_5282);
and U5427 (N_5427,N_5383,N_5349);
nor U5428 (N_5428,N_5389,N_5303);
xnor U5429 (N_5429,N_5285,N_5323);
or U5430 (N_5430,N_5217,N_5392);
or U5431 (N_5431,N_5314,N_5236);
nand U5432 (N_5432,N_5333,N_5342);
nor U5433 (N_5433,N_5215,N_5271);
nand U5434 (N_5434,N_5284,N_5201);
or U5435 (N_5435,N_5288,N_5281);
xor U5436 (N_5436,N_5337,N_5356);
nand U5437 (N_5437,N_5259,N_5385);
xnor U5438 (N_5438,N_5221,N_5367);
and U5439 (N_5439,N_5298,N_5205);
and U5440 (N_5440,N_5353,N_5237);
nor U5441 (N_5441,N_5243,N_5379);
and U5442 (N_5442,N_5289,N_5376);
or U5443 (N_5443,N_5372,N_5343);
nand U5444 (N_5444,N_5213,N_5352);
or U5445 (N_5445,N_5360,N_5265);
or U5446 (N_5446,N_5306,N_5307);
or U5447 (N_5447,N_5209,N_5233);
nor U5448 (N_5448,N_5227,N_5399);
xor U5449 (N_5449,N_5396,N_5338);
nand U5450 (N_5450,N_5348,N_5200);
nand U5451 (N_5451,N_5257,N_5339);
nor U5452 (N_5452,N_5394,N_5340);
nand U5453 (N_5453,N_5212,N_5366);
and U5454 (N_5454,N_5270,N_5228);
nand U5455 (N_5455,N_5224,N_5390);
or U5456 (N_5456,N_5304,N_5369);
nor U5457 (N_5457,N_5355,N_5286);
or U5458 (N_5458,N_5319,N_5207);
nor U5459 (N_5459,N_5283,N_5239);
nand U5460 (N_5460,N_5220,N_5229);
nand U5461 (N_5461,N_5252,N_5295);
xor U5462 (N_5462,N_5251,N_5219);
nand U5463 (N_5463,N_5346,N_5206);
nor U5464 (N_5464,N_5275,N_5313);
or U5465 (N_5465,N_5294,N_5386);
nor U5466 (N_5466,N_5278,N_5354);
nor U5467 (N_5467,N_5391,N_5204);
or U5468 (N_5468,N_5253,N_5345);
nand U5469 (N_5469,N_5393,N_5292);
nand U5470 (N_5470,N_5334,N_5256);
nor U5471 (N_5471,N_5375,N_5358);
and U5472 (N_5472,N_5240,N_5244);
xnor U5473 (N_5473,N_5232,N_5377);
and U5474 (N_5474,N_5318,N_5364);
nand U5475 (N_5475,N_5331,N_5330);
nor U5476 (N_5476,N_5297,N_5249);
and U5477 (N_5477,N_5384,N_5290);
or U5478 (N_5478,N_5381,N_5322);
xnor U5479 (N_5479,N_5241,N_5273);
nor U5480 (N_5480,N_5263,N_5266);
nand U5481 (N_5481,N_5301,N_5250);
or U5482 (N_5482,N_5293,N_5202);
nor U5483 (N_5483,N_5296,N_5350);
nand U5484 (N_5484,N_5234,N_5309);
nand U5485 (N_5485,N_5279,N_5274);
nor U5486 (N_5486,N_5261,N_5268);
nand U5487 (N_5487,N_5226,N_5260);
and U5488 (N_5488,N_5218,N_5351);
nor U5489 (N_5489,N_5254,N_5277);
nand U5490 (N_5490,N_5315,N_5316);
and U5491 (N_5491,N_5312,N_5344);
and U5492 (N_5492,N_5287,N_5223);
nand U5493 (N_5493,N_5347,N_5300);
nand U5494 (N_5494,N_5365,N_5397);
and U5495 (N_5495,N_5247,N_5258);
xor U5496 (N_5496,N_5246,N_5302);
nor U5497 (N_5497,N_5248,N_5361);
or U5498 (N_5498,N_5262,N_5378);
nand U5499 (N_5499,N_5341,N_5231);
nor U5500 (N_5500,N_5342,N_5399);
and U5501 (N_5501,N_5347,N_5250);
nor U5502 (N_5502,N_5359,N_5377);
or U5503 (N_5503,N_5315,N_5323);
nor U5504 (N_5504,N_5295,N_5349);
or U5505 (N_5505,N_5247,N_5376);
nand U5506 (N_5506,N_5216,N_5300);
nand U5507 (N_5507,N_5319,N_5366);
and U5508 (N_5508,N_5285,N_5290);
or U5509 (N_5509,N_5348,N_5373);
nand U5510 (N_5510,N_5338,N_5222);
and U5511 (N_5511,N_5230,N_5250);
nand U5512 (N_5512,N_5391,N_5390);
or U5513 (N_5513,N_5300,N_5346);
or U5514 (N_5514,N_5249,N_5302);
nor U5515 (N_5515,N_5232,N_5372);
xor U5516 (N_5516,N_5351,N_5357);
or U5517 (N_5517,N_5207,N_5217);
and U5518 (N_5518,N_5241,N_5323);
nor U5519 (N_5519,N_5343,N_5354);
nand U5520 (N_5520,N_5311,N_5351);
nor U5521 (N_5521,N_5213,N_5249);
or U5522 (N_5522,N_5290,N_5286);
and U5523 (N_5523,N_5364,N_5281);
nand U5524 (N_5524,N_5337,N_5351);
nand U5525 (N_5525,N_5280,N_5376);
nand U5526 (N_5526,N_5291,N_5372);
and U5527 (N_5527,N_5342,N_5316);
nand U5528 (N_5528,N_5214,N_5334);
or U5529 (N_5529,N_5228,N_5292);
nand U5530 (N_5530,N_5216,N_5243);
nor U5531 (N_5531,N_5304,N_5224);
and U5532 (N_5532,N_5243,N_5309);
and U5533 (N_5533,N_5244,N_5245);
nor U5534 (N_5534,N_5237,N_5250);
or U5535 (N_5535,N_5330,N_5370);
xor U5536 (N_5536,N_5331,N_5283);
nand U5537 (N_5537,N_5352,N_5304);
nand U5538 (N_5538,N_5347,N_5304);
and U5539 (N_5539,N_5278,N_5346);
or U5540 (N_5540,N_5274,N_5351);
nor U5541 (N_5541,N_5322,N_5209);
nor U5542 (N_5542,N_5330,N_5250);
or U5543 (N_5543,N_5325,N_5338);
and U5544 (N_5544,N_5371,N_5235);
and U5545 (N_5545,N_5358,N_5355);
nor U5546 (N_5546,N_5247,N_5286);
or U5547 (N_5547,N_5212,N_5372);
or U5548 (N_5548,N_5399,N_5392);
nand U5549 (N_5549,N_5340,N_5263);
nor U5550 (N_5550,N_5345,N_5326);
xnor U5551 (N_5551,N_5290,N_5216);
nor U5552 (N_5552,N_5333,N_5267);
nand U5553 (N_5553,N_5212,N_5375);
or U5554 (N_5554,N_5383,N_5211);
and U5555 (N_5555,N_5350,N_5374);
or U5556 (N_5556,N_5213,N_5332);
or U5557 (N_5557,N_5216,N_5376);
nor U5558 (N_5558,N_5283,N_5372);
and U5559 (N_5559,N_5215,N_5216);
nand U5560 (N_5560,N_5240,N_5320);
nand U5561 (N_5561,N_5295,N_5350);
and U5562 (N_5562,N_5271,N_5262);
nor U5563 (N_5563,N_5237,N_5321);
and U5564 (N_5564,N_5346,N_5331);
xnor U5565 (N_5565,N_5328,N_5291);
and U5566 (N_5566,N_5251,N_5227);
nor U5567 (N_5567,N_5353,N_5349);
or U5568 (N_5568,N_5291,N_5208);
nor U5569 (N_5569,N_5219,N_5233);
nor U5570 (N_5570,N_5288,N_5248);
nand U5571 (N_5571,N_5372,N_5208);
or U5572 (N_5572,N_5377,N_5264);
and U5573 (N_5573,N_5280,N_5345);
nand U5574 (N_5574,N_5344,N_5214);
nand U5575 (N_5575,N_5312,N_5208);
or U5576 (N_5576,N_5324,N_5202);
nor U5577 (N_5577,N_5302,N_5329);
nand U5578 (N_5578,N_5212,N_5282);
and U5579 (N_5579,N_5335,N_5236);
xnor U5580 (N_5580,N_5207,N_5365);
nand U5581 (N_5581,N_5311,N_5287);
nand U5582 (N_5582,N_5248,N_5250);
nand U5583 (N_5583,N_5391,N_5370);
nor U5584 (N_5584,N_5344,N_5289);
nand U5585 (N_5585,N_5274,N_5215);
or U5586 (N_5586,N_5352,N_5302);
nand U5587 (N_5587,N_5331,N_5296);
nor U5588 (N_5588,N_5368,N_5360);
or U5589 (N_5589,N_5317,N_5313);
and U5590 (N_5590,N_5381,N_5244);
and U5591 (N_5591,N_5335,N_5314);
xnor U5592 (N_5592,N_5352,N_5314);
nor U5593 (N_5593,N_5372,N_5229);
and U5594 (N_5594,N_5298,N_5238);
or U5595 (N_5595,N_5263,N_5377);
nor U5596 (N_5596,N_5367,N_5329);
and U5597 (N_5597,N_5258,N_5262);
nand U5598 (N_5598,N_5308,N_5359);
or U5599 (N_5599,N_5262,N_5264);
or U5600 (N_5600,N_5410,N_5484);
and U5601 (N_5601,N_5446,N_5534);
and U5602 (N_5602,N_5572,N_5432);
or U5603 (N_5603,N_5406,N_5597);
nor U5604 (N_5604,N_5408,N_5434);
nor U5605 (N_5605,N_5591,N_5433);
nand U5606 (N_5606,N_5500,N_5498);
or U5607 (N_5607,N_5416,N_5599);
and U5608 (N_5608,N_5456,N_5424);
nor U5609 (N_5609,N_5515,N_5556);
nand U5610 (N_5610,N_5587,N_5536);
and U5611 (N_5611,N_5481,N_5490);
or U5612 (N_5612,N_5496,N_5524);
or U5613 (N_5613,N_5548,N_5522);
nor U5614 (N_5614,N_5404,N_5480);
and U5615 (N_5615,N_5403,N_5503);
xnor U5616 (N_5616,N_5443,N_5405);
or U5617 (N_5617,N_5499,N_5519);
nand U5618 (N_5618,N_5558,N_5474);
nor U5619 (N_5619,N_5458,N_5575);
and U5620 (N_5620,N_5539,N_5477);
nand U5621 (N_5621,N_5593,N_5582);
nor U5622 (N_5622,N_5584,N_5567);
xnor U5623 (N_5623,N_5566,N_5440);
or U5624 (N_5624,N_5532,N_5400);
xnor U5625 (N_5625,N_5486,N_5520);
or U5626 (N_5626,N_5588,N_5563);
or U5627 (N_5627,N_5576,N_5560);
xnor U5628 (N_5628,N_5493,N_5487);
and U5629 (N_5629,N_5544,N_5527);
nor U5630 (N_5630,N_5421,N_5429);
or U5631 (N_5631,N_5465,N_5444);
nand U5632 (N_5632,N_5451,N_5598);
xor U5633 (N_5633,N_5533,N_5578);
or U5634 (N_5634,N_5547,N_5521);
nand U5635 (N_5635,N_5460,N_5495);
nor U5636 (N_5636,N_5554,N_5531);
nand U5637 (N_5637,N_5482,N_5543);
or U5638 (N_5638,N_5479,N_5426);
xor U5639 (N_5639,N_5549,N_5541);
and U5640 (N_5640,N_5476,N_5555);
and U5641 (N_5641,N_5431,N_5468);
nor U5642 (N_5642,N_5530,N_5430);
nor U5643 (N_5643,N_5436,N_5564);
and U5644 (N_5644,N_5427,N_5497);
nor U5645 (N_5645,N_5573,N_5418);
nor U5646 (N_5646,N_5492,N_5506);
nand U5647 (N_5647,N_5489,N_5469);
or U5648 (N_5648,N_5550,N_5570);
or U5649 (N_5649,N_5442,N_5419);
or U5650 (N_5650,N_5513,N_5420);
nor U5651 (N_5651,N_5449,N_5509);
or U5652 (N_5652,N_5401,N_5594);
and U5653 (N_5653,N_5512,N_5540);
nor U5654 (N_5654,N_5455,N_5445);
nand U5655 (N_5655,N_5413,N_5437);
nor U5656 (N_5656,N_5501,N_5415);
nand U5657 (N_5657,N_5553,N_5485);
nor U5658 (N_5658,N_5467,N_5473);
and U5659 (N_5659,N_5546,N_5529);
nor U5660 (N_5660,N_5414,N_5488);
and U5661 (N_5661,N_5508,N_5470);
nand U5662 (N_5662,N_5459,N_5478);
or U5663 (N_5663,N_5579,N_5528);
nor U5664 (N_5664,N_5526,N_5423);
nand U5665 (N_5665,N_5463,N_5595);
nand U5666 (N_5666,N_5457,N_5464);
nand U5667 (N_5667,N_5590,N_5454);
nor U5668 (N_5668,N_5517,N_5461);
or U5669 (N_5669,N_5422,N_5452);
or U5670 (N_5670,N_5537,N_5583);
or U5671 (N_5671,N_5581,N_5483);
xnor U5672 (N_5672,N_5462,N_5510);
nor U5673 (N_5673,N_5438,N_5557);
nand U5674 (N_5674,N_5523,N_5428);
nand U5675 (N_5675,N_5569,N_5545);
and U5676 (N_5676,N_5542,N_5448);
nand U5677 (N_5677,N_5409,N_5514);
nor U5678 (N_5678,N_5411,N_5402);
or U5679 (N_5679,N_5561,N_5453);
nand U5680 (N_5680,N_5466,N_5435);
nand U5681 (N_5681,N_5425,N_5447);
nor U5682 (N_5682,N_5494,N_5589);
nand U5683 (N_5683,N_5580,N_5450);
nand U5684 (N_5684,N_5574,N_5505);
or U5685 (N_5685,N_5535,N_5407);
or U5686 (N_5686,N_5475,N_5586);
or U5687 (N_5687,N_5417,N_5491);
nand U5688 (N_5688,N_5596,N_5441);
or U5689 (N_5689,N_5592,N_5412);
xor U5690 (N_5690,N_5518,N_5507);
nor U5691 (N_5691,N_5568,N_5471);
nand U5692 (N_5692,N_5504,N_5439);
and U5693 (N_5693,N_5577,N_5472);
or U5694 (N_5694,N_5525,N_5552);
or U5695 (N_5695,N_5565,N_5562);
nor U5696 (N_5696,N_5571,N_5502);
and U5697 (N_5697,N_5559,N_5585);
nand U5698 (N_5698,N_5538,N_5516);
and U5699 (N_5699,N_5551,N_5511);
or U5700 (N_5700,N_5505,N_5514);
nand U5701 (N_5701,N_5529,N_5474);
and U5702 (N_5702,N_5419,N_5535);
xor U5703 (N_5703,N_5485,N_5597);
nor U5704 (N_5704,N_5521,N_5475);
xnor U5705 (N_5705,N_5492,N_5577);
nand U5706 (N_5706,N_5505,N_5467);
and U5707 (N_5707,N_5489,N_5462);
or U5708 (N_5708,N_5505,N_5591);
xnor U5709 (N_5709,N_5516,N_5559);
nor U5710 (N_5710,N_5416,N_5520);
and U5711 (N_5711,N_5473,N_5557);
nor U5712 (N_5712,N_5549,N_5546);
nor U5713 (N_5713,N_5473,N_5527);
and U5714 (N_5714,N_5531,N_5529);
nor U5715 (N_5715,N_5441,N_5495);
nor U5716 (N_5716,N_5574,N_5535);
nor U5717 (N_5717,N_5497,N_5419);
nand U5718 (N_5718,N_5521,N_5400);
xnor U5719 (N_5719,N_5506,N_5586);
nor U5720 (N_5720,N_5540,N_5412);
nor U5721 (N_5721,N_5597,N_5419);
nor U5722 (N_5722,N_5426,N_5515);
or U5723 (N_5723,N_5407,N_5444);
or U5724 (N_5724,N_5401,N_5449);
xor U5725 (N_5725,N_5557,N_5540);
or U5726 (N_5726,N_5445,N_5530);
nor U5727 (N_5727,N_5583,N_5572);
xnor U5728 (N_5728,N_5486,N_5535);
nand U5729 (N_5729,N_5505,N_5477);
nor U5730 (N_5730,N_5503,N_5430);
and U5731 (N_5731,N_5529,N_5499);
nand U5732 (N_5732,N_5450,N_5473);
nand U5733 (N_5733,N_5551,N_5599);
nor U5734 (N_5734,N_5487,N_5507);
and U5735 (N_5735,N_5503,N_5595);
and U5736 (N_5736,N_5496,N_5538);
nor U5737 (N_5737,N_5423,N_5536);
nor U5738 (N_5738,N_5416,N_5465);
nand U5739 (N_5739,N_5410,N_5536);
or U5740 (N_5740,N_5463,N_5418);
and U5741 (N_5741,N_5568,N_5404);
and U5742 (N_5742,N_5517,N_5495);
nor U5743 (N_5743,N_5474,N_5580);
and U5744 (N_5744,N_5521,N_5456);
and U5745 (N_5745,N_5507,N_5585);
and U5746 (N_5746,N_5554,N_5479);
xor U5747 (N_5747,N_5583,N_5518);
nand U5748 (N_5748,N_5425,N_5574);
nand U5749 (N_5749,N_5505,N_5541);
or U5750 (N_5750,N_5430,N_5432);
nand U5751 (N_5751,N_5514,N_5496);
nand U5752 (N_5752,N_5540,N_5443);
nand U5753 (N_5753,N_5546,N_5497);
xnor U5754 (N_5754,N_5421,N_5435);
or U5755 (N_5755,N_5551,N_5543);
and U5756 (N_5756,N_5436,N_5484);
or U5757 (N_5757,N_5457,N_5442);
and U5758 (N_5758,N_5493,N_5410);
or U5759 (N_5759,N_5404,N_5570);
nor U5760 (N_5760,N_5556,N_5529);
nor U5761 (N_5761,N_5553,N_5575);
or U5762 (N_5762,N_5536,N_5407);
nand U5763 (N_5763,N_5595,N_5470);
xor U5764 (N_5764,N_5470,N_5510);
nor U5765 (N_5765,N_5545,N_5436);
or U5766 (N_5766,N_5475,N_5543);
or U5767 (N_5767,N_5548,N_5440);
and U5768 (N_5768,N_5544,N_5412);
nand U5769 (N_5769,N_5596,N_5496);
or U5770 (N_5770,N_5481,N_5586);
nor U5771 (N_5771,N_5410,N_5416);
nand U5772 (N_5772,N_5404,N_5453);
and U5773 (N_5773,N_5598,N_5508);
nand U5774 (N_5774,N_5500,N_5540);
nand U5775 (N_5775,N_5417,N_5501);
or U5776 (N_5776,N_5471,N_5572);
nor U5777 (N_5777,N_5532,N_5594);
nor U5778 (N_5778,N_5441,N_5553);
or U5779 (N_5779,N_5473,N_5549);
xor U5780 (N_5780,N_5449,N_5477);
or U5781 (N_5781,N_5430,N_5439);
nand U5782 (N_5782,N_5510,N_5570);
and U5783 (N_5783,N_5470,N_5552);
xor U5784 (N_5784,N_5591,N_5455);
or U5785 (N_5785,N_5562,N_5408);
nand U5786 (N_5786,N_5516,N_5448);
nand U5787 (N_5787,N_5522,N_5512);
nor U5788 (N_5788,N_5455,N_5430);
or U5789 (N_5789,N_5532,N_5440);
or U5790 (N_5790,N_5543,N_5593);
nand U5791 (N_5791,N_5510,N_5445);
nor U5792 (N_5792,N_5431,N_5503);
nand U5793 (N_5793,N_5480,N_5594);
nor U5794 (N_5794,N_5455,N_5510);
and U5795 (N_5795,N_5509,N_5576);
or U5796 (N_5796,N_5406,N_5564);
nand U5797 (N_5797,N_5528,N_5408);
and U5798 (N_5798,N_5404,N_5544);
and U5799 (N_5799,N_5500,N_5547);
nor U5800 (N_5800,N_5647,N_5779);
or U5801 (N_5801,N_5696,N_5601);
nand U5802 (N_5802,N_5784,N_5756);
xnor U5803 (N_5803,N_5616,N_5698);
nor U5804 (N_5804,N_5678,N_5721);
or U5805 (N_5805,N_5742,N_5798);
nor U5806 (N_5806,N_5791,N_5680);
nand U5807 (N_5807,N_5603,N_5621);
nor U5808 (N_5808,N_5747,N_5645);
or U5809 (N_5809,N_5674,N_5613);
nand U5810 (N_5810,N_5730,N_5725);
nor U5811 (N_5811,N_5775,N_5617);
nor U5812 (N_5812,N_5713,N_5649);
nand U5813 (N_5813,N_5724,N_5711);
nand U5814 (N_5814,N_5728,N_5655);
xor U5815 (N_5815,N_5642,N_5774);
nor U5816 (N_5816,N_5787,N_5703);
or U5817 (N_5817,N_5666,N_5634);
or U5818 (N_5818,N_5644,N_5654);
nand U5819 (N_5819,N_5631,N_5650);
nor U5820 (N_5820,N_5618,N_5785);
or U5821 (N_5821,N_5662,N_5619);
nand U5822 (N_5822,N_5684,N_5770);
nor U5823 (N_5823,N_5738,N_5632);
and U5824 (N_5824,N_5679,N_5754);
nand U5825 (N_5825,N_5729,N_5615);
xnor U5826 (N_5826,N_5608,N_5653);
nand U5827 (N_5827,N_5793,N_5772);
nand U5828 (N_5828,N_5697,N_5646);
nor U5829 (N_5829,N_5715,N_5667);
or U5830 (N_5830,N_5780,N_5665);
and U5831 (N_5831,N_5688,N_5788);
nor U5832 (N_5832,N_5718,N_5760);
nand U5833 (N_5833,N_5658,N_5744);
xnor U5834 (N_5834,N_5630,N_5737);
or U5835 (N_5835,N_5722,N_5694);
and U5836 (N_5836,N_5768,N_5767);
and U5837 (N_5837,N_5799,N_5605);
nor U5838 (N_5838,N_5639,N_5739);
nor U5839 (N_5839,N_5637,N_5704);
and U5840 (N_5840,N_5746,N_5640);
xor U5841 (N_5841,N_5687,N_5607);
or U5842 (N_5842,N_5627,N_5610);
nand U5843 (N_5843,N_5762,N_5755);
nor U5844 (N_5844,N_5781,N_5651);
or U5845 (N_5845,N_5792,N_5782);
nor U5846 (N_5846,N_5714,N_5777);
and U5847 (N_5847,N_5752,N_5604);
nor U5848 (N_5848,N_5691,N_5643);
and U5849 (N_5849,N_5695,N_5789);
and U5850 (N_5850,N_5641,N_5749);
nand U5851 (N_5851,N_5656,N_5638);
or U5852 (N_5852,N_5702,N_5701);
nand U5853 (N_5853,N_5764,N_5740);
nor U5854 (N_5854,N_5668,N_5727);
xnor U5855 (N_5855,N_5622,N_5794);
or U5856 (N_5856,N_5606,N_5612);
nand U5857 (N_5857,N_5685,N_5731);
or U5858 (N_5858,N_5663,N_5693);
and U5859 (N_5859,N_5648,N_5769);
nand U5860 (N_5860,N_5776,N_5705);
nor U5861 (N_5861,N_5602,N_5726);
or U5862 (N_5862,N_5786,N_5690);
nand U5863 (N_5863,N_5797,N_5623);
nand U5864 (N_5864,N_5706,N_5759);
and U5865 (N_5865,N_5635,N_5750);
xor U5866 (N_5866,N_5660,N_5699);
and U5867 (N_5867,N_5710,N_5686);
nand U5868 (N_5868,N_5717,N_5766);
nor U5869 (N_5869,N_5765,N_5745);
or U5870 (N_5870,N_5677,N_5761);
or U5871 (N_5871,N_5748,N_5636);
nor U5872 (N_5872,N_5692,N_5743);
and U5873 (N_5873,N_5669,N_5734);
and U5874 (N_5874,N_5652,N_5609);
nand U5875 (N_5875,N_5720,N_5620);
and U5876 (N_5876,N_5626,N_5682);
xor U5877 (N_5877,N_5757,N_5676);
nand U5878 (N_5878,N_5700,N_5708);
or U5879 (N_5879,N_5670,N_5683);
and U5880 (N_5880,N_5763,N_5751);
nor U5881 (N_5881,N_5795,N_5716);
xnor U5882 (N_5882,N_5771,N_5723);
or U5883 (N_5883,N_5614,N_5629);
nand U5884 (N_5884,N_5709,N_5783);
and U5885 (N_5885,N_5773,N_5657);
nor U5886 (N_5886,N_5753,N_5625);
nand U5887 (N_5887,N_5628,N_5796);
or U5888 (N_5888,N_5707,N_5758);
or U5889 (N_5889,N_5712,N_5600);
nand U5890 (N_5890,N_5778,N_5671);
nand U5891 (N_5891,N_5733,N_5659);
and U5892 (N_5892,N_5719,N_5673);
xnor U5893 (N_5893,N_5790,N_5732);
nor U5894 (N_5894,N_5672,N_5611);
nor U5895 (N_5895,N_5736,N_5681);
nand U5896 (N_5896,N_5735,N_5624);
nand U5897 (N_5897,N_5661,N_5633);
nor U5898 (N_5898,N_5675,N_5741);
or U5899 (N_5899,N_5689,N_5664);
nand U5900 (N_5900,N_5677,N_5783);
nor U5901 (N_5901,N_5723,N_5674);
or U5902 (N_5902,N_5771,N_5701);
nor U5903 (N_5903,N_5607,N_5678);
or U5904 (N_5904,N_5747,N_5782);
nor U5905 (N_5905,N_5717,N_5640);
or U5906 (N_5906,N_5724,N_5701);
nor U5907 (N_5907,N_5666,N_5729);
and U5908 (N_5908,N_5650,N_5692);
nor U5909 (N_5909,N_5784,N_5746);
and U5910 (N_5910,N_5730,N_5628);
and U5911 (N_5911,N_5792,N_5604);
nand U5912 (N_5912,N_5642,N_5701);
nor U5913 (N_5913,N_5724,N_5640);
nand U5914 (N_5914,N_5781,N_5642);
or U5915 (N_5915,N_5643,N_5678);
xor U5916 (N_5916,N_5743,N_5737);
nand U5917 (N_5917,N_5625,N_5646);
or U5918 (N_5918,N_5642,N_5674);
and U5919 (N_5919,N_5688,N_5714);
nor U5920 (N_5920,N_5760,N_5629);
or U5921 (N_5921,N_5741,N_5627);
and U5922 (N_5922,N_5623,N_5741);
nor U5923 (N_5923,N_5790,N_5777);
and U5924 (N_5924,N_5617,N_5606);
xnor U5925 (N_5925,N_5615,N_5753);
and U5926 (N_5926,N_5784,N_5650);
nor U5927 (N_5927,N_5725,N_5706);
nand U5928 (N_5928,N_5784,N_5626);
xnor U5929 (N_5929,N_5631,N_5617);
nor U5930 (N_5930,N_5734,N_5638);
and U5931 (N_5931,N_5693,N_5613);
or U5932 (N_5932,N_5654,N_5720);
nand U5933 (N_5933,N_5730,N_5710);
and U5934 (N_5934,N_5741,N_5727);
nor U5935 (N_5935,N_5719,N_5770);
and U5936 (N_5936,N_5602,N_5763);
nand U5937 (N_5937,N_5623,N_5604);
nand U5938 (N_5938,N_5670,N_5760);
and U5939 (N_5939,N_5684,N_5703);
nand U5940 (N_5940,N_5659,N_5612);
nand U5941 (N_5941,N_5602,N_5728);
and U5942 (N_5942,N_5655,N_5684);
nand U5943 (N_5943,N_5699,N_5695);
nand U5944 (N_5944,N_5726,N_5750);
nand U5945 (N_5945,N_5661,N_5712);
and U5946 (N_5946,N_5635,N_5722);
nand U5947 (N_5947,N_5772,N_5607);
or U5948 (N_5948,N_5633,N_5720);
or U5949 (N_5949,N_5708,N_5711);
nor U5950 (N_5950,N_5737,N_5642);
nand U5951 (N_5951,N_5666,N_5795);
nor U5952 (N_5952,N_5778,N_5674);
and U5953 (N_5953,N_5608,N_5600);
nand U5954 (N_5954,N_5722,N_5669);
and U5955 (N_5955,N_5612,N_5792);
nor U5956 (N_5956,N_5610,N_5721);
or U5957 (N_5957,N_5640,N_5618);
nor U5958 (N_5958,N_5637,N_5671);
or U5959 (N_5959,N_5686,N_5645);
nor U5960 (N_5960,N_5746,N_5631);
nor U5961 (N_5961,N_5621,N_5636);
nand U5962 (N_5962,N_5698,N_5707);
nand U5963 (N_5963,N_5608,N_5759);
nand U5964 (N_5964,N_5621,N_5784);
nand U5965 (N_5965,N_5623,N_5692);
nand U5966 (N_5966,N_5724,N_5741);
nor U5967 (N_5967,N_5782,N_5788);
and U5968 (N_5968,N_5600,N_5783);
and U5969 (N_5969,N_5692,N_5628);
nand U5970 (N_5970,N_5708,N_5703);
nand U5971 (N_5971,N_5635,N_5690);
nor U5972 (N_5972,N_5770,N_5720);
and U5973 (N_5973,N_5760,N_5797);
or U5974 (N_5974,N_5615,N_5750);
nor U5975 (N_5975,N_5689,N_5701);
xnor U5976 (N_5976,N_5717,N_5760);
and U5977 (N_5977,N_5756,N_5723);
or U5978 (N_5978,N_5792,N_5702);
nor U5979 (N_5979,N_5747,N_5638);
nand U5980 (N_5980,N_5731,N_5633);
xor U5981 (N_5981,N_5674,N_5661);
or U5982 (N_5982,N_5640,N_5731);
xnor U5983 (N_5983,N_5639,N_5661);
nor U5984 (N_5984,N_5751,N_5777);
xor U5985 (N_5985,N_5650,N_5660);
or U5986 (N_5986,N_5663,N_5798);
nor U5987 (N_5987,N_5786,N_5681);
or U5988 (N_5988,N_5717,N_5702);
and U5989 (N_5989,N_5766,N_5774);
xor U5990 (N_5990,N_5646,N_5739);
nand U5991 (N_5991,N_5779,N_5786);
or U5992 (N_5992,N_5737,N_5754);
or U5993 (N_5993,N_5793,N_5679);
and U5994 (N_5994,N_5795,N_5622);
or U5995 (N_5995,N_5618,N_5630);
or U5996 (N_5996,N_5713,N_5741);
and U5997 (N_5997,N_5654,N_5698);
nand U5998 (N_5998,N_5613,N_5720);
and U5999 (N_5999,N_5670,N_5743);
nor U6000 (N_6000,N_5808,N_5873);
or U6001 (N_6001,N_5963,N_5970);
or U6002 (N_6002,N_5939,N_5812);
xor U6003 (N_6003,N_5817,N_5904);
and U6004 (N_6004,N_5898,N_5848);
and U6005 (N_6005,N_5885,N_5974);
and U6006 (N_6006,N_5975,N_5907);
and U6007 (N_6007,N_5979,N_5947);
nand U6008 (N_6008,N_5996,N_5805);
or U6009 (N_6009,N_5899,N_5832);
or U6010 (N_6010,N_5825,N_5830);
and U6011 (N_6011,N_5821,N_5870);
and U6012 (N_6012,N_5835,N_5881);
or U6013 (N_6013,N_5890,N_5901);
or U6014 (N_6014,N_5931,N_5920);
nor U6015 (N_6015,N_5822,N_5884);
xor U6016 (N_6016,N_5802,N_5807);
nor U6017 (N_6017,N_5992,N_5871);
nand U6018 (N_6018,N_5876,N_5868);
nand U6019 (N_6019,N_5872,N_5813);
or U6020 (N_6020,N_5980,N_5982);
and U6021 (N_6021,N_5972,N_5999);
xnor U6022 (N_6022,N_5914,N_5809);
nor U6023 (N_6023,N_5858,N_5866);
or U6024 (N_6024,N_5845,N_5895);
or U6025 (N_6025,N_5942,N_5846);
nand U6026 (N_6026,N_5861,N_5935);
and U6027 (N_6027,N_5887,N_5943);
or U6028 (N_6028,N_5915,N_5940);
and U6029 (N_6029,N_5998,N_5806);
nand U6030 (N_6030,N_5838,N_5891);
nand U6031 (N_6031,N_5965,N_5828);
nand U6032 (N_6032,N_5969,N_5928);
and U6033 (N_6033,N_5869,N_5847);
nor U6034 (N_6034,N_5816,N_5993);
and U6035 (N_6035,N_5952,N_5883);
xnor U6036 (N_6036,N_5938,N_5919);
nor U6037 (N_6037,N_5853,N_5867);
or U6038 (N_6038,N_5916,N_5855);
and U6039 (N_6039,N_5836,N_5811);
nand U6040 (N_6040,N_5926,N_5837);
nand U6041 (N_6041,N_5810,N_5893);
nor U6042 (N_6042,N_5878,N_5911);
or U6043 (N_6043,N_5995,N_5864);
nand U6044 (N_6044,N_5909,N_5962);
and U6045 (N_6045,N_5829,N_5981);
nor U6046 (N_6046,N_5964,N_5986);
or U6047 (N_6047,N_5960,N_5906);
or U6048 (N_6048,N_5852,N_5801);
and U6049 (N_6049,N_5921,N_5823);
and U6050 (N_6050,N_5959,N_5875);
nand U6051 (N_6051,N_5857,N_5958);
nor U6052 (N_6052,N_5936,N_5944);
or U6053 (N_6053,N_5840,N_5849);
and U6054 (N_6054,N_5994,N_5957);
nor U6055 (N_6055,N_5833,N_5856);
or U6056 (N_6056,N_5804,N_5976);
and U6057 (N_6057,N_5818,N_5839);
nor U6058 (N_6058,N_5879,N_5984);
nand U6059 (N_6059,N_5886,N_5859);
xnor U6060 (N_6060,N_5929,N_5934);
and U6061 (N_6061,N_5923,N_5800);
or U6062 (N_6062,N_5882,N_5908);
or U6063 (N_6063,N_5930,N_5918);
nand U6064 (N_6064,N_5819,N_5896);
xnor U6065 (N_6065,N_5956,N_5874);
nor U6066 (N_6066,N_5880,N_5925);
or U6067 (N_6067,N_5954,N_5987);
nor U6068 (N_6068,N_5978,N_5903);
or U6069 (N_6069,N_5851,N_5877);
and U6070 (N_6070,N_5951,N_5988);
or U6071 (N_6071,N_5902,N_5961);
or U6072 (N_6072,N_5900,N_5860);
xor U6073 (N_6073,N_5950,N_5888);
and U6074 (N_6074,N_5917,N_5953);
nand U6075 (N_6075,N_5971,N_5933);
and U6076 (N_6076,N_5955,N_5927);
or U6077 (N_6077,N_5941,N_5983);
nand U6078 (N_6078,N_5973,N_5912);
and U6079 (N_6079,N_5863,N_5990);
nor U6080 (N_6080,N_5910,N_5946);
and U6081 (N_6081,N_5826,N_5815);
xor U6082 (N_6082,N_5967,N_5803);
nand U6083 (N_6083,N_5842,N_5968);
or U6084 (N_6084,N_5854,N_5966);
and U6085 (N_6085,N_5824,N_5977);
nor U6086 (N_6086,N_5892,N_5820);
and U6087 (N_6087,N_5932,N_5985);
or U6088 (N_6088,N_5924,N_5844);
nand U6089 (N_6089,N_5894,N_5997);
nor U6090 (N_6090,N_5814,N_5991);
and U6091 (N_6091,N_5889,N_5831);
nand U6092 (N_6092,N_5865,N_5862);
or U6093 (N_6093,N_5827,N_5913);
nand U6094 (N_6094,N_5850,N_5905);
nor U6095 (N_6095,N_5834,N_5948);
or U6096 (N_6096,N_5989,N_5949);
or U6097 (N_6097,N_5945,N_5922);
or U6098 (N_6098,N_5897,N_5937);
xor U6099 (N_6099,N_5843,N_5841);
xnor U6100 (N_6100,N_5897,N_5863);
and U6101 (N_6101,N_5978,N_5858);
nand U6102 (N_6102,N_5899,N_5936);
or U6103 (N_6103,N_5908,N_5833);
and U6104 (N_6104,N_5976,N_5994);
and U6105 (N_6105,N_5983,N_5914);
xnor U6106 (N_6106,N_5908,N_5848);
or U6107 (N_6107,N_5822,N_5853);
nor U6108 (N_6108,N_5924,N_5956);
or U6109 (N_6109,N_5866,N_5946);
or U6110 (N_6110,N_5994,N_5954);
nand U6111 (N_6111,N_5963,N_5911);
and U6112 (N_6112,N_5966,N_5881);
or U6113 (N_6113,N_5807,N_5871);
or U6114 (N_6114,N_5929,N_5801);
and U6115 (N_6115,N_5868,N_5822);
and U6116 (N_6116,N_5813,N_5968);
and U6117 (N_6117,N_5854,N_5863);
and U6118 (N_6118,N_5941,N_5874);
nand U6119 (N_6119,N_5964,N_5889);
nand U6120 (N_6120,N_5885,N_5811);
nor U6121 (N_6121,N_5876,N_5846);
nor U6122 (N_6122,N_5902,N_5964);
nor U6123 (N_6123,N_5845,N_5885);
nor U6124 (N_6124,N_5804,N_5867);
nor U6125 (N_6125,N_5865,N_5804);
nand U6126 (N_6126,N_5867,N_5933);
or U6127 (N_6127,N_5951,N_5963);
xnor U6128 (N_6128,N_5868,N_5983);
nand U6129 (N_6129,N_5848,N_5828);
nor U6130 (N_6130,N_5879,N_5950);
nor U6131 (N_6131,N_5950,N_5805);
nor U6132 (N_6132,N_5933,N_5805);
and U6133 (N_6133,N_5951,N_5975);
nand U6134 (N_6134,N_5804,N_5967);
nor U6135 (N_6135,N_5837,N_5823);
nand U6136 (N_6136,N_5999,N_5801);
nand U6137 (N_6137,N_5869,N_5995);
or U6138 (N_6138,N_5945,N_5866);
nor U6139 (N_6139,N_5886,N_5862);
nor U6140 (N_6140,N_5919,N_5890);
and U6141 (N_6141,N_5949,N_5998);
and U6142 (N_6142,N_5982,N_5935);
nor U6143 (N_6143,N_5937,N_5971);
nand U6144 (N_6144,N_5847,N_5918);
nor U6145 (N_6145,N_5831,N_5979);
or U6146 (N_6146,N_5828,N_5894);
xnor U6147 (N_6147,N_5961,N_5939);
and U6148 (N_6148,N_5954,N_5886);
nand U6149 (N_6149,N_5981,N_5815);
and U6150 (N_6150,N_5953,N_5905);
and U6151 (N_6151,N_5965,N_5810);
nor U6152 (N_6152,N_5874,N_5826);
nor U6153 (N_6153,N_5917,N_5937);
nand U6154 (N_6154,N_5870,N_5969);
and U6155 (N_6155,N_5831,N_5866);
nor U6156 (N_6156,N_5884,N_5881);
nor U6157 (N_6157,N_5906,N_5850);
or U6158 (N_6158,N_5917,N_5973);
or U6159 (N_6159,N_5893,N_5915);
or U6160 (N_6160,N_5815,N_5846);
or U6161 (N_6161,N_5977,N_5804);
and U6162 (N_6162,N_5839,N_5975);
nor U6163 (N_6163,N_5964,N_5916);
nor U6164 (N_6164,N_5878,N_5869);
or U6165 (N_6165,N_5834,N_5839);
nor U6166 (N_6166,N_5991,N_5815);
nor U6167 (N_6167,N_5870,N_5914);
and U6168 (N_6168,N_5990,N_5961);
and U6169 (N_6169,N_5864,N_5982);
and U6170 (N_6170,N_5950,N_5934);
or U6171 (N_6171,N_5962,N_5960);
nor U6172 (N_6172,N_5946,N_5854);
xnor U6173 (N_6173,N_5939,N_5992);
nor U6174 (N_6174,N_5959,N_5907);
and U6175 (N_6175,N_5909,N_5847);
xnor U6176 (N_6176,N_5961,N_5972);
or U6177 (N_6177,N_5971,N_5894);
xnor U6178 (N_6178,N_5840,N_5994);
nor U6179 (N_6179,N_5936,N_5803);
nor U6180 (N_6180,N_5859,N_5826);
and U6181 (N_6181,N_5949,N_5992);
nor U6182 (N_6182,N_5871,N_5912);
and U6183 (N_6183,N_5973,N_5901);
xnor U6184 (N_6184,N_5983,N_5954);
nand U6185 (N_6185,N_5971,N_5881);
nand U6186 (N_6186,N_5946,N_5875);
nor U6187 (N_6187,N_5871,N_5811);
xnor U6188 (N_6188,N_5961,N_5999);
nand U6189 (N_6189,N_5851,N_5827);
or U6190 (N_6190,N_5904,N_5898);
or U6191 (N_6191,N_5854,N_5867);
nor U6192 (N_6192,N_5841,N_5820);
and U6193 (N_6193,N_5929,N_5957);
and U6194 (N_6194,N_5850,N_5857);
nor U6195 (N_6195,N_5961,N_5816);
nor U6196 (N_6196,N_5893,N_5901);
or U6197 (N_6197,N_5885,N_5919);
nor U6198 (N_6198,N_5903,N_5907);
and U6199 (N_6199,N_5809,N_5859);
or U6200 (N_6200,N_6083,N_6012);
or U6201 (N_6201,N_6047,N_6094);
nor U6202 (N_6202,N_6062,N_6178);
nand U6203 (N_6203,N_6115,N_6106);
or U6204 (N_6204,N_6024,N_6150);
or U6205 (N_6205,N_6026,N_6055);
nand U6206 (N_6206,N_6125,N_6086);
or U6207 (N_6207,N_6114,N_6120);
and U6208 (N_6208,N_6173,N_6085);
and U6209 (N_6209,N_6091,N_6021);
and U6210 (N_6210,N_6035,N_6181);
and U6211 (N_6211,N_6102,N_6159);
nor U6212 (N_6212,N_6029,N_6195);
or U6213 (N_6213,N_6148,N_6138);
nand U6214 (N_6214,N_6191,N_6113);
xor U6215 (N_6215,N_6137,N_6103);
or U6216 (N_6216,N_6043,N_6112);
and U6217 (N_6217,N_6053,N_6110);
nand U6218 (N_6218,N_6118,N_6186);
and U6219 (N_6219,N_6171,N_6182);
or U6220 (N_6220,N_6160,N_6071);
or U6221 (N_6221,N_6065,N_6097);
nand U6222 (N_6222,N_6111,N_6005);
nor U6223 (N_6223,N_6072,N_6116);
nor U6224 (N_6224,N_6014,N_6164);
and U6225 (N_6225,N_6064,N_6121);
nand U6226 (N_6226,N_6066,N_6162);
and U6227 (N_6227,N_6156,N_6140);
nand U6228 (N_6228,N_6139,N_6147);
nor U6229 (N_6229,N_6092,N_6036);
or U6230 (N_6230,N_6108,N_6176);
nand U6231 (N_6231,N_6199,N_6002);
nand U6232 (N_6232,N_6197,N_6010);
nand U6233 (N_6233,N_6166,N_6167);
or U6234 (N_6234,N_6135,N_6174);
nand U6235 (N_6235,N_6141,N_6130);
nand U6236 (N_6236,N_6013,N_6009);
nand U6237 (N_6237,N_6152,N_6158);
xor U6238 (N_6238,N_6142,N_6008);
or U6239 (N_6239,N_6104,N_6132);
nand U6240 (N_6240,N_6041,N_6100);
nand U6241 (N_6241,N_6179,N_6196);
nor U6242 (N_6242,N_6081,N_6031);
and U6243 (N_6243,N_6042,N_6190);
or U6244 (N_6244,N_6069,N_6089);
nor U6245 (N_6245,N_6076,N_6122);
or U6246 (N_6246,N_6131,N_6168);
nor U6247 (N_6247,N_6109,N_6101);
nand U6248 (N_6248,N_6063,N_6129);
or U6249 (N_6249,N_6044,N_6022);
nor U6250 (N_6250,N_6049,N_6073);
nand U6251 (N_6251,N_6025,N_6084);
nor U6252 (N_6252,N_6070,N_6032);
and U6253 (N_6253,N_6165,N_6090);
xor U6254 (N_6254,N_6105,N_6144);
and U6255 (N_6255,N_6033,N_6187);
nor U6256 (N_6256,N_6128,N_6019);
or U6257 (N_6257,N_6000,N_6080);
or U6258 (N_6258,N_6037,N_6133);
and U6259 (N_6259,N_6074,N_6058);
nor U6260 (N_6260,N_6119,N_6154);
xnor U6261 (N_6261,N_6050,N_6151);
nand U6262 (N_6262,N_6015,N_6143);
nor U6263 (N_6263,N_6003,N_6077);
xnor U6264 (N_6264,N_6027,N_6180);
nand U6265 (N_6265,N_6146,N_6172);
and U6266 (N_6266,N_6038,N_6059);
nor U6267 (N_6267,N_6061,N_6057);
or U6268 (N_6268,N_6054,N_6126);
or U6269 (N_6269,N_6177,N_6099);
nor U6270 (N_6270,N_6034,N_6136);
nand U6271 (N_6271,N_6123,N_6157);
nor U6272 (N_6272,N_6007,N_6075);
xor U6273 (N_6273,N_6149,N_6161);
nor U6274 (N_6274,N_6006,N_6051);
xor U6275 (N_6275,N_6096,N_6124);
nor U6276 (N_6276,N_6060,N_6134);
nand U6277 (N_6277,N_6056,N_6127);
nand U6278 (N_6278,N_6039,N_6107);
or U6279 (N_6279,N_6078,N_6193);
nor U6280 (N_6280,N_6011,N_6188);
or U6281 (N_6281,N_6082,N_6045);
nor U6282 (N_6282,N_6093,N_6198);
and U6283 (N_6283,N_6163,N_6155);
nand U6284 (N_6284,N_6052,N_6183);
nor U6285 (N_6285,N_6023,N_6145);
nand U6286 (N_6286,N_6194,N_6016);
and U6287 (N_6287,N_6079,N_6192);
xnor U6288 (N_6288,N_6004,N_6153);
xor U6289 (N_6289,N_6185,N_6175);
nor U6290 (N_6290,N_6184,N_6018);
and U6291 (N_6291,N_6028,N_6068);
nor U6292 (N_6292,N_6040,N_6001);
or U6293 (N_6293,N_6030,N_6088);
nor U6294 (N_6294,N_6095,N_6087);
or U6295 (N_6295,N_6020,N_6170);
nand U6296 (N_6296,N_6189,N_6067);
and U6297 (N_6297,N_6046,N_6017);
nand U6298 (N_6298,N_6098,N_6117);
and U6299 (N_6299,N_6048,N_6169);
and U6300 (N_6300,N_6151,N_6149);
and U6301 (N_6301,N_6143,N_6156);
nor U6302 (N_6302,N_6049,N_6179);
nand U6303 (N_6303,N_6187,N_6009);
xor U6304 (N_6304,N_6109,N_6174);
nor U6305 (N_6305,N_6193,N_6050);
nor U6306 (N_6306,N_6016,N_6122);
nand U6307 (N_6307,N_6036,N_6106);
nor U6308 (N_6308,N_6156,N_6125);
or U6309 (N_6309,N_6090,N_6192);
nand U6310 (N_6310,N_6024,N_6079);
nand U6311 (N_6311,N_6155,N_6086);
nand U6312 (N_6312,N_6019,N_6087);
or U6313 (N_6313,N_6050,N_6144);
xor U6314 (N_6314,N_6086,N_6087);
nand U6315 (N_6315,N_6180,N_6186);
or U6316 (N_6316,N_6072,N_6173);
nand U6317 (N_6317,N_6103,N_6008);
nor U6318 (N_6318,N_6015,N_6018);
nor U6319 (N_6319,N_6110,N_6194);
and U6320 (N_6320,N_6023,N_6184);
xor U6321 (N_6321,N_6092,N_6033);
nor U6322 (N_6322,N_6167,N_6122);
or U6323 (N_6323,N_6012,N_6037);
nand U6324 (N_6324,N_6058,N_6198);
xor U6325 (N_6325,N_6081,N_6028);
and U6326 (N_6326,N_6055,N_6156);
or U6327 (N_6327,N_6022,N_6085);
and U6328 (N_6328,N_6115,N_6110);
and U6329 (N_6329,N_6135,N_6021);
nand U6330 (N_6330,N_6027,N_6124);
nand U6331 (N_6331,N_6131,N_6184);
nand U6332 (N_6332,N_6175,N_6044);
xnor U6333 (N_6333,N_6169,N_6060);
nand U6334 (N_6334,N_6078,N_6135);
nand U6335 (N_6335,N_6121,N_6022);
nor U6336 (N_6336,N_6028,N_6082);
nor U6337 (N_6337,N_6159,N_6015);
or U6338 (N_6338,N_6167,N_6194);
and U6339 (N_6339,N_6074,N_6172);
and U6340 (N_6340,N_6187,N_6143);
or U6341 (N_6341,N_6122,N_6043);
or U6342 (N_6342,N_6088,N_6028);
nor U6343 (N_6343,N_6133,N_6127);
nor U6344 (N_6344,N_6171,N_6098);
and U6345 (N_6345,N_6117,N_6140);
nor U6346 (N_6346,N_6073,N_6129);
or U6347 (N_6347,N_6098,N_6139);
nor U6348 (N_6348,N_6013,N_6144);
nor U6349 (N_6349,N_6170,N_6153);
or U6350 (N_6350,N_6191,N_6020);
nor U6351 (N_6351,N_6139,N_6124);
nor U6352 (N_6352,N_6134,N_6169);
and U6353 (N_6353,N_6070,N_6141);
and U6354 (N_6354,N_6023,N_6139);
or U6355 (N_6355,N_6012,N_6043);
xor U6356 (N_6356,N_6099,N_6040);
nand U6357 (N_6357,N_6077,N_6105);
nor U6358 (N_6358,N_6138,N_6195);
nand U6359 (N_6359,N_6075,N_6126);
and U6360 (N_6360,N_6042,N_6069);
and U6361 (N_6361,N_6016,N_6110);
or U6362 (N_6362,N_6151,N_6159);
nand U6363 (N_6363,N_6196,N_6115);
nor U6364 (N_6364,N_6020,N_6056);
nor U6365 (N_6365,N_6046,N_6033);
nand U6366 (N_6366,N_6002,N_6117);
and U6367 (N_6367,N_6134,N_6151);
nand U6368 (N_6368,N_6045,N_6035);
nor U6369 (N_6369,N_6051,N_6177);
nand U6370 (N_6370,N_6125,N_6167);
xor U6371 (N_6371,N_6096,N_6160);
nor U6372 (N_6372,N_6062,N_6196);
or U6373 (N_6373,N_6055,N_6082);
or U6374 (N_6374,N_6063,N_6008);
or U6375 (N_6375,N_6075,N_6185);
nand U6376 (N_6376,N_6070,N_6055);
and U6377 (N_6377,N_6028,N_6173);
and U6378 (N_6378,N_6010,N_6011);
nand U6379 (N_6379,N_6187,N_6072);
nor U6380 (N_6380,N_6114,N_6087);
and U6381 (N_6381,N_6019,N_6014);
and U6382 (N_6382,N_6082,N_6093);
nand U6383 (N_6383,N_6160,N_6001);
and U6384 (N_6384,N_6044,N_6025);
nand U6385 (N_6385,N_6191,N_6197);
xnor U6386 (N_6386,N_6126,N_6010);
or U6387 (N_6387,N_6166,N_6181);
or U6388 (N_6388,N_6078,N_6129);
and U6389 (N_6389,N_6121,N_6173);
nand U6390 (N_6390,N_6028,N_6073);
nor U6391 (N_6391,N_6007,N_6112);
and U6392 (N_6392,N_6103,N_6138);
xor U6393 (N_6393,N_6005,N_6016);
xor U6394 (N_6394,N_6146,N_6176);
nor U6395 (N_6395,N_6172,N_6061);
and U6396 (N_6396,N_6091,N_6024);
nor U6397 (N_6397,N_6070,N_6056);
nand U6398 (N_6398,N_6045,N_6098);
nand U6399 (N_6399,N_6094,N_6191);
nor U6400 (N_6400,N_6335,N_6208);
nor U6401 (N_6401,N_6221,N_6363);
and U6402 (N_6402,N_6298,N_6270);
nor U6403 (N_6403,N_6343,N_6211);
xnor U6404 (N_6404,N_6290,N_6389);
nand U6405 (N_6405,N_6289,N_6231);
nand U6406 (N_6406,N_6253,N_6263);
or U6407 (N_6407,N_6362,N_6313);
nor U6408 (N_6408,N_6275,N_6259);
and U6409 (N_6409,N_6248,N_6318);
and U6410 (N_6410,N_6361,N_6317);
or U6411 (N_6411,N_6203,N_6353);
or U6412 (N_6412,N_6204,N_6288);
or U6413 (N_6413,N_6226,N_6321);
or U6414 (N_6414,N_6356,N_6387);
or U6415 (N_6415,N_6309,N_6252);
and U6416 (N_6416,N_6247,N_6234);
and U6417 (N_6417,N_6314,N_6339);
nand U6418 (N_6418,N_6383,N_6315);
nor U6419 (N_6419,N_6293,N_6341);
nor U6420 (N_6420,N_6281,N_6224);
xnor U6421 (N_6421,N_6254,N_6307);
and U6422 (N_6422,N_6394,N_6225);
and U6423 (N_6423,N_6207,N_6260);
and U6424 (N_6424,N_6265,N_6354);
nor U6425 (N_6425,N_6355,N_6250);
nor U6426 (N_6426,N_6292,N_6351);
and U6427 (N_6427,N_6308,N_6212);
nand U6428 (N_6428,N_6216,N_6337);
nor U6429 (N_6429,N_6230,N_6323);
or U6430 (N_6430,N_6336,N_6338);
nand U6431 (N_6431,N_6302,N_6229);
or U6432 (N_6432,N_6391,N_6306);
nand U6433 (N_6433,N_6373,N_6284);
or U6434 (N_6434,N_6320,N_6379);
xor U6435 (N_6435,N_6255,N_6294);
xor U6436 (N_6436,N_6241,N_6269);
nand U6437 (N_6437,N_6277,N_6228);
and U6438 (N_6438,N_6214,N_6202);
nor U6439 (N_6439,N_6358,N_6276);
nand U6440 (N_6440,N_6227,N_6342);
or U6441 (N_6441,N_6279,N_6310);
and U6442 (N_6442,N_6299,N_6236);
or U6443 (N_6443,N_6380,N_6311);
or U6444 (N_6444,N_6374,N_6328);
and U6445 (N_6445,N_6238,N_6200);
nor U6446 (N_6446,N_6297,N_6364);
and U6447 (N_6447,N_6326,N_6369);
nor U6448 (N_6448,N_6395,N_6392);
or U6449 (N_6449,N_6327,N_6213);
and U6450 (N_6450,N_6257,N_6296);
nand U6451 (N_6451,N_6367,N_6283);
nand U6452 (N_6452,N_6324,N_6390);
and U6453 (N_6453,N_6258,N_6268);
nand U6454 (N_6454,N_6201,N_6271);
and U6455 (N_6455,N_6382,N_6240);
or U6456 (N_6456,N_6376,N_6237);
xnor U6457 (N_6457,N_6377,N_6352);
and U6458 (N_6458,N_6262,N_6386);
or U6459 (N_6459,N_6206,N_6359);
nand U6460 (N_6460,N_6357,N_6267);
nor U6461 (N_6461,N_6329,N_6345);
nand U6462 (N_6462,N_6393,N_6285);
nand U6463 (N_6463,N_6273,N_6397);
and U6464 (N_6464,N_6251,N_6218);
and U6465 (N_6465,N_6233,N_6316);
and U6466 (N_6466,N_6280,N_6372);
nor U6467 (N_6467,N_6340,N_6222);
nand U6468 (N_6468,N_6205,N_6246);
xor U6469 (N_6469,N_6239,N_6223);
or U6470 (N_6470,N_6274,N_6300);
xnor U6471 (N_6471,N_6396,N_6332);
or U6472 (N_6472,N_6245,N_6334);
or U6473 (N_6473,N_6291,N_6325);
nor U6474 (N_6474,N_6312,N_6381);
or U6475 (N_6475,N_6368,N_6278);
or U6476 (N_6476,N_6348,N_6370);
xor U6477 (N_6477,N_6330,N_6232);
nor U6478 (N_6478,N_6384,N_6319);
or U6479 (N_6479,N_6282,N_6371);
or U6480 (N_6480,N_6366,N_6350);
xor U6481 (N_6481,N_6388,N_6242);
xnor U6482 (N_6482,N_6219,N_6261);
and U6483 (N_6483,N_6322,N_6349);
and U6484 (N_6484,N_6399,N_6287);
nand U6485 (N_6485,N_6243,N_6360);
and U6486 (N_6486,N_6331,N_6272);
nand U6487 (N_6487,N_6398,N_6304);
or U6488 (N_6488,N_6286,N_6217);
or U6489 (N_6489,N_6235,N_6365);
nand U6490 (N_6490,N_6244,N_6347);
nand U6491 (N_6491,N_6264,N_6333);
or U6492 (N_6492,N_6220,N_6385);
or U6493 (N_6493,N_6301,N_6346);
or U6494 (N_6494,N_6210,N_6303);
and U6495 (N_6495,N_6378,N_6215);
and U6496 (N_6496,N_6256,N_6209);
nor U6497 (N_6497,N_6305,N_6375);
and U6498 (N_6498,N_6249,N_6295);
nand U6499 (N_6499,N_6344,N_6266);
or U6500 (N_6500,N_6342,N_6245);
and U6501 (N_6501,N_6209,N_6284);
nor U6502 (N_6502,N_6343,N_6262);
xor U6503 (N_6503,N_6388,N_6385);
nand U6504 (N_6504,N_6226,N_6245);
or U6505 (N_6505,N_6253,N_6349);
or U6506 (N_6506,N_6311,N_6262);
nand U6507 (N_6507,N_6203,N_6387);
or U6508 (N_6508,N_6319,N_6345);
nand U6509 (N_6509,N_6272,N_6355);
nand U6510 (N_6510,N_6242,N_6228);
xnor U6511 (N_6511,N_6357,N_6364);
nor U6512 (N_6512,N_6255,N_6259);
nor U6513 (N_6513,N_6366,N_6218);
nor U6514 (N_6514,N_6207,N_6344);
nor U6515 (N_6515,N_6385,N_6395);
or U6516 (N_6516,N_6303,N_6217);
nand U6517 (N_6517,N_6372,N_6237);
and U6518 (N_6518,N_6299,N_6303);
xnor U6519 (N_6519,N_6269,N_6307);
and U6520 (N_6520,N_6346,N_6322);
or U6521 (N_6521,N_6205,N_6320);
or U6522 (N_6522,N_6317,N_6258);
nand U6523 (N_6523,N_6204,N_6211);
nand U6524 (N_6524,N_6210,N_6255);
nor U6525 (N_6525,N_6215,N_6250);
nor U6526 (N_6526,N_6309,N_6349);
nand U6527 (N_6527,N_6363,N_6205);
xor U6528 (N_6528,N_6295,N_6217);
nor U6529 (N_6529,N_6243,N_6251);
or U6530 (N_6530,N_6315,N_6260);
or U6531 (N_6531,N_6205,N_6287);
nand U6532 (N_6532,N_6218,N_6377);
and U6533 (N_6533,N_6232,N_6222);
nand U6534 (N_6534,N_6386,N_6288);
nand U6535 (N_6535,N_6264,N_6341);
and U6536 (N_6536,N_6366,N_6242);
nor U6537 (N_6537,N_6396,N_6228);
and U6538 (N_6538,N_6399,N_6384);
and U6539 (N_6539,N_6354,N_6209);
or U6540 (N_6540,N_6200,N_6311);
xnor U6541 (N_6541,N_6378,N_6377);
or U6542 (N_6542,N_6292,N_6209);
nor U6543 (N_6543,N_6322,N_6393);
nor U6544 (N_6544,N_6205,N_6226);
xnor U6545 (N_6545,N_6219,N_6267);
nor U6546 (N_6546,N_6297,N_6336);
nor U6547 (N_6547,N_6298,N_6267);
and U6548 (N_6548,N_6292,N_6364);
or U6549 (N_6549,N_6342,N_6282);
or U6550 (N_6550,N_6260,N_6359);
nand U6551 (N_6551,N_6296,N_6202);
and U6552 (N_6552,N_6249,N_6293);
nor U6553 (N_6553,N_6355,N_6338);
xor U6554 (N_6554,N_6325,N_6365);
nor U6555 (N_6555,N_6293,N_6318);
and U6556 (N_6556,N_6337,N_6301);
nor U6557 (N_6557,N_6345,N_6310);
nand U6558 (N_6558,N_6276,N_6286);
nand U6559 (N_6559,N_6291,N_6390);
or U6560 (N_6560,N_6399,N_6338);
or U6561 (N_6561,N_6238,N_6218);
and U6562 (N_6562,N_6378,N_6227);
xnor U6563 (N_6563,N_6351,N_6394);
or U6564 (N_6564,N_6254,N_6239);
or U6565 (N_6565,N_6294,N_6340);
nand U6566 (N_6566,N_6217,N_6323);
or U6567 (N_6567,N_6367,N_6291);
or U6568 (N_6568,N_6259,N_6290);
or U6569 (N_6569,N_6253,N_6310);
or U6570 (N_6570,N_6276,N_6333);
or U6571 (N_6571,N_6330,N_6295);
and U6572 (N_6572,N_6313,N_6393);
or U6573 (N_6573,N_6334,N_6325);
nand U6574 (N_6574,N_6376,N_6341);
nand U6575 (N_6575,N_6342,N_6250);
or U6576 (N_6576,N_6367,N_6299);
xnor U6577 (N_6577,N_6362,N_6318);
nand U6578 (N_6578,N_6207,N_6265);
or U6579 (N_6579,N_6271,N_6221);
nand U6580 (N_6580,N_6372,N_6386);
nor U6581 (N_6581,N_6202,N_6278);
nor U6582 (N_6582,N_6259,N_6369);
nand U6583 (N_6583,N_6381,N_6259);
nor U6584 (N_6584,N_6256,N_6364);
or U6585 (N_6585,N_6289,N_6389);
or U6586 (N_6586,N_6230,N_6344);
nand U6587 (N_6587,N_6266,N_6209);
or U6588 (N_6588,N_6343,N_6387);
or U6589 (N_6589,N_6247,N_6250);
or U6590 (N_6590,N_6346,N_6247);
or U6591 (N_6591,N_6246,N_6268);
xnor U6592 (N_6592,N_6281,N_6339);
or U6593 (N_6593,N_6262,N_6255);
nand U6594 (N_6594,N_6220,N_6342);
and U6595 (N_6595,N_6363,N_6200);
or U6596 (N_6596,N_6289,N_6318);
nor U6597 (N_6597,N_6357,N_6231);
nand U6598 (N_6598,N_6361,N_6365);
nand U6599 (N_6599,N_6385,N_6278);
or U6600 (N_6600,N_6588,N_6412);
nand U6601 (N_6601,N_6478,N_6556);
and U6602 (N_6602,N_6469,N_6500);
and U6603 (N_6603,N_6462,N_6404);
nand U6604 (N_6604,N_6484,N_6436);
or U6605 (N_6605,N_6498,N_6593);
nor U6606 (N_6606,N_6485,N_6482);
nand U6607 (N_6607,N_6425,N_6416);
nor U6608 (N_6608,N_6509,N_6580);
or U6609 (N_6609,N_6594,N_6555);
or U6610 (N_6610,N_6584,N_6545);
or U6611 (N_6611,N_6465,N_6502);
nor U6612 (N_6612,N_6558,N_6559);
and U6613 (N_6613,N_6468,N_6449);
and U6614 (N_6614,N_6420,N_6419);
and U6615 (N_6615,N_6493,N_6477);
xnor U6616 (N_6616,N_6583,N_6529);
nor U6617 (N_6617,N_6524,N_6410);
or U6618 (N_6618,N_6541,N_6514);
xor U6619 (N_6619,N_6408,N_6472);
or U6620 (N_6620,N_6494,N_6476);
nor U6621 (N_6621,N_6491,N_6573);
nor U6622 (N_6622,N_6461,N_6553);
or U6623 (N_6623,N_6577,N_6546);
or U6624 (N_6624,N_6532,N_6599);
nor U6625 (N_6625,N_6483,N_6400);
nor U6626 (N_6626,N_6522,N_6411);
nor U6627 (N_6627,N_6505,N_6456);
or U6628 (N_6628,N_6422,N_6525);
nor U6629 (N_6629,N_6473,N_6442);
xor U6630 (N_6630,N_6474,N_6579);
nor U6631 (N_6631,N_6513,N_6592);
nand U6632 (N_6632,N_6459,N_6575);
and U6633 (N_6633,N_6569,N_6572);
nand U6634 (N_6634,N_6551,N_6479);
and U6635 (N_6635,N_6518,N_6512);
nor U6636 (N_6636,N_6455,N_6538);
nand U6637 (N_6637,N_6451,N_6424);
xor U6638 (N_6638,N_6535,N_6453);
or U6639 (N_6639,N_6571,N_6433);
or U6640 (N_6640,N_6450,N_6501);
or U6641 (N_6641,N_6435,N_6519);
and U6642 (N_6642,N_6511,N_6540);
nor U6643 (N_6643,N_6466,N_6417);
or U6644 (N_6644,N_6457,N_6548);
and U6645 (N_6645,N_6527,N_6486);
and U6646 (N_6646,N_6567,N_6507);
nor U6647 (N_6647,N_6533,N_6528);
and U6648 (N_6648,N_6431,N_6531);
nand U6649 (N_6649,N_6570,N_6547);
xnor U6650 (N_6650,N_6402,N_6508);
or U6651 (N_6651,N_6443,N_6550);
nand U6652 (N_6652,N_6510,N_6471);
or U6653 (N_6653,N_6516,N_6564);
nor U6654 (N_6654,N_6418,N_6561);
nand U6655 (N_6655,N_6409,N_6504);
and U6656 (N_6656,N_6576,N_6565);
xor U6657 (N_6657,N_6578,N_6421);
nor U6658 (N_6658,N_6499,N_6446);
and U6659 (N_6659,N_6497,N_6423);
nand U6660 (N_6660,N_6487,N_6568);
and U6661 (N_6661,N_6595,N_6554);
or U6662 (N_6662,N_6429,N_6536);
xnor U6663 (N_6663,N_6523,N_6437);
nor U6664 (N_6664,N_6426,N_6434);
or U6665 (N_6665,N_6539,N_6521);
or U6666 (N_6666,N_6544,N_6585);
nor U6667 (N_6667,N_6481,N_6427);
nor U6668 (N_6668,N_6444,N_6496);
nand U6669 (N_6669,N_6447,N_6587);
nor U6670 (N_6670,N_6440,N_6407);
or U6671 (N_6671,N_6520,N_6537);
or U6672 (N_6672,N_6503,N_6403);
nor U6673 (N_6673,N_6401,N_6489);
nor U6674 (N_6674,N_6432,N_6495);
nor U6675 (N_6675,N_6463,N_6464);
nor U6676 (N_6676,N_6566,N_6530);
nand U6677 (N_6677,N_6598,N_6590);
nand U6678 (N_6678,N_6414,N_6445);
or U6679 (N_6679,N_6470,N_6517);
or U6680 (N_6680,N_6480,N_6492);
nor U6681 (N_6681,N_6439,N_6589);
and U6682 (N_6682,N_6542,N_6441);
and U6683 (N_6683,N_6458,N_6438);
nand U6684 (N_6684,N_6405,N_6581);
nand U6685 (N_6685,N_6582,N_6596);
or U6686 (N_6686,N_6460,N_6591);
or U6687 (N_6687,N_6563,N_6506);
or U6688 (N_6688,N_6475,N_6413);
nor U6689 (N_6689,N_6562,N_6430);
nor U6690 (N_6690,N_6597,N_6549);
nor U6691 (N_6691,N_6448,N_6415);
nand U6692 (N_6692,N_6428,N_6488);
and U6693 (N_6693,N_6534,N_6543);
nor U6694 (N_6694,N_6552,N_6560);
nand U6695 (N_6695,N_6406,N_6515);
nor U6696 (N_6696,N_6574,N_6526);
nor U6697 (N_6697,N_6454,N_6586);
nor U6698 (N_6698,N_6490,N_6467);
nor U6699 (N_6699,N_6557,N_6452);
or U6700 (N_6700,N_6563,N_6590);
xnor U6701 (N_6701,N_6580,N_6586);
or U6702 (N_6702,N_6458,N_6562);
nor U6703 (N_6703,N_6410,N_6549);
and U6704 (N_6704,N_6433,N_6426);
and U6705 (N_6705,N_6519,N_6441);
nand U6706 (N_6706,N_6411,N_6482);
nor U6707 (N_6707,N_6572,N_6495);
nand U6708 (N_6708,N_6403,N_6558);
and U6709 (N_6709,N_6554,N_6580);
xnor U6710 (N_6710,N_6543,N_6560);
or U6711 (N_6711,N_6444,N_6459);
nand U6712 (N_6712,N_6562,N_6456);
nand U6713 (N_6713,N_6437,N_6410);
and U6714 (N_6714,N_6435,N_6464);
and U6715 (N_6715,N_6502,N_6409);
or U6716 (N_6716,N_6539,N_6550);
nand U6717 (N_6717,N_6559,N_6565);
nor U6718 (N_6718,N_6547,N_6459);
nand U6719 (N_6719,N_6456,N_6569);
nand U6720 (N_6720,N_6456,N_6429);
and U6721 (N_6721,N_6473,N_6531);
and U6722 (N_6722,N_6452,N_6432);
and U6723 (N_6723,N_6505,N_6509);
xnor U6724 (N_6724,N_6423,N_6543);
nor U6725 (N_6725,N_6485,N_6481);
nor U6726 (N_6726,N_6539,N_6564);
xnor U6727 (N_6727,N_6548,N_6420);
nor U6728 (N_6728,N_6481,N_6512);
or U6729 (N_6729,N_6420,N_6402);
xnor U6730 (N_6730,N_6488,N_6496);
nand U6731 (N_6731,N_6545,N_6408);
or U6732 (N_6732,N_6582,N_6484);
and U6733 (N_6733,N_6524,N_6470);
xor U6734 (N_6734,N_6454,N_6572);
nand U6735 (N_6735,N_6589,N_6530);
nor U6736 (N_6736,N_6548,N_6462);
or U6737 (N_6737,N_6401,N_6570);
and U6738 (N_6738,N_6517,N_6430);
or U6739 (N_6739,N_6576,N_6445);
nor U6740 (N_6740,N_6480,N_6577);
and U6741 (N_6741,N_6427,N_6585);
nand U6742 (N_6742,N_6490,N_6410);
and U6743 (N_6743,N_6444,N_6466);
nand U6744 (N_6744,N_6490,N_6496);
and U6745 (N_6745,N_6454,N_6485);
nand U6746 (N_6746,N_6511,N_6565);
nor U6747 (N_6747,N_6473,N_6516);
nand U6748 (N_6748,N_6570,N_6420);
nor U6749 (N_6749,N_6582,N_6495);
nor U6750 (N_6750,N_6534,N_6469);
nand U6751 (N_6751,N_6414,N_6420);
or U6752 (N_6752,N_6498,N_6435);
nand U6753 (N_6753,N_6599,N_6566);
nand U6754 (N_6754,N_6580,N_6555);
nand U6755 (N_6755,N_6590,N_6441);
nor U6756 (N_6756,N_6572,N_6500);
nand U6757 (N_6757,N_6589,N_6468);
nor U6758 (N_6758,N_6510,N_6541);
or U6759 (N_6759,N_6531,N_6472);
nand U6760 (N_6760,N_6541,N_6533);
xor U6761 (N_6761,N_6591,N_6459);
or U6762 (N_6762,N_6416,N_6465);
nor U6763 (N_6763,N_6419,N_6535);
nand U6764 (N_6764,N_6543,N_6521);
nand U6765 (N_6765,N_6447,N_6411);
nor U6766 (N_6766,N_6415,N_6499);
or U6767 (N_6767,N_6562,N_6440);
and U6768 (N_6768,N_6488,N_6454);
nor U6769 (N_6769,N_6537,N_6459);
or U6770 (N_6770,N_6451,N_6519);
or U6771 (N_6771,N_6528,N_6547);
and U6772 (N_6772,N_6463,N_6405);
xnor U6773 (N_6773,N_6432,N_6565);
nor U6774 (N_6774,N_6571,N_6577);
nand U6775 (N_6775,N_6434,N_6576);
nor U6776 (N_6776,N_6424,N_6477);
nor U6777 (N_6777,N_6564,N_6509);
or U6778 (N_6778,N_6551,N_6527);
or U6779 (N_6779,N_6551,N_6594);
or U6780 (N_6780,N_6467,N_6423);
nor U6781 (N_6781,N_6403,N_6453);
nand U6782 (N_6782,N_6575,N_6513);
xnor U6783 (N_6783,N_6556,N_6598);
xor U6784 (N_6784,N_6498,N_6580);
and U6785 (N_6785,N_6583,N_6444);
xor U6786 (N_6786,N_6508,N_6580);
or U6787 (N_6787,N_6450,N_6576);
and U6788 (N_6788,N_6549,N_6474);
and U6789 (N_6789,N_6403,N_6588);
and U6790 (N_6790,N_6420,N_6499);
nand U6791 (N_6791,N_6516,N_6551);
xor U6792 (N_6792,N_6529,N_6596);
nor U6793 (N_6793,N_6537,N_6441);
nor U6794 (N_6794,N_6590,N_6455);
and U6795 (N_6795,N_6599,N_6402);
or U6796 (N_6796,N_6449,N_6506);
nor U6797 (N_6797,N_6463,N_6498);
and U6798 (N_6798,N_6403,N_6561);
nand U6799 (N_6799,N_6489,N_6502);
and U6800 (N_6800,N_6679,N_6753);
nand U6801 (N_6801,N_6699,N_6653);
or U6802 (N_6802,N_6621,N_6669);
or U6803 (N_6803,N_6768,N_6761);
and U6804 (N_6804,N_6623,N_6637);
nand U6805 (N_6805,N_6723,N_6718);
nor U6806 (N_6806,N_6703,N_6722);
nand U6807 (N_6807,N_6784,N_6698);
nor U6808 (N_6808,N_6724,N_6656);
and U6809 (N_6809,N_6757,N_6765);
nand U6810 (N_6810,N_6790,N_6687);
nor U6811 (N_6811,N_6631,N_6689);
xor U6812 (N_6812,N_6685,N_6763);
or U6813 (N_6813,N_6683,N_6707);
or U6814 (N_6814,N_6785,N_6636);
and U6815 (N_6815,N_6600,N_6727);
and U6816 (N_6816,N_6728,N_6684);
or U6817 (N_6817,N_6688,N_6791);
xnor U6818 (N_6818,N_6779,N_6759);
and U6819 (N_6819,N_6675,N_6682);
nand U6820 (N_6820,N_6674,N_6788);
nor U6821 (N_6821,N_6767,N_6694);
and U6822 (N_6822,N_6643,N_6617);
nand U6823 (N_6823,N_6787,N_6701);
or U6824 (N_6824,N_6678,N_6601);
nand U6825 (N_6825,N_6622,N_6745);
nand U6826 (N_6826,N_6642,N_6792);
or U6827 (N_6827,N_6746,N_6705);
or U6828 (N_6828,N_6750,N_6664);
nand U6829 (N_6829,N_6609,N_6650);
nor U6830 (N_6830,N_6681,N_6704);
xor U6831 (N_6831,N_6747,N_6624);
nand U6832 (N_6832,N_6794,N_6644);
or U6833 (N_6833,N_6676,N_6645);
nor U6834 (N_6834,N_6696,N_6741);
or U6835 (N_6835,N_6708,N_6630);
or U6836 (N_6836,N_6693,N_6734);
and U6837 (N_6837,N_6690,N_6720);
or U6838 (N_6838,N_6796,N_6719);
nor U6839 (N_6839,N_6615,N_6772);
nand U6840 (N_6840,N_6655,N_6737);
xnor U6841 (N_6841,N_6602,N_6700);
nor U6842 (N_6842,N_6660,N_6668);
or U6843 (N_6843,N_6692,N_6752);
xnor U6844 (N_6844,N_6775,N_6658);
nor U6845 (N_6845,N_6610,N_6786);
and U6846 (N_6846,N_6721,N_6799);
and U6847 (N_6847,N_6716,N_6762);
or U6848 (N_6848,N_6742,N_6638);
nor U6849 (N_6849,N_6639,N_6625);
and U6850 (N_6850,N_6628,N_6611);
or U6851 (N_6851,N_6738,N_6697);
or U6852 (N_6852,N_6773,N_6717);
or U6853 (N_6853,N_6603,N_6733);
nor U6854 (N_6854,N_6735,N_6795);
and U6855 (N_6855,N_6648,N_6783);
and U6856 (N_6856,N_6756,N_6743);
nor U6857 (N_6857,N_6652,N_6782);
nand U6858 (N_6858,N_6758,N_6729);
or U6859 (N_6859,N_6618,N_6730);
and U6860 (N_6860,N_6647,N_6726);
xor U6861 (N_6861,N_6736,N_6793);
nand U6862 (N_6862,N_6691,N_6608);
and U6863 (N_6863,N_6731,N_6654);
or U6864 (N_6864,N_6626,N_6619);
nor U6865 (N_6865,N_6725,N_6633);
nor U6866 (N_6866,N_6777,N_6672);
and U6867 (N_6867,N_6686,N_6641);
or U6868 (N_6868,N_6709,N_6760);
or U6869 (N_6869,N_6706,N_6713);
xnor U6870 (N_6870,N_6635,N_6614);
or U6871 (N_6871,N_6695,N_6661);
nor U6872 (N_6872,N_6606,N_6778);
or U6873 (N_6873,N_6677,N_6646);
nand U6874 (N_6874,N_6616,N_6755);
or U6875 (N_6875,N_6754,N_6680);
nor U6876 (N_6876,N_6774,N_6781);
xor U6877 (N_6877,N_6749,N_6640);
or U6878 (N_6878,N_6673,N_6607);
nand U6879 (N_6879,N_6751,N_6766);
nor U6880 (N_6880,N_6605,N_6780);
nor U6881 (N_6881,N_6659,N_6744);
nor U6882 (N_6882,N_6665,N_6629);
xnor U6883 (N_6883,N_6612,N_6620);
nand U6884 (N_6884,N_6649,N_6667);
nor U6885 (N_6885,N_6702,N_6604);
nand U6886 (N_6886,N_6714,N_6627);
and U6887 (N_6887,N_6613,N_6798);
and U6888 (N_6888,N_6651,N_6634);
nor U6889 (N_6889,N_6764,N_6740);
nor U6890 (N_6890,N_6769,N_6712);
or U6891 (N_6891,N_6770,N_6771);
and U6892 (N_6892,N_6657,N_6748);
nand U6893 (N_6893,N_6739,N_6670);
nor U6894 (N_6894,N_6663,N_6662);
xnor U6895 (N_6895,N_6711,N_6632);
or U6896 (N_6896,N_6797,N_6710);
and U6897 (N_6897,N_6732,N_6776);
nand U6898 (N_6898,N_6671,N_6666);
nor U6899 (N_6899,N_6715,N_6789);
or U6900 (N_6900,N_6637,N_6735);
nor U6901 (N_6901,N_6635,N_6637);
nor U6902 (N_6902,N_6697,N_6764);
xor U6903 (N_6903,N_6641,N_6699);
and U6904 (N_6904,N_6742,N_6619);
xnor U6905 (N_6905,N_6622,N_6609);
or U6906 (N_6906,N_6689,N_6742);
nand U6907 (N_6907,N_6615,N_6725);
and U6908 (N_6908,N_6699,N_6705);
xor U6909 (N_6909,N_6749,N_6618);
and U6910 (N_6910,N_6716,N_6628);
or U6911 (N_6911,N_6742,N_6672);
xor U6912 (N_6912,N_6645,N_6677);
xor U6913 (N_6913,N_6713,N_6649);
or U6914 (N_6914,N_6753,N_6638);
nand U6915 (N_6915,N_6612,N_6763);
and U6916 (N_6916,N_6659,N_6757);
nor U6917 (N_6917,N_6650,N_6664);
or U6918 (N_6918,N_6718,N_6763);
and U6919 (N_6919,N_6686,N_6700);
nand U6920 (N_6920,N_6668,N_6657);
and U6921 (N_6921,N_6746,N_6718);
or U6922 (N_6922,N_6754,N_6747);
and U6923 (N_6923,N_6798,N_6647);
and U6924 (N_6924,N_6731,N_6745);
nor U6925 (N_6925,N_6669,N_6789);
nor U6926 (N_6926,N_6612,N_6648);
or U6927 (N_6927,N_6734,N_6781);
or U6928 (N_6928,N_6643,N_6655);
nor U6929 (N_6929,N_6696,N_6733);
nand U6930 (N_6930,N_6661,N_6787);
and U6931 (N_6931,N_6738,N_6769);
or U6932 (N_6932,N_6791,N_6638);
and U6933 (N_6933,N_6610,N_6717);
or U6934 (N_6934,N_6601,N_6750);
nor U6935 (N_6935,N_6669,N_6746);
nand U6936 (N_6936,N_6793,N_6729);
nand U6937 (N_6937,N_6751,N_6784);
and U6938 (N_6938,N_6616,N_6721);
and U6939 (N_6939,N_6715,N_6637);
nand U6940 (N_6940,N_6679,N_6668);
and U6941 (N_6941,N_6710,N_6685);
nand U6942 (N_6942,N_6654,N_6672);
nor U6943 (N_6943,N_6706,N_6672);
nand U6944 (N_6944,N_6749,N_6677);
nand U6945 (N_6945,N_6725,N_6670);
or U6946 (N_6946,N_6636,N_6655);
and U6947 (N_6947,N_6702,N_6681);
and U6948 (N_6948,N_6641,N_6670);
nand U6949 (N_6949,N_6757,N_6602);
nand U6950 (N_6950,N_6619,N_6715);
nand U6951 (N_6951,N_6663,N_6792);
xnor U6952 (N_6952,N_6765,N_6605);
or U6953 (N_6953,N_6647,N_6707);
nand U6954 (N_6954,N_6614,N_6693);
nand U6955 (N_6955,N_6713,N_6646);
xnor U6956 (N_6956,N_6797,N_6790);
nand U6957 (N_6957,N_6611,N_6691);
nor U6958 (N_6958,N_6719,N_6660);
nand U6959 (N_6959,N_6610,N_6675);
nand U6960 (N_6960,N_6650,N_6639);
and U6961 (N_6961,N_6740,N_6620);
or U6962 (N_6962,N_6764,N_6631);
nand U6963 (N_6963,N_6609,N_6632);
and U6964 (N_6964,N_6780,N_6618);
or U6965 (N_6965,N_6783,N_6754);
and U6966 (N_6966,N_6774,N_6662);
nand U6967 (N_6967,N_6654,N_6734);
nand U6968 (N_6968,N_6753,N_6636);
nor U6969 (N_6969,N_6652,N_6684);
nor U6970 (N_6970,N_6603,N_6624);
nand U6971 (N_6971,N_6770,N_6787);
and U6972 (N_6972,N_6687,N_6749);
or U6973 (N_6973,N_6688,N_6712);
nand U6974 (N_6974,N_6618,N_6770);
and U6975 (N_6975,N_6691,N_6669);
nand U6976 (N_6976,N_6621,N_6741);
xor U6977 (N_6977,N_6671,N_6723);
nor U6978 (N_6978,N_6601,N_6762);
and U6979 (N_6979,N_6635,N_6668);
or U6980 (N_6980,N_6775,N_6608);
or U6981 (N_6981,N_6699,N_6747);
nand U6982 (N_6982,N_6612,N_6757);
and U6983 (N_6983,N_6734,N_6640);
and U6984 (N_6984,N_6743,N_6782);
or U6985 (N_6985,N_6661,N_6649);
nor U6986 (N_6986,N_6744,N_6650);
nand U6987 (N_6987,N_6607,N_6787);
and U6988 (N_6988,N_6622,N_6786);
nor U6989 (N_6989,N_6778,N_6779);
or U6990 (N_6990,N_6625,N_6605);
nand U6991 (N_6991,N_6747,N_6738);
xor U6992 (N_6992,N_6717,N_6619);
or U6993 (N_6993,N_6708,N_6679);
nand U6994 (N_6994,N_6756,N_6779);
and U6995 (N_6995,N_6724,N_6728);
nor U6996 (N_6996,N_6641,N_6630);
nand U6997 (N_6997,N_6646,N_6672);
nand U6998 (N_6998,N_6709,N_6658);
and U6999 (N_6999,N_6700,N_6762);
or U7000 (N_7000,N_6843,N_6897);
or U7001 (N_7001,N_6802,N_6960);
and U7002 (N_7002,N_6906,N_6825);
or U7003 (N_7003,N_6890,N_6929);
and U7004 (N_7004,N_6872,N_6842);
nand U7005 (N_7005,N_6922,N_6923);
or U7006 (N_7006,N_6969,N_6968);
and U7007 (N_7007,N_6862,N_6820);
or U7008 (N_7008,N_6903,N_6954);
nor U7009 (N_7009,N_6803,N_6946);
or U7010 (N_7010,N_6880,N_6902);
and U7011 (N_7011,N_6961,N_6904);
nand U7012 (N_7012,N_6836,N_6984);
and U7013 (N_7013,N_6990,N_6863);
xnor U7014 (N_7014,N_6936,N_6896);
and U7015 (N_7015,N_6943,N_6833);
nor U7016 (N_7016,N_6881,N_6933);
and U7017 (N_7017,N_6875,N_6972);
or U7018 (N_7018,N_6959,N_6870);
xor U7019 (N_7019,N_6938,N_6812);
nand U7020 (N_7020,N_6884,N_6999);
xor U7021 (N_7021,N_6895,N_6966);
or U7022 (N_7022,N_6971,N_6994);
xnor U7023 (N_7023,N_6924,N_6981);
or U7024 (N_7024,N_6908,N_6907);
nor U7025 (N_7025,N_6829,N_6837);
nor U7026 (N_7026,N_6920,N_6914);
and U7027 (N_7027,N_6921,N_6830);
or U7028 (N_7028,N_6822,N_6985);
nor U7029 (N_7029,N_6974,N_6816);
nor U7030 (N_7030,N_6888,N_6934);
nor U7031 (N_7031,N_6909,N_6824);
or U7032 (N_7032,N_6848,N_6819);
nor U7033 (N_7033,N_6901,N_6852);
nand U7034 (N_7034,N_6814,N_6970);
and U7035 (N_7035,N_6905,N_6885);
nor U7036 (N_7036,N_6965,N_6850);
and U7037 (N_7037,N_6804,N_6826);
nor U7038 (N_7038,N_6913,N_6996);
and U7039 (N_7039,N_6982,N_6979);
nor U7040 (N_7040,N_6879,N_6951);
nand U7041 (N_7041,N_6801,N_6918);
nand U7042 (N_7042,N_6853,N_6944);
or U7043 (N_7043,N_6956,N_6932);
and U7044 (N_7044,N_6937,N_6939);
nand U7045 (N_7045,N_6839,N_6856);
or U7046 (N_7046,N_6807,N_6838);
xnor U7047 (N_7047,N_6886,N_6991);
and U7048 (N_7048,N_6935,N_6992);
or U7049 (N_7049,N_6864,N_6846);
and U7050 (N_7050,N_6834,N_6989);
and U7051 (N_7051,N_6827,N_6831);
nor U7052 (N_7052,N_6806,N_6868);
and U7053 (N_7053,N_6894,N_6874);
nor U7054 (N_7054,N_6912,N_6997);
and U7055 (N_7055,N_6917,N_6861);
and U7056 (N_7056,N_6995,N_6947);
or U7057 (N_7057,N_6962,N_6821);
and U7058 (N_7058,N_6915,N_6987);
nor U7059 (N_7059,N_6840,N_6916);
or U7060 (N_7060,N_6805,N_6855);
nor U7061 (N_7061,N_6986,N_6851);
and U7062 (N_7062,N_6873,N_6832);
nor U7063 (N_7063,N_6849,N_6823);
xnor U7064 (N_7064,N_6871,N_6828);
and U7065 (N_7065,N_6898,N_6977);
nand U7066 (N_7066,N_6811,N_6891);
or U7067 (N_7067,N_6931,N_6963);
or U7068 (N_7068,N_6865,N_6930);
or U7069 (N_7069,N_6967,N_6813);
or U7070 (N_7070,N_6877,N_6955);
nor U7071 (N_7071,N_6800,N_6857);
xnor U7072 (N_7072,N_6808,N_6949);
nor U7073 (N_7073,N_6809,N_6998);
nand U7074 (N_7074,N_6940,N_6815);
nand U7075 (N_7075,N_6957,N_6878);
nand U7076 (N_7076,N_6919,N_6844);
xnor U7077 (N_7077,N_6860,N_6818);
or U7078 (N_7078,N_6900,N_6975);
nand U7079 (N_7079,N_6928,N_6942);
or U7080 (N_7080,N_6952,N_6835);
and U7081 (N_7081,N_6953,N_6973);
and U7082 (N_7082,N_6910,N_6950);
nor U7083 (N_7083,N_6887,N_6892);
nand U7084 (N_7084,N_6958,N_6976);
and U7085 (N_7085,N_6927,N_6964);
nor U7086 (N_7086,N_6893,N_6983);
nand U7087 (N_7087,N_6847,N_6876);
nor U7088 (N_7088,N_6926,N_6899);
or U7089 (N_7089,N_6867,N_6945);
or U7090 (N_7090,N_6988,N_6911);
and U7091 (N_7091,N_6980,N_6858);
or U7092 (N_7092,N_6993,N_6882);
nor U7093 (N_7093,N_6854,N_6941);
nand U7094 (N_7094,N_6866,N_6845);
xor U7095 (N_7095,N_6948,N_6841);
and U7096 (N_7096,N_6889,N_6817);
xor U7097 (N_7097,N_6859,N_6883);
and U7098 (N_7098,N_6810,N_6925);
nand U7099 (N_7099,N_6869,N_6978);
or U7100 (N_7100,N_6935,N_6821);
nor U7101 (N_7101,N_6922,N_6970);
nand U7102 (N_7102,N_6946,N_6857);
nor U7103 (N_7103,N_6958,N_6913);
nor U7104 (N_7104,N_6883,N_6981);
or U7105 (N_7105,N_6926,N_6803);
nand U7106 (N_7106,N_6955,N_6950);
nand U7107 (N_7107,N_6930,N_6947);
and U7108 (N_7108,N_6894,N_6896);
nand U7109 (N_7109,N_6943,N_6980);
nand U7110 (N_7110,N_6917,N_6821);
or U7111 (N_7111,N_6965,N_6918);
or U7112 (N_7112,N_6949,N_6859);
and U7113 (N_7113,N_6810,N_6867);
or U7114 (N_7114,N_6864,N_6982);
and U7115 (N_7115,N_6939,N_6867);
and U7116 (N_7116,N_6895,N_6865);
nor U7117 (N_7117,N_6867,N_6898);
and U7118 (N_7118,N_6924,N_6813);
nand U7119 (N_7119,N_6958,N_6827);
nand U7120 (N_7120,N_6948,N_6875);
and U7121 (N_7121,N_6855,N_6916);
and U7122 (N_7122,N_6968,N_6932);
and U7123 (N_7123,N_6884,N_6982);
or U7124 (N_7124,N_6823,N_6992);
or U7125 (N_7125,N_6891,N_6967);
and U7126 (N_7126,N_6924,N_6889);
or U7127 (N_7127,N_6900,N_6904);
nor U7128 (N_7128,N_6880,N_6843);
or U7129 (N_7129,N_6965,N_6969);
or U7130 (N_7130,N_6890,N_6820);
xnor U7131 (N_7131,N_6995,N_6850);
or U7132 (N_7132,N_6974,N_6814);
nand U7133 (N_7133,N_6958,N_6841);
nand U7134 (N_7134,N_6913,N_6995);
nand U7135 (N_7135,N_6971,N_6841);
and U7136 (N_7136,N_6939,N_6922);
and U7137 (N_7137,N_6903,N_6806);
nor U7138 (N_7138,N_6992,N_6885);
nand U7139 (N_7139,N_6974,N_6955);
nand U7140 (N_7140,N_6995,N_6849);
or U7141 (N_7141,N_6868,N_6876);
nor U7142 (N_7142,N_6949,N_6946);
xor U7143 (N_7143,N_6988,N_6953);
or U7144 (N_7144,N_6812,N_6886);
and U7145 (N_7145,N_6957,N_6920);
xnor U7146 (N_7146,N_6934,N_6800);
or U7147 (N_7147,N_6983,N_6895);
nand U7148 (N_7148,N_6819,N_6961);
nor U7149 (N_7149,N_6804,N_6835);
xnor U7150 (N_7150,N_6820,N_6959);
and U7151 (N_7151,N_6989,N_6916);
or U7152 (N_7152,N_6900,N_6960);
or U7153 (N_7153,N_6940,N_6882);
nor U7154 (N_7154,N_6810,N_6923);
and U7155 (N_7155,N_6822,N_6834);
and U7156 (N_7156,N_6927,N_6892);
or U7157 (N_7157,N_6802,N_6886);
and U7158 (N_7158,N_6952,N_6851);
or U7159 (N_7159,N_6920,N_6804);
and U7160 (N_7160,N_6900,N_6952);
nand U7161 (N_7161,N_6940,N_6833);
nor U7162 (N_7162,N_6826,N_6811);
nor U7163 (N_7163,N_6867,N_6845);
nand U7164 (N_7164,N_6905,N_6895);
xnor U7165 (N_7165,N_6926,N_6881);
and U7166 (N_7166,N_6894,N_6910);
or U7167 (N_7167,N_6904,N_6910);
nor U7168 (N_7168,N_6841,N_6801);
nor U7169 (N_7169,N_6853,N_6875);
nor U7170 (N_7170,N_6998,N_6822);
and U7171 (N_7171,N_6902,N_6800);
and U7172 (N_7172,N_6820,N_6844);
or U7173 (N_7173,N_6916,N_6800);
or U7174 (N_7174,N_6802,N_6917);
nand U7175 (N_7175,N_6836,N_6838);
and U7176 (N_7176,N_6862,N_6892);
and U7177 (N_7177,N_6866,N_6900);
and U7178 (N_7178,N_6942,N_6845);
nand U7179 (N_7179,N_6862,N_6897);
nor U7180 (N_7180,N_6961,N_6815);
nor U7181 (N_7181,N_6868,N_6904);
or U7182 (N_7182,N_6875,N_6861);
nand U7183 (N_7183,N_6876,N_6999);
or U7184 (N_7184,N_6820,N_6955);
nor U7185 (N_7185,N_6898,N_6829);
nand U7186 (N_7186,N_6802,N_6928);
and U7187 (N_7187,N_6814,N_6830);
nor U7188 (N_7188,N_6862,N_6902);
and U7189 (N_7189,N_6842,N_6864);
and U7190 (N_7190,N_6899,N_6998);
or U7191 (N_7191,N_6879,N_6825);
and U7192 (N_7192,N_6855,N_6914);
nor U7193 (N_7193,N_6931,N_6955);
nor U7194 (N_7194,N_6928,N_6876);
or U7195 (N_7195,N_6884,N_6890);
xnor U7196 (N_7196,N_6888,N_6986);
nand U7197 (N_7197,N_6878,N_6997);
or U7198 (N_7198,N_6972,N_6954);
nor U7199 (N_7199,N_6978,N_6834);
and U7200 (N_7200,N_7029,N_7100);
nand U7201 (N_7201,N_7015,N_7175);
or U7202 (N_7202,N_7067,N_7050);
and U7203 (N_7203,N_7032,N_7096);
and U7204 (N_7204,N_7031,N_7071);
or U7205 (N_7205,N_7042,N_7075);
xor U7206 (N_7206,N_7064,N_7146);
and U7207 (N_7207,N_7144,N_7035);
and U7208 (N_7208,N_7091,N_7123);
and U7209 (N_7209,N_7151,N_7170);
nand U7210 (N_7210,N_7113,N_7198);
nand U7211 (N_7211,N_7177,N_7078);
and U7212 (N_7212,N_7045,N_7041);
or U7213 (N_7213,N_7109,N_7011);
xnor U7214 (N_7214,N_7187,N_7025);
nand U7215 (N_7215,N_7046,N_7087);
xor U7216 (N_7216,N_7149,N_7010);
nand U7217 (N_7217,N_7199,N_7107);
nand U7218 (N_7218,N_7085,N_7058);
xnor U7219 (N_7219,N_7108,N_7018);
nor U7220 (N_7220,N_7157,N_7000);
or U7221 (N_7221,N_7008,N_7150);
nor U7222 (N_7222,N_7145,N_7083);
and U7223 (N_7223,N_7072,N_7136);
or U7224 (N_7224,N_7047,N_7112);
nor U7225 (N_7225,N_7158,N_7188);
and U7226 (N_7226,N_7094,N_7054);
nor U7227 (N_7227,N_7048,N_7102);
nand U7228 (N_7228,N_7126,N_7111);
nor U7229 (N_7229,N_7160,N_7086);
or U7230 (N_7230,N_7174,N_7081);
or U7231 (N_7231,N_7129,N_7153);
nor U7232 (N_7232,N_7180,N_7004);
nor U7233 (N_7233,N_7074,N_7166);
nand U7234 (N_7234,N_7117,N_7159);
nor U7235 (N_7235,N_7125,N_7131);
or U7236 (N_7236,N_7043,N_7060);
and U7237 (N_7237,N_7140,N_7038);
nor U7238 (N_7238,N_7190,N_7070);
and U7239 (N_7239,N_7089,N_7092);
xor U7240 (N_7240,N_7186,N_7103);
and U7241 (N_7241,N_7055,N_7051);
or U7242 (N_7242,N_7127,N_7168);
and U7243 (N_7243,N_7154,N_7147);
or U7244 (N_7244,N_7104,N_7026);
and U7245 (N_7245,N_7195,N_7196);
and U7246 (N_7246,N_7013,N_7016);
nand U7247 (N_7247,N_7143,N_7114);
xnor U7248 (N_7248,N_7115,N_7155);
nor U7249 (N_7249,N_7057,N_7105);
nand U7250 (N_7250,N_7189,N_7152);
and U7251 (N_7251,N_7193,N_7183);
nand U7252 (N_7252,N_7110,N_7121);
or U7253 (N_7253,N_7028,N_7039);
nand U7254 (N_7254,N_7068,N_7024);
or U7255 (N_7255,N_7095,N_7002);
nand U7256 (N_7256,N_7132,N_7080);
and U7257 (N_7257,N_7098,N_7017);
and U7258 (N_7258,N_7148,N_7012);
xor U7259 (N_7259,N_7137,N_7122);
nor U7260 (N_7260,N_7181,N_7061);
nand U7261 (N_7261,N_7176,N_7101);
nand U7262 (N_7262,N_7118,N_7079);
nor U7263 (N_7263,N_7056,N_7184);
nor U7264 (N_7264,N_7093,N_7178);
xnor U7265 (N_7265,N_7120,N_7073);
or U7266 (N_7266,N_7171,N_7052);
or U7267 (N_7267,N_7116,N_7040);
nand U7268 (N_7268,N_7030,N_7133);
and U7269 (N_7269,N_7049,N_7192);
xnor U7270 (N_7270,N_7169,N_7076);
xnor U7271 (N_7271,N_7006,N_7007);
nor U7272 (N_7272,N_7001,N_7138);
nor U7273 (N_7273,N_7197,N_7179);
nor U7274 (N_7274,N_7097,N_7088);
nor U7275 (N_7275,N_7053,N_7005);
or U7276 (N_7276,N_7161,N_7141);
and U7277 (N_7277,N_7020,N_7191);
nand U7278 (N_7278,N_7065,N_7069);
and U7279 (N_7279,N_7037,N_7156);
nand U7280 (N_7280,N_7062,N_7135);
and U7281 (N_7281,N_7130,N_7139);
nor U7282 (N_7282,N_7082,N_7084);
nand U7283 (N_7283,N_7036,N_7119);
nand U7284 (N_7284,N_7134,N_7090);
or U7285 (N_7285,N_7023,N_7142);
nand U7286 (N_7286,N_7128,N_7167);
and U7287 (N_7287,N_7022,N_7019);
nor U7288 (N_7288,N_7182,N_7194);
nor U7289 (N_7289,N_7014,N_7106);
xnor U7290 (N_7290,N_7063,N_7066);
nor U7291 (N_7291,N_7027,N_7172);
and U7292 (N_7292,N_7124,N_7099);
nand U7293 (N_7293,N_7185,N_7173);
and U7294 (N_7294,N_7163,N_7021);
or U7295 (N_7295,N_7059,N_7009);
and U7296 (N_7296,N_7033,N_7164);
nand U7297 (N_7297,N_7162,N_7165);
and U7298 (N_7298,N_7044,N_7034);
nand U7299 (N_7299,N_7003,N_7077);
xnor U7300 (N_7300,N_7015,N_7174);
xor U7301 (N_7301,N_7129,N_7021);
nor U7302 (N_7302,N_7044,N_7119);
and U7303 (N_7303,N_7145,N_7001);
or U7304 (N_7304,N_7082,N_7168);
or U7305 (N_7305,N_7137,N_7125);
or U7306 (N_7306,N_7044,N_7078);
or U7307 (N_7307,N_7064,N_7112);
or U7308 (N_7308,N_7017,N_7050);
nand U7309 (N_7309,N_7149,N_7067);
nor U7310 (N_7310,N_7124,N_7110);
nand U7311 (N_7311,N_7067,N_7154);
nand U7312 (N_7312,N_7025,N_7193);
nor U7313 (N_7313,N_7130,N_7100);
nor U7314 (N_7314,N_7044,N_7036);
and U7315 (N_7315,N_7025,N_7022);
xor U7316 (N_7316,N_7080,N_7059);
or U7317 (N_7317,N_7031,N_7057);
nor U7318 (N_7318,N_7088,N_7101);
and U7319 (N_7319,N_7170,N_7012);
nor U7320 (N_7320,N_7140,N_7058);
nand U7321 (N_7321,N_7076,N_7070);
nand U7322 (N_7322,N_7064,N_7046);
nor U7323 (N_7323,N_7001,N_7125);
nand U7324 (N_7324,N_7083,N_7059);
nor U7325 (N_7325,N_7097,N_7058);
or U7326 (N_7326,N_7046,N_7133);
and U7327 (N_7327,N_7130,N_7120);
or U7328 (N_7328,N_7070,N_7122);
nor U7329 (N_7329,N_7118,N_7061);
nand U7330 (N_7330,N_7005,N_7021);
or U7331 (N_7331,N_7118,N_7179);
xor U7332 (N_7332,N_7163,N_7169);
or U7333 (N_7333,N_7136,N_7043);
nand U7334 (N_7334,N_7071,N_7151);
or U7335 (N_7335,N_7152,N_7180);
nor U7336 (N_7336,N_7161,N_7102);
xor U7337 (N_7337,N_7032,N_7144);
nor U7338 (N_7338,N_7117,N_7134);
nor U7339 (N_7339,N_7019,N_7182);
nand U7340 (N_7340,N_7025,N_7148);
or U7341 (N_7341,N_7052,N_7035);
nor U7342 (N_7342,N_7009,N_7128);
or U7343 (N_7343,N_7049,N_7012);
nand U7344 (N_7344,N_7123,N_7041);
nand U7345 (N_7345,N_7015,N_7073);
nand U7346 (N_7346,N_7071,N_7022);
and U7347 (N_7347,N_7043,N_7106);
and U7348 (N_7348,N_7028,N_7023);
or U7349 (N_7349,N_7062,N_7019);
nand U7350 (N_7350,N_7171,N_7172);
and U7351 (N_7351,N_7090,N_7045);
and U7352 (N_7352,N_7130,N_7020);
nor U7353 (N_7353,N_7098,N_7149);
nand U7354 (N_7354,N_7027,N_7183);
nor U7355 (N_7355,N_7134,N_7140);
nor U7356 (N_7356,N_7084,N_7113);
nor U7357 (N_7357,N_7046,N_7116);
nor U7358 (N_7358,N_7188,N_7156);
and U7359 (N_7359,N_7171,N_7014);
xor U7360 (N_7360,N_7064,N_7185);
and U7361 (N_7361,N_7158,N_7035);
and U7362 (N_7362,N_7016,N_7080);
and U7363 (N_7363,N_7081,N_7087);
xor U7364 (N_7364,N_7156,N_7116);
nand U7365 (N_7365,N_7087,N_7187);
xor U7366 (N_7366,N_7016,N_7122);
and U7367 (N_7367,N_7075,N_7141);
and U7368 (N_7368,N_7082,N_7095);
nand U7369 (N_7369,N_7008,N_7130);
nor U7370 (N_7370,N_7168,N_7088);
nor U7371 (N_7371,N_7136,N_7156);
nor U7372 (N_7372,N_7064,N_7022);
nand U7373 (N_7373,N_7198,N_7127);
and U7374 (N_7374,N_7090,N_7165);
and U7375 (N_7375,N_7021,N_7102);
and U7376 (N_7376,N_7080,N_7085);
xnor U7377 (N_7377,N_7138,N_7101);
or U7378 (N_7378,N_7196,N_7128);
nor U7379 (N_7379,N_7157,N_7087);
or U7380 (N_7380,N_7139,N_7090);
and U7381 (N_7381,N_7052,N_7199);
nor U7382 (N_7382,N_7036,N_7188);
and U7383 (N_7383,N_7083,N_7198);
nor U7384 (N_7384,N_7100,N_7158);
nor U7385 (N_7385,N_7091,N_7153);
or U7386 (N_7386,N_7062,N_7160);
nor U7387 (N_7387,N_7141,N_7098);
or U7388 (N_7388,N_7153,N_7060);
nand U7389 (N_7389,N_7035,N_7061);
or U7390 (N_7390,N_7053,N_7062);
nor U7391 (N_7391,N_7028,N_7021);
or U7392 (N_7392,N_7169,N_7028);
or U7393 (N_7393,N_7092,N_7137);
and U7394 (N_7394,N_7187,N_7073);
and U7395 (N_7395,N_7191,N_7173);
nand U7396 (N_7396,N_7173,N_7152);
or U7397 (N_7397,N_7032,N_7050);
nand U7398 (N_7398,N_7156,N_7032);
and U7399 (N_7399,N_7137,N_7050);
or U7400 (N_7400,N_7268,N_7387);
or U7401 (N_7401,N_7279,N_7215);
nand U7402 (N_7402,N_7216,N_7208);
and U7403 (N_7403,N_7309,N_7220);
nand U7404 (N_7404,N_7255,N_7316);
or U7405 (N_7405,N_7290,N_7313);
and U7406 (N_7406,N_7291,N_7351);
nand U7407 (N_7407,N_7240,N_7259);
or U7408 (N_7408,N_7314,N_7392);
nand U7409 (N_7409,N_7369,N_7366);
nand U7410 (N_7410,N_7306,N_7218);
nand U7411 (N_7411,N_7329,N_7200);
or U7412 (N_7412,N_7398,N_7379);
and U7413 (N_7413,N_7337,N_7353);
or U7414 (N_7414,N_7211,N_7278);
nor U7415 (N_7415,N_7371,N_7356);
nand U7416 (N_7416,N_7342,N_7222);
or U7417 (N_7417,N_7307,N_7280);
or U7418 (N_7418,N_7370,N_7294);
or U7419 (N_7419,N_7274,N_7385);
or U7420 (N_7420,N_7324,N_7299);
nor U7421 (N_7421,N_7272,N_7281);
nor U7422 (N_7422,N_7263,N_7384);
or U7423 (N_7423,N_7288,N_7372);
nand U7424 (N_7424,N_7249,N_7297);
xor U7425 (N_7425,N_7322,N_7214);
nor U7426 (N_7426,N_7245,N_7204);
nand U7427 (N_7427,N_7336,N_7348);
and U7428 (N_7428,N_7358,N_7357);
or U7429 (N_7429,N_7225,N_7292);
and U7430 (N_7430,N_7381,N_7203);
xor U7431 (N_7431,N_7315,N_7303);
nand U7432 (N_7432,N_7248,N_7285);
xor U7433 (N_7433,N_7333,N_7246);
or U7434 (N_7434,N_7340,N_7394);
and U7435 (N_7435,N_7254,N_7219);
and U7436 (N_7436,N_7266,N_7221);
or U7437 (N_7437,N_7383,N_7232);
nor U7438 (N_7438,N_7344,N_7349);
or U7439 (N_7439,N_7326,N_7239);
nor U7440 (N_7440,N_7304,N_7227);
and U7441 (N_7441,N_7296,N_7258);
or U7442 (N_7442,N_7264,N_7390);
or U7443 (N_7443,N_7275,N_7354);
nand U7444 (N_7444,N_7250,N_7312);
or U7445 (N_7445,N_7260,N_7359);
and U7446 (N_7446,N_7380,N_7375);
nand U7447 (N_7447,N_7267,N_7311);
and U7448 (N_7448,N_7271,N_7223);
nor U7449 (N_7449,N_7210,N_7321);
nor U7450 (N_7450,N_7376,N_7335);
nor U7451 (N_7451,N_7345,N_7319);
or U7452 (N_7452,N_7364,N_7338);
nand U7453 (N_7453,N_7201,N_7212);
nor U7454 (N_7454,N_7256,N_7346);
nor U7455 (N_7455,N_7270,N_7238);
or U7456 (N_7456,N_7362,N_7305);
xnor U7457 (N_7457,N_7341,N_7273);
xor U7458 (N_7458,N_7202,N_7393);
and U7459 (N_7459,N_7209,N_7350);
xnor U7460 (N_7460,N_7388,N_7295);
or U7461 (N_7461,N_7378,N_7284);
and U7462 (N_7462,N_7399,N_7352);
nor U7463 (N_7463,N_7287,N_7343);
nand U7464 (N_7464,N_7365,N_7332);
nor U7465 (N_7465,N_7396,N_7377);
or U7466 (N_7466,N_7247,N_7205);
or U7467 (N_7467,N_7301,N_7241);
nor U7468 (N_7468,N_7234,N_7286);
nand U7469 (N_7469,N_7317,N_7373);
xor U7470 (N_7470,N_7233,N_7213);
nor U7471 (N_7471,N_7374,N_7360);
or U7472 (N_7472,N_7323,N_7327);
nor U7473 (N_7473,N_7265,N_7308);
nand U7474 (N_7474,N_7217,N_7318);
xor U7475 (N_7475,N_7235,N_7236);
nand U7476 (N_7476,N_7328,N_7206);
or U7477 (N_7477,N_7251,N_7325);
nor U7478 (N_7478,N_7389,N_7368);
nor U7479 (N_7479,N_7386,N_7334);
nor U7480 (N_7480,N_7230,N_7257);
nor U7481 (N_7481,N_7331,N_7229);
xor U7482 (N_7482,N_7382,N_7339);
nor U7483 (N_7483,N_7228,N_7361);
or U7484 (N_7484,N_7237,N_7397);
nor U7485 (N_7485,N_7262,N_7289);
or U7486 (N_7486,N_7347,N_7244);
or U7487 (N_7487,N_7253,N_7355);
nand U7488 (N_7488,N_7277,N_7207);
nor U7489 (N_7489,N_7320,N_7261);
or U7490 (N_7490,N_7293,N_7242);
nand U7491 (N_7491,N_7395,N_7283);
and U7492 (N_7492,N_7224,N_7231);
nor U7493 (N_7493,N_7226,N_7269);
or U7494 (N_7494,N_7276,N_7363);
and U7495 (N_7495,N_7310,N_7302);
and U7496 (N_7496,N_7282,N_7243);
nand U7497 (N_7497,N_7330,N_7300);
nand U7498 (N_7498,N_7367,N_7298);
nor U7499 (N_7499,N_7252,N_7391);
or U7500 (N_7500,N_7236,N_7285);
or U7501 (N_7501,N_7334,N_7305);
nor U7502 (N_7502,N_7357,N_7250);
nand U7503 (N_7503,N_7339,N_7310);
xnor U7504 (N_7504,N_7233,N_7372);
xnor U7505 (N_7505,N_7326,N_7265);
or U7506 (N_7506,N_7342,N_7360);
nand U7507 (N_7507,N_7242,N_7334);
or U7508 (N_7508,N_7340,N_7206);
nand U7509 (N_7509,N_7258,N_7208);
and U7510 (N_7510,N_7283,N_7381);
nand U7511 (N_7511,N_7255,N_7229);
or U7512 (N_7512,N_7344,N_7299);
nor U7513 (N_7513,N_7356,N_7201);
and U7514 (N_7514,N_7397,N_7354);
xnor U7515 (N_7515,N_7304,N_7343);
xor U7516 (N_7516,N_7320,N_7209);
xor U7517 (N_7517,N_7348,N_7319);
or U7518 (N_7518,N_7228,N_7354);
or U7519 (N_7519,N_7340,N_7309);
nand U7520 (N_7520,N_7319,N_7218);
and U7521 (N_7521,N_7248,N_7396);
xnor U7522 (N_7522,N_7280,N_7399);
and U7523 (N_7523,N_7336,N_7382);
or U7524 (N_7524,N_7343,N_7333);
and U7525 (N_7525,N_7263,N_7291);
nand U7526 (N_7526,N_7227,N_7325);
and U7527 (N_7527,N_7222,N_7311);
and U7528 (N_7528,N_7326,N_7213);
or U7529 (N_7529,N_7276,N_7391);
nand U7530 (N_7530,N_7225,N_7276);
or U7531 (N_7531,N_7315,N_7389);
and U7532 (N_7532,N_7202,N_7290);
and U7533 (N_7533,N_7288,N_7384);
nand U7534 (N_7534,N_7376,N_7297);
nand U7535 (N_7535,N_7324,N_7336);
and U7536 (N_7536,N_7382,N_7264);
and U7537 (N_7537,N_7364,N_7308);
and U7538 (N_7538,N_7343,N_7212);
nand U7539 (N_7539,N_7285,N_7317);
nor U7540 (N_7540,N_7278,N_7221);
or U7541 (N_7541,N_7298,N_7241);
or U7542 (N_7542,N_7318,N_7255);
and U7543 (N_7543,N_7302,N_7251);
or U7544 (N_7544,N_7280,N_7270);
xnor U7545 (N_7545,N_7395,N_7234);
and U7546 (N_7546,N_7362,N_7216);
and U7547 (N_7547,N_7310,N_7301);
and U7548 (N_7548,N_7304,N_7288);
or U7549 (N_7549,N_7362,N_7377);
and U7550 (N_7550,N_7373,N_7246);
or U7551 (N_7551,N_7397,N_7218);
nor U7552 (N_7552,N_7240,N_7258);
or U7553 (N_7553,N_7347,N_7327);
and U7554 (N_7554,N_7393,N_7251);
nor U7555 (N_7555,N_7279,N_7355);
and U7556 (N_7556,N_7266,N_7296);
or U7557 (N_7557,N_7272,N_7337);
or U7558 (N_7558,N_7228,N_7329);
or U7559 (N_7559,N_7395,N_7352);
and U7560 (N_7560,N_7207,N_7284);
nor U7561 (N_7561,N_7300,N_7288);
or U7562 (N_7562,N_7387,N_7331);
nor U7563 (N_7563,N_7273,N_7250);
and U7564 (N_7564,N_7350,N_7368);
and U7565 (N_7565,N_7315,N_7239);
nor U7566 (N_7566,N_7392,N_7327);
nand U7567 (N_7567,N_7358,N_7331);
or U7568 (N_7568,N_7354,N_7303);
and U7569 (N_7569,N_7279,N_7249);
xnor U7570 (N_7570,N_7393,N_7312);
and U7571 (N_7571,N_7204,N_7332);
nand U7572 (N_7572,N_7223,N_7313);
xor U7573 (N_7573,N_7205,N_7325);
nor U7574 (N_7574,N_7353,N_7399);
or U7575 (N_7575,N_7303,N_7382);
or U7576 (N_7576,N_7241,N_7326);
or U7577 (N_7577,N_7225,N_7239);
nand U7578 (N_7578,N_7247,N_7352);
or U7579 (N_7579,N_7294,N_7285);
or U7580 (N_7580,N_7397,N_7362);
nor U7581 (N_7581,N_7239,N_7378);
xnor U7582 (N_7582,N_7289,N_7290);
and U7583 (N_7583,N_7319,N_7247);
nor U7584 (N_7584,N_7318,N_7264);
and U7585 (N_7585,N_7258,N_7256);
nand U7586 (N_7586,N_7361,N_7364);
or U7587 (N_7587,N_7286,N_7260);
and U7588 (N_7588,N_7217,N_7317);
or U7589 (N_7589,N_7257,N_7365);
nand U7590 (N_7590,N_7361,N_7221);
nor U7591 (N_7591,N_7360,N_7317);
or U7592 (N_7592,N_7398,N_7317);
and U7593 (N_7593,N_7313,N_7285);
or U7594 (N_7594,N_7379,N_7202);
nand U7595 (N_7595,N_7233,N_7298);
and U7596 (N_7596,N_7230,N_7261);
nand U7597 (N_7597,N_7315,N_7282);
nor U7598 (N_7598,N_7359,N_7308);
nor U7599 (N_7599,N_7206,N_7230);
nand U7600 (N_7600,N_7483,N_7436);
or U7601 (N_7601,N_7443,N_7509);
and U7602 (N_7602,N_7441,N_7474);
xor U7603 (N_7603,N_7584,N_7404);
xnor U7604 (N_7604,N_7554,N_7477);
xor U7605 (N_7605,N_7530,N_7598);
xor U7606 (N_7606,N_7550,N_7578);
nor U7607 (N_7607,N_7406,N_7416);
or U7608 (N_7608,N_7494,N_7545);
and U7609 (N_7609,N_7505,N_7454);
and U7610 (N_7610,N_7446,N_7570);
xor U7611 (N_7611,N_7587,N_7520);
and U7612 (N_7612,N_7444,N_7486);
or U7613 (N_7613,N_7424,N_7585);
and U7614 (N_7614,N_7596,N_7498);
xor U7615 (N_7615,N_7423,N_7482);
or U7616 (N_7616,N_7496,N_7525);
nand U7617 (N_7617,N_7572,N_7490);
and U7618 (N_7618,N_7588,N_7434);
or U7619 (N_7619,N_7507,N_7410);
or U7620 (N_7620,N_7564,N_7546);
and U7621 (N_7621,N_7593,N_7480);
or U7622 (N_7622,N_7568,N_7499);
nor U7623 (N_7623,N_7468,N_7551);
or U7624 (N_7624,N_7521,N_7582);
xor U7625 (N_7625,N_7552,N_7581);
and U7626 (N_7626,N_7532,N_7466);
nor U7627 (N_7627,N_7426,N_7541);
nand U7628 (N_7628,N_7481,N_7467);
nor U7629 (N_7629,N_7594,N_7591);
or U7630 (N_7630,N_7538,N_7575);
and U7631 (N_7631,N_7514,N_7543);
nand U7632 (N_7632,N_7409,N_7403);
and U7633 (N_7633,N_7500,N_7449);
xnor U7634 (N_7634,N_7513,N_7430);
nand U7635 (N_7635,N_7524,N_7492);
or U7636 (N_7636,N_7528,N_7579);
or U7637 (N_7637,N_7448,N_7461);
and U7638 (N_7638,N_7501,N_7464);
xor U7639 (N_7639,N_7457,N_7590);
or U7640 (N_7640,N_7566,N_7460);
nand U7641 (N_7641,N_7439,N_7401);
and U7642 (N_7642,N_7567,N_7465);
xnor U7643 (N_7643,N_7418,N_7517);
nor U7644 (N_7644,N_7537,N_7438);
and U7645 (N_7645,N_7479,N_7476);
nor U7646 (N_7646,N_7452,N_7435);
or U7647 (N_7647,N_7565,N_7548);
and U7648 (N_7648,N_7455,N_7447);
or U7649 (N_7649,N_7561,N_7506);
xnor U7650 (N_7650,N_7470,N_7489);
or U7651 (N_7651,N_7433,N_7408);
nand U7652 (N_7652,N_7487,N_7450);
or U7653 (N_7653,N_7415,N_7592);
and U7654 (N_7654,N_7508,N_7456);
nor U7655 (N_7655,N_7534,N_7471);
or U7656 (N_7656,N_7458,N_7493);
and U7657 (N_7657,N_7419,N_7549);
nand U7658 (N_7658,N_7539,N_7445);
nor U7659 (N_7659,N_7533,N_7407);
nor U7660 (N_7660,N_7432,N_7511);
or U7661 (N_7661,N_7428,N_7442);
xor U7662 (N_7662,N_7555,N_7597);
nor U7663 (N_7663,N_7519,N_7557);
and U7664 (N_7664,N_7523,N_7485);
or U7665 (N_7665,N_7580,N_7472);
xor U7666 (N_7666,N_7413,N_7402);
or U7667 (N_7667,N_7583,N_7421);
or U7668 (N_7668,N_7469,N_7558);
xor U7669 (N_7669,N_7497,N_7531);
and U7670 (N_7670,N_7462,N_7495);
and U7671 (N_7671,N_7412,N_7427);
xnor U7672 (N_7672,N_7562,N_7475);
and U7673 (N_7673,N_7518,N_7556);
or U7674 (N_7674,N_7559,N_7515);
nor U7675 (N_7675,N_7414,N_7535);
xnor U7676 (N_7676,N_7503,N_7437);
nand U7677 (N_7677,N_7527,N_7451);
nor U7678 (N_7678,N_7459,N_7573);
nand U7679 (N_7679,N_7577,N_7595);
nor U7680 (N_7680,N_7431,N_7502);
xnor U7681 (N_7681,N_7599,N_7571);
and U7682 (N_7682,N_7512,N_7522);
and U7683 (N_7683,N_7560,N_7488);
nor U7684 (N_7684,N_7422,N_7400);
nand U7685 (N_7685,N_7542,N_7536);
nor U7686 (N_7686,N_7586,N_7491);
nor U7687 (N_7687,N_7510,N_7425);
nand U7688 (N_7688,N_7563,N_7589);
and U7689 (N_7689,N_7405,N_7463);
xnor U7690 (N_7690,N_7553,N_7529);
and U7691 (N_7691,N_7478,N_7473);
xnor U7692 (N_7692,N_7516,N_7417);
or U7693 (N_7693,N_7569,N_7504);
nor U7694 (N_7694,N_7484,N_7411);
or U7695 (N_7695,N_7429,N_7526);
xor U7696 (N_7696,N_7440,N_7544);
or U7697 (N_7697,N_7453,N_7576);
nor U7698 (N_7698,N_7420,N_7547);
nor U7699 (N_7699,N_7574,N_7540);
nand U7700 (N_7700,N_7446,N_7594);
nor U7701 (N_7701,N_7594,N_7538);
nand U7702 (N_7702,N_7569,N_7471);
nand U7703 (N_7703,N_7482,N_7465);
nand U7704 (N_7704,N_7540,N_7584);
and U7705 (N_7705,N_7590,N_7468);
nand U7706 (N_7706,N_7424,N_7512);
xor U7707 (N_7707,N_7431,N_7549);
nand U7708 (N_7708,N_7491,N_7590);
nor U7709 (N_7709,N_7573,N_7470);
xor U7710 (N_7710,N_7564,N_7410);
nand U7711 (N_7711,N_7571,N_7565);
and U7712 (N_7712,N_7560,N_7578);
nor U7713 (N_7713,N_7454,N_7483);
nor U7714 (N_7714,N_7592,N_7499);
nor U7715 (N_7715,N_7413,N_7555);
nor U7716 (N_7716,N_7510,N_7524);
nor U7717 (N_7717,N_7446,N_7533);
xor U7718 (N_7718,N_7431,N_7523);
xor U7719 (N_7719,N_7433,N_7520);
or U7720 (N_7720,N_7482,N_7555);
and U7721 (N_7721,N_7524,N_7462);
nand U7722 (N_7722,N_7509,N_7537);
and U7723 (N_7723,N_7570,N_7415);
and U7724 (N_7724,N_7504,N_7548);
nand U7725 (N_7725,N_7443,N_7480);
or U7726 (N_7726,N_7505,N_7597);
xor U7727 (N_7727,N_7532,N_7436);
nor U7728 (N_7728,N_7552,N_7481);
or U7729 (N_7729,N_7447,N_7488);
nor U7730 (N_7730,N_7403,N_7560);
nand U7731 (N_7731,N_7547,N_7588);
or U7732 (N_7732,N_7456,N_7419);
nor U7733 (N_7733,N_7579,N_7436);
nor U7734 (N_7734,N_7552,N_7572);
nand U7735 (N_7735,N_7433,N_7598);
nor U7736 (N_7736,N_7500,N_7591);
xnor U7737 (N_7737,N_7537,N_7450);
or U7738 (N_7738,N_7513,N_7449);
nand U7739 (N_7739,N_7422,N_7412);
and U7740 (N_7740,N_7564,N_7569);
nor U7741 (N_7741,N_7524,N_7587);
and U7742 (N_7742,N_7552,N_7430);
or U7743 (N_7743,N_7467,N_7447);
or U7744 (N_7744,N_7437,N_7460);
nor U7745 (N_7745,N_7497,N_7532);
nor U7746 (N_7746,N_7544,N_7557);
nor U7747 (N_7747,N_7483,N_7402);
and U7748 (N_7748,N_7508,N_7475);
nand U7749 (N_7749,N_7584,N_7468);
xnor U7750 (N_7750,N_7577,N_7544);
and U7751 (N_7751,N_7520,N_7477);
xnor U7752 (N_7752,N_7499,N_7503);
xnor U7753 (N_7753,N_7507,N_7411);
and U7754 (N_7754,N_7562,N_7414);
nand U7755 (N_7755,N_7467,N_7542);
nand U7756 (N_7756,N_7573,N_7577);
and U7757 (N_7757,N_7425,N_7423);
nor U7758 (N_7758,N_7430,N_7572);
nor U7759 (N_7759,N_7530,N_7428);
nor U7760 (N_7760,N_7483,N_7508);
xor U7761 (N_7761,N_7529,N_7413);
nand U7762 (N_7762,N_7429,N_7452);
or U7763 (N_7763,N_7437,N_7568);
and U7764 (N_7764,N_7423,N_7525);
nand U7765 (N_7765,N_7456,N_7451);
nor U7766 (N_7766,N_7521,N_7502);
or U7767 (N_7767,N_7591,N_7420);
and U7768 (N_7768,N_7481,N_7497);
nand U7769 (N_7769,N_7539,N_7428);
nand U7770 (N_7770,N_7595,N_7587);
nand U7771 (N_7771,N_7447,N_7590);
and U7772 (N_7772,N_7496,N_7481);
xor U7773 (N_7773,N_7486,N_7544);
nor U7774 (N_7774,N_7417,N_7532);
and U7775 (N_7775,N_7584,N_7587);
and U7776 (N_7776,N_7482,N_7494);
nand U7777 (N_7777,N_7550,N_7498);
nor U7778 (N_7778,N_7472,N_7526);
nand U7779 (N_7779,N_7440,N_7528);
nand U7780 (N_7780,N_7529,N_7423);
or U7781 (N_7781,N_7424,N_7562);
or U7782 (N_7782,N_7512,N_7511);
nor U7783 (N_7783,N_7417,N_7422);
or U7784 (N_7784,N_7549,N_7500);
or U7785 (N_7785,N_7409,N_7587);
nand U7786 (N_7786,N_7457,N_7461);
nor U7787 (N_7787,N_7482,N_7492);
or U7788 (N_7788,N_7532,N_7520);
or U7789 (N_7789,N_7574,N_7597);
xor U7790 (N_7790,N_7568,N_7406);
xor U7791 (N_7791,N_7476,N_7420);
nand U7792 (N_7792,N_7527,N_7513);
or U7793 (N_7793,N_7493,N_7567);
and U7794 (N_7794,N_7586,N_7566);
nor U7795 (N_7795,N_7409,N_7432);
and U7796 (N_7796,N_7406,N_7549);
nand U7797 (N_7797,N_7587,N_7582);
nor U7798 (N_7798,N_7458,N_7594);
and U7799 (N_7799,N_7452,N_7570);
or U7800 (N_7800,N_7665,N_7747);
and U7801 (N_7801,N_7709,N_7748);
nand U7802 (N_7802,N_7668,N_7751);
and U7803 (N_7803,N_7698,N_7754);
and U7804 (N_7804,N_7659,N_7601);
or U7805 (N_7805,N_7615,N_7777);
nor U7806 (N_7806,N_7781,N_7727);
or U7807 (N_7807,N_7732,N_7787);
or U7808 (N_7808,N_7684,N_7688);
xnor U7809 (N_7809,N_7768,N_7609);
nand U7810 (N_7810,N_7794,N_7696);
xnor U7811 (N_7811,N_7648,N_7756);
nor U7812 (N_7812,N_7753,N_7765);
nand U7813 (N_7813,N_7715,N_7743);
nand U7814 (N_7814,N_7625,N_7626);
nor U7815 (N_7815,N_7633,N_7735);
nor U7816 (N_7816,N_7785,N_7602);
nand U7817 (N_7817,N_7640,N_7676);
nand U7818 (N_7818,N_7632,N_7677);
xor U7819 (N_7819,N_7651,N_7667);
nor U7820 (N_7820,N_7690,N_7619);
nand U7821 (N_7821,N_7796,N_7728);
nand U7822 (N_7822,N_7742,N_7663);
and U7823 (N_7823,N_7786,N_7737);
nor U7824 (N_7824,N_7702,N_7711);
nand U7825 (N_7825,N_7661,N_7726);
or U7826 (N_7826,N_7712,N_7789);
nor U7827 (N_7827,N_7731,N_7631);
nand U7828 (N_7828,N_7622,N_7760);
xor U7829 (N_7829,N_7607,N_7681);
and U7830 (N_7830,N_7611,N_7618);
nand U7831 (N_7831,N_7750,N_7657);
xnor U7832 (N_7832,N_7795,N_7713);
or U7833 (N_7833,N_7654,N_7788);
nor U7834 (N_7834,N_7630,N_7687);
and U7835 (N_7835,N_7738,N_7606);
and U7836 (N_7836,N_7784,N_7790);
nand U7837 (N_7837,N_7730,N_7699);
nand U7838 (N_7838,N_7758,N_7704);
and U7839 (N_7839,N_7718,N_7741);
or U7840 (N_7840,N_7761,N_7764);
or U7841 (N_7841,N_7736,N_7733);
nor U7842 (N_7842,N_7766,N_7639);
and U7843 (N_7843,N_7664,N_7683);
and U7844 (N_7844,N_7769,N_7762);
or U7845 (N_7845,N_7649,N_7636);
and U7846 (N_7846,N_7637,N_7608);
nor U7847 (N_7847,N_7617,N_7703);
or U7848 (N_7848,N_7641,N_7674);
nand U7849 (N_7849,N_7746,N_7624);
or U7850 (N_7850,N_7798,N_7644);
nor U7851 (N_7851,N_7685,N_7791);
or U7852 (N_7852,N_7604,N_7623);
nand U7853 (N_7853,N_7686,N_7744);
nand U7854 (N_7854,N_7759,N_7675);
nor U7855 (N_7855,N_7603,N_7638);
and U7856 (N_7856,N_7714,N_7679);
nand U7857 (N_7857,N_7778,N_7749);
and U7858 (N_7858,N_7776,N_7745);
nor U7859 (N_7859,N_7629,N_7628);
and U7860 (N_7860,N_7650,N_7783);
nand U7861 (N_7861,N_7647,N_7720);
nor U7862 (N_7862,N_7763,N_7614);
and U7863 (N_7863,N_7610,N_7772);
and U7864 (N_7864,N_7627,N_7701);
and U7865 (N_7865,N_7656,N_7616);
nor U7866 (N_7866,N_7672,N_7620);
and U7867 (N_7867,N_7717,N_7613);
nand U7868 (N_7868,N_7666,N_7682);
nor U7869 (N_7869,N_7605,N_7646);
nor U7870 (N_7870,N_7634,N_7643);
nor U7871 (N_7871,N_7792,N_7678);
xor U7872 (N_7872,N_7775,N_7734);
nand U7873 (N_7873,N_7774,N_7721);
and U7874 (N_7874,N_7621,N_7692);
and U7875 (N_7875,N_7705,N_7653);
or U7876 (N_7876,N_7671,N_7680);
nor U7877 (N_7877,N_7767,N_7773);
nor U7878 (N_7878,N_7706,N_7693);
nor U7879 (N_7879,N_7652,N_7710);
xor U7880 (N_7880,N_7725,N_7642);
nand U7881 (N_7881,N_7799,N_7752);
or U7882 (N_7882,N_7779,N_7770);
nor U7883 (N_7883,N_7662,N_7755);
nor U7884 (N_7884,N_7612,N_7635);
nor U7885 (N_7885,N_7695,N_7700);
and U7886 (N_7886,N_7739,N_7797);
nor U7887 (N_7887,N_7670,N_7716);
or U7888 (N_7888,N_7655,N_7673);
xor U7889 (N_7889,N_7669,N_7708);
or U7890 (N_7890,N_7658,N_7757);
nor U7891 (N_7891,N_7782,N_7719);
or U7892 (N_7892,N_7729,N_7697);
or U7893 (N_7893,N_7689,N_7645);
and U7894 (N_7894,N_7600,N_7707);
nor U7895 (N_7895,N_7723,N_7771);
nand U7896 (N_7896,N_7793,N_7724);
nand U7897 (N_7897,N_7780,N_7691);
nand U7898 (N_7898,N_7722,N_7740);
nor U7899 (N_7899,N_7694,N_7660);
and U7900 (N_7900,N_7607,N_7750);
nand U7901 (N_7901,N_7603,N_7704);
nor U7902 (N_7902,N_7718,N_7761);
nand U7903 (N_7903,N_7693,N_7757);
nand U7904 (N_7904,N_7637,N_7696);
nand U7905 (N_7905,N_7620,N_7705);
nor U7906 (N_7906,N_7603,N_7622);
or U7907 (N_7907,N_7711,N_7668);
nor U7908 (N_7908,N_7770,N_7725);
or U7909 (N_7909,N_7607,N_7741);
xor U7910 (N_7910,N_7637,N_7740);
xnor U7911 (N_7911,N_7750,N_7707);
or U7912 (N_7912,N_7763,N_7699);
xor U7913 (N_7913,N_7628,N_7775);
nand U7914 (N_7914,N_7783,N_7763);
nor U7915 (N_7915,N_7738,N_7620);
nand U7916 (N_7916,N_7621,N_7769);
or U7917 (N_7917,N_7759,N_7784);
xnor U7918 (N_7918,N_7732,N_7681);
nand U7919 (N_7919,N_7604,N_7754);
nor U7920 (N_7920,N_7625,N_7776);
nor U7921 (N_7921,N_7672,N_7622);
nand U7922 (N_7922,N_7738,N_7657);
nand U7923 (N_7923,N_7622,N_7786);
or U7924 (N_7924,N_7791,N_7659);
nor U7925 (N_7925,N_7611,N_7685);
xnor U7926 (N_7926,N_7647,N_7607);
xor U7927 (N_7927,N_7622,N_7655);
nor U7928 (N_7928,N_7749,N_7795);
or U7929 (N_7929,N_7601,N_7708);
xnor U7930 (N_7930,N_7626,N_7609);
or U7931 (N_7931,N_7634,N_7797);
and U7932 (N_7932,N_7649,N_7696);
or U7933 (N_7933,N_7650,N_7683);
nor U7934 (N_7934,N_7747,N_7666);
nand U7935 (N_7935,N_7779,N_7745);
and U7936 (N_7936,N_7717,N_7601);
or U7937 (N_7937,N_7797,N_7766);
or U7938 (N_7938,N_7668,N_7659);
or U7939 (N_7939,N_7630,N_7654);
nand U7940 (N_7940,N_7685,N_7651);
and U7941 (N_7941,N_7794,N_7622);
nor U7942 (N_7942,N_7709,N_7774);
nand U7943 (N_7943,N_7763,N_7753);
nor U7944 (N_7944,N_7705,N_7792);
nor U7945 (N_7945,N_7649,N_7702);
or U7946 (N_7946,N_7672,N_7751);
or U7947 (N_7947,N_7721,N_7708);
and U7948 (N_7948,N_7638,N_7736);
and U7949 (N_7949,N_7615,N_7787);
xor U7950 (N_7950,N_7786,N_7642);
nand U7951 (N_7951,N_7793,N_7784);
nand U7952 (N_7952,N_7687,N_7648);
and U7953 (N_7953,N_7696,N_7745);
and U7954 (N_7954,N_7609,N_7617);
xnor U7955 (N_7955,N_7656,N_7768);
or U7956 (N_7956,N_7764,N_7720);
nand U7957 (N_7957,N_7730,N_7661);
xnor U7958 (N_7958,N_7683,N_7737);
or U7959 (N_7959,N_7771,N_7718);
nor U7960 (N_7960,N_7655,N_7737);
nor U7961 (N_7961,N_7697,N_7763);
or U7962 (N_7962,N_7693,N_7644);
and U7963 (N_7963,N_7796,N_7660);
and U7964 (N_7964,N_7638,N_7611);
nor U7965 (N_7965,N_7646,N_7684);
or U7966 (N_7966,N_7694,N_7725);
nor U7967 (N_7967,N_7615,N_7679);
nand U7968 (N_7968,N_7604,N_7756);
nand U7969 (N_7969,N_7748,N_7786);
or U7970 (N_7970,N_7632,N_7772);
nand U7971 (N_7971,N_7659,N_7769);
or U7972 (N_7972,N_7668,N_7625);
nor U7973 (N_7973,N_7604,N_7651);
or U7974 (N_7974,N_7676,N_7716);
nand U7975 (N_7975,N_7694,N_7610);
nand U7976 (N_7976,N_7721,N_7775);
nor U7977 (N_7977,N_7763,N_7662);
and U7978 (N_7978,N_7643,N_7776);
nor U7979 (N_7979,N_7688,N_7796);
or U7980 (N_7980,N_7629,N_7745);
nor U7981 (N_7981,N_7713,N_7779);
nand U7982 (N_7982,N_7763,N_7622);
nand U7983 (N_7983,N_7650,N_7687);
and U7984 (N_7984,N_7742,N_7701);
and U7985 (N_7985,N_7756,N_7793);
and U7986 (N_7986,N_7687,N_7776);
and U7987 (N_7987,N_7687,N_7731);
and U7988 (N_7988,N_7762,N_7618);
nand U7989 (N_7989,N_7685,N_7786);
and U7990 (N_7990,N_7722,N_7664);
nor U7991 (N_7991,N_7700,N_7653);
and U7992 (N_7992,N_7636,N_7612);
nand U7993 (N_7993,N_7706,N_7696);
or U7994 (N_7994,N_7666,N_7768);
and U7995 (N_7995,N_7611,N_7783);
nand U7996 (N_7996,N_7746,N_7780);
and U7997 (N_7997,N_7730,N_7608);
nand U7998 (N_7998,N_7752,N_7798);
nand U7999 (N_7999,N_7612,N_7634);
and U8000 (N_8000,N_7925,N_7902);
or U8001 (N_8001,N_7882,N_7830);
and U8002 (N_8002,N_7912,N_7889);
and U8003 (N_8003,N_7805,N_7847);
and U8004 (N_8004,N_7972,N_7890);
nand U8005 (N_8005,N_7992,N_7899);
or U8006 (N_8006,N_7822,N_7933);
nand U8007 (N_8007,N_7873,N_7875);
nor U8008 (N_8008,N_7924,N_7807);
and U8009 (N_8009,N_7802,N_7950);
nand U8010 (N_8010,N_7834,N_7947);
and U8011 (N_8011,N_7987,N_7817);
nand U8012 (N_8012,N_7978,N_7975);
nand U8013 (N_8013,N_7918,N_7981);
nand U8014 (N_8014,N_7880,N_7877);
and U8015 (N_8015,N_7839,N_7881);
nor U8016 (N_8016,N_7943,N_7980);
nor U8017 (N_8017,N_7852,N_7908);
or U8018 (N_8018,N_7824,N_7879);
nor U8019 (N_8019,N_7958,N_7961);
and U8020 (N_8020,N_7888,N_7838);
and U8021 (N_8021,N_7966,N_7968);
nand U8022 (N_8022,N_7809,N_7867);
and U8023 (N_8023,N_7938,N_7960);
nand U8024 (N_8024,N_7808,N_7853);
nand U8025 (N_8025,N_7923,N_7855);
nand U8026 (N_8026,N_7917,N_7970);
and U8027 (N_8027,N_7862,N_7914);
nand U8028 (N_8028,N_7840,N_7894);
or U8029 (N_8029,N_7955,N_7998);
or U8030 (N_8030,N_7928,N_7836);
nor U8031 (N_8031,N_7982,N_7874);
nor U8032 (N_8032,N_7878,N_7926);
and U8033 (N_8033,N_7940,N_7921);
nor U8034 (N_8034,N_7833,N_7850);
or U8035 (N_8035,N_7945,N_7871);
and U8036 (N_8036,N_7997,N_7962);
and U8037 (N_8037,N_7870,N_7896);
or U8038 (N_8038,N_7930,N_7971);
and U8039 (N_8039,N_7932,N_7976);
nand U8040 (N_8040,N_7964,N_7984);
xor U8041 (N_8041,N_7967,N_7897);
and U8042 (N_8042,N_7952,N_7919);
nor U8043 (N_8043,N_7910,N_7835);
and U8044 (N_8044,N_7861,N_7973);
and U8045 (N_8045,N_7946,N_7898);
nor U8046 (N_8046,N_7996,N_7883);
nor U8047 (N_8047,N_7885,N_7869);
xor U8048 (N_8048,N_7956,N_7988);
xnor U8049 (N_8049,N_7904,N_7866);
nor U8050 (N_8050,N_7893,N_7991);
and U8051 (N_8051,N_7963,N_7815);
nor U8052 (N_8052,N_7806,N_7920);
nand U8053 (N_8053,N_7985,N_7849);
or U8054 (N_8054,N_7977,N_7915);
nor U8055 (N_8055,N_7829,N_7845);
or U8056 (N_8056,N_7842,N_7927);
and U8057 (N_8057,N_7954,N_7911);
and U8058 (N_8058,N_7837,N_7937);
nor U8059 (N_8059,N_7993,N_7944);
and U8060 (N_8060,N_7990,N_7851);
or U8061 (N_8061,N_7819,N_7941);
nand U8062 (N_8062,N_7999,N_7931);
nand U8063 (N_8063,N_7872,N_7865);
nor U8064 (N_8064,N_7826,N_7939);
or U8065 (N_8065,N_7922,N_7953);
and U8066 (N_8066,N_7936,N_7856);
nor U8067 (N_8067,N_7827,N_7816);
or U8068 (N_8068,N_7823,N_7951);
and U8069 (N_8069,N_7994,N_7965);
or U8070 (N_8070,N_7863,N_7846);
or U8071 (N_8071,N_7906,N_7986);
nand U8072 (N_8072,N_7957,N_7989);
and U8073 (N_8073,N_7909,N_7995);
nand U8074 (N_8074,N_7887,N_7859);
nor U8075 (N_8075,N_7907,N_7929);
and U8076 (N_8076,N_7828,N_7983);
and U8077 (N_8077,N_7803,N_7804);
nor U8078 (N_8078,N_7886,N_7858);
xnor U8079 (N_8079,N_7820,N_7974);
or U8080 (N_8080,N_7864,N_7900);
xnor U8081 (N_8081,N_7969,N_7844);
or U8082 (N_8082,N_7935,N_7843);
or U8083 (N_8083,N_7854,N_7831);
xor U8084 (N_8084,N_7818,N_7812);
or U8085 (N_8085,N_7916,N_7895);
or U8086 (N_8086,N_7942,N_7810);
nor U8087 (N_8087,N_7868,N_7979);
or U8088 (N_8088,N_7913,N_7959);
nor U8089 (N_8089,N_7876,N_7800);
nor U8090 (N_8090,N_7949,N_7841);
and U8091 (N_8091,N_7811,N_7825);
and U8092 (N_8092,N_7901,N_7948);
nor U8093 (N_8093,N_7884,N_7814);
xor U8094 (N_8094,N_7905,N_7857);
xnor U8095 (N_8095,N_7821,N_7813);
nor U8096 (N_8096,N_7934,N_7860);
and U8097 (N_8097,N_7832,N_7801);
and U8098 (N_8098,N_7903,N_7892);
nor U8099 (N_8099,N_7891,N_7848);
nor U8100 (N_8100,N_7996,N_7991);
or U8101 (N_8101,N_7876,N_7980);
and U8102 (N_8102,N_7977,N_7995);
nand U8103 (N_8103,N_7986,N_7810);
nand U8104 (N_8104,N_7892,N_7896);
or U8105 (N_8105,N_7857,N_7957);
nand U8106 (N_8106,N_7833,N_7836);
and U8107 (N_8107,N_7869,N_7838);
nand U8108 (N_8108,N_7822,N_7864);
or U8109 (N_8109,N_7901,N_7903);
nand U8110 (N_8110,N_7829,N_7866);
and U8111 (N_8111,N_7898,N_7987);
nor U8112 (N_8112,N_7931,N_7982);
nor U8113 (N_8113,N_7803,N_7976);
and U8114 (N_8114,N_7891,N_7999);
or U8115 (N_8115,N_7956,N_7835);
nor U8116 (N_8116,N_7837,N_7865);
nor U8117 (N_8117,N_7947,N_7827);
nor U8118 (N_8118,N_7944,N_7873);
nor U8119 (N_8119,N_7947,N_7875);
nand U8120 (N_8120,N_7826,N_7964);
nand U8121 (N_8121,N_7946,N_7834);
and U8122 (N_8122,N_7834,N_7968);
xor U8123 (N_8123,N_7996,N_7871);
or U8124 (N_8124,N_7878,N_7877);
and U8125 (N_8125,N_7816,N_7829);
nor U8126 (N_8126,N_7813,N_7872);
and U8127 (N_8127,N_7994,N_7926);
xnor U8128 (N_8128,N_7969,N_7843);
nand U8129 (N_8129,N_7928,N_7930);
nor U8130 (N_8130,N_7926,N_7808);
nand U8131 (N_8131,N_7876,N_7909);
or U8132 (N_8132,N_7904,N_7820);
nor U8133 (N_8133,N_7869,N_7981);
nor U8134 (N_8134,N_7959,N_7967);
nand U8135 (N_8135,N_7945,N_7853);
nor U8136 (N_8136,N_7845,N_7927);
or U8137 (N_8137,N_7821,N_7851);
or U8138 (N_8138,N_7974,N_7863);
nor U8139 (N_8139,N_7922,N_7987);
and U8140 (N_8140,N_7886,N_7902);
and U8141 (N_8141,N_7883,N_7953);
and U8142 (N_8142,N_7816,N_7881);
nand U8143 (N_8143,N_7808,N_7892);
nand U8144 (N_8144,N_7960,N_7925);
and U8145 (N_8145,N_7905,N_7803);
or U8146 (N_8146,N_7877,N_7862);
or U8147 (N_8147,N_7831,N_7982);
or U8148 (N_8148,N_7986,N_7958);
or U8149 (N_8149,N_7973,N_7847);
or U8150 (N_8150,N_7805,N_7885);
and U8151 (N_8151,N_7811,N_7901);
and U8152 (N_8152,N_7807,N_7915);
xnor U8153 (N_8153,N_7920,N_7984);
nand U8154 (N_8154,N_7961,N_7808);
or U8155 (N_8155,N_7926,N_7979);
or U8156 (N_8156,N_7989,N_7804);
nor U8157 (N_8157,N_7896,N_7940);
or U8158 (N_8158,N_7984,N_7930);
and U8159 (N_8159,N_7809,N_7851);
or U8160 (N_8160,N_7954,N_7958);
nor U8161 (N_8161,N_7839,N_7806);
nand U8162 (N_8162,N_7899,N_7988);
or U8163 (N_8163,N_7814,N_7858);
xnor U8164 (N_8164,N_7902,N_7933);
or U8165 (N_8165,N_7889,N_7983);
or U8166 (N_8166,N_7969,N_7897);
nor U8167 (N_8167,N_7944,N_7991);
or U8168 (N_8168,N_7804,N_7940);
xnor U8169 (N_8169,N_7827,N_7933);
nand U8170 (N_8170,N_7893,N_7826);
xnor U8171 (N_8171,N_7835,N_7947);
nand U8172 (N_8172,N_7938,N_7899);
and U8173 (N_8173,N_7872,N_7974);
or U8174 (N_8174,N_7910,N_7844);
nor U8175 (N_8175,N_7807,N_7935);
xnor U8176 (N_8176,N_7984,N_7857);
and U8177 (N_8177,N_7877,N_7820);
nor U8178 (N_8178,N_7862,N_7825);
nand U8179 (N_8179,N_7815,N_7920);
and U8180 (N_8180,N_7829,N_7909);
nor U8181 (N_8181,N_7862,N_7873);
and U8182 (N_8182,N_7924,N_7838);
or U8183 (N_8183,N_7963,N_7899);
nor U8184 (N_8184,N_7960,N_7844);
or U8185 (N_8185,N_7885,N_7979);
nor U8186 (N_8186,N_7906,N_7814);
nor U8187 (N_8187,N_7885,N_7895);
and U8188 (N_8188,N_7881,N_7921);
nand U8189 (N_8189,N_7897,N_7894);
nor U8190 (N_8190,N_7900,N_7838);
nor U8191 (N_8191,N_7878,N_7979);
and U8192 (N_8192,N_7951,N_7892);
and U8193 (N_8193,N_7855,N_7868);
nand U8194 (N_8194,N_7960,N_7803);
nor U8195 (N_8195,N_7999,N_7975);
xnor U8196 (N_8196,N_7975,N_7887);
and U8197 (N_8197,N_7996,N_7811);
or U8198 (N_8198,N_7952,N_7901);
or U8199 (N_8199,N_7867,N_7880);
and U8200 (N_8200,N_8021,N_8022);
or U8201 (N_8201,N_8005,N_8141);
and U8202 (N_8202,N_8092,N_8152);
nand U8203 (N_8203,N_8115,N_8184);
or U8204 (N_8204,N_8043,N_8017);
nand U8205 (N_8205,N_8137,N_8151);
nor U8206 (N_8206,N_8166,N_8102);
xor U8207 (N_8207,N_8170,N_8051);
and U8208 (N_8208,N_8155,N_8087);
xor U8209 (N_8209,N_8003,N_8072);
nand U8210 (N_8210,N_8150,N_8073);
nand U8211 (N_8211,N_8113,N_8065);
xnor U8212 (N_8212,N_8035,N_8082);
xnor U8213 (N_8213,N_8000,N_8078);
and U8214 (N_8214,N_8168,N_8160);
xnor U8215 (N_8215,N_8156,N_8176);
nor U8216 (N_8216,N_8131,N_8054);
and U8217 (N_8217,N_8091,N_8061);
nor U8218 (N_8218,N_8041,N_8026);
or U8219 (N_8219,N_8085,N_8178);
nor U8220 (N_8220,N_8192,N_8145);
nand U8221 (N_8221,N_8097,N_8023);
nand U8222 (N_8222,N_8029,N_8121);
xor U8223 (N_8223,N_8187,N_8019);
nand U8224 (N_8224,N_8118,N_8039);
nor U8225 (N_8225,N_8134,N_8001);
nor U8226 (N_8226,N_8090,N_8095);
nand U8227 (N_8227,N_8159,N_8196);
nand U8228 (N_8228,N_8175,N_8044);
and U8229 (N_8229,N_8074,N_8112);
and U8230 (N_8230,N_8071,N_8030);
xor U8231 (N_8231,N_8181,N_8167);
or U8232 (N_8232,N_8109,N_8114);
and U8233 (N_8233,N_8047,N_8182);
and U8234 (N_8234,N_8098,N_8125);
nand U8235 (N_8235,N_8117,N_8110);
nand U8236 (N_8236,N_8049,N_8094);
nand U8237 (N_8237,N_8127,N_8066);
and U8238 (N_8238,N_8008,N_8009);
and U8239 (N_8239,N_8052,N_8136);
nand U8240 (N_8240,N_8174,N_8036);
and U8241 (N_8241,N_8055,N_8033);
nor U8242 (N_8242,N_8165,N_8086);
nand U8243 (N_8243,N_8111,N_8011);
and U8244 (N_8244,N_8037,N_8056);
nand U8245 (N_8245,N_8116,N_8190);
or U8246 (N_8246,N_8018,N_8154);
and U8247 (N_8247,N_8139,N_8169);
nor U8248 (N_8248,N_8157,N_8040);
or U8249 (N_8249,N_8031,N_8162);
or U8250 (N_8250,N_8140,N_8084);
nor U8251 (N_8251,N_8158,N_8130);
nand U8252 (N_8252,N_8058,N_8057);
nand U8253 (N_8253,N_8068,N_8002);
nand U8254 (N_8254,N_8173,N_8053);
or U8255 (N_8255,N_8194,N_8006);
nor U8256 (N_8256,N_8010,N_8186);
nand U8257 (N_8257,N_8171,N_8120);
nand U8258 (N_8258,N_8089,N_8042);
or U8259 (N_8259,N_8107,N_8147);
or U8260 (N_8260,N_8063,N_8079);
or U8261 (N_8261,N_8088,N_8148);
xor U8262 (N_8262,N_8067,N_8126);
xnor U8263 (N_8263,N_8142,N_8199);
nor U8264 (N_8264,N_8062,N_8195);
or U8265 (N_8265,N_8138,N_8004);
nor U8266 (N_8266,N_8185,N_8027);
nor U8267 (N_8267,N_8104,N_8164);
and U8268 (N_8268,N_8024,N_8163);
or U8269 (N_8269,N_8193,N_8077);
nor U8270 (N_8270,N_8135,N_8128);
nand U8271 (N_8271,N_8096,N_8197);
nor U8272 (N_8272,N_8119,N_8014);
or U8273 (N_8273,N_8038,N_8070);
nand U8274 (N_8274,N_8132,N_8076);
xor U8275 (N_8275,N_8179,N_8198);
and U8276 (N_8276,N_8191,N_8028);
and U8277 (N_8277,N_8123,N_8101);
nand U8278 (N_8278,N_8149,N_8081);
or U8279 (N_8279,N_8032,N_8100);
nand U8280 (N_8280,N_8188,N_8144);
nand U8281 (N_8281,N_8013,N_8106);
xor U8282 (N_8282,N_8016,N_8069);
xnor U8283 (N_8283,N_8059,N_8133);
nand U8284 (N_8284,N_8105,N_8161);
or U8285 (N_8285,N_8189,N_8080);
or U8286 (N_8286,N_8046,N_8064);
and U8287 (N_8287,N_8007,N_8099);
xor U8288 (N_8288,N_8129,N_8075);
or U8289 (N_8289,N_8012,N_8172);
xor U8290 (N_8290,N_8034,N_8108);
or U8291 (N_8291,N_8180,N_8093);
nor U8292 (N_8292,N_8124,N_8103);
nand U8293 (N_8293,N_8050,N_8177);
nor U8294 (N_8294,N_8122,N_8153);
nand U8295 (N_8295,N_8183,N_8060);
nand U8296 (N_8296,N_8045,N_8146);
and U8297 (N_8297,N_8020,N_8015);
nand U8298 (N_8298,N_8083,N_8025);
nor U8299 (N_8299,N_8048,N_8143);
nand U8300 (N_8300,N_8057,N_8159);
and U8301 (N_8301,N_8161,N_8032);
nand U8302 (N_8302,N_8120,N_8152);
or U8303 (N_8303,N_8081,N_8137);
or U8304 (N_8304,N_8041,N_8121);
nor U8305 (N_8305,N_8003,N_8012);
nand U8306 (N_8306,N_8025,N_8116);
or U8307 (N_8307,N_8113,N_8022);
nor U8308 (N_8308,N_8071,N_8145);
or U8309 (N_8309,N_8190,N_8103);
nand U8310 (N_8310,N_8183,N_8021);
or U8311 (N_8311,N_8011,N_8151);
nand U8312 (N_8312,N_8049,N_8051);
xnor U8313 (N_8313,N_8054,N_8116);
nor U8314 (N_8314,N_8163,N_8011);
nand U8315 (N_8315,N_8056,N_8177);
and U8316 (N_8316,N_8175,N_8084);
or U8317 (N_8317,N_8141,N_8021);
and U8318 (N_8318,N_8057,N_8168);
or U8319 (N_8319,N_8030,N_8007);
or U8320 (N_8320,N_8159,N_8114);
nor U8321 (N_8321,N_8103,N_8130);
and U8322 (N_8322,N_8037,N_8189);
or U8323 (N_8323,N_8163,N_8111);
or U8324 (N_8324,N_8189,N_8023);
or U8325 (N_8325,N_8165,N_8125);
and U8326 (N_8326,N_8128,N_8140);
xnor U8327 (N_8327,N_8170,N_8141);
nor U8328 (N_8328,N_8151,N_8111);
and U8329 (N_8329,N_8152,N_8124);
and U8330 (N_8330,N_8135,N_8044);
or U8331 (N_8331,N_8102,N_8177);
nor U8332 (N_8332,N_8131,N_8060);
xor U8333 (N_8333,N_8068,N_8001);
nand U8334 (N_8334,N_8123,N_8167);
nor U8335 (N_8335,N_8142,N_8021);
nand U8336 (N_8336,N_8055,N_8030);
and U8337 (N_8337,N_8113,N_8096);
and U8338 (N_8338,N_8181,N_8002);
and U8339 (N_8339,N_8115,N_8089);
and U8340 (N_8340,N_8186,N_8130);
nor U8341 (N_8341,N_8141,N_8115);
or U8342 (N_8342,N_8009,N_8192);
and U8343 (N_8343,N_8101,N_8018);
or U8344 (N_8344,N_8119,N_8091);
and U8345 (N_8345,N_8085,N_8191);
nor U8346 (N_8346,N_8155,N_8167);
and U8347 (N_8347,N_8138,N_8043);
xnor U8348 (N_8348,N_8023,N_8154);
or U8349 (N_8349,N_8181,N_8127);
nand U8350 (N_8350,N_8176,N_8002);
and U8351 (N_8351,N_8149,N_8132);
nand U8352 (N_8352,N_8122,N_8072);
nand U8353 (N_8353,N_8061,N_8056);
or U8354 (N_8354,N_8047,N_8004);
nand U8355 (N_8355,N_8139,N_8111);
nand U8356 (N_8356,N_8185,N_8161);
and U8357 (N_8357,N_8198,N_8025);
and U8358 (N_8358,N_8038,N_8086);
nand U8359 (N_8359,N_8181,N_8149);
or U8360 (N_8360,N_8112,N_8095);
or U8361 (N_8361,N_8190,N_8039);
and U8362 (N_8362,N_8199,N_8081);
nor U8363 (N_8363,N_8008,N_8189);
or U8364 (N_8364,N_8050,N_8027);
nor U8365 (N_8365,N_8116,N_8098);
or U8366 (N_8366,N_8103,N_8072);
or U8367 (N_8367,N_8108,N_8075);
nand U8368 (N_8368,N_8195,N_8043);
nand U8369 (N_8369,N_8059,N_8021);
nor U8370 (N_8370,N_8195,N_8152);
nand U8371 (N_8371,N_8189,N_8087);
or U8372 (N_8372,N_8026,N_8001);
or U8373 (N_8373,N_8029,N_8055);
nand U8374 (N_8374,N_8087,N_8003);
or U8375 (N_8375,N_8023,N_8176);
and U8376 (N_8376,N_8011,N_8175);
or U8377 (N_8377,N_8108,N_8145);
or U8378 (N_8378,N_8156,N_8072);
nor U8379 (N_8379,N_8012,N_8167);
and U8380 (N_8380,N_8123,N_8113);
nor U8381 (N_8381,N_8035,N_8079);
and U8382 (N_8382,N_8015,N_8171);
nor U8383 (N_8383,N_8030,N_8082);
nand U8384 (N_8384,N_8014,N_8162);
and U8385 (N_8385,N_8008,N_8196);
and U8386 (N_8386,N_8101,N_8075);
or U8387 (N_8387,N_8083,N_8096);
or U8388 (N_8388,N_8146,N_8054);
and U8389 (N_8389,N_8119,N_8045);
nand U8390 (N_8390,N_8060,N_8130);
or U8391 (N_8391,N_8089,N_8059);
nand U8392 (N_8392,N_8007,N_8145);
and U8393 (N_8393,N_8064,N_8122);
nand U8394 (N_8394,N_8193,N_8150);
or U8395 (N_8395,N_8101,N_8194);
or U8396 (N_8396,N_8066,N_8195);
and U8397 (N_8397,N_8010,N_8077);
nor U8398 (N_8398,N_8068,N_8171);
and U8399 (N_8399,N_8113,N_8180);
xnor U8400 (N_8400,N_8262,N_8223);
or U8401 (N_8401,N_8302,N_8216);
nor U8402 (N_8402,N_8363,N_8272);
and U8403 (N_8403,N_8229,N_8230);
or U8404 (N_8404,N_8389,N_8362);
or U8405 (N_8405,N_8207,N_8331);
xor U8406 (N_8406,N_8398,N_8211);
and U8407 (N_8407,N_8317,N_8399);
nand U8408 (N_8408,N_8328,N_8383);
nand U8409 (N_8409,N_8313,N_8382);
xnor U8410 (N_8410,N_8357,N_8254);
and U8411 (N_8411,N_8256,N_8310);
nand U8412 (N_8412,N_8245,N_8220);
or U8413 (N_8413,N_8227,N_8283);
xor U8414 (N_8414,N_8319,N_8228);
and U8415 (N_8415,N_8321,N_8213);
or U8416 (N_8416,N_8322,N_8369);
and U8417 (N_8417,N_8205,N_8329);
nand U8418 (N_8418,N_8351,N_8294);
nand U8419 (N_8419,N_8247,N_8252);
nor U8420 (N_8420,N_8333,N_8242);
or U8421 (N_8421,N_8366,N_8299);
nand U8422 (N_8422,N_8244,N_8232);
or U8423 (N_8423,N_8275,N_8343);
nand U8424 (N_8424,N_8268,N_8209);
xnor U8425 (N_8425,N_8392,N_8217);
nand U8426 (N_8426,N_8296,N_8312);
xnor U8427 (N_8427,N_8231,N_8249);
xnor U8428 (N_8428,N_8314,N_8277);
or U8429 (N_8429,N_8270,N_8251);
and U8430 (N_8430,N_8340,N_8222);
xnor U8431 (N_8431,N_8326,N_8352);
and U8432 (N_8432,N_8241,N_8334);
nor U8433 (N_8433,N_8237,N_8315);
nor U8434 (N_8434,N_8248,N_8287);
nor U8435 (N_8435,N_8236,N_8370);
nor U8436 (N_8436,N_8218,N_8293);
and U8437 (N_8437,N_8298,N_8238);
or U8438 (N_8438,N_8320,N_8279);
nand U8439 (N_8439,N_8282,N_8311);
or U8440 (N_8440,N_8365,N_8267);
and U8441 (N_8441,N_8304,N_8381);
nor U8442 (N_8442,N_8271,N_8323);
and U8443 (N_8443,N_8342,N_8206);
nor U8444 (N_8444,N_8316,N_8212);
or U8445 (N_8445,N_8221,N_8373);
and U8446 (N_8446,N_8204,N_8301);
nand U8447 (N_8447,N_8393,N_8219);
nand U8448 (N_8448,N_8263,N_8318);
or U8449 (N_8449,N_8388,N_8233);
nand U8450 (N_8450,N_8258,N_8337);
nor U8451 (N_8451,N_8397,N_8264);
nand U8452 (N_8452,N_8280,N_8353);
nor U8453 (N_8453,N_8305,N_8261);
and U8454 (N_8454,N_8346,N_8274);
nor U8455 (N_8455,N_8390,N_8200);
nor U8456 (N_8456,N_8203,N_8341);
nand U8457 (N_8457,N_8276,N_8377);
nor U8458 (N_8458,N_8288,N_8234);
xor U8459 (N_8459,N_8385,N_8307);
and U8460 (N_8460,N_8210,N_8384);
or U8461 (N_8461,N_8350,N_8345);
and U8462 (N_8462,N_8344,N_8356);
and U8463 (N_8463,N_8269,N_8335);
nand U8464 (N_8464,N_8284,N_8224);
nand U8465 (N_8465,N_8368,N_8285);
nand U8466 (N_8466,N_8201,N_8265);
nand U8467 (N_8467,N_8376,N_8250);
and U8468 (N_8468,N_8303,N_8348);
nor U8469 (N_8469,N_8281,N_8300);
nand U8470 (N_8470,N_8215,N_8354);
xnor U8471 (N_8471,N_8255,N_8309);
nand U8472 (N_8472,N_8360,N_8208);
or U8473 (N_8473,N_8332,N_8286);
or U8474 (N_8474,N_8225,N_8214);
or U8475 (N_8475,N_8297,N_8386);
or U8476 (N_8476,N_8327,N_8355);
xor U8477 (N_8477,N_8273,N_8290);
nand U8478 (N_8478,N_8339,N_8260);
nor U8479 (N_8479,N_8240,N_8349);
and U8480 (N_8480,N_8259,N_8375);
or U8481 (N_8481,N_8239,N_8396);
nand U8482 (N_8482,N_8235,N_8324);
and U8483 (N_8483,N_8336,N_8278);
and U8484 (N_8484,N_8202,N_8330);
xnor U8485 (N_8485,N_8306,N_8367);
nand U8486 (N_8486,N_8380,N_8243);
nand U8487 (N_8487,N_8371,N_8289);
or U8488 (N_8488,N_8394,N_8253);
and U8489 (N_8489,N_8266,N_8374);
nor U8490 (N_8490,N_8295,N_8308);
or U8491 (N_8491,N_8372,N_8391);
and U8492 (N_8492,N_8226,N_8379);
nor U8493 (N_8493,N_8338,N_8395);
nor U8494 (N_8494,N_8364,N_8246);
nand U8495 (N_8495,N_8292,N_8291);
nand U8496 (N_8496,N_8378,N_8361);
or U8497 (N_8497,N_8387,N_8325);
xnor U8498 (N_8498,N_8359,N_8347);
nand U8499 (N_8499,N_8257,N_8358);
xnor U8500 (N_8500,N_8246,N_8284);
or U8501 (N_8501,N_8324,N_8236);
nand U8502 (N_8502,N_8324,N_8206);
nand U8503 (N_8503,N_8262,N_8338);
or U8504 (N_8504,N_8267,N_8281);
nand U8505 (N_8505,N_8246,N_8395);
nor U8506 (N_8506,N_8380,N_8353);
nand U8507 (N_8507,N_8351,N_8245);
xnor U8508 (N_8508,N_8333,N_8255);
or U8509 (N_8509,N_8347,N_8396);
nand U8510 (N_8510,N_8397,N_8331);
nand U8511 (N_8511,N_8276,N_8233);
nand U8512 (N_8512,N_8356,N_8274);
or U8513 (N_8513,N_8375,N_8254);
nor U8514 (N_8514,N_8305,N_8310);
and U8515 (N_8515,N_8372,N_8256);
or U8516 (N_8516,N_8208,N_8273);
nor U8517 (N_8517,N_8347,N_8233);
nor U8518 (N_8518,N_8300,N_8299);
nor U8519 (N_8519,N_8332,N_8380);
or U8520 (N_8520,N_8228,N_8375);
or U8521 (N_8521,N_8204,N_8281);
nor U8522 (N_8522,N_8372,N_8359);
nor U8523 (N_8523,N_8382,N_8391);
nand U8524 (N_8524,N_8275,N_8352);
and U8525 (N_8525,N_8363,N_8237);
nand U8526 (N_8526,N_8297,N_8304);
and U8527 (N_8527,N_8329,N_8272);
and U8528 (N_8528,N_8310,N_8235);
or U8529 (N_8529,N_8362,N_8315);
nor U8530 (N_8530,N_8240,N_8205);
nand U8531 (N_8531,N_8233,N_8311);
nor U8532 (N_8532,N_8269,N_8294);
nand U8533 (N_8533,N_8264,N_8284);
xnor U8534 (N_8534,N_8316,N_8255);
nor U8535 (N_8535,N_8287,N_8280);
and U8536 (N_8536,N_8237,N_8223);
nand U8537 (N_8537,N_8318,N_8289);
and U8538 (N_8538,N_8258,N_8274);
or U8539 (N_8539,N_8289,N_8363);
or U8540 (N_8540,N_8249,N_8205);
or U8541 (N_8541,N_8361,N_8258);
nand U8542 (N_8542,N_8224,N_8237);
or U8543 (N_8543,N_8376,N_8324);
and U8544 (N_8544,N_8394,N_8263);
or U8545 (N_8545,N_8212,N_8339);
or U8546 (N_8546,N_8361,N_8244);
nor U8547 (N_8547,N_8202,N_8245);
nor U8548 (N_8548,N_8345,N_8305);
or U8549 (N_8549,N_8340,N_8266);
nor U8550 (N_8550,N_8213,N_8330);
and U8551 (N_8551,N_8303,N_8207);
or U8552 (N_8552,N_8312,N_8234);
nor U8553 (N_8553,N_8234,N_8229);
or U8554 (N_8554,N_8389,N_8242);
nor U8555 (N_8555,N_8246,N_8294);
xor U8556 (N_8556,N_8335,N_8215);
or U8557 (N_8557,N_8283,N_8356);
or U8558 (N_8558,N_8391,N_8240);
xor U8559 (N_8559,N_8218,N_8219);
nor U8560 (N_8560,N_8385,N_8252);
and U8561 (N_8561,N_8223,N_8342);
nand U8562 (N_8562,N_8231,N_8347);
nor U8563 (N_8563,N_8228,N_8391);
nor U8564 (N_8564,N_8340,N_8318);
and U8565 (N_8565,N_8389,N_8249);
or U8566 (N_8566,N_8308,N_8294);
xnor U8567 (N_8567,N_8388,N_8229);
xor U8568 (N_8568,N_8369,N_8325);
xor U8569 (N_8569,N_8271,N_8389);
nand U8570 (N_8570,N_8299,N_8340);
and U8571 (N_8571,N_8342,N_8318);
and U8572 (N_8572,N_8348,N_8344);
or U8573 (N_8573,N_8298,N_8257);
nor U8574 (N_8574,N_8248,N_8278);
nand U8575 (N_8575,N_8252,N_8240);
nand U8576 (N_8576,N_8210,N_8368);
nand U8577 (N_8577,N_8342,N_8300);
or U8578 (N_8578,N_8283,N_8218);
or U8579 (N_8579,N_8318,N_8381);
nor U8580 (N_8580,N_8251,N_8378);
xnor U8581 (N_8581,N_8351,N_8250);
and U8582 (N_8582,N_8245,N_8285);
or U8583 (N_8583,N_8202,N_8397);
or U8584 (N_8584,N_8306,N_8260);
and U8585 (N_8585,N_8343,N_8269);
or U8586 (N_8586,N_8392,N_8276);
xor U8587 (N_8587,N_8384,N_8212);
nand U8588 (N_8588,N_8251,N_8328);
and U8589 (N_8589,N_8347,N_8217);
nand U8590 (N_8590,N_8268,N_8355);
xor U8591 (N_8591,N_8273,N_8243);
nor U8592 (N_8592,N_8378,N_8366);
and U8593 (N_8593,N_8271,N_8381);
nand U8594 (N_8594,N_8222,N_8253);
nor U8595 (N_8595,N_8341,N_8274);
nor U8596 (N_8596,N_8229,N_8393);
nor U8597 (N_8597,N_8342,N_8367);
and U8598 (N_8598,N_8393,N_8225);
nor U8599 (N_8599,N_8267,N_8321);
nor U8600 (N_8600,N_8436,N_8411);
nor U8601 (N_8601,N_8459,N_8435);
or U8602 (N_8602,N_8506,N_8432);
nor U8603 (N_8603,N_8545,N_8467);
and U8604 (N_8604,N_8541,N_8422);
nor U8605 (N_8605,N_8447,N_8589);
and U8606 (N_8606,N_8542,N_8554);
nor U8607 (N_8607,N_8492,N_8441);
and U8608 (N_8608,N_8553,N_8413);
nand U8609 (N_8609,N_8527,N_8585);
xnor U8610 (N_8610,N_8513,N_8455);
and U8611 (N_8611,N_8480,N_8466);
nor U8612 (N_8612,N_8535,N_8590);
and U8613 (N_8613,N_8409,N_8454);
xor U8614 (N_8614,N_8517,N_8504);
nand U8615 (N_8615,N_8579,N_8534);
and U8616 (N_8616,N_8568,N_8404);
and U8617 (N_8617,N_8563,N_8428);
nor U8618 (N_8618,N_8514,N_8482);
nand U8619 (N_8619,N_8452,N_8471);
nand U8620 (N_8620,N_8421,N_8418);
or U8621 (N_8621,N_8543,N_8414);
and U8622 (N_8622,N_8412,N_8434);
nand U8623 (N_8623,N_8566,N_8594);
and U8624 (N_8624,N_8401,N_8475);
nor U8625 (N_8625,N_8509,N_8445);
and U8626 (N_8626,N_8481,N_8438);
or U8627 (N_8627,N_8552,N_8575);
or U8628 (N_8628,N_8463,N_8495);
and U8629 (N_8629,N_8551,N_8430);
and U8630 (N_8630,N_8581,N_8596);
nor U8631 (N_8631,N_8582,N_8460);
nor U8632 (N_8632,N_8538,N_8577);
nand U8633 (N_8633,N_8571,N_8451);
nand U8634 (N_8634,N_8501,N_8427);
and U8635 (N_8635,N_8415,N_8464);
or U8636 (N_8636,N_8499,N_8556);
or U8637 (N_8637,N_8448,N_8567);
nor U8638 (N_8638,N_8530,N_8494);
nand U8639 (N_8639,N_8592,N_8505);
nor U8640 (N_8640,N_8423,N_8518);
or U8641 (N_8641,N_8457,N_8419);
nor U8642 (N_8642,N_8531,N_8400);
nand U8643 (N_8643,N_8580,N_8444);
nand U8644 (N_8644,N_8520,N_8511);
or U8645 (N_8645,N_8476,N_8485);
or U8646 (N_8646,N_8473,N_8420);
nand U8647 (N_8647,N_8570,N_8562);
or U8648 (N_8648,N_8524,N_8472);
and U8649 (N_8649,N_8521,N_8458);
and U8650 (N_8650,N_8437,N_8493);
and U8651 (N_8651,N_8496,N_8561);
nor U8652 (N_8652,N_8565,N_8417);
or U8653 (N_8653,N_8453,N_8573);
nand U8654 (N_8654,N_8489,N_8512);
and U8655 (N_8655,N_8508,N_8555);
nor U8656 (N_8656,N_8503,N_8569);
nand U8657 (N_8657,N_8431,N_8597);
or U8658 (N_8658,N_8442,N_8449);
and U8659 (N_8659,N_8502,N_8591);
or U8660 (N_8660,N_8572,N_8558);
or U8661 (N_8661,N_8510,N_8516);
nor U8662 (N_8662,N_8539,N_8544);
nand U8663 (N_8663,N_8497,N_8507);
and U8664 (N_8664,N_8528,N_8470);
and U8665 (N_8665,N_8576,N_8429);
or U8666 (N_8666,N_8461,N_8578);
nor U8667 (N_8667,N_8462,N_8443);
or U8668 (N_8668,N_8557,N_8598);
xnor U8669 (N_8669,N_8456,N_8450);
nand U8670 (N_8670,N_8440,N_8533);
nand U8671 (N_8671,N_8407,N_8525);
nor U8672 (N_8672,N_8586,N_8488);
nor U8673 (N_8673,N_8587,N_8479);
nand U8674 (N_8674,N_8410,N_8491);
nor U8675 (N_8675,N_8406,N_8477);
nand U8676 (N_8676,N_8532,N_8583);
nor U8677 (N_8677,N_8446,N_8515);
and U8678 (N_8678,N_8564,N_8519);
and U8679 (N_8679,N_8424,N_8593);
nor U8680 (N_8680,N_8478,N_8500);
or U8681 (N_8681,N_8469,N_8433);
or U8682 (N_8682,N_8588,N_8523);
and U8683 (N_8683,N_8574,N_8522);
nor U8684 (N_8684,N_8584,N_8465);
and U8685 (N_8685,N_8484,N_8559);
or U8686 (N_8686,N_8474,N_8483);
and U8687 (N_8687,N_8403,N_8408);
and U8688 (N_8688,N_8487,N_8490);
or U8689 (N_8689,N_8402,N_8550);
nor U8690 (N_8690,N_8546,N_8595);
or U8691 (N_8691,N_8526,N_8599);
nor U8692 (N_8692,N_8486,N_8425);
or U8693 (N_8693,N_8548,N_8540);
nor U8694 (N_8694,N_8560,N_8549);
xor U8695 (N_8695,N_8405,N_8468);
and U8696 (N_8696,N_8547,N_8439);
nor U8697 (N_8697,N_8498,N_8536);
or U8698 (N_8698,N_8537,N_8416);
or U8699 (N_8699,N_8529,N_8426);
nor U8700 (N_8700,N_8598,N_8594);
nor U8701 (N_8701,N_8428,N_8539);
and U8702 (N_8702,N_8431,N_8411);
or U8703 (N_8703,N_8419,N_8435);
or U8704 (N_8704,N_8427,N_8410);
or U8705 (N_8705,N_8493,N_8588);
nand U8706 (N_8706,N_8403,N_8515);
xnor U8707 (N_8707,N_8496,N_8539);
or U8708 (N_8708,N_8474,N_8462);
nand U8709 (N_8709,N_8507,N_8452);
and U8710 (N_8710,N_8535,N_8554);
and U8711 (N_8711,N_8458,N_8588);
nor U8712 (N_8712,N_8502,N_8457);
nor U8713 (N_8713,N_8461,N_8488);
nand U8714 (N_8714,N_8520,N_8582);
and U8715 (N_8715,N_8527,N_8447);
nor U8716 (N_8716,N_8539,N_8525);
nand U8717 (N_8717,N_8588,N_8490);
or U8718 (N_8718,N_8446,N_8448);
and U8719 (N_8719,N_8409,N_8532);
xnor U8720 (N_8720,N_8449,N_8597);
or U8721 (N_8721,N_8589,N_8412);
nor U8722 (N_8722,N_8580,N_8589);
and U8723 (N_8723,N_8470,N_8568);
and U8724 (N_8724,N_8407,N_8420);
and U8725 (N_8725,N_8417,N_8443);
nand U8726 (N_8726,N_8590,N_8457);
and U8727 (N_8727,N_8531,N_8453);
nand U8728 (N_8728,N_8402,N_8490);
nand U8729 (N_8729,N_8406,N_8413);
nand U8730 (N_8730,N_8433,N_8541);
nand U8731 (N_8731,N_8511,N_8440);
nor U8732 (N_8732,N_8442,N_8425);
and U8733 (N_8733,N_8458,N_8439);
nor U8734 (N_8734,N_8506,N_8408);
or U8735 (N_8735,N_8529,N_8542);
and U8736 (N_8736,N_8406,N_8508);
or U8737 (N_8737,N_8480,N_8519);
xor U8738 (N_8738,N_8595,N_8563);
nand U8739 (N_8739,N_8565,N_8408);
nor U8740 (N_8740,N_8457,N_8541);
nand U8741 (N_8741,N_8530,N_8412);
or U8742 (N_8742,N_8573,N_8516);
xnor U8743 (N_8743,N_8592,N_8442);
and U8744 (N_8744,N_8502,N_8445);
or U8745 (N_8745,N_8410,N_8540);
and U8746 (N_8746,N_8487,N_8429);
nand U8747 (N_8747,N_8435,N_8440);
and U8748 (N_8748,N_8484,N_8566);
and U8749 (N_8749,N_8408,N_8564);
and U8750 (N_8750,N_8540,N_8502);
nand U8751 (N_8751,N_8578,N_8522);
nand U8752 (N_8752,N_8583,N_8579);
nor U8753 (N_8753,N_8485,N_8434);
nor U8754 (N_8754,N_8545,N_8536);
nor U8755 (N_8755,N_8515,N_8547);
and U8756 (N_8756,N_8451,N_8416);
or U8757 (N_8757,N_8465,N_8566);
and U8758 (N_8758,N_8555,N_8493);
nor U8759 (N_8759,N_8515,N_8538);
nand U8760 (N_8760,N_8553,N_8513);
nor U8761 (N_8761,N_8461,N_8536);
nor U8762 (N_8762,N_8420,N_8539);
xnor U8763 (N_8763,N_8588,N_8530);
or U8764 (N_8764,N_8430,N_8438);
nor U8765 (N_8765,N_8466,N_8425);
nand U8766 (N_8766,N_8593,N_8470);
nor U8767 (N_8767,N_8469,N_8511);
and U8768 (N_8768,N_8427,N_8494);
or U8769 (N_8769,N_8592,N_8482);
or U8770 (N_8770,N_8576,N_8580);
and U8771 (N_8771,N_8528,N_8537);
or U8772 (N_8772,N_8416,N_8596);
or U8773 (N_8773,N_8529,N_8565);
or U8774 (N_8774,N_8444,N_8567);
or U8775 (N_8775,N_8532,N_8530);
or U8776 (N_8776,N_8596,N_8582);
and U8777 (N_8777,N_8545,N_8560);
and U8778 (N_8778,N_8547,N_8406);
nand U8779 (N_8779,N_8565,N_8506);
nor U8780 (N_8780,N_8433,N_8498);
and U8781 (N_8781,N_8533,N_8545);
and U8782 (N_8782,N_8533,N_8414);
and U8783 (N_8783,N_8540,N_8453);
nand U8784 (N_8784,N_8551,N_8588);
and U8785 (N_8785,N_8598,N_8456);
and U8786 (N_8786,N_8463,N_8487);
or U8787 (N_8787,N_8491,N_8564);
or U8788 (N_8788,N_8551,N_8526);
or U8789 (N_8789,N_8425,N_8532);
or U8790 (N_8790,N_8573,N_8410);
nor U8791 (N_8791,N_8435,N_8574);
or U8792 (N_8792,N_8409,N_8499);
nand U8793 (N_8793,N_8550,N_8444);
and U8794 (N_8794,N_8454,N_8423);
and U8795 (N_8795,N_8461,N_8432);
or U8796 (N_8796,N_8510,N_8419);
nand U8797 (N_8797,N_8595,N_8421);
and U8798 (N_8798,N_8510,N_8455);
xor U8799 (N_8799,N_8548,N_8564);
xor U8800 (N_8800,N_8655,N_8746);
nor U8801 (N_8801,N_8664,N_8780);
nor U8802 (N_8802,N_8745,N_8641);
nand U8803 (N_8803,N_8677,N_8744);
xnor U8804 (N_8804,N_8785,N_8720);
nor U8805 (N_8805,N_8615,N_8635);
nand U8806 (N_8806,N_8680,N_8600);
nand U8807 (N_8807,N_8732,N_8630);
or U8808 (N_8808,N_8726,N_8658);
or U8809 (N_8809,N_8652,N_8647);
or U8810 (N_8810,N_8638,N_8793);
nor U8811 (N_8811,N_8642,N_8712);
nor U8812 (N_8812,N_8684,N_8792);
nand U8813 (N_8813,N_8775,N_8737);
or U8814 (N_8814,N_8645,N_8715);
and U8815 (N_8815,N_8742,N_8623);
or U8816 (N_8816,N_8603,N_8781);
and U8817 (N_8817,N_8694,N_8782);
nor U8818 (N_8818,N_8665,N_8673);
or U8819 (N_8819,N_8735,N_8768);
nand U8820 (N_8820,N_8753,N_8749);
nand U8821 (N_8821,N_8707,N_8730);
nand U8822 (N_8822,N_8686,N_8788);
nor U8823 (N_8823,N_8644,N_8795);
nor U8824 (N_8824,N_8731,N_8696);
and U8825 (N_8825,N_8646,N_8692);
or U8826 (N_8826,N_8724,N_8794);
or U8827 (N_8827,N_8670,N_8761);
nor U8828 (N_8828,N_8725,N_8675);
xor U8829 (N_8829,N_8700,N_8659);
and U8830 (N_8830,N_8783,N_8637);
nor U8831 (N_8831,N_8769,N_8755);
or U8832 (N_8832,N_8619,N_8682);
nor U8833 (N_8833,N_8653,N_8657);
xor U8834 (N_8834,N_8674,N_8617);
and U8835 (N_8835,N_8727,N_8690);
nor U8836 (N_8836,N_8639,N_8671);
xnor U8837 (N_8837,N_8634,N_8743);
or U8838 (N_8838,N_8713,N_8602);
nand U8839 (N_8839,N_8799,N_8734);
nor U8840 (N_8840,N_8767,N_8778);
nor U8841 (N_8841,N_8679,N_8708);
nand U8842 (N_8842,N_8620,N_8625);
or U8843 (N_8843,N_8606,N_8758);
xor U8844 (N_8844,N_8759,N_8748);
nor U8845 (N_8845,N_8757,N_8672);
and U8846 (N_8846,N_8704,N_8756);
and U8847 (N_8847,N_8640,N_8777);
and U8848 (N_8848,N_8666,N_8702);
nor U8849 (N_8849,N_8669,N_8774);
or U8850 (N_8850,N_8699,N_8733);
or U8851 (N_8851,N_8689,N_8668);
nor U8852 (N_8852,N_8622,N_8791);
nand U8853 (N_8853,N_8698,N_8651);
nand U8854 (N_8854,N_8687,N_8693);
and U8855 (N_8855,N_8739,N_8604);
or U8856 (N_8856,N_8771,N_8648);
nand U8857 (N_8857,N_8628,N_8740);
and U8858 (N_8858,N_8701,N_8797);
or U8859 (N_8859,N_8705,N_8626);
nor U8860 (N_8860,N_8751,N_8773);
or U8861 (N_8861,N_8754,N_8770);
nand U8862 (N_8862,N_8656,N_8786);
nand U8863 (N_8863,N_8798,N_8632);
nor U8864 (N_8864,N_8613,N_8611);
and U8865 (N_8865,N_8681,N_8636);
nand U8866 (N_8866,N_8765,N_8661);
nand U8867 (N_8867,N_8763,N_8631);
and U8868 (N_8868,N_8663,N_8789);
xor U8869 (N_8869,N_8691,N_8633);
nand U8870 (N_8870,N_8752,N_8678);
nor U8871 (N_8871,N_8750,N_8784);
or U8872 (N_8872,N_8779,N_8710);
or U8873 (N_8873,N_8716,N_8790);
and U8874 (N_8874,N_8723,N_8612);
xnor U8875 (N_8875,N_8762,N_8736);
or U8876 (N_8876,N_8660,N_8741);
and U8877 (N_8877,N_8618,N_8719);
nand U8878 (N_8878,N_8711,N_8703);
or U8879 (N_8879,N_8697,N_8605);
and U8880 (N_8880,N_8721,N_8650);
or U8881 (N_8881,N_8614,N_8610);
or U8882 (N_8882,N_8616,N_8718);
and U8883 (N_8883,N_8760,N_8695);
or U8884 (N_8884,N_8621,N_8714);
nor U8885 (N_8885,N_8676,N_8683);
nor U8886 (N_8886,N_8609,N_8738);
and U8887 (N_8887,N_8772,N_8728);
nand U8888 (N_8888,N_8662,N_8688);
and U8889 (N_8889,N_8796,N_8729);
and U8890 (N_8890,N_8649,N_8627);
and U8891 (N_8891,N_8654,N_8764);
nand U8892 (N_8892,N_8776,N_8624);
and U8893 (N_8893,N_8601,N_8722);
nor U8894 (N_8894,N_8685,N_8747);
nor U8895 (N_8895,N_8706,N_8787);
nor U8896 (N_8896,N_8709,N_8608);
or U8897 (N_8897,N_8766,N_8667);
nor U8898 (N_8898,N_8643,N_8717);
and U8899 (N_8899,N_8629,N_8607);
xor U8900 (N_8900,N_8707,N_8608);
nand U8901 (N_8901,N_8736,N_8624);
nand U8902 (N_8902,N_8705,N_8718);
nor U8903 (N_8903,N_8702,N_8783);
or U8904 (N_8904,N_8625,N_8730);
nor U8905 (N_8905,N_8632,N_8721);
nor U8906 (N_8906,N_8718,N_8637);
or U8907 (N_8907,N_8655,N_8776);
and U8908 (N_8908,N_8756,N_8614);
or U8909 (N_8909,N_8664,N_8669);
xnor U8910 (N_8910,N_8778,N_8606);
or U8911 (N_8911,N_8659,N_8773);
and U8912 (N_8912,N_8741,N_8635);
nand U8913 (N_8913,N_8786,N_8611);
and U8914 (N_8914,N_8709,N_8630);
nand U8915 (N_8915,N_8791,N_8636);
nor U8916 (N_8916,N_8698,N_8619);
and U8917 (N_8917,N_8761,N_8783);
nor U8918 (N_8918,N_8758,N_8616);
nor U8919 (N_8919,N_8625,N_8609);
or U8920 (N_8920,N_8755,N_8648);
or U8921 (N_8921,N_8678,N_8699);
or U8922 (N_8922,N_8798,N_8688);
nand U8923 (N_8923,N_8723,N_8613);
xor U8924 (N_8924,N_8657,N_8608);
or U8925 (N_8925,N_8678,N_8672);
xor U8926 (N_8926,N_8733,N_8707);
and U8927 (N_8927,N_8689,N_8664);
nand U8928 (N_8928,N_8658,N_8651);
or U8929 (N_8929,N_8751,N_8775);
nor U8930 (N_8930,N_8754,N_8602);
nor U8931 (N_8931,N_8669,N_8670);
nand U8932 (N_8932,N_8634,N_8655);
or U8933 (N_8933,N_8631,N_8717);
nor U8934 (N_8934,N_8625,N_8715);
and U8935 (N_8935,N_8700,N_8738);
or U8936 (N_8936,N_8662,N_8628);
and U8937 (N_8937,N_8694,N_8745);
nor U8938 (N_8938,N_8718,N_8735);
or U8939 (N_8939,N_8759,N_8798);
nand U8940 (N_8940,N_8777,N_8753);
nor U8941 (N_8941,N_8690,N_8678);
and U8942 (N_8942,N_8794,N_8657);
nor U8943 (N_8943,N_8665,N_8751);
nor U8944 (N_8944,N_8776,N_8723);
nor U8945 (N_8945,N_8635,N_8629);
nor U8946 (N_8946,N_8711,N_8779);
nand U8947 (N_8947,N_8755,N_8763);
or U8948 (N_8948,N_8695,N_8691);
nor U8949 (N_8949,N_8794,N_8620);
and U8950 (N_8950,N_8797,N_8671);
and U8951 (N_8951,N_8675,N_8695);
nand U8952 (N_8952,N_8624,N_8716);
or U8953 (N_8953,N_8652,N_8602);
nor U8954 (N_8954,N_8767,N_8663);
nor U8955 (N_8955,N_8650,N_8722);
and U8956 (N_8956,N_8653,N_8680);
nand U8957 (N_8957,N_8625,N_8756);
nor U8958 (N_8958,N_8664,N_8760);
or U8959 (N_8959,N_8673,N_8725);
and U8960 (N_8960,N_8766,N_8683);
nand U8961 (N_8961,N_8623,N_8615);
nand U8962 (N_8962,N_8730,N_8757);
and U8963 (N_8963,N_8609,N_8662);
and U8964 (N_8964,N_8669,N_8642);
and U8965 (N_8965,N_8761,N_8679);
or U8966 (N_8966,N_8604,N_8767);
nor U8967 (N_8967,N_8695,N_8677);
xor U8968 (N_8968,N_8783,N_8669);
nor U8969 (N_8969,N_8798,N_8742);
xnor U8970 (N_8970,N_8741,N_8602);
or U8971 (N_8971,N_8664,N_8750);
and U8972 (N_8972,N_8608,N_8673);
and U8973 (N_8973,N_8613,N_8753);
or U8974 (N_8974,N_8603,N_8648);
nor U8975 (N_8975,N_8721,N_8607);
and U8976 (N_8976,N_8744,N_8664);
or U8977 (N_8977,N_8649,N_8776);
and U8978 (N_8978,N_8791,N_8650);
nor U8979 (N_8979,N_8619,N_8642);
xnor U8980 (N_8980,N_8640,N_8643);
and U8981 (N_8981,N_8769,N_8659);
nor U8982 (N_8982,N_8652,N_8731);
nor U8983 (N_8983,N_8725,N_8702);
nand U8984 (N_8984,N_8718,N_8714);
or U8985 (N_8985,N_8660,N_8702);
and U8986 (N_8986,N_8630,N_8658);
and U8987 (N_8987,N_8740,N_8677);
or U8988 (N_8988,N_8716,N_8660);
or U8989 (N_8989,N_8797,N_8608);
nand U8990 (N_8990,N_8719,N_8721);
or U8991 (N_8991,N_8758,N_8607);
nor U8992 (N_8992,N_8677,N_8647);
nand U8993 (N_8993,N_8775,N_8628);
nor U8994 (N_8994,N_8781,N_8645);
nand U8995 (N_8995,N_8780,N_8653);
nor U8996 (N_8996,N_8632,N_8614);
xor U8997 (N_8997,N_8678,N_8731);
nor U8998 (N_8998,N_8623,N_8782);
nor U8999 (N_8999,N_8649,N_8630);
or U9000 (N_9000,N_8961,N_8843);
or U9001 (N_9001,N_8975,N_8823);
nand U9002 (N_9002,N_8923,N_8864);
or U9003 (N_9003,N_8841,N_8996);
nor U9004 (N_9004,N_8819,N_8862);
nor U9005 (N_9005,N_8997,N_8908);
nor U9006 (N_9006,N_8968,N_8880);
or U9007 (N_9007,N_8884,N_8994);
and U9008 (N_9008,N_8954,N_8831);
nor U9009 (N_9009,N_8984,N_8826);
nor U9010 (N_9010,N_8910,N_8838);
or U9011 (N_9011,N_8893,N_8845);
and U9012 (N_9012,N_8883,N_8955);
nor U9013 (N_9013,N_8999,N_8947);
nor U9014 (N_9014,N_8974,N_8851);
and U9015 (N_9015,N_8988,N_8861);
and U9016 (N_9016,N_8816,N_8906);
and U9017 (N_9017,N_8922,N_8888);
nor U9018 (N_9018,N_8897,N_8875);
or U9019 (N_9019,N_8869,N_8813);
nor U9020 (N_9020,N_8944,N_8825);
xnor U9021 (N_9021,N_8927,N_8860);
xor U9022 (N_9022,N_8802,N_8980);
xnor U9023 (N_9023,N_8953,N_8806);
or U9024 (N_9024,N_8989,N_8842);
nand U9025 (N_9025,N_8814,N_8914);
or U9026 (N_9026,N_8858,N_8963);
and U9027 (N_9027,N_8801,N_8878);
or U9028 (N_9028,N_8934,N_8859);
and U9029 (N_9029,N_8931,N_8967);
nand U9030 (N_9030,N_8871,N_8949);
nor U9031 (N_9031,N_8853,N_8977);
nand U9032 (N_9032,N_8918,N_8822);
nand U9033 (N_9033,N_8900,N_8958);
and U9034 (N_9034,N_8857,N_8892);
nand U9035 (N_9035,N_8846,N_8965);
xor U9036 (N_9036,N_8956,N_8852);
or U9037 (N_9037,N_8925,N_8990);
nor U9038 (N_9038,N_8946,N_8948);
xor U9039 (N_9039,N_8837,N_8902);
nand U9040 (N_9040,N_8898,N_8836);
nand U9041 (N_9041,N_8926,N_8879);
or U9042 (N_9042,N_8964,N_8986);
or U9043 (N_9043,N_8848,N_8932);
and U9044 (N_9044,N_8978,N_8886);
xor U9045 (N_9045,N_8877,N_8920);
and U9046 (N_9046,N_8928,N_8889);
nor U9047 (N_9047,N_8844,N_8936);
xnor U9048 (N_9048,N_8976,N_8894);
xor U9049 (N_9049,N_8933,N_8809);
and U9050 (N_9050,N_8807,N_8921);
or U9051 (N_9051,N_8824,N_8873);
and U9052 (N_9052,N_8828,N_8972);
nand U9053 (N_9053,N_8985,N_8820);
nand U9054 (N_9054,N_8827,N_8973);
nand U9055 (N_9055,N_8867,N_8992);
nand U9056 (N_9056,N_8850,N_8830);
nand U9057 (N_9057,N_8885,N_8890);
and U9058 (N_9058,N_8959,N_8939);
nand U9059 (N_9059,N_8919,N_8821);
or U9060 (N_9060,N_8876,N_8929);
xnor U9061 (N_9061,N_8950,N_8901);
nand U9062 (N_9062,N_8833,N_8943);
and U9063 (N_9063,N_8941,N_8800);
and U9064 (N_9064,N_8979,N_8911);
xnor U9065 (N_9065,N_8991,N_8969);
xnor U9066 (N_9066,N_8863,N_8872);
and U9067 (N_9067,N_8896,N_8839);
nand U9068 (N_9068,N_8832,N_8812);
nor U9069 (N_9069,N_8811,N_8835);
nor U9070 (N_9070,N_8856,N_8993);
or U9071 (N_9071,N_8870,N_8840);
and U9072 (N_9072,N_8895,N_8935);
xnor U9073 (N_9073,N_8940,N_8909);
and U9074 (N_9074,N_8913,N_8887);
or U9075 (N_9075,N_8849,N_8881);
nor U9076 (N_9076,N_8866,N_8891);
or U9077 (N_9077,N_8907,N_8966);
nor U9078 (N_9078,N_8865,N_8915);
or U9079 (N_9079,N_8960,N_8882);
or U9080 (N_9080,N_8938,N_8981);
nor U9081 (N_9081,N_8904,N_8951);
and U9082 (N_9082,N_8957,N_8970);
nand U9083 (N_9083,N_8952,N_8905);
and U9084 (N_9084,N_8855,N_8818);
and U9085 (N_9085,N_8912,N_8810);
xnor U9086 (N_9086,N_8917,N_8803);
nand U9087 (N_9087,N_8916,N_8987);
nand U9088 (N_9088,N_8995,N_8930);
nand U9089 (N_9089,N_8924,N_8829);
nand U9090 (N_9090,N_8942,N_8983);
and U9091 (N_9091,N_8805,N_8971);
and U9092 (N_9092,N_8962,N_8854);
nand U9093 (N_9093,N_8903,N_8817);
or U9094 (N_9094,N_8847,N_8874);
or U9095 (N_9095,N_8982,N_8998);
nor U9096 (N_9096,N_8937,N_8808);
and U9097 (N_9097,N_8815,N_8899);
or U9098 (N_9098,N_8945,N_8834);
xnor U9099 (N_9099,N_8804,N_8868);
nor U9100 (N_9100,N_8893,N_8930);
and U9101 (N_9101,N_8996,N_8849);
xnor U9102 (N_9102,N_8942,N_8832);
nand U9103 (N_9103,N_8866,N_8832);
nand U9104 (N_9104,N_8838,N_8967);
nor U9105 (N_9105,N_8930,N_8950);
nand U9106 (N_9106,N_8843,N_8844);
nor U9107 (N_9107,N_8943,N_8843);
and U9108 (N_9108,N_8805,N_8825);
nand U9109 (N_9109,N_8963,N_8928);
nor U9110 (N_9110,N_8968,N_8917);
nand U9111 (N_9111,N_8948,N_8960);
nand U9112 (N_9112,N_8829,N_8904);
or U9113 (N_9113,N_8912,N_8821);
and U9114 (N_9114,N_8970,N_8865);
and U9115 (N_9115,N_8800,N_8963);
or U9116 (N_9116,N_8891,N_8997);
nor U9117 (N_9117,N_8971,N_8943);
nor U9118 (N_9118,N_8998,N_8988);
xnor U9119 (N_9119,N_8818,N_8995);
and U9120 (N_9120,N_8805,N_8816);
nand U9121 (N_9121,N_8899,N_8963);
nor U9122 (N_9122,N_8859,N_8920);
or U9123 (N_9123,N_8924,N_8989);
nor U9124 (N_9124,N_8873,N_8867);
nand U9125 (N_9125,N_8923,N_8947);
or U9126 (N_9126,N_8974,N_8924);
nand U9127 (N_9127,N_8943,N_8886);
nor U9128 (N_9128,N_8946,N_8813);
and U9129 (N_9129,N_8837,N_8938);
and U9130 (N_9130,N_8974,N_8840);
or U9131 (N_9131,N_8815,N_8895);
nand U9132 (N_9132,N_8859,N_8994);
nand U9133 (N_9133,N_8928,N_8824);
xnor U9134 (N_9134,N_8831,N_8988);
or U9135 (N_9135,N_8856,N_8965);
nand U9136 (N_9136,N_8803,N_8975);
and U9137 (N_9137,N_8956,N_8958);
nor U9138 (N_9138,N_8855,N_8951);
xor U9139 (N_9139,N_8817,N_8994);
and U9140 (N_9140,N_8949,N_8996);
or U9141 (N_9141,N_8876,N_8915);
nand U9142 (N_9142,N_8922,N_8865);
xnor U9143 (N_9143,N_8960,N_8929);
or U9144 (N_9144,N_8964,N_8880);
or U9145 (N_9145,N_8964,N_8953);
nor U9146 (N_9146,N_8969,N_8840);
xnor U9147 (N_9147,N_8958,N_8994);
and U9148 (N_9148,N_8883,N_8950);
and U9149 (N_9149,N_8908,N_8840);
or U9150 (N_9150,N_8826,N_8848);
xnor U9151 (N_9151,N_8925,N_8891);
nor U9152 (N_9152,N_8838,N_8994);
nand U9153 (N_9153,N_8818,N_8810);
or U9154 (N_9154,N_8800,N_8880);
or U9155 (N_9155,N_8875,N_8937);
or U9156 (N_9156,N_8967,N_8827);
and U9157 (N_9157,N_8807,N_8987);
and U9158 (N_9158,N_8991,N_8955);
or U9159 (N_9159,N_8918,N_8925);
xnor U9160 (N_9160,N_8859,N_8927);
nand U9161 (N_9161,N_8806,N_8907);
nor U9162 (N_9162,N_8885,N_8864);
and U9163 (N_9163,N_8905,N_8802);
or U9164 (N_9164,N_8852,N_8889);
or U9165 (N_9165,N_8999,N_8967);
nor U9166 (N_9166,N_8875,N_8976);
nand U9167 (N_9167,N_8899,N_8985);
nor U9168 (N_9168,N_8902,N_8921);
xnor U9169 (N_9169,N_8833,N_8812);
or U9170 (N_9170,N_8807,N_8931);
or U9171 (N_9171,N_8996,N_8872);
xor U9172 (N_9172,N_8957,N_8827);
nand U9173 (N_9173,N_8931,N_8802);
and U9174 (N_9174,N_8960,N_8858);
and U9175 (N_9175,N_8926,N_8866);
or U9176 (N_9176,N_8857,N_8928);
nor U9177 (N_9177,N_8902,N_8911);
or U9178 (N_9178,N_8930,N_8966);
nor U9179 (N_9179,N_8836,N_8913);
xnor U9180 (N_9180,N_8977,N_8800);
nand U9181 (N_9181,N_8997,N_8974);
xnor U9182 (N_9182,N_8977,N_8803);
nor U9183 (N_9183,N_8826,N_8836);
or U9184 (N_9184,N_8849,N_8913);
or U9185 (N_9185,N_8962,N_8803);
nor U9186 (N_9186,N_8897,N_8836);
or U9187 (N_9187,N_8889,N_8845);
nand U9188 (N_9188,N_8995,N_8806);
and U9189 (N_9189,N_8923,N_8983);
nand U9190 (N_9190,N_8902,N_8842);
and U9191 (N_9191,N_8905,N_8913);
nor U9192 (N_9192,N_8879,N_8809);
and U9193 (N_9193,N_8985,N_8916);
and U9194 (N_9194,N_8838,N_8807);
xor U9195 (N_9195,N_8954,N_8967);
nand U9196 (N_9196,N_8859,N_8851);
and U9197 (N_9197,N_8974,N_8915);
xor U9198 (N_9198,N_8901,N_8939);
nand U9199 (N_9199,N_8895,N_8831);
and U9200 (N_9200,N_9145,N_9031);
or U9201 (N_9201,N_9149,N_9192);
nor U9202 (N_9202,N_9148,N_9179);
nand U9203 (N_9203,N_9075,N_9073);
nor U9204 (N_9204,N_9110,N_9000);
and U9205 (N_9205,N_9109,N_9135);
xnor U9206 (N_9206,N_9144,N_9166);
xnor U9207 (N_9207,N_9060,N_9199);
or U9208 (N_9208,N_9159,N_9011);
or U9209 (N_9209,N_9175,N_9098);
and U9210 (N_9210,N_9133,N_9162);
or U9211 (N_9211,N_9029,N_9112);
and U9212 (N_9212,N_9102,N_9129);
or U9213 (N_9213,N_9055,N_9045);
and U9214 (N_9214,N_9051,N_9044);
nand U9215 (N_9215,N_9082,N_9131);
nand U9216 (N_9216,N_9089,N_9063);
or U9217 (N_9217,N_9189,N_9118);
or U9218 (N_9218,N_9081,N_9009);
nand U9219 (N_9219,N_9168,N_9076);
nor U9220 (N_9220,N_9190,N_9062);
or U9221 (N_9221,N_9172,N_9163);
nand U9222 (N_9222,N_9068,N_9121);
or U9223 (N_9223,N_9003,N_9173);
xor U9224 (N_9224,N_9197,N_9174);
nand U9225 (N_9225,N_9128,N_9139);
nand U9226 (N_9226,N_9085,N_9065);
or U9227 (N_9227,N_9191,N_9117);
and U9228 (N_9228,N_9134,N_9050);
xnor U9229 (N_9229,N_9052,N_9100);
nand U9230 (N_9230,N_9183,N_9024);
nor U9231 (N_9231,N_9083,N_9171);
and U9232 (N_9232,N_9026,N_9103);
or U9233 (N_9233,N_9164,N_9165);
or U9234 (N_9234,N_9027,N_9104);
nor U9235 (N_9235,N_9157,N_9080);
nor U9236 (N_9236,N_9049,N_9096);
and U9237 (N_9237,N_9125,N_9116);
or U9238 (N_9238,N_9167,N_9105);
or U9239 (N_9239,N_9115,N_9039);
xnor U9240 (N_9240,N_9095,N_9037);
nor U9241 (N_9241,N_9023,N_9017);
nor U9242 (N_9242,N_9016,N_9067);
or U9243 (N_9243,N_9053,N_9072);
nand U9244 (N_9244,N_9140,N_9180);
nand U9245 (N_9245,N_9176,N_9142);
or U9246 (N_9246,N_9113,N_9141);
or U9247 (N_9247,N_9119,N_9152);
nand U9248 (N_9248,N_9097,N_9106);
and U9249 (N_9249,N_9021,N_9198);
or U9250 (N_9250,N_9187,N_9136);
and U9251 (N_9251,N_9132,N_9182);
nand U9252 (N_9252,N_9070,N_9127);
or U9253 (N_9253,N_9040,N_9099);
nand U9254 (N_9254,N_9043,N_9177);
or U9255 (N_9255,N_9087,N_9086);
and U9256 (N_9256,N_9146,N_9126);
nand U9257 (N_9257,N_9088,N_9046);
and U9258 (N_9258,N_9057,N_9091);
and U9259 (N_9259,N_9158,N_9169);
nand U9260 (N_9260,N_9194,N_9147);
xnor U9261 (N_9261,N_9001,N_9004);
xnor U9262 (N_9262,N_9150,N_9079);
and U9263 (N_9263,N_9008,N_9030);
nor U9264 (N_9264,N_9005,N_9094);
and U9265 (N_9265,N_9042,N_9059);
nor U9266 (N_9266,N_9090,N_9074);
nand U9267 (N_9267,N_9114,N_9036);
nor U9268 (N_9268,N_9012,N_9120);
xnor U9269 (N_9269,N_9041,N_9122);
xor U9270 (N_9270,N_9178,N_9066);
and U9271 (N_9271,N_9124,N_9056);
or U9272 (N_9272,N_9108,N_9064);
xor U9273 (N_9273,N_9123,N_9002);
nand U9274 (N_9274,N_9181,N_9020);
or U9275 (N_9275,N_9032,N_9084);
xnor U9276 (N_9276,N_9093,N_9019);
and U9277 (N_9277,N_9170,N_9156);
nor U9278 (N_9278,N_9022,N_9058);
or U9279 (N_9279,N_9061,N_9015);
and U9280 (N_9280,N_9138,N_9054);
or U9281 (N_9281,N_9101,N_9048);
and U9282 (N_9282,N_9107,N_9196);
xor U9283 (N_9283,N_9137,N_9078);
nand U9284 (N_9284,N_9155,N_9014);
or U9285 (N_9285,N_9035,N_9033);
and U9286 (N_9286,N_9007,N_9153);
or U9287 (N_9287,N_9186,N_9034);
and U9288 (N_9288,N_9111,N_9013);
or U9289 (N_9289,N_9151,N_9071);
or U9290 (N_9290,N_9193,N_9195);
nor U9291 (N_9291,N_9092,N_9047);
and U9292 (N_9292,N_9161,N_9160);
and U9293 (N_9293,N_9010,N_9130);
nand U9294 (N_9294,N_9028,N_9069);
xor U9295 (N_9295,N_9077,N_9188);
and U9296 (N_9296,N_9143,N_9185);
nand U9297 (N_9297,N_9006,N_9025);
nand U9298 (N_9298,N_9154,N_9184);
or U9299 (N_9299,N_9018,N_9038);
xor U9300 (N_9300,N_9139,N_9195);
xnor U9301 (N_9301,N_9073,N_9109);
and U9302 (N_9302,N_9059,N_9108);
and U9303 (N_9303,N_9005,N_9110);
xor U9304 (N_9304,N_9117,N_9034);
nand U9305 (N_9305,N_9083,N_9178);
and U9306 (N_9306,N_9001,N_9082);
and U9307 (N_9307,N_9076,N_9173);
xor U9308 (N_9308,N_9181,N_9006);
and U9309 (N_9309,N_9027,N_9008);
and U9310 (N_9310,N_9099,N_9069);
nand U9311 (N_9311,N_9149,N_9027);
and U9312 (N_9312,N_9155,N_9075);
and U9313 (N_9313,N_9188,N_9034);
nand U9314 (N_9314,N_9049,N_9005);
and U9315 (N_9315,N_9063,N_9114);
nand U9316 (N_9316,N_9011,N_9186);
and U9317 (N_9317,N_9001,N_9085);
or U9318 (N_9318,N_9186,N_9055);
or U9319 (N_9319,N_9074,N_9024);
and U9320 (N_9320,N_9012,N_9160);
xnor U9321 (N_9321,N_9026,N_9176);
xor U9322 (N_9322,N_9054,N_9096);
nor U9323 (N_9323,N_9044,N_9156);
and U9324 (N_9324,N_9056,N_9122);
or U9325 (N_9325,N_9119,N_9076);
and U9326 (N_9326,N_9109,N_9115);
nand U9327 (N_9327,N_9127,N_9094);
xor U9328 (N_9328,N_9122,N_9177);
and U9329 (N_9329,N_9056,N_9119);
and U9330 (N_9330,N_9189,N_9193);
nor U9331 (N_9331,N_9096,N_9061);
xor U9332 (N_9332,N_9130,N_9071);
nand U9333 (N_9333,N_9138,N_9101);
or U9334 (N_9334,N_9025,N_9131);
xnor U9335 (N_9335,N_9057,N_9077);
and U9336 (N_9336,N_9152,N_9110);
nor U9337 (N_9337,N_9039,N_9145);
nor U9338 (N_9338,N_9111,N_9099);
and U9339 (N_9339,N_9176,N_9173);
or U9340 (N_9340,N_9016,N_9178);
and U9341 (N_9341,N_9082,N_9009);
nor U9342 (N_9342,N_9108,N_9096);
or U9343 (N_9343,N_9180,N_9056);
and U9344 (N_9344,N_9173,N_9063);
nand U9345 (N_9345,N_9042,N_9076);
and U9346 (N_9346,N_9047,N_9024);
nor U9347 (N_9347,N_9112,N_9110);
nor U9348 (N_9348,N_9094,N_9178);
nor U9349 (N_9349,N_9017,N_9185);
nor U9350 (N_9350,N_9091,N_9151);
and U9351 (N_9351,N_9148,N_9168);
nor U9352 (N_9352,N_9088,N_9018);
nor U9353 (N_9353,N_9040,N_9160);
nor U9354 (N_9354,N_9119,N_9187);
nand U9355 (N_9355,N_9025,N_9031);
or U9356 (N_9356,N_9198,N_9178);
nor U9357 (N_9357,N_9107,N_9147);
nor U9358 (N_9358,N_9006,N_9051);
and U9359 (N_9359,N_9136,N_9019);
and U9360 (N_9360,N_9169,N_9054);
nand U9361 (N_9361,N_9160,N_9137);
nand U9362 (N_9362,N_9116,N_9141);
or U9363 (N_9363,N_9022,N_9017);
or U9364 (N_9364,N_9199,N_9155);
xnor U9365 (N_9365,N_9041,N_9018);
nor U9366 (N_9366,N_9030,N_9095);
and U9367 (N_9367,N_9119,N_9191);
or U9368 (N_9368,N_9169,N_9044);
and U9369 (N_9369,N_9074,N_9089);
nor U9370 (N_9370,N_9141,N_9175);
nor U9371 (N_9371,N_9146,N_9086);
or U9372 (N_9372,N_9059,N_9048);
or U9373 (N_9373,N_9136,N_9064);
nand U9374 (N_9374,N_9031,N_9055);
and U9375 (N_9375,N_9064,N_9094);
or U9376 (N_9376,N_9051,N_9071);
or U9377 (N_9377,N_9170,N_9040);
nor U9378 (N_9378,N_9136,N_9038);
or U9379 (N_9379,N_9036,N_9055);
and U9380 (N_9380,N_9086,N_9017);
nor U9381 (N_9381,N_9074,N_9009);
nand U9382 (N_9382,N_9168,N_9005);
or U9383 (N_9383,N_9081,N_9189);
and U9384 (N_9384,N_9140,N_9045);
or U9385 (N_9385,N_9018,N_9188);
nor U9386 (N_9386,N_9082,N_9088);
nand U9387 (N_9387,N_9112,N_9184);
or U9388 (N_9388,N_9014,N_9066);
and U9389 (N_9389,N_9009,N_9127);
nand U9390 (N_9390,N_9059,N_9175);
or U9391 (N_9391,N_9040,N_9103);
or U9392 (N_9392,N_9141,N_9197);
xor U9393 (N_9393,N_9161,N_9019);
or U9394 (N_9394,N_9078,N_9161);
nand U9395 (N_9395,N_9191,N_9187);
and U9396 (N_9396,N_9001,N_9047);
nor U9397 (N_9397,N_9148,N_9087);
and U9398 (N_9398,N_9127,N_9004);
and U9399 (N_9399,N_9086,N_9149);
and U9400 (N_9400,N_9288,N_9374);
nor U9401 (N_9401,N_9232,N_9264);
nor U9402 (N_9402,N_9315,N_9205);
or U9403 (N_9403,N_9281,N_9202);
xnor U9404 (N_9404,N_9214,N_9295);
and U9405 (N_9405,N_9370,N_9316);
nor U9406 (N_9406,N_9361,N_9268);
nor U9407 (N_9407,N_9274,N_9373);
nor U9408 (N_9408,N_9320,N_9350);
or U9409 (N_9409,N_9228,N_9211);
nor U9410 (N_9410,N_9207,N_9297);
or U9411 (N_9411,N_9254,N_9203);
or U9412 (N_9412,N_9383,N_9356);
or U9413 (N_9413,N_9218,N_9200);
and U9414 (N_9414,N_9275,N_9349);
and U9415 (N_9415,N_9330,N_9221);
or U9416 (N_9416,N_9265,N_9319);
nor U9417 (N_9417,N_9276,N_9352);
nor U9418 (N_9418,N_9227,N_9266);
xor U9419 (N_9419,N_9269,N_9306);
and U9420 (N_9420,N_9393,N_9236);
nand U9421 (N_9421,N_9229,N_9286);
and U9422 (N_9422,N_9395,N_9251);
nor U9423 (N_9423,N_9230,N_9293);
nor U9424 (N_9424,N_9308,N_9325);
xnor U9425 (N_9425,N_9209,N_9382);
nand U9426 (N_9426,N_9327,N_9260);
nor U9427 (N_9427,N_9380,N_9307);
and U9428 (N_9428,N_9305,N_9240);
or U9429 (N_9429,N_9375,N_9273);
nand U9430 (N_9430,N_9242,N_9311);
and U9431 (N_9431,N_9348,N_9280);
nand U9432 (N_9432,N_9359,N_9290);
or U9433 (N_9433,N_9289,N_9340);
or U9434 (N_9434,N_9335,N_9398);
nor U9435 (N_9435,N_9353,N_9285);
and U9436 (N_9436,N_9296,N_9376);
or U9437 (N_9437,N_9368,N_9313);
nor U9438 (N_9438,N_9371,N_9256);
nand U9439 (N_9439,N_9241,N_9360);
nor U9440 (N_9440,N_9392,N_9252);
nor U9441 (N_9441,N_9381,N_9329);
and U9442 (N_9442,N_9226,N_9346);
and U9443 (N_9443,N_9345,N_9364);
nand U9444 (N_9444,N_9238,N_9250);
nand U9445 (N_9445,N_9336,N_9222);
and U9446 (N_9446,N_9337,N_9271);
and U9447 (N_9447,N_9219,N_9216);
or U9448 (N_9448,N_9323,N_9237);
and U9449 (N_9449,N_9302,N_9261);
and U9450 (N_9450,N_9235,N_9388);
nand U9451 (N_9451,N_9365,N_9326);
and U9452 (N_9452,N_9386,N_9262);
nor U9453 (N_9453,N_9298,N_9201);
or U9454 (N_9454,N_9246,N_9377);
xor U9455 (N_9455,N_9332,N_9304);
or U9456 (N_9456,N_9292,N_9247);
nand U9457 (N_9457,N_9355,N_9314);
nand U9458 (N_9458,N_9263,N_9391);
nor U9459 (N_9459,N_9249,N_9294);
nand U9460 (N_9460,N_9309,N_9328);
nor U9461 (N_9461,N_9378,N_9284);
and U9462 (N_9462,N_9253,N_9208);
nor U9463 (N_9463,N_9317,N_9367);
nand U9464 (N_9464,N_9257,N_9267);
and U9465 (N_9465,N_9372,N_9341);
and U9466 (N_9466,N_9212,N_9239);
nand U9467 (N_9467,N_9389,N_9301);
or U9468 (N_9468,N_9343,N_9399);
nor U9469 (N_9469,N_9344,N_9258);
nor U9470 (N_9470,N_9390,N_9234);
or U9471 (N_9471,N_9259,N_9223);
nor U9472 (N_9472,N_9366,N_9397);
or U9473 (N_9473,N_9231,N_9333);
and U9474 (N_9474,N_9217,N_9233);
and U9475 (N_9475,N_9358,N_9282);
and U9476 (N_9476,N_9255,N_9324);
nor U9477 (N_9477,N_9322,N_9387);
xor U9478 (N_9478,N_9351,N_9342);
xnor U9479 (N_9479,N_9334,N_9379);
nand U9480 (N_9480,N_9303,N_9204);
xnor U9481 (N_9481,N_9243,N_9300);
xor U9482 (N_9482,N_9287,N_9225);
nor U9483 (N_9483,N_9385,N_9278);
or U9484 (N_9484,N_9394,N_9310);
or U9485 (N_9485,N_9396,N_9210);
nand U9486 (N_9486,N_9384,N_9248);
or U9487 (N_9487,N_9279,N_9299);
and U9488 (N_9488,N_9318,N_9272);
and U9489 (N_9489,N_9224,N_9220);
or U9490 (N_9490,N_9213,N_9244);
xnor U9491 (N_9491,N_9331,N_9321);
nor U9492 (N_9492,N_9277,N_9357);
nand U9493 (N_9493,N_9363,N_9339);
nor U9494 (N_9494,N_9283,N_9354);
nand U9495 (N_9495,N_9206,N_9270);
or U9496 (N_9496,N_9245,N_9347);
xor U9497 (N_9497,N_9291,N_9338);
and U9498 (N_9498,N_9362,N_9215);
nor U9499 (N_9499,N_9312,N_9369);
nand U9500 (N_9500,N_9214,N_9284);
and U9501 (N_9501,N_9378,N_9330);
xor U9502 (N_9502,N_9291,N_9205);
and U9503 (N_9503,N_9238,N_9209);
and U9504 (N_9504,N_9202,N_9323);
nand U9505 (N_9505,N_9298,N_9282);
nand U9506 (N_9506,N_9335,N_9278);
and U9507 (N_9507,N_9220,N_9262);
nand U9508 (N_9508,N_9370,N_9360);
or U9509 (N_9509,N_9379,N_9204);
nand U9510 (N_9510,N_9366,N_9208);
and U9511 (N_9511,N_9246,N_9382);
nand U9512 (N_9512,N_9397,N_9340);
or U9513 (N_9513,N_9291,N_9361);
nor U9514 (N_9514,N_9284,N_9250);
or U9515 (N_9515,N_9208,N_9254);
or U9516 (N_9516,N_9236,N_9368);
nand U9517 (N_9517,N_9304,N_9212);
nand U9518 (N_9518,N_9364,N_9293);
or U9519 (N_9519,N_9210,N_9233);
nor U9520 (N_9520,N_9204,N_9201);
and U9521 (N_9521,N_9356,N_9359);
or U9522 (N_9522,N_9304,N_9247);
nor U9523 (N_9523,N_9322,N_9278);
nand U9524 (N_9524,N_9243,N_9340);
or U9525 (N_9525,N_9359,N_9355);
nor U9526 (N_9526,N_9309,N_9369);
and U9527 (N_9527,N_9293,N_9277);
nor U9528 (N_9528,N_9236,N_9311);
nand U9529 (N_9529,N_9395,N_9236);
nor U9530 (N_9530,N_9340,N_9219);
nand U9531 (N_9531,N_9215,N_9308);
nand U9532 (N_9532,N_9343,N_9285);
and U9533 (N_9533,N_9345,N_9220);
or U9534 (N_9534,N_9280,N_9282);
nor U9535 (N_9535,N_9345,N_9335);
and U9536 (N_9536,N_9336,N_9367);
nor U9537 (N_9537,N_9341,N_9208);
or U9538 (N_9538,N_9298,N_9398);
nor U9539 (N_9539,N_9310,N_9214);
nor U9540 (N_9540,N_9353,N_9281);
and U9541 (N_9541,N_9253,N_9320);
or U9542 (N_9542,N_9355,N_9213);
nand U9543 (N_9543,N_9321,N_9327);
nor U9544 (N_9544,N_9271,N_9345);
and U9545 (N_9545,N_9214,N_9228);
nand U9546 (N_9546,N_9261,N_9373);
nand U9547 (N_9547,N_9340,N_9309);
nor U9548 (N_9548,N_9363,N_9245);
nand U9549 (N_9549,N_9369,N_9224);
nor U9550 (N_9550,N_9337,N_9322);
nand U9551 (N_9551,N_9221,N_9383);
nor U9552 (N_9552,N_9282,N_9350);
or U9553 (N_9553,N_9297,N_9283);
nor U9554 (N_9554,N_9339,N_9347);
or U9555 (N_9555,N_9390,N_9278);
or U9556 (N_9556,N_9230,N_9302);
or U9557 (N_9557,N_9378,N_9295);
nand U9558 (N_9558,N_9204,N_9275);
nor U9559 (N_9559,N_9321,N_9360);
or U9560 (N_9560,N_9319,N_9311);
nand U9561 (N_9561,N_9371,N_9253);
xnor U9562 (N_9562,N_9396,N_9360);
or U9563 (N_9563,N_9378,N_9230);
or U9564 (N_9564,N_9234,N_9237);
nand U9565 (N_9565,N_9252,N_9312);
nand U9566 (N_9566,N_9372,N_9220);
or U9567 (N_9567,N_9305,N_9332);
and U9568 (N_9568,N_9373,N_9211);
nor U9569 (N_9569,N_9281,N_9265);
and U9570 (N_9570,N_9286,N_9215);
and U9571 (N_9571,N_9344,N_9219);
nand U9572 (N_9572,N_9227,N_9282);
or U9573 (N_9573,N_9316,N_9234);
and U9574 (N_9574,N_9228,N_9343);
nor U9575 (N_9575,N_9239,N_9208);
xor U9576 (N_9576,N_9378,N_9345);
nor U9577 (N_9577,N_9292,N_9251);
nor U9578 (N_9578,N_9214,N_9392);
nor U9579 (N_9579,N_9263,N_9393);
nand U9580 (N_9580,N_9233,N_9317);
nand U9581 (N_9581,N_9356,N_9398);
nand U9582 (N_9582,N_9244,N_9338);
nand U9583 (N_9583,N_9307,N_9250);
and U9584 (N_9584,N_9341,N_9248);
nor U9585 (N_9585,N_9363,N_9322);
nor U9586 (N_9586,N_9228,N_9346);
nor U9587 (N_9587,N_9388,N_9253);
or U9588 (N_9588,N_9329,N_9355);
nor U9589 (N_9589,N_9390,N_9305);
nand U9590 (N_9590,N_9271,N_9280);
or U9591 (N_9591,N_9333,N_9338);
nand U9592 (N_9592,N_9381,N_9264);
and U9593 (N_9593,N_9332,N_9338);
nand U9594 (N_9594,N_9286,N_9214);
nor U9595 (N_9595,N_9386,N_9350);
or U9596 (N_9596,N_9223,N_9209);
nand U9597 (N_9597,N_9261,N_9307);
or U9598 (N_9598,N_9373,N_9267);
and U9599 (N_9599,N_9381,N_9368);
nor U9600 (N_9600,N_9481,N_9480);
and U9601 (N_9601,N_9556,N_9502);
or U9602 (N_9602,N_9414,N_9529);
nand U9603 (N_9603,N_9458,N_9571);
nor U9604 (N_9604,N_9585,N_9555);
and U9605 (N_9605,N_9425,N_9479);
and U9606 (N_9606,N_9440,N_9509);
or U9607 (N_9607,N_9558,N_9421);
nor U9608 (N_9608,N_9550,N_9514);
nor U9609 (N_9609,N_9415,N_9438);
nand U9610 (N_9610,N_9590,N_9548);
xnor U9611 (N_9611,N_9586,N_9576);
or U9612 (N_9612,N_9431,N_9582);
nand U9613 (N_9613,N_9460,N_9557);
nor U9614 (N_9614,N_9504,N_9473);
nor U9615 (N_9615,N_9450,N_9443);
nand U9616 (N_9616,N_9523,N_9562);
xnor U9617 (N_9617,N_9467,N_9498);
nor U9618 (N_9618,N_9553,N_9537);
or U9619 (N_9619,N_9486,N_9488);
or U9620 (N_9620,N_9566,N_9567);
xor U9621 (N_9621,N_9409,N_9511);
nor U9622 (N_9622,N_9494,N_9452);
or U9623 (N_9623,N_9500,N_9598);
nor U9624 (N_9624,N_9591,N_9441);
and U9625 (N_9625,N_9540,N_9516);
nor U9626 (N_9626,N_9515,N_9564);
nor U9627 (N_9627,N_9594,N_9573);
nor U9628 (N_9628,N_9401,N_9593);
or U9629 (N_9629,N_9413,N_9448);
or U9630 (N_9630,N_9539,N_9536);
nor U9631 (N_9631,N_9478,N_9424);
nor U9632 (N_9632,N_9459,N_9496);
or U9633 (N_9633,N_9457,N_9595);
and U9634 (N_9634,N_9545,N_9422);
and U9635 (N_9635,N_9597,N_9417);
and U9636 (N_9636,N_9411,N_9507);
nand U9637 (N_9637,N_9531,N_9577);
and U9638 (N_9638,N_9472,N_9474);
nand U9639 (N_9639,N_9569,N_9489);
nand U9640 (N_9640,N_9400,N_9455);
or U9641 (N_9641,N_9527,N_9596);
nand U9642 (N_9642,N_9552,N_9461);
nand U9643 (N_9643,N_9407,N_9532);
nand U9644 (N_9644,N_9416,N_9547);
or U9645 (N_9645,N_9512,N_9442);
xnor U9646 (N_9646,N_9477,N_9549);
xnor U9647 (N_9647,N_9592,N_9575);
or U9648 (N_9648,N_9476,N_9538);
nand U9649 (N_9649,N_9439,N_9453);
nand U9650 (N_9650,N_9517,N_9454);
nor U9651 (N_9651,N_9584,N_9587);
xor U9652 (N_9652,N_9521,N_9470);
and U9653 (N_9653,N_9526,N_9497);
nor U9654 (N_9654,N_9519,N_9508);
nor U9655 (N_9655,N_9465,N_9463);
xor U9656 (N_9656,N_9501,N_9492);
or U9657 (N_9657,N_9551,N_9403);
or U9658 (N_9658,N_9433,N_9530);
and U9659 (N_9659,N_9437,N_9589);
nor U9660 (N_9660,N_9543,N_9542);
or U9661 (N_9661,N_9466,N_9432);
nand U9662 (N_9662,N_9434,N_9491);
xor U9663 (N_9663,N_9580,N_9525);
or U9664 (N_9664,N_9588,N_9565);
xnor U9665 (N_9665,N_9462,N_9449);
nor U9666 (N_9666,N_9469,N_9471);
or U9667 (N_9667,N_9495,N_9524);
nor U9668 (N_9668,N_9546,N_9563);
nand U9669 (N_9669,N_9499,N_9483);
and U9670 (N_9670,N_9485,N_9554);
and U9671 (N_9671,N_9406,N_9518);
nor U9672 (N_9672,N_9419,N_9506);
nor U9673 (N_9673,N_9559,N_9560);
nand U9674 (N_9674,N_9599,N_9578);
or U9675 (N_9675,N_9446,N_9544);
and U9676 (N_9676,N_9445,N_9534);
nand U9677 (N_9677,N_9561,N_9484);
nor U9678 (N_9678,N_9493,N_9570);
nand U9679 (N_9679,N_9513,N_9475);
and U9680 (N_9680,N_9420,N_9429);
or U9681 (N_9681,N_9505,N_9487);
or U9682 (N_9682,N_9541,N_9444);
and U9683 (N_9683,N_9410,N_9581);
nor U9684 (N_9684,N_9412,N_9418);
xnor U9685 (N_9685,N_9456,N_9535);
and U9686 (N_9686,N_9436,N_9464);
xnor U9687 (N_9687,N_9579,N_9528);
and U9688 (N_9688,N_9405,N_9574);
xor U9689 (N_9689,N_9426,N_9522);
nor U9690 (N_9690,N_9490,N_9451);
nand U9691 (N_9691,N_9428,N_9468);
or U9692 (N_9692,N_9402,N_9568);
or U9693 (N_9693,N_9447,N_9533);
xnor U9694 (N_9694,N_9583,N_9520);
nor U9695 (N_9695,N_9408,N_9404);
or U9696 (N_9696,N_9572,N_9430);
nor U9697 (N_9697,N_9423,N_9510);
nand U9698 (N_9698,N_9482,N_9427);
and U9699 (N_9699,N_9435,N_9503);
nand U9700 (N_9700,N_9520,N_9481);
nor U9701 (N_9701,N_9534,N_9458);
nand U9702 (N_9702,N_9471,N_9523);
nand U9703 (N_9703,N_9464,N_9493);
nand U9704 (N_9704,N_9524,N_9579);
nand U9705 (N_9705,N_9481,N_9446);
nor U9706 (N_9706,N_9465,N_9575);
and U9707 (N_9707,N_9519,N_9576);
and U9708 (N_9708,N_9514,N_9433);
and U9709 (N_9709,N_9496,N_9544);
nand U9710 (N_9710,N_9564,N_9506);
or U9711 (N_9711,N_9584,N_9541);
and U9712 (N_9712,N_9582,N_9548);
or U9713 (N_9713,N_9446,N_9422);
or U9714 (N_9714,N_9572,N_9442);
xnor U9715 (N_9715,N_9599,N_9593);
nor U9716 (N_9716,N_9430,N_9427);
or U9717 (N_9717,N_9480,N_9554);
nor U9718 (N_9718,N_9580,N_9478);
nor U9719 (N_9719,N_9551,N_9552);
and U9720 (N_9720,N_9533,N_9584);
xnor U9721 (N_9721,N_9567,N_9559);
or U9722 (N_9722,N_9458,N_9489);
nor U9723 (N_9723,N_9495,N_9480);
nand U9724 (N_9724,N_9430,N_9406);
nor U9725 (N_9725,N_9450,N_9531);
nand U9726 (N_9726,N_9548,N_9500);
and U9727 (N_9727,N_9566,N_9596);
xor U9728 (N_9728,N_9403,N_9503);
nand U9729 (N_9729,N_9569,N_9460);
nor U9730 (N_9730,N_9559,N_9517);
nor U9731 (N_9731,N_9491,N_9587);
nand U9732 (N_9732,N_9546,N_9540);
nor U9733 (N_9733,N_9524,N_9443);
nor U9734 (N_9734,N_9490,N_9487);
nand U9735 (N_9735,N_9437,N_9577);
and U9736 (N_9736,N_9573,N_9414);
or U9737 (N_9737,N_9403,N_9495);
nor U9738 (N_9738,N_9437,N_9554);
and U9739 (N_9739,N_9548,N_9449);
nor U9740 (N_9740,N_9406,N_9482);
xnor U9741 (N_9741,N_9579,N_9527);
nand U9742 (N_9742,N_9561,N_9480);
nor U9743 (N_9743,N_9559,N_9490);
nor U9744 (N_9744,N_9443,N_9422);
nor U9745 (N_9745,N_9555,N_9460);
nor U9746 (N_9746,N_9439,N_9518);
and U9747 (N_9747,N_9466,N_9520);
or U9748 (N_9748,N_9506,N_9502);
and U9749 (N_9749,N_9588,N_9572);
nor U9750 (N_9750,N_9596,N_9554);
or U9751 (N_9751,N_9495,N_9450);
and U9752 (N_9752,N_9415,N_9595);
nand U9753 (N_9753,N_9403,N_9519);
nor U9754 (N_9754,N_9437,N_9542);
xor U9755 (N_9755,N_9484,N_9582);
or U9756 (N_9756,N_9572,N_9414);
and U9757 (N_9757,N_9452,N_9438);
nor U9758 (N_9758,N_9552,N_9579);
and U9759 (N_9759,N_9588,N_9472);
and U9760 (N_9760,N_9454,N_9584);
nand U9761 (N_9761,N_9465,N_9511);
nand U9762 (N_9762,N_9507,N_9559);
nand U9763 (N_9763,N_9575,N_9423);
and U9764 (N_9764,N_9407,N_9549);
and U9765 (N_9765,N_9580,N_9545);
or U9766 (N_9766,N_9489,N_9466);
and U9767 (N_9767,N_9561,N_9412);
or U9768 (N_9768,N_9491,N_9507);
and U9769 (N_9769,N_9559,N_9479);
xnor U9770 (N_9770,N_9534,N_9515);
and U9771 (N_9771,N_9583,N_9427);
xnor U9772 (N_9772,N_9486,N_9561);
or U9773 (N_9773,N_9574,N_9518);
or U9774 (N_9774,N_9579,N_9438);
nand U9775 (N_9775,N_9545,N_9513);
and U9776 (N_9776,N_9589,N_9449);
or U9777 (N_9777,N_9493,N_9402);
nand U9778 (N_9778,N_9512,N_9428);
xnor U9779 (N_9779,N_9502,N_9581);
nor U9780 (N_9780,N_9479,N_9428);
nor U9781 (N_9781,N_9418,N_9503);
nand U9782 (N_9782,N_9416,N_9566);
nand U9783 (N_9783,N_9450,N_9573);
nand U9784 (N_9784,N_9491,N_9479);
and U9785 (N_9785,N_9430,N_9447);
nand U9786 (N_9786,N_9469,N_9456);
nor U9787 (N_9787,N_9431,N_9518);
and U9788 (N_9788,N_9591,N_9501);
and U9789 (N_9789,N_9591,N_9404);
or U9790 (N_9790,N_9587,N_9413);
xor U9791 (N_9791,N_9554,N_9515);
and U9792 (N_9792,N_9573,N_9474);
and U9793 (N_9793,N_9550,N_9546);
nor U9794 (N_9794,N_9480,N_9585);
or U9795 (N_9795,N_9588,N_9583);
nand U9796 (N_9796,N_9426,N_9501);
nand U9797 (N_9797,N_9544,N_9412);
and U9798 (N_9798,N_9508,N_9440);
xor U9799 (N_9799,N_9588,N_9495);
or U9800 (N_9800,N_9693,N_9710);
nor U9801 (N_9801,N_9662,N_9624);
or U9802 (N_9802,N_9762,N_9752);
nand U9803 (N_9803,N_9640,N_9749);
nor U9804 (N_9804,N_9653,N_9705);
or U9805 (N_9805,N_9697,N_9727);
and U9806 (N_9806,N_9639,N_9698);
or U9807 (N_9807,N_9751,N_9729);
or U9808 (N_9808,N_9670,N_9789);
nor U9809 (N_9809,N_9621,N_9606);
or U9810 (N_9810,N_9676,N_9793);
nor U9811 (N_9811,N_9700,N_9766);
nand U9812 (N_9812,N_9768,N_9753);
nor U9813 (N_9813,N_9742,N_9612);
nand U9814 (N_9814,N_9786,N_9649);
nor U9815 (N_9815,N_9661,N_9652);
or U9816 (N_9816,N_9772,N_9763);
and U9817 (N_9817,N_9758,N_9782);
or U9818 (N_9818,N_9761,N_9701);
nor U9819 (N_9819,N_9778,N_9680);
nand U9820 (N_9820,N_9643,N_9694);
nor U9821 (N_9821,N_9739,N_9745);
nor U9822 (N_9822,N_9605,N_9699);
or U9823 (N_9823,N_9725,N_9607);
xnor U9824 (N_9824,N_9783,N_9666);
nand U9825 (N_9825,N_9792,N_9618);
xnor U9826 (N_9826,N_9733,N_9647);
and U9827 (N_9827,N_9628,N_9634);
nor U9828 (N_9828,N_9728,N_9794);
nor U9829 (N_9829,N_9630,N_9719);
and U9830 (N_9830,N_9717,N_9600);
xnor U9831 (N_9831,N_9735,N_9608);
and U9832 (N_9832,N_9686,N_9620);
nand U9833 (N_9833,N_9642,N_9748);
xor U9834 (N_9834,N_9711,N_9734);
and U9835 (N_9835,N_9707,N_9648);
nand U9836 (N_9836,N_9626,N_9689);
nor U9837 (N_9837,N_9613,N_9685);
nand U9838 (N_9838,N_9740,N_9646);
and U9839 (N_9839,N_9712,N_9784);
or U9840 (N_9840,N_9674,N_9704);
nand U9841 (N_9841,N_9737,N_9682);
nand U9842 (N_9842,N_9775,N_9769);
or U9843 (N_9843,N_9681,N_9691);
or U9844 (N_9844,N_9622,N_9785);
nand U9845 (N_9845,N_9799,N_9790);
and U9846 (N_9846,N_9774,N_9603);
and U9847 (N_9847,N_9629,N_9668);
xor U9848 (N_9848,N_9779,N_9696);
nand U9849 (N_9849,N_9732,N_9747);
and U9850 (N_9850,N_9619,N_9736);
or U9851 (N_9851,N_9754,N_9695);
and U9852 (N_9852,N_9746,N_9636);
and U9853 (N_9853,N_9756,N_9780);
nor U9854 (N_9854,N_9687,N_9675);
nand U9855 (N_9855,N_9669,N_9770);
and U9856 (N_9856,N_9655,N_9767);
nor U9857 (N_9857,N_9708,N_9798);
nor U9858 (N_9858,N_9667,N_9760);
nand U9859 (N_9859,N_9611,N_9617);
nor U9860 (N_9860,N_9721,N_9637);
or U9861 (N_9861,N_9602,N_9664);
nor U9862 (N_9862,N_9632,N_9773);
nand U9863 (N_9863,N_9658,N_9663);
and U9864 (N_9864,N_9609,N_9764);
or U9865 (N_9865,N_9679,N_9788);
nor U9866 (N_9866,N_9627,N_9615);
and U9867 (N_9867,N_9703,N_9677);
or U9868 (N_9868,N_9616,N_9731);
nor U9869 (N_9869,N_9795,N_9610);
nor U9870 (N_9870,N_9777,N_9715);
or U9871 (N_9871,N_9645,N_9771);
and U9872 (N_9872,N_9730,N_9631);
nor U9873 (N_9873,N_9671,N_9623);
xor U9874 (N_9874,N_9713,N_9744);
xnor U9875 (N_9875,N_9601,N_9716);
nor U9876 (N_9876,N_9741,N_9641);
nor U9877 (N_9877,N_9755,N_9723);
and U9878 (N_9878,N_9750,N_9722);
nand U9879 (N_9879,N_9660,N_9656);
and U9880 (N_9880,N_9638,N_9709);
nor U9881 (N_9881,N_9673,N_9659);
nor U9882 (N_9882,N_9692,N_9657);
nor U9883 (N_9883,N_9625,N_9724);
and U9884 (N_9884,N_9720,N_9759);
or U9885 (N_9885,N_9604,N_9787);
nand U9886 (N_9886,N_9757,N_9644);
or U9887 (N_9887,N_9678,N_9738);
or U9888 (N_9888,N_9672,N_9796);
nand U9889 (N_9889,N_9684,N_9683);
or U9890 (N_9890,N_9635,N_9688);
nand U9891 (N_9891,N_9614,N_9650);
or U9892 (N_9892,N_9791,N_9726);
xnor U9893 (N_9893,N_9706,N_9781);
nand U9894 (N_9894,N_9690,N_9633);
or U9895 (N_9895,N_9797,N_9714);
nand U9896 (N_9896,N_9665,N_9702);
nand U9897 (N_9897,N_9654,N_9651);
or U9898 (N_9898,N_9765,N_9743);
xor U9899 (N_9899,N_9776,N_9718);
nor U9900 (N_9900,N_9713,N_9625);
nand U9901 (N_9901,N_9709,N_9722);
xor U9902 (N_9902,N_9767,N_9694);
xor U9903 (N_9903,N_9657,N_9634);
xor U9904 (N_9904,N_9669,N_9615);
xor U9905 (N_9905,N_9781,N_9783);
and U9906 (N_9906,N_9687,N_9780);
xor U9907 (N_9907,N_9709,N_9752);
and U9908 (N_9908,N_9797,N_9618);
and U9909 (N_9909,N_9723,N_9720);
nor U9910 (N_9910,N_9626,N_9658);
and U9911 (N_9911,N_9703,N_9605);
nand U9912 (N_9912,N_9712,N_9610);
and U9913 (N_9913,N_9624,N_9716);
or U9914 (N_9914,N_9791,N_9664);
nand U9915 (N_9915,N_9733,N_9627);
and U9916 (N_9916,N_9768,N_9635);
xor U9917 (N_9917,N_9737,N_9768);
nor U9918 (N_9918,N_9640,N_9718);
xnor U9919 (N_9919,N_9680,N_9751);
nor U9920 (N_9920,N_9735,N_9771);
xor U9921 (N_9921,N_9639,N_9772);
xor U9922 (N_9922,N_9662,N_9646);
or U9923 (N_9923,N_9630,N_9725);
or U9924 (N_9924,N_9764,N_9687);
nand U9925 (N_9925,N_9783,N_9678);
xnor U9926 (N_9926,N_9779,N_9768);
nor U9927 (N_9927,N_9705,N_9606);
xnor U9928 (N_9928,N_9612,N_9670);
and U9929 (N_9929,N_9771,N_9615);
nand U9930 (N_9930,N_9757,N_9722);
xor U9931 (N_9931,N_9755,N_9628);
or U9932 (N_9932,N_9711,N_9775);
and U9933 (N_9933,N_9682,N_9604);
and U9934 (N_9934,N_9658,N_9758);
xnor U9935 (N_9935,N_9768,N_9662);
or U9936 (N_9936,N_9643,N_9756);
nand U9937 (N_9937,N_9798,N_9636);
nand U9938 (N_9938,N_9700,N_9792);
and U9939 (N_9939,N_9773,N_9616);
and U9940 (N_9940,N_9794,N_9617);
nand U9941 (N_9941,N_9659,N_9730);
nor U9942 (N_9942,N_9727,N_9769);
nand U9943 (N_9943,N_9799,N_9644);
and U9944 (N_9944,N_9704,N_9656);
nand U9945 (N_9945,N_9687,N_9643);
and U9946 (N_9946,N_9785,N_9659);
nor U9947 (N_9947,N_9705,N_9721);
and U9948 (N_9948,N_9798,N_9722);
or U9949 (N_9949,N_9789,N_9686);
xnor U9950 (N_9950,N_9729,N_9774);
nor U9951 (N_9951,N_9709,N_9606);
or U9952 (N_9952,N_9724,N_9728);
nor U9953 (N_9953,N_9738,N_9763);
or U9954 (N_9954,N_9677,N_9775);
or U9955 (N_9955,N_9653,N_9601);
nand U9956 (N_9956,N_9701,N_9715);
and U9957 (N_9957,N_9789,N_9600);
nand U9958 (N_9958,N_9617,N_9677);
nand U9959 (N_9959,N_9721,N_9798);
xnor U9960 (N_9960,N_9754,N_9698);
and U9961 (N_9961,N_9711,N_9612);
nor U9962 (N_9962,N_9637,N_9624);
and U9963 (N_9963,N_9618,N_9636);
or U9964 (N_9964,N_9783,N_9650);
and U9965 (N_9965,N_9773,N_9664);
nand U9966 (N_9966,N_9766,N_9672);
nor U9967 (N_9967,N_9703,N_9771);
nor U9968 (N_9968,N_9623,N_9736);
and U9969 (N_9969,N_9780,N_9683);
xor U9970 (N_9970,N_9733,N_9695);
nor U9971 (N_9971,N_9768,N_9690);
xor U9972 (N_9972,N_9778,N_9715);
and U9973 (N_9973,N_9669,N_9625);
or U9974 (N_9974,N_9766,N_9749);
and U9975 (N_9975,N_9613,N_9729);
nand U9976 (N_9976,N_9706,N_9704);
nor U9977 (N_9977,N_9606,N_9631);
or U9978 (N_9978,N_9750,N_9610);
nor U9979 (N_9979,N_9646,N_9737);
nor U9980 (N_9980,N_9708,N_9715);
or U9981 (N_9981,N_9638,N_9769);
xnor U9982 (N_9982,N_9723,N_9668);
nand U9983 (N_9983,N_9792,N_9785);
or U9984 (N_9984,N_9765,N_9612);
or U9985 (N_9985,N_9647,N_9716);
nand U9986 (N_9986,N_9616,N_9719);
nand U9987 (N_9987,N_9719,N_9779);
or U9988 (N_9988,N_9766,N_9684);
nor U9989 (N_9989,N_9775,N_9624);
xnor U9990 (N_9990,N_9648,N_9612);
nand U9991 (N_9991,N_9622,N_9655);
nor U9992 (N_9992,N_9664,N_9772);
nand U9993 (N_9993,N_9720,N_9784);
and U9994 (N_9994,N_9723,N_9776);
nand U9995 (N_9995,N_9714,N_9758);
xnor U9996 (N_9996,N_9796,N_9703);
nor U9997 (N_9997,N_9694,N_9789);
xnor U9998 (N_9998,N_9700,N_9753);
or U9999 (N_9999,N_9769,N_9753);
nand UO_0 (O_0,N_9874,N_9915);
nand UO_1 (O_1,N_9876,N_9818);
or UO_2 (O_2,N_9990,N_9880);
nor UO_3 (O_3,N_9961,N_9815);
and UO_4 (O_4,N_9803,N_9847);
nor UO_5 (O_5,N_9948,N_9875);
nor UO_6 (O_6,N_9844,N_9907);
and UO_7 (O_7,N_9871,N_9826);
nor UO_8 (O_8,N_9920,N_9986);
nor UO_9 (O_9,N_9861,N_9902);
and UO_10 (O_10,N_9996,N_9938);
nor UO_11 (O_11,N_9936,N_9912);
nand UO_12 (O_12,N_9831,N_9893);
nand UO_13 (O_13,N_9879,N_9979);
nor UO_14 (O_14,N_9819,N_9901);
nand UO_15 (O_15,N_9835,N_9957);
or UO_16 (O_16,N_9987,N_9897);
nor UO_17 (O_17,N_9993,N_9995);
nor UO_18 (O_18,N_9949,N_9945);
and UO_19 (O_19,N_9944,N_9852);
and UO_20 (O_20,N_9841,N_9825);
nand UO_21 (O_21,N_9867,N_9959);
nor UO_22 (O_22,N_9952,N_9821);
and UO_23 (O_23,N_9923,N_9994);
or UO_24 (O_24,N_9911,N_9917);
nor UO_25 (O_25,N_9909,N_9805);
nor UO_26 (O_26,N_9962,N_9977);
and UO_27 (O_27,N_9943,N_9982);
or UO_28 (O_28,N_9854,N_9814);
or UO_29 (O_29,N_9946,N_9882);
nand UO_30 (O_30,N_9878,N_9817);
and UO_31 (O_31,N_9981,N_9836);
or UO_32 (O_32,N_9864,N_9964);
and UO_33 (O_33,N_9892,N_9856);
or UO_34 (O_34,N_9937,N_9884);
or UO_35 (O_35,N_9984,N_9886);
or UO_36 (O_36,N_9809,N_9906);
nand UO_37 (O_37,N_9860,N_9839);
nor UO_38 (O_38,N_9992,N_9843);
or UO_39 (O_39,N_9968,N_9833);
or UO_40 (O_40,N_9830,N_9868);
nand UO_41 (O_41,N_9919,N_9850);
nand UO_42 (O_42,N_9940,N_9980);
nor UO_43 (O_43,N_9922,N_9908);
nor UO_44 (O_44,N_9820,N_9804);
or UO_45 (O_45,N_9877,N_9932);
and UO_46 (O_46,N_9991,N_9828);
nor UO_47 (O_47,N_9842,N_9966);
and UO_48 (O_48,N_9972,N_9941);
nor UO_49 (O_49,N_9812,N_9971);
xnor UO_50 (O_50,N_9913,N_9975);
and UO_51 (O_51,N_9898,N_9929);
or UO_52 (O_52,N_9978,N_9899);
nand UO_53 (O_53,N_9811,N_9960);
nor UO_54 (O_54,N_9905,N_9851);
xnor UO_55 (O_55,N_9885,N_9985);
and UO_56 (O_56,N_9837,N_9808);
and UO_57 (O_57,N_9862,N_9806);
xnor UO_58 (O_58,N_9849,N_9965);
nand UO_59 (O_59,N_9933,N_9883);
and UO_60 (O_60,N_9895,N_9935);
nor UO_61 (O_61,N_9910,N_9976);
nor UO_62 (O_62,N_9918,N_9869);
or UO_63 (O_63,N_9950,N_9924);
or UO_64 (O_64,N_9958,N_9865);
nand UO_65 (O_65,N_9840,N_9858);
or UO_66 (O_66,N_9872,N_9953);
xnor UO_67 (O_67,N_9823,N_9816);
or UO_68 (O_68,N_9989,N_9827);
nor UO_69 (O_69,N_9866,N_9925);
nor UO_70 (O_70,N_9926,N_9914);
xnor UO_71 (O_71,N_9999,N_9921);
xnor UO_72 (O_72,N_9870,N_9970);
or UO_73 (O_73,N_9954,N_9846);
and UO_74 (O_74,N_9887,N_9927);
nand UO_75 (O_75,N_9988,N_9942);
or UO_76 (O_76,N_9916,N_9983);
nor UO_77 (O_77,N_9813,N_9807);
nand UO_78 (O_78,N_9881,N_9896);
and UO_79 (O_79,N_9888,N_9963);
and UO_80 (O_80,N_9939,N_9801);
or UO_81 (O_81,N_9969,N_9894);
and UO_82 (O_82,N_9931,N_9873);
nand UO_83 (O_83,N_9810,N_9973);
and UO_84 (O_84,N_9834,N_9967);
xnor UO_85 (O_85,N_9848,N_9890);
and UO_86 (O_86,N_9974,N_9859);
and UO_87 (O_87,N_9930,N_9802);
nor UO_88 (O_88,N_9855,N_9951);
or UO_89 (O_89,N_9934,N_9829);
nor UO_90 (O_90,N_9863,N_9832);
nor UO_91 (O_91,N_9891,N_9903);
and UO_92 (O_92,N_9800,N_9824);
xnor UO_93 (O_93,N_9997,N_9853);
nand UO_94 (O_94,N_9928,N_9998);
nor UO_95 (O_95,N_9955,N_9956);
nand UO_96 (O_96,N_9857,N_9889);
or UO_97 (O_97,N_9900,N_9822);
and UO_98 (O_98,N_9838,N_9845);
or UO_99 (O_99,N_9904,N_9947);
nor UO_100 (O_100,N_9962,N_9825);
or UO_101 (O_101,N_9998,N_9975);
xnor UO_102 (O_102,N_9942,N_9878);
or UO_103 (O_103,N_9961,N_9863);
xor UO_104 (O_104,N_9838,N_9961);
and UO_105 (O_105,N_9958,N_9890);
or UO_106 (O_106,N_9869,N_9954);
or UO_107 (O_107,N_9850,N_9909);
nor UO_108 (O_108,N_9947,N_9867);
and UO_109 (O_109,N_9976,N_9803);
or UO_110 (O_110,N_9968,N_9902);
or UO_111 (O_111,N_9817,N_9944);
nand UO_112 (O_112,N_9843,N_9868);
nor UO_113 (O_113,N_9862,N_9831);
or UO_114 (O_114,N_9869,N_9958);
and UO_115 (O_115,N_9846,N_9822);
xor UO_116 (O_116,N_9900,N_9863);
and UO_117 (O_117,N_9817,N_9845);
or UO_118 (O_118,N_9977,N_9906);
or UO_119 (O_119,N_9809,N_9975);
xnor UO_120 (O_120,N_9835,N_9961);
nor UO_121 (O_121,N_9890,N_9967);
nand UO_122 (O_122,N_9826,N_9944);
or UO_123 (O_123,N_9957,N_9935);
nand UO_124 (O_124,N_9969,N_9974);
nor UO_125 (O_125,N_9817,N_9921);
and UO_126 (O_126,N_9918,N_9902);
or UO_127 (O_127,N_9998,N_9958);
nand UO_128 (O_128,N_9857,N_9933);
nor UO_129 (O_129,N_9928,N_9875);
nor UO_130 (O_130,N_9905,N_9939);
and UO_131 (O_131,N_9943,N_9954);
or UO_132 (O_132,N_9837,N_9893);
nand UO_133 (O_133,N_9943,N_9904);
nor UO_134 (O_134,N_9823,N_9919);
nand UO_135 (O_135,N_9861,N_9918);
or UO_136 (O_136,N_9955,N_9868);
and UO_137 (O_137,N_9902,N_9814);
or UO_138 (O_138,N_9904,N_9863);
nand UO_139 (O_139,N_9852,N_9824);
nor UO_140 (O_140,N_9979,N_9978);
or UO_141 (O_141,N_9814,N_9895);
nor UO_142 (O_142,N_9947,N_9931);
nand UO_143 (O_143,N_9825,N_9826);
or UO_144 (O_144,N_9817,N_9871);
and UO_145 (O_145,N_9922,N_9884);
and UO_146 (O_146,N_9913,N_9813);
or UO_147 (O_147,N_9873,N_9894);
and UO_148 (O_148,N_9937,N_9942);
or UO_149 (O_149,N_9906,N_9919);
and UO_150 (O_150,N_9925,N_9888);
or UO_151 (O_151,N_9843,N_9890);
nand UO_152 (O_152,N_9927,N_9959);
xnor UO_153 (O_153,N_9838,N_9826);
nand UO_154 (O_154,N_9921,N_9986);
nand UO_155 (O_155,N_9959,N_9966);
nand UO_156 (O_156,N_9817,N_9873);
nor UO_157 (O_157,N_9895,N_9916);
or UO_158 (O_158,N_9967,N_9946);
nor UO_159 (O_159,N_9841,N_9911);
or UO_160 (O_160,N_9927,N_9922);
nand UO_161 (O_161,N_9956,N_9873);
and UO_162 (O_162,N_9975,N_9860);
nand UO_163 (O_163,N_9979,N_9918);
nor UO_164 (O_164,N_9965,N_9868);
and UO_165 (O_165,N_9942,N_9998);
nor UO_166 (O_166,N_9904,N_9940);
and UO_167 (O_167,N_9955,N_9996);
nor UO_168 (O_168,N_9889,N_9897);
nor UO_169 (O_169,N_9987,N_9905);
or UO_170 (O_170,N_9948,N_9852);
nor UO_171 (O_171,N_9902,N_9943);
or UO_172 (O_172,N_9801,N_9853);
nor UO_173 (O_173,N_9904,N_9996);
and UO_174 (O_174,N_9819,N_9816);
or UO_175 (O_175,N_9927,N_9807);
nand UO_176 (O_176,N_9850,N_9868);
or UO_177 (O_177,N_9996,N_9945);
nor UO_178 (O_178,N_9801,N_9980);
nand UO_179 (O_179,N_9959,N_9815);
nor UO_180 (O_180,N_9801,N_9876);
nand UO_181 (O_181,N_9980,N_9993);
xor UO_182 (O_182,N_9821,N_9899);
nor UO_183 (O_183,N_9972,N_9985);
nor UO_184 (O_184,N_9885,N_9835);
xor UO_185 (O_185,N_9853,N_9934);
nand UO_186 (O_186,N_9981,N_9833);
nor UO_187 (O_187,N_9992,N_9933);
nor UO_188 (O_188,N_9974,N_9992);
nand UO_189 (O_189,N_9961,N_9867);
nor UO_190 (O_190,N_9970,N_9901);
or UO_191 (O_191,N_9849,N_9981);
or UO_192 (O_192,N_9997,N_9806);
nand UO_193 (O_193,N_9909,N_9904);
nor UO_194 (O_194,N_9913,N_9989);
and UO_195 (O_195,N_9906,N_9816);
nand UO_196 (O_196,N_9947,N_9841);
nand UO_197 (O_197,N_9958,N_9889);
nand UO_198 (O_198,N_9924,N_9912);
nand UO_199 (O_199,N_9965,N_9872);
or UO_200 (O_200,N_9947,N_9982);
and UO_201 (O_201,N_9868,N_9902);
and UO_202 (O_202,N_9953,N_9827);
and UO_203 (O_203,N_9878,N_9956);
nor UO_204 (O_204,N_9884,N_9857);
or UO_205 (O_205,N_9860,N_9897);
nor UO_206 (O_206,N_9936,N_9867);
nor UO_207 (O_207,N_9834,N_9864);
and UO_208 (O_208,N_9804,N_9931);
and UO_209 (O_209,N_9955,N_9899);
or UO_210 (O_210,N_9824,N_9968);
and UO_211 (O_211,N_9890,N_9996);
and UO_212 (O_212,N_9956,N_9830);
nand UO_213 (O_213,N_9945,N_9870);
and UO_214 (O_214,N_9947,N_9977);
or UO_215 (O_215,N_9863,N_9816);
and UO_216 (O_216,N_9938,N_9963);
and UO_217 (O_217,N_9978,N_9859);
xnor UO_218 (O_218,N_9937,N_9910);
xnor UO_219 (O_219,N_9844,N_9815);
nor UO_220 (O_220,N_9899,N_9989);
and UO_221 (O_221,N_9888,N_9833);
and UO_222 (O_222,N_9915,N_9951);
nand UO_223 (O_223,N_9895,N_9820);
nand UO_224 (O_224,N_9915,N_9879);
xor UO_225 (O_225,N_9941,N_9902);
and UO_226 (O_226,N_9898,N_9842);
nand UO_227 (O_227,N_9863,N_9805);
and UO_228 (O_228,N_9853,N_9818);
nand UO_229 (O_229,N_9956,N_9925);
nand UO_230 (O_230,N_9971,N_9912);
nand UO_231 (O_231,N_9813,N_9846);
and UO_232 (O_232,N_9880,N_9970);
nand UO_233 (O_233,N_9806,N_9832);
nor UO_234 (O_234,N_9980,N_9893);
or UO_235 (O_235,N_9812,N_9835);
nor UO_236 (O_236,N_9916,N_9939);
xnor UO_237 (O_237,N_9874,N_9926);
or UO_238 (O_238,N_9976,N_9847);
xor UO_239 (O_239,N_9969,N_9975);
nand UO_240 (O_240,N_9923,N_9818);
and UO_241 (O_241,N_9967,N_9971);
or UO_242 (O_242,N_9963,N_9854);
nand UO_243 (O_243,N_9885,N_9973);
and UO_244 (O_244,N_9989,N_9931);
and UO_245 (O_245,N_9830,N_9879);
nor UO_246 (O_246,N_9832,N_9877);
nand UO_247 (O_247,N_9876,N_9857);
or UO_248 (O_248,N_9930,N_9990);
nor UO_249 (O_249,N_9927,N_9916);
and UO_250 (O_250,N_9921,N_9806);
or UO_251 (O_251,N_9805,N_9905);
or UO_252 (O_252,N_9867,N_9919);
and UO_253 (O_253,N_9985,N_9925);
or UO_254 (O_254,N_9924,N_9831);
nor UO_255 (O_255,N_9960,N_9852);
nor UO_256 (O_256,N_9997,N_9874);
xnor UO_257 (O_257,N_9973,N_9942);
xor UO_258 (O_258,N_9947,N_9923);
or UO_259 (O_259,N_9986,N_9988);
or UO_260 (O_260,N_9995,N_9883);
or UO_261 (O_261,N_9905,N_9902);
or UO_262 (O_262,N_9840,N_9877);
nor UO_263 (O_263,N_9940,N_9876);
and UO_264 (O_264,N_9846,N_9972);
or UO_265 (O_265,N_9835,N_9865);
nand UO_266 (O_266,N_9982,N_9973);
nor UO_267 (O_267,N_9938,N_9847);
nand UO_268 (O_268,N_9970,N_9825);
xnor UO_269 (O_269,N_9839,N_9871);
and UO_270 (O_270,N_9985,N_9829);
or UO_271 (O_271,N_9858,N_9910);
nand UO_272 (O_272,N_9966,N_9894);
nand UO_273 (O_273,N_9909,N_9898);
and UO_274 (O_274,N_9922,N_9917);
or UO_275 (O_275,N_9871,N_9914);
nor UO_276 (O_276,N_9877,N_9962);
nor UO_277 (O_277,N_9806,N_9903);
xor UO_278 (O_278,N_9898,N_9923);
or UO_279 (O_279,N_9843,N_9918);
nand UO_280 (O_280,N_9961,N_9976);
or UO_281 (O_281,N_9990,N_9989);
and UO_282 (O_282,N_9979,N_9810);
or UO_283 (O_283,N_9825,N_9896);
nor UO_284 (O_284,N_9972,N_9967);
or UO_285 (O_285,N_9961,N_9850);
nand UO_286 (O_286,N_9879,N_9948);
xnor UO_287 (O_287,N_9835,N_9813);
nand UO_288 (O_288,N_9995,N_9994);
xnor UO_289 (O_289,N_9870,N_9965);
nor UO_290 (O_290,N_9910,N_9802);
nor UO_291 (O_291,N_9888,N_9815);
and UO_292 (O_292,N_9957,N_9964);
or UO_293 (O_293,N_9927,N_9987);
or UO_294 (O_294,N_9892,N_9912);
nand UO_295 (O_295,N_9987,N_9983);
nand UO_296 (O_296,N_9802,N_9983);
nand UO_297 (O_297,N_9804,N_9935);
nor UO_298 (O_298,N_9935,N_9904);
or UO_299 (O_299,N_9953,N_9821);
nor UO_300 (O_300,N_9881,N_9901);
xnor UO_301 (O_301,N_9831,N_9847);
nand UO_302 (O_302,N_9934,N_9802);
nand UO_303 (O_303,N_9954,N_9808);
and UO_304 (O_304,N_9826,N_9801);
and UO_305 (O_305,N_9948,N_9977);
nor UO_306 (O_306,N_9998,N_9880);
and UO_307 (O_307,N_9886,N_9870);
and UO_308 (O_308,N_9996,N_9829);
nor UO_309 (O_309,N_9951,N_9903);
nand UO_310 (O_310,N_9833,N_9860);
or UO_311 (O_311,N_9976,N_9887);
xor UO_312 (O_312,N_9959,N_9985);
nor UO_313 (O_313,N_9990,N_9857);
nand UO_314 (O_314,N_9927,N_9881);
and UO_315 (O_315,N_9930,N_9879);
nor UO_316 (O_316,N_9992,N_9817);
nor UO_317 (O_317,N_9964,N_9904);
nor UO_318 (O_318,N_9951,N_9822);
and UO_319 (O_319,N_9893,N_9928);
or UO_320 (O_320,N_9978,N_9874);
and UO_321 (O_321,N_9900,N_9824);
or UO_322 (O_322,N_9965,N_9947);
and UO_323 (O_323,N_9802,N_9809);
and UO_324 (O_324,N_9813,N_9817);
nand UO_325 (O_325,N_9964,N_9930);
and UO_326 (O_326,N_9892,N_9957);
or UO_327 (O_327,N_9947,N_9911);
nand UO_328 (O_328,N_9817,N_9838);
or UO_329 (O_329,N_9946,N_9962);
or UO_330 (O_330,N_9833,N_9984);
nor UO_331 (O_331,N_9836,N_9878);
and UO_332 (O_332,N_9924,N_9800);
nor UO_333 (O_333,N_9968,N_9815);
or UO_334 (O_334,N_9948,N_9933);
or UO_335 (O_335,N_9892,N_9886);
or UO_336 (O_336,N_9981,N_9934);
or UO_337 (O_337,N_9864,N_9805);
nor UO_338 (O_338,N_9956,N_9876);
nor UO_339 (O_339,N_9887,N_9944);
nand UO_340 (O_340,N_9980,N_9971);
nor UO_341 (O_341,N_9967,N_9968);
or UO_342 (O_342,N_9934,N_9808);
nor UO_343 (O_343,N_9924,N_9932);
xnor UO_344 (O_344,N_9816,N_9904);
and UO_345 (O_345,N_9860,N_9837);
or UO_346 (O_346,N_9886,N_9926);
xor UO_347 (O_347,N_9940,N_9955);
nor UO_348 (O_348,N_9928,N_9804);
nor UO_349 (O_349,N_9937,N_9993);
and UO_350 (O_350,N_9963,N_9809);
xnor UO_351 (O_351,N_9991,N_9817);
or UO_352 (O_352,N_9980,N_9873);
nor UO_353 (O_353,N_9880,N_9968);
and UO_354 (O_354,N_9853,N_9828);
nand UO_355 (O_355,N_9857,N_9899);
or UO_356 (O_356,N_9962,N_9994);
xor UO_357 (O_357,N_9972,N_9962);
and UO_358 (O_358,N_9867,N_9823);
nor UO_359 (O_359,N_9906,N_9984);
nand UO_360 (O_360,N_9966,N_9898);
and UO_361 (O_361,N_9957,N_9975);
xnor UO_362 (O_362,N_9972,N_9965);
nor UO_363 (O_363,N_9971,N_9817);
nand UO_364 (O_364,N_9987,N_9824);
and UO_365 (O_365,N_9888,N_9947);
or UO_366 (O_366,N_9971,N_9858);
and UO_367 (O_367,N_9979,N_9833);
and UO_368 (O_368,N_9966,N_9963);
and UO_369 (O_369,N_9820,N_9954);
and UO_370 (O_370,N_9939,N_9956);
nand UO_371 (O_371,N_9894,N_9838);
xnor UO_372 (O_372,N_9868,N_9990);
nor UO_373 (O_373,N_9858,N_9917);
or UO_374 (O_374,N_9926,N_9991);
xor UO_375 (O_375,N_9914,N_9835);
or UO_376 (O_376,N_9819,N_9890);
nand UO_377 (O_377,N_9935,N_9848);
and UO_378 (O_378,N_9953,N_9995);
xor UO_379 (O_379,N_9846,N_9939);
and UO_380 (O_380,N_9893,N_9815);
and UO_381 (O_381,N_9981,N_9855);
nand UO_382 (O_382,N_9914,N_9809);
and UO_383 (O_383,N_9925,N_9969);
or UO_384 (O_384,N_9947,N_9817);
and UO_385 (O_385,N_9910,N_9957);
and UO_386 (O_386,N_9814,N_9878);
and UO_387 (O_387,N_9998,N_9837);
or UO_388 (O_388,N_9864,N_9846);
or UO_389 (O_389,N_9936,N_9993);
nand UO_390 (O_390,N_9875,N_9890);
nor UO_391 (O_391,N_9880,N_9947);
and UO_392 (O_392,N_9941,N_9932);
nand UO_393 (O_393,N_9893,N_9902);
and UO_394 (O_394,N_9816,N_9884);
or UO_395 (O_395,N_9820,N_9986);
nand UO_396 (O_396,N_9935,N_9887);
nand UO_397 (O_397,N_9858,N_9832);
xnor UO_398 (O_398,N_9926,N_9960);
and UO_399 (O_399,N_9864,N_9875);
and UO_400 (O_400,N_9833,N_9805);
nand UO_401 (O_401,N_9945,N_9932);
and UO_402 (O_402,N_9895,N_9989);
xnor UO_403 (O_403,N_9801,N_9992);
or UO_404 (O_404,N_9844,N_9855);
nor UO_405 (O_405,N_9855,N_9867);
nand UO_406 (O_406,N_9975,N_9990);
or UO_407 (O_407,N_9836,N_9879);
and UO_408 (O_408,N_9979,N_9968);
nand UO_409 (O_409,N_9890,N_9931);
or UO_410 (O_410,N_9945,N_9834);
or UO_411 (O_411,N_9864,N_9960);
or UO_412 (O_412,N_9948,N_9822);
nand UO_413 (O_413,N_9844,N_9969);
and UO_414 (O_414,N_9906,N_9852);
nand UO_415 (O_415,N_9820,N_9930);
nand UO_416 (O_416,N_9966,N_9968);
and UO_417 (O_417,N_9981,N_9856);
nor UO_418 (O_418,N_9901,N_9979);
and UO_419 (O_419,N_9884,N_9966);
nor UO_420 (O_420,N_9886,N_9913);
and UO_421 (O_421,N_9886,N_9954);
nand UO_422 (O_422,N_9949,N_9929);
and UO_423 (O_423,N_9934,N_9862);
and UO_424 (O_424,N_9991,N_9918);
and UO_425 (O_425,N_9928,N_9865);
nor UO_426 (O_426,N_9964,N_9998);
or UO_427 (O_427,N_9907,N_9816);
nand UO_428 (O_428,N_9994,N_9859);
or UO_429 (O_429,N_9800,N_9813);
nor UO_430 (O_430,N_9824,N_9907);
nand UO_431 (O_431,N_9888,N_9851);
nand UO_432 (O_432,N_9868,N_9862);
and UO_433 (O_433,N_9996,N_9823);
or UO_434 (O_434,N_9842,N_9816);
xor UO_435 (O_435,N_9892,N_9930);
or UO_436 (O_436,N_9945,N_9922);
and UO_437 (O_437,N_9800,N_9951);
or UO_438 (O_438,N_9831,N_9921);
nand UO_439 (O_439,N_9850,N_9862);
nand UO_440 (O_440,N_9891,N_9849);
nand UO_441 (O_441,N_9955,N_9913);
nand UO_442 (O_442,N_9902,N_9904);
or UO_443 (O_443,N_9959,N_9938);
nor UO_444 (O_444,N_9802,N_9940);
xnor UO_445 (O_445,N_9858,N_9887);
and UO_446 (O_446,N_9873,N_9904);
nand UO_447 (O_447,N_9914,N_9843);
and UO_448 (O_448,N_9828,N_9925);
xor UO_449 (O_449,N_9935,N_9997);
and UO_450 (O_450,N_9847,N_9914);
xnor UO_451 (O_451,N_9916,N_9886);
nand UO_452 (O_452,N_9801,N_9989);
or UO_453 (O_453,N_9861,N_9860);
nor UO_454 (O_454,N_9867,N_9897);
xor UO_455 (O_455,N_9887,N_9932);
or UO_456 (O_456,N_9989,N_9921);
and UO_457 (O_457,N_9850,N_9942);
or UO_458 (O_458,N_9806,N_9898);
nand UO_459 (O_459,N_9848,N_9876);
nor UO_460 (O_460,N_9858,N_9853);
nor UO_461 (O_461,N_9886,N_9844);
and UO_462 (O_462,N_9933,N_9817);
nand UO_463 (O_463,N_9850,N_9929);
nor UO_464 (O_464,N_9872,N_9903);
or UO_465 (O_465,N_9909,N_9955);
or UO_466 (O_466,N_9805,N_9894);
and UO_467 (O_467,N_9916,N_9890);
or UO_468 (O_468,N_9901,N_9886);
nand UO_469 (O_469,N_9963,N_9896);
nand UO_470 (O_470,N_9928,N_9800);
xnor UO_471 (O_471,N_9959,N_9844);
nor UO_472 (O_472,N_9821,N_9881);
xor UO_473 (O_473,N_9910,N_9934);
nor UO_474 (O_474,N_9902,N_9907);
or UO_475 (O_475,N_9907,N_9948);
nand UO_476 (O_476,N_9901,N_9909);
and UO_477 (O_477,N_9903,N_9962);
xor UO_478 (O_478,N_9954,N_9902);
nand UO_479 (O_479,N_9942,N_9912);
and UO_480 (O_480,N_9837,N_9807);
nor UO_481 (O_481,N_9985,N_9961);
nand UO_482 (O_482,N_9995,N_9989);
and UO_483 (O_483,N_9881,N_9861);
nand UO_484 (O_484,N_9932,N_9870);
xor UO_485 (O_485,N_9973,N_9922);
xor UO_486 (O_486,N_9810,N_9872);
nand UO_487 (O_487,N_9901,N_9844);
nor UO_488 (O_488,N_9978,N_9883);
nor UO_489 (O_489,N_9977,N_9974);
nand UO_490 (O_490,N_9913,N_9884);
nor UO_491 (O_491,N_9860,N_9997);
nor UO_492 (O_492,N_9905,N_9990);
nor UO_493 (O_493,N_9800,N_9860);
nor UO_494 (O_494,N_9829,N_9915);
or UO_495 (O_495,N_9990,N_9882);
nand UO_496 (O_496,N_9971,N_9859);
nand UO_497 (O_497,N_9981,N_9820);
or UO_498 (O_498,N_9990,N_9831);
and UO_499 (O_499,N_9834,N_9909);
nand UO_500 (O_500,N_9887,N_9946);
nor UO_501 (O_501,N_9903,N_9853);
nand UO_502 (O_502,N_9925,N_9918);
and UO_503 (O_503,N_9920,N_9941);
nor UO_504 (O_504,N_9934,N_9999);
nand UO_505 (O_505,N_9839,N_9857);
nor UO_506 (O_506,N_9888,N_9813);
xnor UO_507 (O_507,N_9930,N_9839);
and UO_508 (O_508,N_9897,N_9970);
nand UO_509 (O_509,N_9854,N_9855);
nand UO_510 (O_510,N_9831,N_9933);
or UO_511 (O_511,N_9812,N_9905);
nor UO_512 (O_512,N_9817,N_9844);
and UO_513 (O_513,N_9881,N_9966);
and UO_514 (O_514,N_9990,N_9826);
xor UO_515 (O_515,N_9927,N_9911);
nor UO_516 (O_516,N_9888,N_9967);
xnor UO_517 (O_517,N_9975,N_9918);
nand UO_518 (O_518,N_9954,N_9810);
or UO_519 (O_519,N_9913,N_9803);
and UO_520 (O_520,N_9969,N_9937);
or UO_521 (O_521,N_9923,N_9874);
nor UO_522 (O_522,N_9896,N_9807);
nand UO_523 (O_523,N_9859,N_9879);
and UO_524 (O_524,N_9835,N_9884);
or UO_525 (O_525,N_9821,N_9927);
and UO_526 (O_526,N_9969,N_9942);
and UO_527 (O_527,N_9846,N_9925);
and UO_528 (O_528,N_9966,N_9804);
or UO_529 (O_529,N_9816,N_9828);
or UO_530 (O_530,N_9996,N_9991);
nand UO_531 (O_531,N_9862,N_9893);
nor UO_532 (O_532,N_9892,N_9822);
and UO_533 (O_533,N_9960,N_9869);
and UO_534 (O_534,N_9890,N_9980);
and UO_535 (O_535,N_9889,N_9821);
nand UO_536 (O_536,N_9894,N_9851);
and UO_537 (O_537,N_9937,N_9863);
or UO_538 (O_538,N_9873,N_9861);
and UO_539 (O_539,N_9818,N_9954);
nor UO_540 (O_540,N_9828,N_9852);
xor UO_541 (O_541,N_9864,N_9858);
or UO_542 (O_542,N_9897,N_9962);
nor UO_543 (O_543,N_9915,N_9891);
xnor UO_544 (O_544,N_9956,N_9944);
xnor UO_545 (O_545,N_9845,N_9810);
xnor UO_546 (O_546,N_9834,N_9896);
and UO_547 (O_547,N_9979,N_9984);
nor UO_548 (O_548,N_9830,N_9957);
or UO_549 (O_549,N_9974,N_9807);
nor UO_550 (O_550,N_9957,N_9951);
nand UO_551 (O_551,N_9830,N_9872);
and UO_552 (O_552,N_9923,N_9936);
nand UO_553 (O_553,N_9811,N_9929);
xnor UO_554 (O_554,N_9931,N_9885);
or UO_555 (O_555,N_9848,N_9844);
nand UO_556 (O_556,N_9974,N_9813);
nand UO_557 (O_557,N_9858,N_9916);
or UO_558 (O_558,N_9815,N_9973);
and UO_559 (O_559,N_9901,N_9866);
nor UO_560 (O_560,N_9872,N_9889);
and UO_561 (O_561,N_9979,N_9845);
nand UO_562 (O_562,N_9961,N_9869);
and UO_563 (O_563,N_9803,N_9960);
nand UO_564 (O_564,N_9996,N_9920);
nand UO_565 (O_565,N_9948,N_9873);
xor UO_566 (O_566,N_9907,N_9959);
nor UO_567 (O_567,N_9922,N_9823);
nor UO_568 (O_568,N_9879,N_9860);
and UO_569 (O_569,N_9958,N_9841);
xor UO_570 (O_570,N_9946,N_9894);
xnor UO_571 (O_571,N_9843,N_9825);
and UO_572 (O_572,N_9903,N_9923);
nor UO_573 (O_573,N_9836,N_9984);
nand UO_574 (O_574,N_9906,N_9976);
and UO_575 (O_575,N_9901,N_9975);
nor UO_576 (O_576,N_9847,N_9885);
nand UO_577 (O_577,N_9823,N_9872);
xnor UO_578 (O_578,N_9852,N_9914);
nand UO_579 (O_579,N_9972,N_9885);
nand UO_580 (O_580,N_9874,N_9907);
xor UO_581 (O_581,N_9816,N_9937);
or UO_582 (O_582,N_9865,N_9859);
or UO_583 (O_583,N_9984,N_9988);
nor UO_584 (O_584,N_9970,N_9999);
nand UO_585 (O_585,N_9958,N_9805);
xor UO_586 (O_586,N_9905,N_9977);
xnor UO_587 (O_587,N_9918,N_9874);
nand UO_588 (O_588,N_9876,N_9855);
xnor UO_589 (O_589,N_9929,N_9862);
or UO_590 (O_590,N_9872,N_9803);
and UO_591 (O_591,N_9870,N_9930);
or UO_592 (O_592,N_9896,N_9942);
or UO_593 (O_593,N_9820,N_9891);
nand UO_594 (O_594,N_9885,N_9944);
nor UO_595 (O_595,N_9838,N_9850);
nor UO_596 (O_596,N_9800,N_9980);
and UO_597 (O_597,N_9994,N_9903);
or UO_598 (O_598,N_9969,N_9808);
nand UO_599 (O_599,N_9910,N_9966);
nand UO_600 (O_600,N_9951,N_9900);
nor UO_601 (O_601,N_9883,N_9854);
nor UO_602 (O_602,N_9827,N_9981);
nand UO_603 (O_603,N_9943,N_9905);
and UO_604 (O_604,N_9863,N_9844);
xor UO_605 (O_605,N_9871,N_9906);
nor UO_606 (O_606,N_9909,N_9883);
nand UO_607 (O_607,N_9997,N_9988);
and UO_608 (O_608,N_9935,N_9909);
nand UO_609 (O_609,N_9934,N_9883);
nor UO_610 (O_610,N_9937,N_9953);
or UO_611 (O_611,N_9880,N_9978);
nor UO_612 (O_612,N_9990,N_9948);
and UO_613 (O_613,N_9818,N_9979);
nand UO_614 (O_614,N_9997,N_9810);
nor UO_615 (O_615,N_9875,N_9871);
nor UO_616 (O_616,N_9863,N_9975);
or UO_617 (O_617,N_9928,N_9902);
xor UO_618 (O_618,N_9930,N_9987);
nor UO_619 (O_619,N_9826,N_9897);
and UO_620 (O_620,N_9934,N_9837);
and UO_621 (O_621,N_9874,N_9848);
or UO_622 (O_622,N_9836,N_9828);
nand UO_623 (O_623,N_9855,N_9933);
or UO_624 (O_624,N_9923,N_9931);
and UO_625 (O_625,N_9824,N_9940);
and UO_626 (O_626,N_9938,N_9880);
and UO_627 (O_627,N_9813,N_9801);
xor UO_628 (O_628,N_9973,N_9937);
nor UO_629 (O_629,N_9998,N_9907);
nor UO_630 (O_630,N_9955,N_9840);
nor UO_631 (O_631,N_9979,N_9950);
nor UO_632 (O_632,N_9876,N_9917);
or UO_633 (O_633,N_9805,N_9945);
nand UO_634 (O_634,N_9916,N_9962);
nor UO_635 (O_635,N_9864,N_9990);
or UO_636 (O_636,N_9925,N_9980);
and UO_637 (O_637,N_9911,N_9816);
nor UO_638 (O_638,N_9964,N_9809);
or UO_639 (O_639,N_9983,N_9970);
nand UO_640 (O_640,N_9817,N_9862);
and UO_641 (O_641,N_9929,N_9928);
nor UO_642 (O_642,N_9961,N_9974);
nand UO_643 (O_643,N_9999,N_9889);
and UO_644 (O_644,N_9823,N_9977);
nor UO_645 (O_645,N_9877,N_9917);
nand UO_646 (O_646,N_9800,N_9945);
or UO_647 (O_647,N_9941,N_9966);
xor UO_648 (O_648,N_9823,N_9881);
and UO_649 (O_649,N_9991,N_9938);
nor UO_650 (O_650,N_9889,N_9855);
nor UO_651 (O_651,N_9924,N_9895);
or UO_652 (O_652,N_9843,N_9907);
nand UO_653 (O_653,N_9923,N_9840);
or UO_654 (O_654,N_9951,N_9879);
or UO_655 (O_655,N_9866,N_9826);
or UO_656 (O_656,N_9825,N_9862);
nor UO_657 (O_657,N_9805,N_9984);
and UO_658 (O_658,N_9969,N_9837);
and UO_659 (O_659,N_9880,N_9999);
nand UO_660 (O_660,N_9963,N_9801);
nand UO_661 (O_661,N_9967,N_9978);
nor UO_662 (O_662,N_9836,N_9933);
and UO_663 (O_663,N_9990,N_9870);
nand UO_664 (O_664,N_9814,N_9990);
nor UO_665 (O_665,N_9999,N_9954);
and UO_666 (O_666,N_9904,N_9896);
nor UO_667 (O_667,N_9858,N_9865);
and UO_668 (O_668,N_9914,N_9902);
nor UO_669 (O_669,N_9994,N_9884);
nand UO_670 (O_670,N_9899,N_9967);
nor UO_671 (O_671,N_9882,N_9954);
nand UO_672 (O_672,N_9990,N_9961);
or UO_673 (O_673,N_9816,N_9939);
nand UO_674 (O_674,N_9821,N_9824);
xor UO_675 (O_675,N_9908,N_9900);
nand UO_676 (O_676,N_9949,N_9850);
xor UO_677 (O_677,N_9833,N_9842);
nand UO_678 (O_678,N_9811,N_9974);
nor UO_679 (O_679,N_9860,N_9976);
nand UO_680 (O_680,N_9994,N_9861);
nor UO_681 (O_681,N_9910,N_9983);
and UO_682 (O_682,N_9927,N_9931);
and UO_683 (O_683,N_9969,N_9949);
xnor UO_684 (O_684,N_9867,N_9875);
xnor UO_685 (O_685,N_9889,N_9925);
or UO_686 (O_686,N_9875,N_9981);
or UO_687 (O_687,N_9957,N_9885);
nor UO_688 (O_688,N_9842,N_9856);
and UO_689 (O_689,N_9900,N_9980);
or UO_690 (O_690,N_9893,N_9989);
nor UO_691 (O_691,N_9943,N_9822);
nor UO_692 (O_692,N_9971,N_9876);
xor UO_693 (O_693,N_9949,N_9907);
nand UO_694 (O_694,N_9880,N_9922);
xor UO_695 (O_695,N_9882,N_9955);
or UO_696 (O_696,N_9916,N_9848);
nand UO_697 (O_697,N_9811,N_9864);
xnor UO_698 (O_698,N_9983,N_9833);
nor UO_699 (O_699,N_9887,N_9938);
nor UO_700 (O_700,N_9988,N_9893);
nand UO_701 (O_701,N_9831,N_9926);
nor UO_702 (O_702,N_9822,N_9886);
nand UO_703 (O_703,N_9981,N_9889);
and UO_704 (O_704,N_9941,N_9866);
nor UO_705 (O_705,N_9846,N_9868);
nor UO_706 (O_706,N_9927,N_9850);
nor UO_707 (O_707,N_9905,N_9901);
nand UO_708 (O_708,N_9887,N_9952);
nor UO_709 (O_709,N_9886,N_9934);
nand UO_710 (O_710,N_9898,N_9921);
xnor UO_711 (O_711,N_9901,N_9832);
nor UO_712 (O_712,N_9838,N_9877);
or UO_713 (O_713,N_9819,N_9804);
nor UO_714 (O_714,N_9815,N_9824);
or UO_715 (O_715,N_9934,N_9994);
and UO_716 (O_716,N_9926,N_9978);
or UO_717 (O_717,N_9985,N_9853);
nand UO_718 (O_718,N_9989,N_9979);
or UO_719 (O_719,N_9956,N_9866);
nor UO_720 (O_720,N_9932,N_9834);
nor UO_721 (O_721,N_9887,N_9820);
nand UO_722 (O_722,N_9869,N_9985);
or UO_723 (O_723,N_9996,N_9867);
nand UO_724 (O_724,N_9811,N_9927);
and UO_725 (O_725,N_9978,N_9817);
nand UO_726 (O_726,N_9821,N_9811);
or UO_727 (O_727,N_9806,N_9955);
and UO_728 (O_728,N_9822,N_9974);
xor UO_729 (O_729,N_9894,N_9932);
nand UO_730 (O_730,N_9893,N_9941);
xnor UO_731 (O_731,N_9894,N_9807);
and UO_732 (O_732,N_9926,N_9948);
or UO_733 (O_733,N_9928,N_9900);
nand UO_734 (O_734,N_9919,N_9880);
nand UO_735 (O_735,N_9812,N_9947);
nor UO_736 (O_736,N_9936,N_9966);
xor UO_737 (O_737,N_9999,N_9815);
and UO_738 (O_738,N_9979,N_9816);
nor UO_739 (O_739,N_9921,N_9903);
and UO_740 (O_740,N_9904,N_9923);
nand UO_741 (O_741,N_9824,N_9823);
or UO_742 (O_742,N_9913,N_9912);
and UO_743 (O_743,N_9989,N_9912);
or UO_744 (O_744,N_9902,N_9837);
or UO_745 (O_745,N_9830,N_9832);
nor UO_746 (O_746,N_9912,N_9809);
nand UO_747 (O_747,N_9932,N_9835);
or UO_748 (O_748,N_9840,N_9804);
nand UO_749 (O_749,N_9940,N_9805);
xnor UO_750 (O_750,N_9890,N_9801);
nor UO_751 (O_751,N_9818,N_9889);
nor UO_752 (O_752,N_9848,N_9954);
nor UO_753 (O_753,N_9857,N_9914);
or UO_754 (O_754,N_9898,N_9908);
and UO_755 (O_755,N_9965,N_9967);
nor UO_756 (O_756,N_9836,N_9945);
and UO_757 (O_757,N_9899,N_9942);
and UO_758 (O_758,N_9913,N_9974);
nor UO_759 (O_759,N_9975,N_9965);
nand UO_760 (O_760,N_9836,N_9963);
xnor UO_761 (O_761,N_9965,N_9841);
or UO_762 (O_762,N_9892,N_9853);
or UO_763 (O_763,N_9982,N_9800);
xnor UO_764 (O_764,N_9945,N_9958);
or UO_765 (O_765,N_9870,N_9810);
and UO_766 (O_766,N_9870,N_9872);
and UO_767 (O_767,N_9970,N_9888);
or UO_768 (O_768,N_9807,N_9956);
xnor UO_769 (O_769,N_9995,N_9973);
or UO_770 (O_770,N_9972,N_9988);
nor UO_771 (O_771,N_9890,N_9891);
or UO_772 (O_772,N_9958,N_9850);
nor UO_773 (O_773,N_9953,N_9992);
nand UO_774 (O_774,N_9926,N_9845);
or UO_775 (O_775,N_9918,N_9987);
nand UO_776 (O_776,N_9899,N_9869);
nand UO_777 (O_777,N_9817,N_9814);
nand UO_778 (O_778,N_9812,N_9856);
nand UO_779 (O_779,N_9963,N_9993);
or UO_780 (O_780,N_9919,N_9970);
nand UO_781 (O_781,N_9979,N_9885);
nor UO_782 (O_782,N_9855,N_9905);
nor UO_783 (O_783,N_9907,N_9880);
nand UO_784 (O_784,N_9972,N_9815);
and UO_785 (O_785,N_9923,N_9962);
nand UO_786 (O_786,N_9873,N_9820);
and UO_787 (O_787,N_9904,N_9832);
and UO_788 (O_788,N_9998,N_9875);
or UO_789 (O_789,N_9864,N_9900);
and UO_790 (O_790,N_9851,N_9992);
and UO_791 (O_791,N_9880,N_9963);
and UO_792 (O_792,N_9801,N_9996);
or UO_793 (O_793,N_9943,N_9963);
nand UO_794 (O_794,N_9863,N_9856);
xor UO_795 (O_795,N_9829,N_9943);
and UO_796 (O_796,N_9839,N_9965);
nor UO_797 (O_797,N_9920,N_9952);
or UO_798 (O_798,N_9878,N_9863);
and UO_799 (O_799,N_9842,N_9802);
and UO_800 (O_800,N_9849,N_9908);
or UO_801 (O_801,N_9938,N_9932);
and UO_802 (O_802,N_9991,N_9874);
and UO_803 (O_803,N_9967,N_9920);
and UO_804 (O_804,N_9891,N_9897);
nand UO_805 (O_805,N_9950,N_9833);
or UO_806 (O_806,N_9821,N_9841);
and UO_807 (O_807,N_9877,N_9923);
nor UO_808 (O_808,N_9905,N_9864);
nor UO_809 (O_809,N_9945,N_9936);
nand UO_810 (O_810,N_9915,N_9909);
nor UO_811 (O_811,N_9818,N_9830);
or UO_812 (O_812,N_9857,N_9929);
or UO_813 (O_813,N_9841,N_9916);
nor UO_814 (O_814,N_9951,N_9913);
and UO_815 (O_815,N_9926,N_9945);
nor UO_816 (O_816,N_9920,N_9969);
nand UO_817 (O_817,N_9805,N_9950);
nor UO_818 (O_818,N_9932,N_9975);
xnor UO_819 (O_819,N_9973,N_9821);
nor UO_820 (O_820,N_9866,N_9840);
and UO_821 (O_821,N_9805,N_9936);
and UO_822 (O_822,N_9905,N_9868);
and UO_823 (O_823,N_9851,N_9876);
nand UO_824 (O_824,N_9959,N_9944);
nand UO_825 (O_825,N_9881,N_9806);
and UO_826 (O_826,N_9994,N_9897);
nor UO_827 (O_827,N_9855,N_9924);
nor UO_828 (O_828,N_9911,N_9915);
and UO_829 (O_829,N_9819,N_9861);
nor UO_830 (O_830,N_9896,N_9976);
or UO_831 (O_831,N_9919,N_9806);
nor UO_832 (O_832,N_9999,N_9997);
nand UO_833 (O_833,N_9831,N_9876);
xnor UO_834 (O_834,N_9818,N_9915);
and UO_835 (O_835,N_9858,N_9878);
and UO_836 (O_836,N_9847,N_9806);
or UO_837 (O_837,N_9829,N_9983);
or UO_838 (O_838,N_9999,N_9976);
nor UO_839 (O_839,N_9852,N_9836);
nand UO_840 (O_840,N_9891,N_9951);
and UO_841 (O_841,N_9820,N_9939);
and UO_842 (O_842,N_9973,N_9850);
or UO_843 (O_843,N_9804,N_9894);
nand UO_844 (O_844,N_9823,N_9842);
nor UO_845 (O_845,N_9834,N_9981);
nand UO_846 (O_846,N_9857,N_9831);
xnor UO_847 (O_847,N_9830,N_9933);
or UO_848 (O_848,N_9858,N_9960);
and UO_849 (O_849,N_9885,N_9888);
nand UO_850 (O_850,N_9849,N_9860);
and UO_851 (O_851,N_9973,N_9928);
nand UO_852 (O_852,N_9874,N_9958);
nor UO_853 (O_853,N_9965,N_9999);
nor UO_854 (O_854,N_9887,N_9980);
and UO_855 (O_855,N_9818,N_9994);
nor UO_856 (O_856,N_9825,N_9972);
nor UO_857 (O_857,N_9983,N_9869);
and UO_858 (O_858,N_9864,N_9817);
or UO_859 (O_859,N_9936,N_9989);
or UO_860 (O_860,N_9899,N_9964);
nor UO_861 (O_861,N_9868,N_9816);
or UO_862 (O_862,N_9964,N_9917);
nand UO_863 (O_863,N_9977,N_9967);
nor UO_864 (O_864,N_9952,N_9884);
nor UO_865 (O_865,N_9820,N_9867);
and UO_866 (O_866,N_9949,N_9966);
or UO_867 (O_867,N_9914,N_9813);
or UO_868 (O_868,N_9908,N_9817);
nand UO_869 (O_869,N_9868,N_9827);
and UO_870 (O_870,N_9878,N_9825);
nor UO_871 (O_871,N_9844,N_9832);
and UO_872 (O_872,N_9923,N_9885);
and UO_873 (O_873,N_9985,N_9997);
xor UO_874 (O_874,N_9811,N_9862);
nand UO_875 (O_875,N_9829,N_9825);
and UO_876 (O_876,N_9941,N_9910);
or UO_877 (O_877,N_9929,N_9986);
or UO_878 (O_878,N_9954,N_9807);
xnor UO_879 (O_879,N_9807,N_9988);
nor UO_880 (O_880,N_9983,N_9972);
or UO_881 (O_881,N_9871,N_9935);
xnor UO_882 (O_882,N_9971,N_9875);
and UO_883 (O_883,N_9913,N_9869);
nor UO_884 (O_884,N_9961,N_9829);
nor UO_885 (O_885,N_9914,N_9916);
or UO_886 (O_886,N_9921,N_9865);
and UO_887 (O_887,N_9958,N_9856);
and UO_888 (O_888,N_9983,N_9858);
or UO_889 (O_889,N_9965,N_9888);
nor UO_890 (O_890,N_9862,N_9939);
xnor UO_891 (O_891,N_9855,N_9977);
nand UO_892 (O_892,N_9886,N_9904);
nor UO_893 (O_893,N_9861,N_9893);
xor UO_894 (O_894,N_9884,N_9920);
xor UO_895 (O_895,N_9816,N_9876);
or UO_896 (O_896,N_9935,N_9817);
nand UO_897 (O_897,N_9886,N_9977);
nor UO_898 (O_898,N_9858,N_9919);
nand UO_899 (O_899,N_9904,N_9838);
or UO_900 (O_900,N_9865,N_9984);
nand UO_901 (O_901,N_9890,N_9968);
or UO_902 (O_902,N_9844,N_9813);
and UO_903 (O_903,N_9951,N_9922);
or UO_904 (O_904,N_9810,N_9912);
and UO_905 (O_905,N_9987,N_9945);
or UO_906 (O_906,N_9961,N_9995);
nor UO_907 (O_907,N_9807,N_9976);
nand UO_908 (O_908,N_9971,N_9874);
and UO_909 (O_909,N_9944,N_9968);
or UO_910 (O_910,N_9996,N_9903);
or UO_911 (O_911,N_9985,N_9895);
xnor UO_912 (O_912,N_9971,N_9897);
nor UO_913 (O_913,N_9822,N_9859);
nor UO_914 (O_914,N_9866,N_9991);
or UO_915 (O_915,N_9994,N_9991);
nand UO_916 (O_916,N_9960,N_9994);
and UO_917 (O_917,N_9975,N_9862);
nand UO_918 (O_918,N_9880,N_9835);
nand UO_919 (O_919,N_9869,N_9933);
xnor UO_920 (O_920,N_9836,N_9943);
nor UO_921 (O_921,N_9839,N_9870);
and UO_922 (O_922,N_9975,N_9943);
or UO_923 (O_923,N_9837,N_9924);
nor UO_924 (O_924,N_9839,N_9836);
xor UO_925 (O_925,N_9825,N_9943);
or UO_926 (O_926,N_9835,N_9883);
nand UO_927 (O_927,N_9899,N_9856);
nand UO_928 (O_928,N_9849,N_9862);
nand UO_929 (O_929,N_9885,N_9816);
nand UO_930 (O_930,N_9848,N_9882);
nor UO_931 (O_931,N_9912,N_9991);
and UO_932 (O_932,N_9990,N_9867);
nand UO_933 (O_933,N_9856,N_9879);
nand UO_934 (O_934,N_9846,N_9950);
or UO_935 (O_935,N_9883,N_9829);
and UO_936 (O_936,N_9880,N_9845);
nor UO_937 (O_937,N_9820,N_9935);
nor UO_938 (O_938,N_9986,N_9815);
nor UO_939 (O_939,N_9909,N_9872);
xnor UO_940 (O_940,N_9812,N_9868);
and UO_941 (O_941,N_9989,N_9980);
nor UO_942 (O_942,N_9971,N_9915);
and UO_943 (O_943,N_9896,N_9880);
nand UO_944 (O_944,N_9869,N_9808);
nand UO_945 (O_945,N_9901,N_9860);
and UO_946 (O_946,N_9853,N_9907);
and UO_947 (O_947,N_9843,N_9808);
or UO_948 (O_948,N_9913,N_9937);
xnor UO_949 (O_949,N_9920,N_9874);
nand UO_950 (O_950,N_9887,N_9918);
nor UO_951 (O_951,N_9836,N_9809);
or UO_952 (O_952,N_9984,N_9954);
nand UO_953 (O_953,N_9927,N_9993);
nand UO_954 (O_954,N_9890,N_9807);
xor UO_955 (O_955,N_9976,N_9948);
and UO_956 (O_956,N_9835,N_9917);
nor UO_957 (O_957,N_9923,N_9895);
xnor UO_958 (O_958,N_9918,N_9894);
or UO_959 (O_959,N_9993,N_9952);
and UO_960 (O_960,N_9949,N_9845);
and UO_961 (O_961,N_9818,N_9891);
nand UO_962 (O_962,N_9910,N_9872);
xnor UO_963 (O_963,N_9963,N_9870);
xor UO_964 (O_964,N_9918,N_9944);
nor UO_965 (O_965,N_9823,N_9968);
xor UO_966 (O_966,N_9999,N_9953);
xor UO_967 (O_967,N_9844,N_9870);
or UO_968 (O_968,N_9997,N_9990);
and UO_969 (O_969,N_9917,N_9973);
xor UO_970 (O_970,N_9995,N_9934);
or UO_971 (O_971,N_9834,N_9808);
nor UO_972 (O_972,N_9820,N_9963);
nor UO_973 (O_973,N_9814,N_9816);
nand UO_974 (O_974,N_9937,N_9895);
or UO_975 (O_975,N_9832,N_9958);
nor UO_976 (O_976,N_9952,N_9880);
or UO_977 (O_977,N_9972,N_9808);
nor UO_978 (O_978,N_9963,N_9996);
and UO_979 (O_979,N_9831,N_9845);
nor UO_980 (O_980,N_9901,N_9840);
or UO_981 (O_981,N_9889,N_9913);
nor UO_982 (O_982,N_9914,N_9920);
nand UO_983 (O_983,N_9901,N_9891);
and UO_984 (O_984,N_9923,N_9920);
nor UO_985 (O_985,N_9971,N_9800);
nor UO_986 (O_986,N_9821,N_9946);
or UO_987 (O_987,N_9999,N_9902);
nor UO_988 (O_988,N_9934,N_9848);
nor UO_989 (O_989,N_9923,N_9856);
or UO_990 (O_990,N_9972,N_9854);
nor UO_991 (O_991,N_9856,N_9936);
or UO_992 (O_992,N_9902,N_9911);
nand UO_993 (O_993,N_9862,N_9845);
and UO_994 (O_994,N_9811,N_9893);
xnor UO_995 (O_995,N_9882,N_9956);
nor UO_996 (O_996,N_9876,N_9819);
or UO_997 (O_997,N_9885,N_9801);
xnor UO_998 (O_998,N_9848,N_9817);
and UO_999 (O_999,N_9929,N_9924);
and UO_1000 (O_1000,N_9992,N_9981);
nand UO_1001 (O_1001,N_9967,N_9990);
or UO_1002 (O_1002,N_9954,N_9936);
xnor UO_1003 (O_1003,N_9878,N_9998);
and UO_1004 (O_1004,N_9898,N_9991);
or UO_1005 (O_1005,N_9890,N_9838);
nand UO_1006 (O_1006,N_9933,N_9971);
nand UO_1007 (O_1007,N_9932,N_9937);
and UO_1008 (O_1008,N_9854,N_9853);
nor UO_1009 (O_1009,N_9956,N_9845);
nand UO_1010 (O_1010,N_9806,N_9975);
nand UO_1011 (O_1011,N_9927,N_9978);
nand UO_1012 (O_1012,N_9901,N_9816);
nand UO_1013 (O_1013,N_9925,N_9872);
nand UO_1014 (O_1014,N_9853,N_9918);
nand UO_1015 (O_1015,N_9857,N_9826);
nor UO_1016 (O_1016,N_9893,N_9982);
nand UO_1017 (O_1017,N_9808,N_9984);
nand UO_1018 (O_1018,N_9874,N_9994);
or UO_1019 (O_1019,N_9923,N_9841);
nor UO_1020 (O_1020,N_9987,N_9982);
or UO_1021 (O_1021,N_9882,N_9864);
xnor UO_1022 (O_1022,N_9818,N_9981);
and UO_1023 (O_1023,N_9888,N_9889);
xor UO_1024 (O_1024,N_9853,N_9931);
nand UO_1025 (O_1025,N_9970,N_9850);
nor UO_1026 (O_1026,N_9927,N_9964);
and UO_1027 (O_1027,N_9900,N_9929);
nor UO_1028 (O_1028,N_9919,N_9924);
or UO_1029 (O_1029,N_9992,N_9852);
xnor UO_1030 (O_1030,N_9829,N_9843);
nor UO_1031 (O_1031,N_9890,N_9803);
or UO_1032 (O_1032,N_9899,N_9969);
and UO_1033 (O_1033,N_9871,N_9829);
nor UO_1034 (O_1034,N_9991,N_9863);
or UO_1035 (O_1035,N_9997,N_9930);
and UO_1036 (O_1036,N_9836,N_9803);
and UO_1037 (O_1037,N_9815,N_9976);
and UO_1038 (O_1038,N_9927,N_9970);
xnor UO_1039 (O_1039,N_9822,N_9915);
nand UO_1040 (O_1040,N_9918,N_9886);
and UO_1041 (O_1041,N_9940,N_9898);
xnor UO_1042 (O_1042,N_9994,N_9831);
and UO_1043 (O_1043,N_9900,N_9916);
nor UO_1044 (O_1044,N_9904,N_9864);
or UO_1045 (O_1045,N_9999,N_9837);
nor UO_1046 (O_1046,N_9920,N_9895);
nor UO_1047 (O_1047,N_9934,N_9979);
xor UO_1048 (O_1048,N_9832,N_9995);
nor UO_1049 (O_1049,N_9878,N_9895);
nand UO_1050 (O_1050,N_9972,N_9817);
xnor UO_1051 (O_1051,N_9833,N_9955);
and UO_1052 (O_1052,N_9962,N_9812);
nand UO_1053 (O_1053,N_9825,N_9828);
nand UO_1054 (O_1054,N_9835,N_9993);
nor UO_1055 (O_1055,N_9905,N_9978);
xor UO_1056 (O_1056,N_9812,N_9800);
nor UO_1057 (O_1057,N_9850,N_9926);
xnor UO_1058 (O_1058,N_9999,N_9928);
xnor UO_1059 (O_1059,N_9861,N_9899);
nor UO_1060 (O_1060,N_9831,N_9860);
nand UO_1061 (O_1061,N_9911,N_9808);
nand UO_1062 (O_1062,N_9968,N_9915);
or UO_1063 (O_1063,N_9930,N_9937);
and UO_1064 (O_1064,N_9891,N_9888);
and UO_1065 (O_1065,N_9931,N_9955);
xnor UO_1066 (O_1066,N_9910,N_9927);
and UO_1067 (O_1067,N_9939,N_9967);
nor UO_1068 (O_1068,N_9934,N_9949);
nor UO_1069 (O_1069,N_9894,N_9859);
and UO_1070 (O_1070,N_9879,N_9853);
xnor UO_1071 (O_1071,N_9853,N_9947);
nor UO_1072 (O_1072,N_9830,N_9952);
and UO_1073 (O_1073,N_9908,N_9914);
and UO_1074 (O_1074,N_9997,N_9944);
and UO_1075 (O_1075,N_9823,N_9869);
or UO_1076 (O_1076,N_9929,N_9913);
nor UO_1077 (O_1077,N_9825,N_9954);
nand UO_1078 (O_1078,N_9932,N_9991);
and UO_1079 (O_1079,N_9811,N_9851);
and UO_1080 (O_1080,N_9804,N_9876);
or UO_1081 (O_1081,N_9862,N_9801);
nor UO_1082 (O_1082,N_9969,N_9849);
nand UO_1083 (O_1083,N_9928,N_9831);
and UO_1084 (O_1084,N_9941,N_9812);
nor UO_1085 (O_1085,N_9929,N_9882);
and UO_1086 (O_1086,N_9805,N_9980);
nor UO_1087 (O_1087,N_9919,N_9876);
nand UO_1088 (O_1088,N_9826,N_9867);
nand UO_1089 (O_1089,N_9977,N_9876);
or UO_1090 (O_1090,N_9847,N_9878);
or UO_1091 (O_1091,N_9831,N_9841);
xor UO_1092 (O_1092,N_9830,N_9986);
and UO_1093 (O_1093,N_9939,N_9853);
nor UO_1094 (O_1094,N_9868,N_9858);
and UO_1095 (O_1095,N_9949,N_9910);
nor UO_1096 (O_1096,N_9866,N_9912);
and UO_1097 (O_1097,N_9887,N_9973);
nand UO_1098 (O_1098,N_9985,N_9946);
and UO_1099 (O_1099,N_9800,N_9919);
or UO_1100 (O_1100,N_9946,N_9993);
or UO_1101 (O_1101,N_9956,N_9843);
or UO_1102 (O_1102,N_9930,N_9844);
nand UO_1103 (O_1103,N_9840,N_9928);
nor UO_1104 (O_1104,N_9853,N_9927);
xor UO_1105 (O_1105,N_9912,N_9825);
and UO_1106 (O_1106,N_9816,N_9827);
and UO_1107 (O_1107,N_9995,N_9947);
and UO_1108 (O_1108,N_9990,N_9885);
nand UO_1109 (O_1109,N_9916,N_9845);
and UO_1110 (O_1110,N_9992,N_9990);
or UO_1111 (O_1111,N_9882,N_9898);
nand UO_1112 (O_1112,N_9919,N_9957);
or UO_1113 (O_1113,N_9925,N_9818);
and UO_1114 (O_1114,N_9983,N_9868);
and UO_1115 (O_1115,N_9936,N_9888);
nor UO_1116 (O_1116,N_9841,N_9979);
or UO_1117 (O_1117,N_9842,N_9934);
or UO_1118 (O_1118,N_9929,N_9890);
or UO_1119 (O_1119,N_9820,N_9910);
and UO_1120 (O_1120,N_9902,N_9986);
or UO_1121 (O_1121,N_9898,N_9975);
nor UO_1122 (O_1122,N_9893,N_9839);
nand UO_1123 (O_1123,N_9818,N_9921);
and UO_1124 (O_1124,N_9999,N_9980);
nand UO_1125 (O_1125,N_9890,N_9938);
nor UO_1126 (O_1126,N_9910,N_9929);
nor UO_1127 (O_1127,N_9983,N_9899);
and UO_1128 (O_1128,N_9859,N_9979);
or UO_1129 (O_1129,N_9800,N_9911);
nand UO_1130 (O_1130,N_9815,N_9998);
xnor UO_1131 (O_1131,N_9837,N_9967);
and UO_1132 (O_1132,N_9846,N_9924);
nor UO_1133 (O_1133,N_9831,N_9888);
xnor UO_1134 (O_1134,N_9866,N_9952);
xnor UO_1135 (O_1135,N_9926,N_9985);
and UO_1136 (O_1136,N_9925,N_9995);
nor UO_1137 (O_1137,N_9969,N_9930);
nand UO_1138 (O_1138,N_9895,N_9973);
nor UO_1139 (O_1139,N_9844,N_9846);
nor UO_1140 (O_1140,N_9813,N_9902);
nor UO_1141 (O_1141,N_9845,N_9854);
or UO_1142 (O_1142,N_9981,N_9869);
nor UO_1143 (O_1143,N_9916,N_9987);
nor UO_1144 (O_1144,N_9939,N_9983);
xor UO_1145 (O_1145,N_9938,N_9838);
or UO_1146 (O_1146,N_9899,N_9879);
nand UO_1147 (O_1147,N_9881,N_9851);
and UO_1148 (O_1148,N_9902,N_9971);
xor UO_1149 (O_1149,N_9896,N_9911);
and UO_1150 (O_1150,N_9960,N_9948);
and UO_1151 (O_1151,N_9827,N_9845);
nand UO_1152 (O_1152,N_9971,N_9842);
and UO_1153 (O_1153,N_9956,N_9985);
nor UO_1154 (O_1154,N_9924,N_9984);
nand UO_1155 (O_1155,N_9837,N_9813);
nor UO_1156 (O_1156,N_9930,N_9983);
nand UO_1157 (O_1157,N_9822,N_9808);
or UO_1158 (O_1158,N_9825,N_9882);
xnor UO_1159 (O_1159,N_9950,N_9902);
nor UO_1160 (O_1160,N_9896,N_9802);
nand UO_1161 (O_1161,N_9835,N_9872);
nor UO_1162 (O_1162,N_9892,N_9994);
nor UO_1163 (O_1163,N_9839,N_9994);
or UO_1164 (O_1164,N_9966,N_9844);
nor UO_1165 (O_1165,N_9941,N_9891);
nand UO_1166 (O_1166,N_9899,N_9875);
nor UO_1167 (O_1167,N_9858,N_9923);
nor UO_1168 (O_1168,N_9867,N_9970);
nor UO_1169 (O_1169,N_9917,N_9916);
and UO_1170 (O_1170,N_9912,N_9861);
and UO_1171 (O_1171,N_9892,N_9937);
xor UO_1172 (O_1172,N_9873,N_9918);
or UO_1173 (O_1173,N_9839,N_9979);
and UO_1174 (O_1174,N_9985,N_9991);
nand UO_1175 (O_1175,N_9871,N_9995);
nand UO_1176 (O_1176,N_9875,N_9855);
and UO_1177 (O_1177,N_9993,N_9827);
and UO_1178 (O_1178,N_9855,N_9953);
nand UO_1179 (O_1179,N_9836,N_9907);
or UO_1180 (O_1180,N_9919,N_9923);
and UO_1181 (O_1181,N_9820,N_9933);
nand UO_1182 (O_1182,N_9847,N_9921);
xnor UO_1183 (O_1183,N_9812,N_9955);
nor UO_1184 (O_1184,N_9858,N_9825);
or UO_1185 (O_1185,N_9839,N_9903);
or UO_1186 (O_1186,N_9844,N_9971);
nand UO_1187 (O_1187,N_9949,N_9860);
nand UO_1188 (O_1188,N_9947,N_9816);
and UO_1189 (O_1189,N_9905,N_9960);
xnor UO_1190 (O_1190,N_9896,N_9912);
and UO_1191 (O_1191,N_9935,N_9972);
and UO_1192 (O_1192,N_9988,N_9973);
nor UO_1193 (O_1193,N_9894,N_9967);
nor UO_1194 (O_1194,N_9909,N_9959);
or UO_1195 (O_1195,N_9807,N_9907);
nand UO_1196 (O_1196,N_9944,N_9936);
nand UO_1197 (O_1197,N_9923,N_9817);
or UO_1198 (O_1198,N_9959,N_9824);
and UO_1199 (O_1199,N_9880,N_9939);
and UO_1200 (O_1200,N_9866,N_9888);
nand UO_1201 (O_1201,N_9916,N_9837);
nand UO_1202 (O_1202,N_9906,N_9924);
nand UO_1203 (O_1203,N_9987,N_9869);
xor UO_1204 (O_1204,N_9966,N_9802);
or UO_1205 (O_1205,N_9858,N_9877);
nor UO_1206 (O_1206,N_9845,N_9853);
nand UO_1207 (O_1207,N_9812,N_9950);
nand UO_1208 (O_1208,N_9852,N_9800);
and UO_1209 (O_1209,N_9884,N_9992);
nand UO_1210 (O_1210,N_9845,N_9843);
or UO_1211 (O_1211,N_9879,N_9902);
and UO_1212 (O_1212,N_9991,N_9931);
xor UO_1213 (O_1213,N_9843,N_9903);
nand UO_1214 (O_1214,N_9930,N_9853);
nor UO_1215 (O_1215,N_9809,N_9996);
or UO_1216 (O_1216,N_9991,N_9907);
nand UO_1217 (O_1217,N_9955,N_9836);
nor UO_1218 (O_1218,N_9909,N_9981);
xor UO_1219 (O_1219,N_9977,N_9969);
xnor UO_1220 (O_1220,N_9871,N_9854);
xnor UO_1221 (O_1221,N_9957,N_9843);
nand UO_1222 (O_1222,N_9913,N_9877);
xor UO_1223 (O_1223,N_9932,N_9955);
or UO_1224 (O_1224,N_9883,N_9906);
and UO_1225 (O_1225,N_9859,N_9898);
nand UO_1226 (O_1226,N_9905,N_9830);
or UO_1227 (O_1227,N_9804,N_9910);
or UO_1228 (O_1228,N_9961,N_9914);
and UO_1229 (O_1229,N_9963,N_9903);
and UO_1230 (O_1230,N_9915,N_9887);
and UO_1231 (O_1231,N_9961,N_9902);
nor UO_1232 (O_1232,N_9973,N_9951);
and UO_1233 (O_1233,N_9937,N_9846);
nand UO_1234 (O_1234,N_9841,N_9878);
nand UO_1235 (O_1235,N_9966,N_9917);
and UO_1236 (O_1236,N_9810,N_9880);
xnor UO_1237 (O_1237,N_9826,N_9893);
and UO_1238 (O_1238,N_9830,N_9885);
nand UO_1239 (O_1239,N_9848,N_9860);
or UO_1240 (O_1240,N_9918,N_9940);
or UO_1241 (O_1241,N_9923,N_9879);
nand UO_1242 (O_1242,N_9975,N_9955);
or UO_1243 (O_1243,N_9987,N_9941);
and UO_1244 (O_1244,N_9906,N_9911);
and UO_1245 (O_1245,N_9889,N_9864);
nand UO_1246 (O_1246,N_9976,N_9917);
nand UO_1247 (O_1247,N_9921,N_9864);
nor UO_1248 (O_1248,N_9858,N_9903);
nor UO_1249 (O_1249,N_9884,N_9845);
nand UO_1250 (O_1250,N_9923,N_9944);
nand UO_1251 (O_1251,N_9893,N_9879);
or UO_1252 (O_1252,N_9873,N_9830);
or UO_1253 (O_1253,N_9848,N_9883);
nor UO_1254 (O_1254,N_9921,N_9952);
or UO_1255 (O_1255,N_9913,N_9843);
or UO_1256 (O_1256,N_9841,N_9922);
nand UO_1257 (O_1257,N_9833,N_9909);
nor UO_1258 (O_1258,N_9939,N_9906);
xor UO_1259 (O_1259,N_9957,N_9928);
nand UO_1260 (O_1260,N_9855,N_9908);
and UO_1261 (O_1261,N_9969,N_9994);
nor UO_1262 (O_1262,N_9934,N_9830);
nand UO_1263 (O_1263,N_9804,N_9862);
nand UO_1264 (O_1264,N_9869,N_9834);
nor UO_1265 (O_1265,N_9995,N_9837);
nand UO_1266 (O_1266,N_9904,N_9956);
or UO_1267 (O_1267,N_9873,N_9924);
or UO_1268 (O_1268,N_9950,N_9863);
or UO_1269 (O_1269,N_9815,N_9971);
nor UO_1270 (O_1270,N_9950,N_9890);
nand UO_1271 (O_1271,N_9825,N_9997);
nand UO_1272 (O_1272,N_9898,N_9861);
nand UO_1273 (O_1273,N_9960,N_9954);
and UO_1274 (O_1274,N_9953,N_9860);
nor UO_1275 (O_1275,N_9898,N_9855);
or UO_1276 (O_1276,N_9920,N_9980);
nand UO_1277 (O_1277,N_9964,N_9965);
xnor UO_1278 (O_1278,N_9846,N_9801);
nand UO_1279 (O_1279,N_9915,N_9952);
nand UO_1280 (O_1280,N_9822,N_9911);
nor UO_1281 (O_1281,N_9983,N_9991);
nand UO_1282 (O_1282,N_9882,N_9908);
nor UO_1283 (O_1283,N_9965,N_9963);
and UO_1284 (O_1284,N_9990,N_9846);
and UO_1285 (O_1285,N_9963,N_9927);
or UO_1286 (O_1286,N_9846,N_9922);
nand UO_1287 (O_1287,N_9966,N_9869);
xor UO_1288 (O_1288,N_9820,N_9992);
and UO_1289 (O_1289,N_9865,N_9884);
nor UO_1290 (O_1290,N_9833,N_9989);
xnor UO_1291 (O_1291,N_9913,N_9961);
nor UO_1292 (O_1292,N_9980,N_9970);
nand UO_1293 (O_1293,N_9985,N_9808);
nor UO_1294 (O_1294,N_9914,N_9899);
and UO_1295 (O_1295,N_9953,N_9869);
nand UO_1296 (O_1296,N_9843,N_9984);
xor UO_1297 (O_1297,N_9879,N_9968);
nand UO_1298 (O_1298,N_9812,N_9877);
nor UO_1299 (O_1299,N_9971,N_9822);
nand UO_1300 (O_1300,N_9823,N_9885);
and UO_1301 (O_1301,N_9969,N_9889);
or UO_1302 (O_1302,N_9950,N_9994);
nor UO_1303 (O_1303,N_9811,N_9842);
nor UO_1304 (O_1304,N_9951,N_9885);
nor UO_1305 (O_1305,N_9979,N_9862);
or UO_1306 (O_1306,N_9934,N_9911);
nor UO_1307 (O_1307,N_9834,N_9968);
nand UO_1308 (O_1308,N_9927,N_9877);
nor UO_1309 (O_1309,N_9971,N_9805);
nand UO_1310 (O_1310,N_9906,N_9858);
xnor UO_1311 (O_1311,N_9917,N_9851);
and UO_1312 (O_1312,N_9910,N_9876);
and UO_1313 (O_1313,N_9879,N_9928);
nor UO_1314 (O_1314,N_9833,N_9926);
nor UO_1315 (O_1315,N_9846,N_9891);
nor UO_1316 (O_1316,N_9915,N_9953);
or UO_1317 (O_1317,N_9914,N_9993);
nor UO_1318 (O_1318,N_9906,N_9933);
and UO_1319 (O_1319,N_9909,N_9870);
nor UO_1320 (O_1320,N_9945,N_9843);
nand UO_1321 (O_1321,N_9851,N_9895);
and UO_1322 (O_1322,N_9988,N_9949);
xor UO_1323 (O_1323,N_9989,N_9853);
and UO_1324 (O_1324,N_9974,N_9943);
nor UO_1325 (O_1325,N_9933,N_9915);
nand UO_1326 (O_1326,N_9834,N_9975);
or UO_1327 (O_1327,N_9949,N_9897);
nor UO_1328 (O_1328,N_9982,N_9959);
or UO_1329 (O_1329,N_9832,N_9908);
or UO_1330 (O_1330,N_9829,N_9910);
and UO_1331 (O_1331,N_9876,N_9968);
and UO_1332 (O_1332,N_9992,N_9954);
or UO_1333 (O_1333,N_9920,N_9829);
and UO_1334 (O_1334,N_9979,N_9940);
nor UO_1335 (O_1335,N_9818,N_9829);
nand UO_1336 (O_1336,N_9861,N_9826);
and UO_1337 (O_1337,N_9979,N_9967);
nand UO_1338 (O_1338,N_9809,N_9834);
nor UO_1339 (O_1339,N_9806,N_9960);
and UO_1340 (O_1340,N_9978,N_9886);
nand UO_1341 (O_1341,N_9980,N_9960);
nor UO_1342 (O_1342,N_9992,N_9910);
nand UO_1343 (O_1343,N_9882,N_9899);
nand UO_1344 (O_1344,N_9918,N_9890);
nand UO_1345 (O_1345,N_9885,N_9845);
or UO_1346 (O_1346,N_9903,N_9957);
or UO_1347 (O_1347,N_9821,N_9872);
xnor UO_1348 (O_1348,N_9846,N_9845);
and UO_1349 (O_1349,N_9910,N_9995);
nand UO_1350 (O_1350,N_9917,N_9870);
nor UO_1351 (O_1351,N_9918,N_9826);
nand UO_1352 (O_1352,N_9800,N_9893);
and UO_1353 (O_1353,N_9961,N_9841);
or UO_1354 (O_1354,N_9944,N_9935);
or UO_1355 (O_1355,N_9884,N_9969);
and UO_1356 (O_1356,N_9905,N_9979);
xnor UO_1357 (O_1357,N_9929,N_9911);
nor UO_1358 (O_1358,N_9979,N_9869);
nor UO_1359 (O_1359,N_9915,N_9867);
nor UO_1360 (O_1360,N_9967,N_9806);
xnor UO_1361 (O_1361,N_9841,N_9845);
xnor UO_1362 (O_1362,N_9875,N_9895);
nand UO_1363 (O_1363,N_9953,N_9912);
and UO_1364 (O_1364,N_9903,N_9822);
nor UO_1365 (O_1365,N_9955,N_9900);
or UO_1366 (O_1366,N_9859,N_9863);
or UO_1367 (O_1367,N_9904,N_9995);
nor UO_1368 (O_1368,N_9894,N_9898);
or UO_1369 (O_1369,N_9954,N_9830);
or UO_1370 (O_1370,N_9962,N_9979);
and UO_1371 (O_1371,N_9888,N_9862);
nor UO_1372 (O_1372,N_9864,N_9952);
or UO_1373 (O_1373,N_9880,N_9916);
xnor UO_1374 (O_1374,N_9845,N_9815);
and UO_1375 (O_1375,N_9961,N_9971);
and UO_1376 (O_1376,N_9906,N_9995);
nand UO_1377 (O_1377,N_9938,N_9993);
nand UO_1378 (O_1378,N_9815,N_9994);
nand UO_1379 (O_1379,N_9851,N_9899);
and UO_1380 (O_1380,N_9811,N_9952);
nor UO_1381 (O_1381,N_9884,N_9860);
and UO_1382 (O_1382,N_9961,N_9813);
nand UO_1383 (O_1383,N_9928,N_9851);
nand UO_1384 (O_1384,N_9812,N_9867);
or UO_1385 (O_1385,N_9831,N_9896);
xor UO_1386 (O_1386,N_9943,N_9937);
and UO_1387 (O_1387,N_9899,N_9905);
or UO_1388 (O_1388,N_9817,N_9998);
or UO_1389 (O_1389,N_9981,N_9928);
xor UO_1390 (O_1390,N_9976,N_9882);
nor UO_1391 (O_1391,N_9886,N_9859);
nor UO_1392 (O_1392,N_9862,N_9843);
and UO_1393 (O_1393,N_9830,N_9856);
and UO_1394 (O_1394,N_9803,N_9868);
nor UO_1395 (O_1395,N_9808,N_9930);
and UO_1396 (O_1396,N_9931,N_9907);
nand UO_1397 (O_1397,N_9958,N_9928);
and UO_1398 (O_1398,N_9931,N_9921);
or UO_1399 (O_1399,N_9898,N_9886);
nand UO_1400 (O_1400,N_9848,N_9949);
nor UO_1401 (O_1401,N_9978,N_9930);
nor UO_1402 (O_1402,N_9878,N_9910);
xnor UO_1403 (O_1403,N_9977,N_9853);
nor UO_1404 (O_1404,N_9848,N_9957);
and UO_1405 (O_1405,N_9857,N_9841);
nor UO_1406 (O_1406,N_9852,N_9945);
nor UO_1407 (O_1407,N_9930,N_9828);
or UO_1408 (O_1408,N_9836,N_9835);
and UO_1409 (O_1409,N_9902,N_9860);
or UO_1410 (O_1410,N_9895,N_9929);
and UO_1411 (O_1411,N_9865,N_9910);
nor UO_1412 (O_1412,N_9802,N_9887);
or UO_1413 (O_1413,N_9891,N_9877);
nand UO_1414 (O_1414,N_9990,N_9887);
or UO_1415 (O_1415,N_9819,N_9962);
or UO_1416 (O_1416,N_9926,N_9813);
or UO_1417 (O_1417,N_9864,N_9922);
and UO_1418 (O_1418,N_9835,N_9803);
nor UO_1419 (O_1419,N_9980,N_9870);
nand UO_1420 (O_1420,N_9804,N_9849);
nand UO_1421 (O_1421,N_9964,N_9970);
nand UO_1422 (O_1422,N_9984,N_9917);
or UO_1423 (O_1423,N_9895,N_9932);
nor UO_1424 (O_1424,N_9820,N_9975);
or UO_1425 (O_1425,N_9814,N_9948);
nand UO_1426 (O_1426,N_9875,N_9990);
nor UO_1427 (O_1427,N_9973,N_9800);
xor UO_1428 (O_1428,N_9862,N_9953);
or UO_1429 (O_1429,N_9900,N_9966);
or UO_1430 (O_1430,N_9933,N_9880);
or UO_1431 (O_1431,N_9843,N_9946);
nor UO_1432 (O_1432,N_9846,N_9913);
and UO_1433 (O_1433,N_9921,N_9939);
nor UO_1434 (O_1434,N_9811,N_9925);
xnor UO_1435 (O_1435,N_9803,N_9808);
and UO_1436 (O_1436,N_9854,N_9864);
and UO_1437 (O_1437,N_9981,N_9956);
or UO_1438 (O_1438,N_9976,N_9987);
nor UO_1439 (O_1439,N_9981,N_9896);
nor UO_1440 (O_1440,N_9994,N_9803);
or UO_1441 (O_1441,N_9894,N_9822);
and UO_1442 (O_1442,N_9942,N_9978);
nor UO_1443 (O_1443,N_9831,N_9850);
nand UO_1444 (O_1444,N_9974,N_9975);
and UO_1445 (O_1445,N_9952,N_9879);
nor UO_1446 (O_1446,N_9831,N_9835);
or UO_1447 (O_1447,N_9831,N_9877);
or UO_1448 (O_1448,N_9928,N_9819);
nand UO_1449 (O_1449,N_9917,N_9882);
or UO_1450 (O_1450,N_9954,N_9970);
or UO_1451 (O_1451,N_9916,N_9821);
nand UO_1452 (O_1452,N_9927,N_9923);
or UO_1453 (O_1453,N_9896,N_9805);
or UO_1454 (O_1454,N_9963,N_9876);
or UO_1455 (O_1455,N_9924,N_9968);
nor UO_1456 (O_1456,N_9999,N_9927);
xnor UO_1457 (O_1457,N_9871,N_9981);
and UO_1458 (O_1458,N_9870,N_9923);
or UO_1459 (O_1459,N_9911,N_9852);
nand UO_1460 (O_1460,N_9988,N_9873);
nand UO_1461 (O_1461,N_9806,N_9828);
nor UO_1462 (O_1462,N_9962,N_9861);
or UO_1463 (O_1463,N_9987,N_9861);
or UO_1464 (O_1464,N_9858,N_9933);
and UO_1465 (O_1465,N_9910,N_9971);
and UO_1466 (O_1466,N_9885,N_9858);
nand UO_1467 (O_1467,N_9883,N_9805);
or UO_1468 (O_1468,N_9863,N_9984);
nor UO_1469 (O_1469,N_9973,N_9996);
nor UO_1470 (O_1470,N_9945,N_9846);
nand UO_1471 (O_1471,N_9900,N_9840);
and UO_1472 (O_1472,N_9903,N_9814);
or UO_1473 (O_1473,N_9999,N_9966);
nand UO_1474 (O_1474,N_9945,N_9858);
nor UO_1475 (O_1475,N_9937,N_9843);
and UO_1476 (O_1476,N_9919,N_9885);
or UO_1477 (O_1477,N_9849,N_9974);
or UO_1478 (O_1478,N_9923,N_9811);
nor UO_1479 (O_1479,N_9919,N_9977);
nor UO_1480 (O_1480,N_9814,N_9851);
and UO_1481 (O_1481,N_9991,N_9965);
nand UO_1482 (O_1482,N_9838,N_9955);
or UO_1483 (O_1483,N_9977,N_9873);
xor UO_1484 (O_1484,N_9931,N_9889);
and UO_1485 (O_1485,N_9927,N_9836);
and UO_1486 (O_1486,N_9880,N_9886);
xor UO_1487 (O_1487,N_9810,N_9836);
or UO_1488 (O_1488,N_9956,N_9805);
and UO_1489 (O_1489,N_9823,N_9831);
or UO_1490 (O_1490,N_9803,N_9992);
nor UO_1491 (O_1491,N_9907,N_9911);
and UO_1492 (O_1492,N_9821,N_9951);
nand UO_1493 (O_1493,N_9985,N_9845);
or UO_1494 (O_1494,N_9927,N_9825);
nor UO_1495 (O_1495,N_9829,N_9979);
and UO_1496 (O_1496,N_9831,N_9895);
nand UO_1497 (O_1497,N_9819,N_9887);
or UO_1498 (O_1498,N_9937,N_9821);
or UO_1499 (O_1499,N_9932,N_9836);
endmodule