module basic_500_3000_500_6_levels_2xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_222,In_7);
nor U1 (N_1,In_328,In_322);
nor U2 (N_2,In_339,In_400);
nor U3 (N_3,In_173,In_426);
nor U4 (N_4,In_141,In_406);
and U5 (N_5,In_410,In_289);
and U6 (N_6,In_464,In_110);
nor U7 (N_7,In_143,In_350);
and U8 (N_8,In_261,In_437);
nand U9 (N_9,In_139,In_6);
or U10 (N_10,In_4,In_147);
nand U11 (N_11,In_208,In_156);
nand U12 (N_12,In_272,In_308);
or U13 (N_13,In_335,In_362);
nand U14 (N_14,In_378,In_342);
and U15 (N_15,In_303,In_405);
or U16 (N_16,In_470,In_346);
and U17 (N_17,In_461,In_51);
and U18 (N_18,In_411,In_217);
nor U19 (N_19,In_469,In_178);
and U20 (N_20,In_353,In_41);
and U21 (N_21,In_284,In_34);
or U22 (N_22,In_356,In_279);
nor U23 (N_23,In_103,In_455);
nor U24 (N_24,In_389,In_466);
and U25 (N_25,In_358,In_334);
xnor U26 (N_26,In_17,In_452);
or U27 (N_27,In_204,In_338);
or U28 (N_28,In_499,In_226);
and U29 (N_29,In_319,In_218);
or U30 (N_30,In_55,In_122);
or U31 (N_31,In_314,In_65);
xnor U32 (N_32,In_463,In_417);
nor U33 (N_33,In_93,In_31);
nor U34 (N_34,In_359,In_121);
or U35 (N_35,In_256,In_113);
or U36 (N_36,In_223,In_393);
nand U37 (N_37,In_23,In_128);
or U38 (N_38,In_37,In_131);
nand U39 (N_39,In_453,In_236);
or U40 (N_40,In_440,In_50);
or U41 (N_41,In_89,In_465);
nand U42 (N_42,In_48,In_152);
nor U43 (N_43,In_233,In_396);
and U44 (N_44,In_340,In_162);
and U45 (N_45,In_416,In_214);
nand U46 (N_46,In_354,In_336);
nor U47 (N_47,In_305,In_395);
nand U48 (N_48,In_247,In_387);
nor U49 (N_49,In_420,In_9);
or U50 (N_50,In_313,In_35);
and U51 (N_51,In_375,In_77);
or U52 (N_52,In_443,In_150);
or U53 (N_53,In_133,In_282);
nor U54 (N_54,In_228,In_138);
or U55 (N_55,In_298,In_476);
or U56 (N_56,In_10,In_429);
nand U57 (N_57,In_70,In_300);
nand U58 (N_58,In_490,In_116);
and U59 (N_59,In_459,In_191);
and U60 (N_60,In_449,In_172);
or U61 (N_61,In_215,In_203);
nor U62 (N_62,In_489,In_211);
nand U63 (N_63,In_190,In_45);
or U64 (N_64,In_98,In_49);
or U65 (N_65,In_245,In_183);
or U66 (N_66,In_482,In_188);
or U67 (N_67,In_164,In_423);
nand U68 (N_68,In_158,In_159);
nand U69 (N_69,In_61,In_419);
nand U70 (N_70,In_95,In_132);
and U71 (N_71,In_382,In_104);
and U72 (N_72,In_343,In_281);
nor U73 (N_73,In_360,In_309);
xnor U74 (N_74,In_14,In_324);
and U75 (N_75,In_265,In_192);
and U76 (N_76,In_331,In_404);
and U77 (N_77,In_462,In_287);
xnor U78 (N_78,In_487,In_210);
or U79 (N_79,In_255,In_82);
and U80 (N_80,In_352,In_80);
nor U81 (N_81,In_175,In_398);
or U82 (N_82,In_52,In_205);
nand U83 (N_83,In_428,In_182);
nand U84 (N_84,In_125,In_383);
xor U85 (N_85,In_137,In_28);
nand U86 (N_86,In_126,In_301);
nor U87 (N_87,In_425,In_15);
nand U88 (N_88,In_363,In_0);
nor U89 (N_89,In_239,In_136);
or U90 (N_90,In_240,In_107);
nor U91 (N_91,In_269,In_69);
and U92 (N_92,In_224,In_181);
nor U93 (N_93,In_479,In_492);
nand U94 (N_94,In_421,In_106);
and U95 (N_95,In_250,In_268);
nand U96 (N_96,In_169,In_170);
and U97 (N_97,In_373,In_195);
or U98 (N_98,In_371,In_71);
or U99 (N_99,In_273,In_456);
nor U100 (N_100,In_290,In_366);
or U101 (N_101,In_263,In_196);
and U102 (N_102,In_326,In_227);
nand U103 (N_103,In_96,In_495);
or U104 (N_104,In_193,In_73);
nand U105 (N_105,In_67,In_36);
or U106 (N_106,In_439,In_63);
or U107 (N_107,In_381,In_311);
or U108 (N_108,In_480,In_262);
or U109 (N_109,In_177,In_32);
nand U110 (N_110,In_414,In_212);
or U111 (N_111,In_11,In_86);
and U112 (N_112,In_140,In_40);
nor U113 (N_113,In_307,In_471);
nand U114 (N_114,In_2,In_20);
nand U115 (N_115,In_127,In_16);
nand U116 (N_116,In_22,In_248);
nor U117 (N_117,In_179,In_488);
and U118 (N_118,In_33,In_241);
nand U119 (N_119,In_266,In_18);
or U120 (N_120,In_312,In_385);
nand U121 (N_121,In_286,In_124);
or U122 (N_122,In_430,In_388);
nand U123 (N_123,In_12,In_76);
nor U124 (N_124,In_253,In_75);
nand U125 (N_125,In_165,In_92);
and U126 (N_126,In_333,In_243);
nor U127 (N_127,In_415,In_280);
nor U128 (N_128,In_315,In_294);
or U129 (N_129,In_441,In_90);
xor U130 (N_130,In_30,In_408);
nand U131 (N_131,In_102,In_201);
or U132 (N_132,In_60,In_148);
nor U133 (N_133,In_186,In_392);
and U134 (N_134,In_329,In_99);
and U135 (N_135,In_115,In_232);
and U136 (N_136,In_384,In_142);
nor U137 (N_137,In_88,In_157);
or U138 (N_138,In_259,In_468);
nor U139 (N_139,In_260,In_153);
and U140 (N_140,In_422,In_278);
and U141 (N_141,In_8,In_213);
or U142 (N_142,In_361,In_101);
nand U143 (N_143,In_187,In_364);
nor U144 (N_144,In_87,In_118);
and U145 (N_145,In_344,In_450);
nor U146 (N_146,In_486,In_221);
nor U147 (N_147,In_84,In_166);
or U148 (N_148,In_59,In_238);
nor U149 (N_149,In_401,In_174);
and U150 (N_150,In_380,In_254);
or U151 (N_151,In_317,In_168);
and U152 (N_152,In_83,In_200);
nand U153 (N_153,In_171,In_270);
and U154 (N_154,In_413,In_407);
nand U155 (N_155,In_185,In_38);
nor U156 (N_156,In_206,In_368);
nand U157 (N_157,In_94,In_402);
nand U158 (N_158,In_267,In_299);
nand U159 (N_159,In_1,In_374);
nand U160 (N_160,In_390,In_249);
nand U161 (N_161,In_424,In_438);
nand U162 (N_162,In_473,In_478);
or U163 (N_163,In_78,In_120);
nor U164 (N_164,In_271,In_283);
and U165 (N_165,In_231,In_3);
and U166 (N_166,In_444,In_54);
and U167 (N_167,In_347,In_24);
nand U168 (N_168,In_377,In_306);
or U169 (N_169,In_225,In_318);
or U170 (N_170,In_276,In_467);
nor U171 (N_171,In_100,In_348);
and U172 (N_172,In_19,In_62);
or U173 (N_173,In_246,In_234);
and U174 (N_174,In_337,In_130);
and U175 (N_175,In_197,In_494);
or U176 (N_176,In_341,In_292);
nand U177 (N_177,In_167,In_105);
and U178 (N_178,In_42,In_230);
nor U179 (N_179,In_251,In_258);
and U180 (N_180,In_370,In_27);
nor U181 (N_181,In_295,In_129);
and U182 (N_182,In_448,In_117);
and U183 (N_183,In_144,In_13);
nor U184 (N_184,In_275,In_285);
nand U185 (N_185,In_297,In_330);
or U186 (N_186,In_372,In_433);
or U187 (N_187,In_109,In_26);
nand U188 (N_188,In_367,In_57);
or U189 (N_189,In_446,In_202);
or U190 (N_190,In_293,In_198);
or U191 (N_191,In_394,In_154);
and U192 (N_192,In_119,In_155);
nand U193 (N_193,In_351,In_161);
nor U194 (N_194,In_498,In_345);
nor U195 (N_195,In_209,In_44);
or U196 (N_196,In_349,In_79);
or U197 (N_197,In_123,In_25);
and U198 (N_198,In_474,In_111);
nor U199 (N_199,In_160,In_244);
nor U200 (N_200,In_386,In_145);
and U201 (N_201,In_66,In_485);
or U202 (N_202,In_237,In_68);
and U203 (N_203,In_242,In_151);
nand U204 (N_204,In_445,In_97);
and U205 (N_205,In_323,In_219);
and U206 (N_206,In_458,In_176);
nand U207 (N_207,In_316,In_481);
or U208 (N_208,In_134,In_365);
and U209 (N_209,In_397,In_403);
nor U210 (N_210,In_264,In_108);
nand U211 (N_211,In_332,In_457);
or U212 (N_212,In_277,In_447);
and U213 (N_213,In_475,In_29);
nor U214 (N_214,In_376,In_207);
or U215 (N_215,In_296,In_288);
and U216 (N_216,In_369,In_497);
xnor U217 (N_217,In_43,In_85);
and U218 (N_218,In_435,In_58);
nor U219 (N_219,In_220,In_21);
nand U220 (N_220,In_432,In_72);
nor U221 (N_221,In_53,In_149);
nand U222 (N_222,In_291,In_39);
nor U223 (N_223,In_321,In_252);
and U224 (N_224,In_442,In_493);
nor U225 (N_225,In_163,In_229);
and U226 (N_226,In_418,In_47);
xor U227 (N_227,In_114,In_379);
nand U228 (N_228,In_427,In_460);
and U229 (N_229,In_180,In_216);
nand U230 (N_230,In_355,In_274);
and U231 (N_231,In_436,In_472);
nor U232 (N_232,In_496,In_46);
or U233 (N_233,In_357,In_491);
or U234 (N_234,In_325,In_5);
or U235 (N_235,In_112,In_146);
and U236 (N_236,In_74,In_310);
and U237 (N_237,In_484,In_189);
and U238 (N_238,In_235,In_81);
nand U239 (N_239,In_477,In_184);
or U240 (N_240,In_302,In_64);
nand U241 (N_241,In_451,In_434);
nand U242 (N_242,In_412,In_304);
and U243 (N_243,In_194,In_327);
and U244 (N_244,In_56,In_199);
xnor U245 (N_245,In_454,In_135);
and U246 (N_246,In_91,In_257);
and U247 (N_247,In_409,In_391);
or U248 (N_248,In_320,In_483);
nor U249 (N_249,In_399,In_431);
xnor U250 (N_250,In_273,In_35);
nor U251 (N_251,In_49,In_258);
nand U252 (N_252,In_76,In_445);
nor U253 (N_253,In_21,In_177);
nand U254 (N_254,In_351,In_220);
or U255 (N_255,In_365,In_138);
and U256 (N_256,In_129,In_134);
nand U257 (N_257,In_190,In_438);
or U258 (N_258,In_433,In_238);
nand U259 (N_259,In_385,In_477);
nand U260 (N_260,In_428,In_464);
and U261 (N_261,In_38,In_397);
nand U262 (N_262,In_433,In_363);
and U263 (N_263,In_106,In_245);
xor U264 (N_264,In_433,In_286);
and U265 (N_265,In_266,In_85);
and U266 (N_266,In_293,In_240);
xnor U267 (N_267,In_384,In_151);
and U268 (N_268,In_452,In_268);
nor U269 (N_269,In_34,In_56);
or U270 (N_270,In_10,In_318);
nor U271 (N_271,In_334,In_183);
nand U272 (N_272,In_186,In_369);
or U273 (N_273,In_397,In_229);
and U274 (N_274,In_60,In_251);
nand U275 (N_275,In_274,In_66);
nor U276 (N_276,In_1,In_414);
and U277 (N_277,In_59,In_307);
nor U278 (N_278,In_322,In_16);
or U279 (N_279,In_249,In_169);
nand U280 (N_280,In_340,In_271);
nand U281 (N_281,In_35,In_160);
nor U282 (N_282,In_33,In_279);
or U283 (N_283,In_167,In_85);
and U284 (N_284,In_340,In_280);
or U285 (N_285,In_463,In_263);
nand U286 (N_286,In_143,In_277);
and U287 (N_287,In_321,In_283);
and U288 (N_288,In_444,In_368);
nand U289 (N_289,In_338,In_142);
or U290 (N_290,In_431,In_476);
nor U291 (N_291,In_204,In_371);
nor U292 (N_292,In_133,In_321);
nor U293 (N_293,In_76,In_462);
and U294 (N_294,In_481,In_118);
and U295 (N_295,In_193,In_215);
or U296 (N_296,In_305,In_254);
or U297 (N_297,In_40,In_28);
and U298 (N_298,In_354,In_153);
nand U299 (N_299,In_289,In_149);
or U300 (N_300,In_367,In_423);
xnor U301 (N_301,In_126,In_92);
nand U302 (N_302,In_70,In_434);
or U303 (N_303,In_2,In_139);
and U304 (N_304,In_254,In_144);
or U305 (N_305,In_158,In_320);
or U306 (N_306,In_87,In_260);
and U307 (N_307,In_381,In_12);
or U308 (N_308,In_205,In_353);
nand U309 (N_309,In_498,In_276);
or U310 (N_310,In_81,In_489);
nand U311 (N_311,In_189,In_222);
and U312 (N_312,In_362,In_210);
nand U313 (N_313,In_275,In_450);
and U314 (N_314,In_291,In_398);
and U315 (N_315,In_126,In_146);
nand U316 (N_316,In_30,In_470);
or U317 (N_317,In_304,In_193);
nor U318 (N_318,In_291,In_25);
nand U319 (N_319,In_370,In_373);
and U320 (N_320,In_464,In_183);
nor U321 (N_321,In_251,In_65);
nor U322 (N_322,In_255,In_491);
nand U323 (N_323,In_485,In_129);
nand U324 (N_324,In_224,In_244);
nand U325 (N_325,In_15,In_267);
nor U326 (N_326,In_268,In_112);
nor U327 (N_327,In_384,In_258);
nor U328 (N_328,In_197,In_285);
and U329 (N_329,In_474,In_138);
or U330 (N_330,In_440,In_230);
and U331 (N_331,In_146,In_324);
or U332 (N_332,In_453,In_13);
nor U333 (N_333,In_493,In_167);
or U334 (N_334,In_260,In_390);
and U335 (N_335,In_194,In_120);
and U336 (N_336,In_489,In_361);
nor U337 (N_337,In_255,In_438);
nand U338 (N_338,In_364,In_368);
and U339 (N_339,In_437,In_410);
nand U340 (N_340,In_130,In_421);
nand U341 (N_341,In_422,In_214);
nand U342 (N_342,In_372,In_40);
xnor U343 (N_343,In_223,In_147);
nand U344 (N_344,In_170,In_112);
and U345 (N_345,In_449,In_86);
or U346 (N_346,In_448,In_18);
and U347 (N_347,In_204,In_347);
and U348 (N_348,In_148,In_337);
or U349 (N_349,In_405,In_112);
and U350 (N_350,In_305,In_189);
nand U351 (N_351,In_211,In_8);
and U352 (N_352,In_149,In_111);
or U353 (N_353,In_422,In_201);
nor U354 (N_354,In_419,In_425);
or U355 (N_355,In_261,In_149);
nor U356 (N_356,In_480,In_453);
nor U357 (N_357,In_198,In_262);
nor U358 (N_358,In_275,In_94);
and U359 (N_359,In_287,In_234);
nand U360 (N_360,In_472,In_48);
and U361 (N_361,In_459,In_227);
nand U362 (N_362,In_379,In_181);
xnor U363 (N_363,In_395,In_373);
nand U364 (N_364,In_354,In_10);
or U365 (N_365,In_368,In_363);
nand U366 (N_366,In_166,In_115);
nand U367 (N_367,In_70,In_315);
and U368 (N_368,In_357,In_309);
and U369 (N_369,In_112,In_474);
nor U370 (N_370,In_285,In_376);
nand U371 (N_371,In_27,In_431);
nor U372 (N_372,In_258,In_372);
and U373 (N_373,In_104,In_207);
xnor U374 (N_374,In_486,In_101);
and U375 (N_375,In_162,In_150);
and U376 (N_376,In_399,In_469);
or U377 (N_377,In_336,In_21);
nor U378 (N_378,In_199,In_402);
and U379 (N_379,In_263,In_127);
and U380 (N_380,In_235,In_271);
nand U381 (N_381,In_123,In_210);
and U382 (N_382,In_487,In_176);
nor U383 (N_383,In_0,In_186);
and U384 (N_384,In_68,In_181);
nand U385 (N_385,In_477,In_10);
and U386 (N_386,In_100,In_263);
and U387 (N_387,In_350,In_5);
or U388 (N_388,In_362,In_421);
nor U389 (N_389,In_308,In_420);
nor U390 (N_390,In_36,In_0);
nand U391 (N_391,In_423,In_434);
nor U392 (N_392,In_389,In_80);
and U393 (N_393,In_20,In_337);
and U394 (N_394,In_81,In_348);
or U395 (N_395,In_372,In_290);
or U396 (N_396,In_44,In_197);
or U397 (N_397,In_77,In_373);
and U398 (N_398,In_178,In_270);
or U399 (N_399,In_285,In_463);
nand U400 (N_400,In_483,In_33);
and U401 (N_401,In_109,In_276);
nand U402 (N_402,In_237,In_226);
or U403 (N_403,In_370,In_240);
nor U404 (N_404,In_360,In_277);
nand U405 (N_405,In_158,In_265);
nand U406 (N_406,In_164,In_47);
and U407 (N_407,In_422,In_132);
nor U408 (N_408,In_245,In_147);
nand U409 (N_409,In_398,In_127);
and U410 (N_410,In_241,In_356);
or U411 (N_411,In_493,In_205);
and U412 (N_412,In_207,In_345);
or U413 (N_413,In_411,In_78);
nand U414 (N_414,In_333,In_385);
and U415 (N_415,In_22,In_33);
xnor U416 (N_416,In_379,In_464);
nor U417 (N_417,In_406,In_453);
nor U418 (N_418,In_312,In_302);
or U419 (N_419,In_139,In_91);
nand U420 (N_420,In_419,In_200);
nor U421 (N_421,In_428,In_330);
and U422 (N_422,In_178,In_151);
nor U423 (N_423,In_241,In_221);
nand U424 (N_424,In_128,In_52);
and U425 (N_425,In_91,In_168);
nor U426 (N_426,In_290,In_350);
or U427 (N_427,In_414,In_111);
nand U428 (N_428,In_376,In_433);
and U429 (N_429,In_203,In_415);
and U430 (N_430,In_456,In_397);
nand U431 (N_431,In_103,In_469);
nand U432 (N_432,In_263,In_173);
nor U433 (N_433,In_245,In_429);
or U434 (N_434,In_422,In_341);
nor U435 (N_435,In_214,In_448);
and U436 (N_436,In_229,In_199);
or U437 (N_437,In_276,In_178);
or U438 (N_438,In_90,In_177);
nand U439 (N_439,In_39,In_230);
nand U440 (N_440,In_185,In_301);
and U441 (N_441,In_454,In_5);
and U442 (N_442,In_376,In_409);
nand U443 (N_443,In_330,In_156);
nand U444 (N_444,In_274,In_336);
nor U445 (N_445,In_151,In_161);
and U446 (N_446,In_242,In_124);
or U447 (N_447,In_422,In_228);
nand U448 (N_448,In_491,In_186);
or U449 (N_449,In_460,In_88);
and U450 (N_450,In_413,In_358);
nor U451 (N_451,In_163,In_34);
and U452 (N_452,In_90,In_179);
or U453 (N_453,In_147,In_375);
nor U454 (N_454,In_357,In_131);
nor U455 (N_455,In_61,In_11);
nor U456 (N_456,In_3,In_275);
nand U457 (N_457,In_53,In_471);
or U458 (N_458,In_230,In_352);
and U459 (N_459,In_437,In_242);
or U460 (N_460,In_455,In_248);
or U461 (N_461,In_312,In_300);
nand U462 (N_462,In_158,In_432);
or U463 (N_463,In_237,In_385);
or U464 (N_464,In_278,In_350);
and U465 (N_465,In_288,In_350);
and U466 (N_466,In_294,In_74);
nor U467 (N_467,In_343,In_0);
nand U468 (N_468,In_42,In_413);
nand U469 (N_469,In_426,In_416);
or U470 (N_470,In_468,In_276);
or U471 (N_471,In_274,In_163);
nor U472 (N_472,In_116,In_151);
or U473 (N_473,In_427,In_420);
nand U474 (N_474,In_443,In_496);
nand U475 (N_475,In_91,In_454);
and U476 (N_476,In_142,In_110);
or U477 (N_477,In_384,In_351);
and U478 (N_478,In_334,In_84);
and U479 (N_479,In_368,In_300);
nand U480 (N_480,In_285,In_400);
nand U481 (N_481,In_157,In_211);
or U482 (N_482,In_114,In_346);
nand U483 (N_483,In_56,In_475);
xnor U484 (N_484,In_85,In_25);
and U485 (N_485,In_356,In_381);
and U486 (N_486,In_308,In_459);
or U487 (N_487,In_42,In_43);
or U488 (N_488,In_238,In_402);
nor U489 (N_489,In_84,In_422);
nor U490 (N_490,In_442,In_430);
nor U491 (N_491,In_478,In_62);
or U492 (N_492,In_153,In_107);
and U493 (N_493,In_368,In_359);
and U494 (N_494,In_90,In_103);
nand U495 (N_495,In_402,In_350);
and U496 (N_496,In_485,In_282);
or U497 (N_497,In_154,In_331);
nand U498 (N_498,In_343,In_330);
nand U499 (N_499,In_251,In_26);
nand U500 (N_500,N_61,N_426);
or U501 (N_501,N_442,N_323);
or U502 (N_502,N_321,N_295);
nand U503 (N_503,N_160,N_367);
nor U504 (N_504,N_141,N_66);
nand U505 (N_505,N_2,N_288);
and U506 (N_506,N_98,N_440);
or U507 (N_507,N_252,N_207);
nand U508 (N_508,N_450,N_37);
nand U509 (N_509,N_76,N_162);
and U510 (N_510,N_53,N_497);
or U511 (N_511,N_276,N_153);
nand U512 (N_512,N_167,N_366);
or U513 (N_513,N_372,N_472);
and U514 (N_514,N_401,N_30);
nand U515 (N_515,N_104,N_460);
nand U516 (N_516,N_226,N_130);
or U517 (N_517,N_181,N_376);
nor U518 (N_518,N_95,N_265);
nor U519 (N_519,N_468,N_356);
nor U520 (N_520,N_424,N_240);
nor U521 (N_521,N_57,N_304);
nand U522 (N_522,N_337,N_13);
nor U523 (N_523,N_229,N_219);
nand U524 (N_524,N_488,N_224);
or U525 (N_525,N_112,N_329);
nor U526 (N_526,N_209,N_354);
nand U527 (N_527,N_370,N_218);
nand U528 (N_528,N_429,N_319);
nor U529 (N_529,N_467,N_179);
and U530 (N_530,N_42,N_186);
and U531 (N_531,N_231,N_176);
and U532 (N_532,N_23,N_481);
nor U533 (N_533,N_341,N_109);
nor U534 (N_534,N_364,N_325);
nand U535 (N_535,N_308,N_234);
nor U536 (N_536,N_486,N_458);
or U537 (N_537,N_39,N_375);
or U538 (N_538,N_421,N_430);
nand U539 (N_539,N_236,N_123);
and U540 (N_540,N_335,N_330);
nand U541 (N_541,N_355,N_54);
and U542 (N_542,N_15,N_137);
and U543 (N_543,N_485,N_21);
nor U544 (N_544,N_177,N_267);
nor U545 (N_545,N_345,N_106);
or U546 (N_546,N_79,N_299);
or U547 (N_547,N_48,N_230);
and U548 (N_548,N_483,N_408);
and U549 (N_549,N_175,N_403);
nand U550 (N_550,N_263,N_365);
and U551 (N_551,N_427,N_250);
and U552 (N_552,N_262,N_38);
and U553 (N_553,N_373,N_74);
nor U554 (N_554,N_269,N_397);
and U555 (N_555,N_119,N_285);
nor U556 (N_556,N_145,N_161);
or U557 (N_557,N_72,N_443);
and U558 (N_558,N_261,N_12);
or U559 (N_559,N_422,N_88);
nand U560 (N_560,N_482,N_111);
or U561 (N_561,N_155,N_96);
and U562 (N_562,N_107,N_462);
nor U563 (N_563,N_152,N_143);
and U564 (N_564,N_441,N_16);
or U565 (N_565,N_292,N_447);
nand U566 (N_566,N_147,N_333);
xnor U567 (N_567,N_127,N_387);
or U568 (N_568,N_182,N_245);
nor U569 (N_569,N_60,N_40);
and U570 (N_570,N_383,N_310);
and U571 (N_571,N_394,N_19);
or U572 (N_572,N_85,N_92);
nand U573 (N_573,N_431,N_17);
nand U574 (N_574,N_348,N_69);
and U575 (N_575,N_277,N_469);
nand U576 (N_576,N_433,N_62);
nor U577 (N_577,N_411,N_158);
and U578 (N_578,N_291,N_20);
nand U579 (N_579,N_339,N_289);
nand U580 (N_580,N_18,N_172);
nand U581 (N_581,N_243,N_78);
and U582 (N_582,N_150,N_41);
nand U583 (N_583,N_84,N_228);
or U584 (N_584,N_82,N_75);
nand U585 (N_585,N_331,N_453);
or U586 (N_586,N_242,N_413);
nand U587 (N_587,N_259,N_196);
nor U588 (N_588,N_416,N_379);
or U589 (N_589,N_32,N_210);
nand U590 (N_590,N_398,N_284);
nor U591 (N_591,N_24,N_390);
or U592 (N_592,N_399,N_33);
or U593 (N_593,N_105,N_169);
and U594 (N_594,N_336,N_43);
and U595 (N_595,N_233,N_352);
and U596 (N_596,N_184,N_378);
or U597 (N_597,N_223,N_326);
or U598 (N_598,N_216,N_1);
and U599 (N_599,N_148,N_342);
nand U600 (N_600,N_268,N_139);
or U601 (N_601,N_253,N_102);
nand U602 (N_602,N_126,N_385);
or U603 (N_603,N_165,N_464);
and U604 (N_604,N_118,N_206);
or U605 (N_605,N_166,N_65);
or U606 (N_606,N_451,N_314);
and U607 (N_607,N_97,N_180);
nor U608 (N_608,N_56,N_215);
and U609 (N_609,N_100,N_414);
and U610 (N_610,N_410,N_480);
or U611 (N_611,N_93,N_412);
nor U612 (N_612,N_301,N_396);
nor U613 (N_613,N_437,N_129);
and U614 (N_614,N_183,N_322);
or U615 (N_615,N_131,N_340);
or U616 (N_616,N_34,N_272);
or U617 (N_617,N_374,N_211);
or U618 (N_618,N_492,N_311);
or U619 (N_619,N_212,N_247);
nand U620 (N_620,N_132,N_478);
or U621 (N_621,N_201,N_25);
nor U622 (N_622,N_27,N_439);
and U623 (N_623,N_8,N_257);
nor U624 (N_624,N_280,N_122);
nor U625 (N_625,N_476,N_275);
nor U626 (N_626,N_248,N_477);
or U627 (N_627,N_125,N_22);
or U628 (N_628,N_237,N_448);
and U629 (N_629,N_395,N_94);
nor U630 (N_630,N_349,N_347);
or U631 (N_631,N_296,N_498);
xor U632 (N_632,N_381,N_279);
and U633 (N_633,N_168,N_473);
nand U634 (N_634,N_204,N_353);
nor U635 (N_635,N_116,N_91);
or U636 (N_636,N_121,N_281);
and U637 (N_637,N_222,N_446);
nor U638 (N_638,N_317,N_52);
and U639 (N_639,N_271,N_73);
nand U640 (N_640,N_293,N_404);
nand U641 (N_641,N_418,N_51);
and U642 (N_642,N_178,N_278);
nand U643 (N_643,N_192,N_140);
and U644 (N_644,N_435,N_297);
and U645 (N_645,N_260,N_344);
nor U646 (N_646,N_380,N_157);
nand U647 (N_647,N_4,N_309);
nor U648 (N_648,N_189,N_171);
nand U649 (N_649,N_400,N_273);
nor U650 (N_650,N_244,N_386);
or U651 (N_651,N_235,N_452);
nor U652 (N_652,N_357,N_159);
nor U653 (N_653,N_423,N_164);
or U654 (N_654,N_246,N_313);
xor U655 (N_655,N_101,N_264);
nand U656 (N_656,N_238,N_220);
and U657 (N_657,N_149,N_5);
nand U658 (N_658,N_362,N_203);
or U659 (N_659,N_99,N_493);
and U660 (N_660,N_489,N_46);
or U661 (N_661,N_350,N_459);
nor U662 (N_662,N_146,N_417);
xor U663 (N_663,N_270,N_438);
and U664 (N_664,N_334,N_256);
nor U665 (N_665,N_484,N_205);
or U666 (N_666,N_457,N_0);
xnor U667 (N_667,N_454,N_315);
and U668 (N_668,N_103,N_194);
nor U669 (N_669,N_283,N_202);
or U670 (N_670,N_117,N_120);
and U671 (N_671,N_445,N_318);
nor U672 (N_672,N_64,N_405);
or U673 (N_673,N_346,N_68);
nor U674 (N_674,N_185,N_327);
nand U675 (N_675,N_163,N_81);
nor U676 (N_676,N_108,N_303);
nand U677 (N_677,N_463,N_36);
nor U678 (N_678,N_351,N_298);
nor U679 (N_679,N_343,N_55);
or U680 (N_680,N_9,N_361);
and U681 (N_681,N_136,N_384);
nand U682 (N_682,N_50,N_144);
or U683 (N_683,N_151,N_282);
nand U684 (N_684,N_499,N_409);
nand U685 (N_685,N_225,N_174);
nand U686 (N_686,N_449,N_3);
nor U687 (N_687,N_47,N_360);
nor U688 (N_688,N_113,N_406);
nand U689 (N_689,N_425,N_138);
nor U690 (N_690,N_305,N_11);
nand U691 (N_691,N_474,N_227);
or U692 (N_692,N_191,N_455);
or U693 (N_693,N_491,N_392);
nor U694 (N_694,N_239,N_142);
xor U695 (N_695,N_199,N_221);
nand U696 (N_696,N_6,N_302);
nor U697 (N_697,N_475,N_266);
nand U698 (N_698,N_31,N_35);
nand U699 (N_699,N_110,N_371);
nor U700 (N_700,N_420,N_434);
and U701 (N_701,N_133,N_154);
xor U702 (N_702,N_456,N_290);
or U703 (N_703,N_407,N_432);
nor U704 (N_704,N_419,N_67);
nor U705 (N_705,N_70,N_369);
nor U706 (N_706,N_428,N_26);
or U707 (N_707,N_255,N_294);
and U708 (N_708,N_307,N_134);
nor U709 (N_709,N_382,N_241);
nand U710 (N_710,N_217,N_197);
nor U711 (N_711,N_200,N_389);
nor U712 (N_712,N_258,N_80);
and U713 (N_713,N_358,N_115);
or U714 (N_714,N_135,N_63);
nor U715 (N_715,N_71,N_444);
nand U716 (N_716,N_14,N_466);
or U717 (N_717,N_287,N_436);
nand U718 (N_718,N_208,N_190);
and U719 (N_719,N_286,N_306);
or U720 (N_720,N_391,N_124);
nor U721 (N_721,N_90,N_58);
nor U722 (N_722,N_87,N_312);
nor U723 (N_723,N_232,N_470);
nand U724 (N_724,N_114,N_490);
nand U725 (N_725,N_83,N_393);
or U726 (N_726,N_128,N_368);
or U727 (N_727,N_465,N_316);
or U728 (N_728,N_300,N_187);
nor U729 (N_729,N_10,N_328);
or U730 (N_730,N_487,N_363);
nand U731 (N_731,N_254,N_59);
xnor U732 (N_732,N_198,N_49);
nor U733 (N_733,N_338,N_213);
nor U734 (N_734,N_249,N_388);
or U735 (N_735,N_494,N_332);
or U736 (N_736,N_188,N_320);
nor U737 (N_737,N_193,N_44);
and U738 (N_738,N_45,N_89);
or U739 (N_739,N_274,N_86);
or U740 (N_740,N_471,N_496);
and U741 (N_741,N_77,N_324);
nand U742 (N_742,N_251,N_359);
xor U743 (N_743,N_214,N_156);
and U744 (N_744,N_29,N_28);
nand U745 (N_745,N_495,N_170);
or U746 (N_746,N_195,N_461);
nor U747 (N_747,N_415,N_402);
nor U748 (N_748,N_479,N_173);
xor U749 (N_749,N_7,N_377);
nand U750 (N_750,N_462,N_148);
or U751 (N_751,N_357,N_371);
or U752 (N_752,N_244,N_379);
or U753 (N_753,N_416,N_300);
or U754 (N_754,N_288,N_416);
nand U755 (N_755,N_279,N_201);
nor U756 (N_756,N_15,N_68);
nor U757 (N_757,N_205,N_395);
and U758 (N_758,N_133,N_248);
nand U759 (N_759,N_181,N_480);
and U760 (N_760,N_490,N_388);
xor U761 (N_761,N_32,N_135);
and U762 (N_762,N_107,N_266);
and U763 (N_763,N_296,N_77);
and U764 (N_764,N_61,N_170);
and U765 (N_765,N_197,N_123);
nand U766 (N_766,N_257,N_210);
or U767 (N_767,N_301,N_117);
and U768 (N_768,N_384,N_223);
nand U769 (N_769,N_333,N_44);
or U770 (N_770,N_204,N_159);
xor U771 (N_771,N_5,N_410);
xnor U772 (N_772,N_411,N_259);
nand U773 (N_773,N_431,N_384);
xor U774 (N_774,N_314,N_156);
nor U775 (N_775,N_253,N_331);
or U776 (N_776,N_228,N_37);
nor U777 (N_777,N_495,N_211);
nand U778 (N_778,N_301,N_492);
nand U779 (N_779,N_145,N_400);
and U780 (N_780,N_229,N_133);
and U781 (N_781,N_145,N_337);
or U782 (N_782,N_432,N_96);
or U783 (N_783,N_126,N_290);
and U784 (N_784,N_434,N_51);
or U785 (N_785,N_29,N_402);
and U786 (N_786,N_35,N_246);
or U787 (N_787,N_324,N_58);
or U788 (N_788,N_63,N_421);
nand U789 (N_789,N_186,N_198);
nor U790 (N_790,N_435,N_382);
nand U791 (N_791,N_40,N_47);
nand U792 (N_792,N_282,N_192);
nor U793 (N_793,N_252,N_435);
nand U794 (N_794,N_133,N_367);
nor U795 (N_795,N_484,N_52);
nand U796 (N_796,N_464,N_113);
nor U797 (N_797,N_243,N_79);
or U798 (N_798,N_118,N_78);
xnor U799 (N_799,N_344,N_78);
nor U800 (N_800,N_10,N_402);
and U801 (N_801,N_127,N_490);
nand U802 (N_802,N_213,N_364);
nand U803 (N_803,N_371,N_407);
nor U804 (N_804,N_221,N_394);
and U805 (N_805,N_170,N_91);
nor U806 (N_806,N_482,N_281);
or U807 (N_807,N_298,N_431);
and U808 (N_808,N_474,N_374);
nor U809 (N_809,N_489,N_196);
and U810 (N_810,N_480,N_160);
or U811 (N_811,N_129,N_359);
and U812 (N_812,N_141,N_460);
and U813 (N_813,N_34,N_459);
and U814 (N_814,N_394,N_117);
nand U815 (N_815,N_378,N_445);
or U816 (N_816,N_189,N_191);
nand U817 (N_817,N_276,N_231);
nor U818 (N_818,N_206,N_299);
nand U819 (N_819,N_458,N_111);
and U820 (N_820,N_495,N_53);
nand U821 (N_821,N_474,N_86);
nand U822 (N_822,N_156,N_293);
and U823 (N_823,N_89,N_188);
nand U824 (N_824,N_269,N_2);
nor U825 (N_825,N_300,N_451);
or U826 (N_826,N_452,N_379);
or U827 (N_827,N_156,N_429);
nor U828 (N_828,N_419,N_101);
nor U829 (N_829,N_300,N_333);
nand U830 (N_830,N_350,N_334);
nor U831 (N_831,N_162,N_20);
and U832 (N_832,N_68,N_263);
or U833 (N_833,N_341,N_464);
or U834 (N_834,N_183,N_50);
and U835 (N_835,N_128,N_390);
nor U836 (N_836,N_175,N_89);
nor U837 (N_837,N_294,N_394);
xnor U838 (N_838,N_238,N_217);
nor U839 (N_839,N_462,N_49);
and U840 (N_840,N_128,N_156);
or U841 (N_841,N_220,N_233);
nor U842 (N_842,N_192,N_454);
or U843 (N_843,N_439,N_267);
nand U844 (N_844,N_156,N_68);
nand U845 (N_845,N_238,N_289);
xor U846 (N_846,N_119,N_397);
nor U847 (N_847,N_492,N_19);
and U848 (N_848,N_425,N_205);
and U849 (N_849,N_101,N_299);
nor U850 (N_850,N_421,N_121);
nand U851 (N_851,N_133,N_179);
nor U852 (N_852,N_72,N_32);
nand U853 (N_853,N_135,N_415);
and U854 (N_854,N_124,N_146);
nand U855 (N_855,N_266,N_320);
and U856 (N_856,N_493,N_221);
nand U857 (N_857,N_287,N_329);
or U858 (N_858,N_436,N_134);
or U859 (N_859,N_263,N_112);
nor U860 (N_860,N_130,N_345);
or U861 (N_861,N_4,N_134);
and U862 (N_862,N_72,N_22);
nor U863 (N_863,N_59,N_287);
nand U864 (N_864,N_382,N_354);
nand U865 (N_865,N_88,N_354);
or U866 (N_866,N_83,N_465);
or U867 (N_867,N_252,N_180);
or U868 (N_868,N_168,N_92);
or U869 (N_869,N_42,N_201);
and U870 (N_870,N_85,N_288);
nor U871 (N_871,N_343,N_91);
or U872 (N_872,N_471,N_468);
nand U873 (N_873,N_215,N_53);
or U874 (N_874,N_380,N_339);
nand U875 (N_875,N_345,N_25);
and U876 (N_876,N_295,N_104);
or U877 (N_877,N_422,N_241);
nand U878 (N_878,N_188,N_279);
nor U879 (N_879,N_336,N_393);
and U880 (N_880,N_185,N_418);
or U881 (N_881,N_113,N_474);
nor U882 (N_882,N_72,N_240);
nand U883 (N_883,N_349,N_56);
and U884 (N_884,N_15,N_4);
nand U885 (N_885,N_210,N_168);
nand U886 (N_886,N_475,N_389);
nand U887 (N_887,N_382,N_173);
and U888 (N_888,N_314,N_249);
nand U889 (N_889,N_9,N_438);
nand U890 (N_890,N_356,N_138);
or U891 (N_891,N_19,N_345);
or U892 (N_892,N_96,N_247);
nor U893 (N_893,N_395,N_218);
nand U894 (N_894,N_261,N_255);
nor U895 (N_895,N_152,N_261);
and U896 (N_896,N_50,N_268);
nor U897 (N_897,N_364,N_248);
nor U898 (N_898,N_284,N_82);
nand U899 (N_899,N_462,N_53);
or U900 (N_900,N_453,N_57);
and U901 (N_901,N_188,N_300);
nand U902 (N_902,N_439,N_432);
and U903 (N_903,N_208,N_30);
or U904 (N_904,N_390,N_174);
and U905 (N_905,N_362,N_49);
nor U906 (N_906,N_21,N_334);
nand U907 (N_907,N_147,N_307);
nand U908 (N_908,N_243,N_366);
nand U909 (N_909,N_398,N_176);
or U910 (N_910,N_344,N_444);
nand U911 (N_911,N_24,N_220);
nor U912 (N_912,N_435,N_69);
and U913 (N_913,N_287,N_81);
or U914 (N_914,N_225,N_464);
nor U915 (N_915,N_283,N_316);
or U916 (N_916,N_459,N_205);
and U917 (N_917,N_366,N_140);
and U918 (N_918,N_416,N_96);
and U919 (N_919,N_292,N_401);
or U920 (N_920,N_46,N_327);
nor U921 (N_921,N_83,N_17);
or U922 (N_922,N_315,N_449);
or U923 (N_923,N_140,N_473);
nand U924 (N_924,N_234,N_258);
nor U925 (N_925,N_122,N_348);
nand U926 (N_926,N_452,N_132);
and U927 (N_927,N_82,N_97);
nand U928 (N_928,N_413,N_153);
or U929 (N_929,N_438,N_59);
nor U930 (N_930,N_30,N_257);
or U931 (N_931,N_350,N_417);
or U932 (N_932,N_198,N_81);
xnor U933 (N_933,N_197,N_485);
or U934 (N_934,N_433,N_98);
nand U935 (N_935,N_49,N_179);
nand U936 (N_936,N_281,N_387);
nor U937 (N_937,N_334,N_458);
and U938 (N_938,N_423,N_324);
and U939 (N_939,N_420,N_101);
nand U940 (N_940,N_91,N_20);
nor U941 (N_941,N_149,N_165);
nand U942 (N_942,N_95,N_350);
nand U943 (N_943,N_397,N_6);
nand U944 (N_944,N_219,N_497);
nor U945 (N_945,N_295,N_1);
and U946 (N_946,N_361,N_362);
and U947 (N_947,N_182,N_426);
and U948 (N_948,N_91,N_43);
nand U949 (N_949,N_261,N_38);
or U950 (N_950,N_428,N_460);
or U951 (N_951,N_375,N_220);
or U952 (N_952,N_448,N_17);
nand U953 (N_953,N_187,N_286);
and U954 (N_954,N_202,N_299);
nand U955 (N_955,N_497,N_406);
and U956 (N_956,N_435,N_346);
nand U957 (N_957,N_23,N_488);
and U958 (N_958,N_334,N_71);
and U959 (N_959,N_260,N_411);
nor U960 (N_960,N_301,N_92);
and U961 (N_961,N_474,N_19);
nand U962 (N_962,N_156,N_92);
or U963 (N_963,N_322,N_251);
and U964 (N_964,N_427,N_486);
or U965 (N_965,N_265,N_280);
and U966 (N_966,N_386,N_327);
nor U967 (N_967,N_166,N_11);
nand U968 (N_968,N_199,N_218);
xnor U969 (N_969,N_183,N_15);
nor U970 (N_970,N_385,N_326);
nand U971 (N_971,N_467,N_124);
nand U972 (N_972,N_357,N_456);
and U973 (N_973,N_277,N_488);
and U974 (N_974,N_435,N_132);
or U975 (N_975,N_496,N_314);
and U976 (N_976,N_160,N_6);
or U977 (N_977,N_223,N_177);
or U978 (N_978,N_128,N_246);
and U979 (N_979,N_411,N_242);
or U980 (N_980,N_306,N_298);
nand U981 (N_981,N_491,N_317);
nor U982 (N_982,N_101,N_413);
nand U983 (N_983,N_285,N_191);
nor U984 (N_984,N_25,N_198);
or U985 (N_985,N_169,N_62);
nand U986 (N_986,N_143,N_380);
nand U987 (N_987,N_405,N_402);
nand U988 (N_988,N_95,N_322);
xnor U989 (N_989,N_278,N_174);
nor U990 (N_990,N_133,N_25);
nor U991 (N_991,N_224,N_87);
and U992 (N_992,N_32,N_122);
nor U993 (N_993,N_62,N_201);
nand U994 (N_994,N_57,N_459);
nor U995 (N_995,N_244,N_280);
nor U996 (N_996,N_184,N_193);
nand U997 (N_997,N_0,N_283);
nand U998 (N_998,N_424,N_318);
nand U999 (N_999,N_107,N_207);
and U1000 (N_1000,N_841,N_522);
nand U1001 (N_1001,N_627,N_687);
and U1002 (N_1002,N_840,N_541);
nand U1003 (N_1003,N_760,N_565);
xor U1004 (N_1004,N_692,N_720);
and U1005 (N_1005,N_726,N_976);
and U1006 (N_1006,N_994,N_543);
nand U1007 (N_1007,N_756,N_701);
or U1008 (N_1008,N_509,N_540);
or U1009 (N_1009,N_733,N_981);
or U1010 (N_1010,N_822,N_659);
and U1011 (N_1011,N_949,N_597);
or U1012 (N_1012,N_859,N_698);
xnor U1013 (N_1013,N_853,N_854);
and U1014 (N_1014,N_860,N_801);
or U1015 (N_1015,N_505,N_915);
and U1016 (N_1016,N_845,N_761);
or U1017 (N_1017,N_521,N_638);
nor U1018 (N_1018,N_717,N_777);
nor U1019 (N_1019,N_803,N_811);
or U1020 (N_1020,N_572,N_616);
nor U1021 (N_1021,N_790,N_930);
and U1022 (N_1022,N_762,N_977);
nor U1023 (N_1023,N_747,N_830);
or U1024 (N_1024,N_635,N_922);
nand U1025 (N_1025,N_598,N_754);
nor U1026 (N_1026,N_675,N_604);
or U1027 (N_1027,N_580,N_856);
or U1028 (N_1028,N_574,N_836);
nor U1029 (N_1029,N_834,N_998);
and U1030 (N_1030,N_558,N_883);
and U1031 (N_1031,N_871,N_719);
nand U1032 (N_1032,N_932,N_723);
nor U1033 (N_1033,N_937,N_559);
nand U1034 (N_1034,N_648,N_991);
or U1035 (N_1035,N_749,N_831);
nor U1036 (N_1036,N_557,N_787);
or U1037 (N_1037,N_795,N_984);
nor U1038 (N_1038,N_561,N_780);
nand U1039 (N_1039,N_870,N_705);
nand U1040 (N_1040,N_781,N_877);
nand U1041 (N_1041,N_944,N_872);
nand U1042 (N_1042,N_958,N_992);
nor U1043 (N_1043,N_775,N_700);
nand U1044 (N_1044,N_511,N_562);
nor U1045 (N_1045,N_904,N_873);
nand U1046 (N_1046,N_900,N_793);
nand U1047 (N_1047,N_925,N_690);
and U1048 (N_1048,N_956,N_953);
and U1049 (N_1049,N_670,N_674);
xor U1050 (N_1050,N_539,N_971);
and U1051 (N_1051,N_528,N_600);
and U1052 (N_1052,N_798,N_544);
nand U1053 (N_1053,N_917,N_907);
nand U1054 (N_1054,N_997,N_709);
or U1055 (N_1055,N_563,N_536);
and U1056 (N_1056,N_879,N_661);
or U1057 (N_1057,N_848,N_750);
and U1058 (N_1058,N_636,N_718);
and U1059 (N_1059,N_752,N_551);
or U1060 (N_1060,N_520,N_812);
or U1061 (N_1061,N_951,N_802);
and U1062 (N_1062,N_874,N_881);
nor U1063 (N_1063,N_913,N_791);
or U1064 (N_1064,N_861,N_927);
nand U1065 (N_1065,N_772,N_818);
nor U1066 (N_1066,N_782,N_855);
or U1067 (N_1067,N_882,N_525);
or U1068 (N_1068,N_919,N_739);
and U1069 (N_1069,N_866,N_898);
nor U1070 (N_1070,N_989,N_758);
nor U1071 (N_1071,N_869,N_685);
nand U1072 (N_1072,N_972,N_553);
or U1073 (N_1073,N_918,N_610);
nor U1074 (N_1074,N_732,N_606);
and U1075 (N_1075,N_846,N_897);
and U1076 (N_1076,N_970,N_625);
and U1077 (N_1077,N_658,N_943);
xor U1078 (N_1078,N_864,N_619);
nand U1079 (N_1079,N_626,N_706);
or U1080 (N_1080,N_755,N_671);
xor U1081 (N_1081,N_714,N_783);
or U1082 (N_1082,N_813,N_697);
nor U1083 (N_1083,N_642,N_929);
or U1084 (N_1084,N_885,N_768);
and U1085 (N_1085,N_906,N_650);
nor U1086 (N_1086,N_693,N_672);
and U1087 (N_1087,N_639,N_974);
nor U1088 (N_1088,N_815,N_605);
and U1089 (N_1089,N_660,N_502);
nand U1090 (N_1090,N_538,N_896);
or U1091 (N_1091,N_570,N_542);
nor U1092 (N_1092,N_529,N_601);
and U1093 (N_1093,N_792,N_684);
nor U1094 (N_1094,N_679,N_503);
nand U1095 (N_1095,N_832,N_603);
and U1096 (N_1096,N_620,N_980);
and U1097 (N_1097,N_647,N_916);
nor U1098 (N_1098,N_590,N_569);
xnor U1099 (N_1099,N_887,N_657);
nand U1100 (N_1100,N_865,N_631);
or U1101 (N_1101,N_910,N_985);
or U1102 (N_1102,N_770,N_725);
or U1103 (N_1103,N_945,N_512);
nand U1104 (N_1104,N_796,N_982);
and U1105 (N_1105,N_568,N_814);
or U1106 (N_1106,N_646,N_545);
nand U1107 (N_1107,N_615,N_708);
or U1108 (N_1108,N_892,N_596);
or U1109 (N_1109,N_948,N_594);
xor U1110 (N_1110,N_537,N_954);
nor U1111 (N_1111,N_893,N_794);
nor U1112 (N_1112,N_595,N_552);
nor U1113 (N_1113,N_621,N_788);
nor U1114 (N_1114,N_583,N_979);
and U1115 (N_1115,N_546,N_547);
or U1116 (N_1116,N_681,N_926);
nand U1117 (N_1117,N_664,N_808);
nor U1118 (N_1118,N_576,N_535);
and U1119 (N_1119,N_727,N_931);
nor U1120 (N_1120,N_765,N_902);
and U1121 (N_1121,N_938,N_899);
and U1122 (N_1122,N_805,N_748);
and U1123 (N_1123,N_886,N_969);
nor U1124 (N_1124,N_644,N_584);
nor U1125 (N_1125,N_680,N_963);
nand U1126 (N_1126,N_513,N_618);
nor U1127 (N_1127,N_995,N_599);
nor U1128 (N_1128,N_908,N_738);
nor U1129 (N_1129,N_530,N_939);
or U1130 (N_1130,N_890,N_524);
nor U1131 (N_1131,N_960,N_878);
nor U1132 (N_1132,N_577,N_843);
and U1133 (N_1133,N_724,N_891);
nor U1134 (N_1134,N_523,N_592);
nand U1135 (N_1135,N_767,N_952);
or U1136 (N_1136,N_663,N_966);
nand U1137 (N_1137,N_689,N_667);
nor U1138 (N_1138,N_909,N_729);
and U1139 (N_1139,N_555,N_716);
or U1140 (N_1140,N_810,N_799);
and U1141 (N_1141,N_757,N_500);
nor U1142 (N_1142,N_515,N_769);
and U1143 (N_1143,N_959,N_571);
or U1144 (N_1144,N_624,N_715);
nor U1145 (N_1145,N_589,N_517);
nor U1146 (N_1146,N_912,N_686);
and U1147 (N_1147,N_819,N_759);
or U1148 (N_1148,N_973,N_779);
and U1149 (N_1149,N_634,N_629);
nand U1150 (N_1150,N_921,N_614);
and U1151 (N_1151,N_746,N_514);
nor U1152 (N_1152,N_827,N_633);
and U1153 (N_1153,N_764,N_607);
nand U1154 (N_1154,N_722,N_695);
nand U1155 (N_1155,N_957,N_823);
nor U1156 (N_1156,N_741,N_628);
or U1157 (N_1157,N_842,N_591);
or U1158 (N_1158,N_532,N_721);
nor U1159 (N_1159,N_911,N_742);
or U1160 (N_1160,N_773,N_850);
or U1161 (N_1161,N_575,N_809);
nand U1162 (N_1162,N_554,N_662);
and U1163 (N_1163,N_751,N_645);
nor U1164 (N_1164,N_829,N_778);
nor U1165 (N_1165,N_987,N_946);
xnor U1166 (N_1166,N_924,N_851);
nor U1167 (N_1167,N_875,N_835);
and U1168 (N_1168,N_582,N_964);
and U1169 (N_1169,N_838,N_655);
nor U1170 (N_1170,N_880,N_578);
and U1171 (N_1171,N_707,N_579);
nand U1172 (N_1172,N_978,N_804);
nand U1173 (N_1173,N_612,N_888);
nor U1174 (N_1174,N_797,N_656);
nand U1175 (N_1175,N_609,N_940);
or U1176 (N_1176,N_863,N_825);
nor U1177 (N_1177,N_766,N_611);
and U1178 (N_1178,N_800,N_699);
nand U1179 (N_1179,N_665,N_683);
and U1180 (N_1180,N_771,N_858);
nor U1181 (N_1181,N_999,N_868);
or U1182 (N_1182,N_730,N_857);
or U1183 (N_1183,N_753,N_519);
and U1184 (N_1184,N_548,N_510);
or U1185 (N_1185,N_833,N_824);
or U1186 (N_1186,N_550,N_955);
and U1187 (N_1187,N_744,N_928);
and U1188 (N_1188,N_731,N_901);
nor U1189 (N_1189,N_965,N_622);
nand U1190 (N_1190,N_507,N_527);
and U1191 (N_1191,N_501,N_867);
nor U1192 (N_1192,N_533,N_852);
nor U1193 (N_1193,N_564,N_942);
and U1194 (N_1194,N_806,N_816);
nor U1195 (N_1195,N_711,N_643);
nand U1196 (N_1196,N_704,N_837);
nor U1197 (N_1197,N_807,N_640);
and U1198 (N_1198,N_673,N_641);
or U1199 (N_1199,N_923,N_933);
nand U1200 (N_1200,N_632,N_993);
and U1201 (N_1201,N_996,N_581);
nand U1202 (N_1202,N_986,N_763);
or U1203 (N_1203,N_920,N_531);
nand U1204 (N_1204,N_821,N_735);
or U1205 (N_1205,N_737,N_566);
or U1206 (N_1206,N_950,N_903);
nor U1207 (N_1207,N_968,N_947);
nor U1208 (N_1208,N_593,N_786);
nand U1209 (N_1209,N_703,N_630);
and U1210 (N_1210,N_676,N_588);
or U1211 (N_1211,N_914,N_962);
nand U1212 (N_1212,N_666,N_740);
and U1213 (N_1213,N_560,N_817);
nand U1214 (N_1214,N_862,N_573);
and U1215 (N_1215,N_884,N_934);
or U1216 (N_1216,N_696,N_668);
nand U1217 (N_1217,N_691,N_587);
or U1218 (N_1218,N_549,N_710);
or U1219 (N_1219,N_669,N_975);
xor U1220 (N_1220,N_876,N_905);
and U1221 (N_1221,N_774,N_608);
nand U1222 (N_1222,N_734,N_847);
nor U1223 (N_1223,N_988,N_826);
and U1224 (N_1224,N_623,N_516);
nor U1225 (N_1225,N_567,N_526);
and U1226 (N_1226,N_789,N_990);
and U1227 (N_1227,N_702,N_534);
nor U1228 (N_1228,N_776,N_586);
and U1229 (N_1229,N_743,N_895);
nor U1230 (N_1230,N_694,N_652);
nor U1231 (N_1231,N_518,N_712);
and U1232 (N_1232,N_820,N_936);
or U1233 (N_1233,N_983,N_967);
and U1234 (N_1234,N_784,N_894);
nand U1235 (N_1235,N_935,N_651);
and U1236 (N_1236,N_613,N_828);
xor U1237 (N_1237,N_649,N_682);
and U1238 (N_1238,N_688,N_889);
and U1239 (N_1239,N_736,N_713);
nor U1240 (N_1240,N_602,N_745);
nor U1241 (N_1241,N_504,N_654);
nor U1242 (N_1242,N_941,N_839);
or U1243 (N_1243,N_506,N_637);
or U1244 (N_1244,N_653,N_785);
or U1245 (N_1245,N_508,N_961);
and U1246 (N_1246,N_678,N_677);
and U1247 (N_1247,N_556,N_728);
and U1248 (N_1248,N_849,N_617);
xnor U1249 (N_1249,N_844,N_585);
or U1250 (N_1250,N_774,N_671);
or U1251 (N_1251,N_837,N_848);
nand U1252 (N_1252,N_941,N_821);
or U1253 (N_1253,N_826,N_526);
nand U1254 (N_1254,N_618,N_816);
and U1255 (N_1255,N_814,N_949);
or U1256 (N_1256,N_658,N_981);
nand U1257 (N_1257,N_962,N_660);
xnor U1258 (N_1258,N_696,N_955);
nand U1259 (N_1259,N_614,N_637);
nand U1260 (N_1260,N_655,N_551);
nor U1261 (N_1261,N_561,N_530);
and U1262 (N_1262,N_772,N_689);
or U1263 (N_1263,N_613,N_592);
nand U1264 (N_1264,N_753,N_633);
nand U1265 (N_1265,N_646,N_845);
nand U1266 (N_1266,N_789,N_646);
or U1267 (N_1267,N_637,N_740);
or U1268 (N_1268,N_670,N_731);
nand U1269 (N_1269,N_563,N_739);
or U1270 (N_1270,N_693,N_807);
xor U1271 (N_1271,N_623,N_530);
or U1272 (N_1272,N_954,N_612);
and U1273 (N_1273,N_691,N_542);
nand U1274 (N_1274,N_553,N_827);
nor U1275 (N_1275,N_689,N_709);
or U1276 (N_1276,N_810,N_934);
nor U1277 (N_1277,N_774,N_685);
nor U1278 (N_1278,N_697,N_775);
and U1279 (N_1279,N_854,N_742);
and U1280 (N_1280,N_796,N_503);
nand U1281 (N_1281,N_569,N_789);
nand U1282 (N_1282,N_888,N_637);
nand U1283 (N_1283,N_652,N_856);
or U1284 (N_1284,N_709,N_599);
or U1285 (N_1285,N_992,N_675);
and U1286 (N_1286,N_869,N_820);
and U1287 (N_1287,N_737,N_574);
and U1288 (N_1288,N_961,N_918);
and U1289 (N_1289,N_810,N_961);
nor U1290 (N_1290,N_874,N_787);
nor U1291 (N_1291,N_889,N_602);
nor U1292 (N_1292,N_620,N_628);
nand U1293 (N_1293,N_700,N_763);
nand U1294 (N_1294,N_560,N_709);
nand U1295 (N_1295,N_659,N_739);
or U1296 (N_1296,N_850,N_514);
xor U1297 (N_1297,N_673,N_930);
or U1298 (N_1298,N_764,N_901);
or U1299 (N_1299,N_825,N_616);
nand U1300 (N_1300,N_567,N_589);
nand U1301 (N_1301,N_881,N_923);
and U1302 (N_1302,N_989,N_890);
nand U1303 (N_1303,N_820,N_990);
nand U1304 (N_1304,N_503,N_752);
nor U1305 (N_1305,N_852,N_999);
nor U1306 (N_1306,N_786,N_978);
nor U1307 (N_1307,N_814,N_817);
nor U1308 (N_1308,N_693,N_866);
nor U1309 (N_1309,N_780,N_987);
and U1310 (N_1310,N_953,N_569);
nor U1311 (N_1311,N_703,N_850);
and U1312 (N_1312,N_538,N_852);
nor U1313 (N_1313,N_548,N_511);
or U1314 (N_1314,N_965,N_779);
or U1315 (N_1315,N_519,N_678);
or U1316 (N_1316,N_565,N_654);
or U1317 (N_1317,N_894,N_762);
nand U1318 (N_1318,N_687,N_876);
or U1319 (N_1319,N_846,N_639);
or U1320 (N_1320,N_526,N_708);
and U1321 (N_1321,N_559,N_936);
and U1322 (N_1322,N_641,N_756);
nand U1323 (N_1323,N_938,N_839);
or U1324 (N_1324,N_882,N_605);
or U1325 (N_1325,N_590,N_748);
or U1326 (N_1326,N_635,N_766);
nor U1327 (N_1327,N_574,N_573);
and U1328 (N_1328,N_674,N_662);
or U1329 (N_1329,N_992,N_956);
or U1330 (N_1330,N_710,N_886);
nor U1331 (N_1331,N_947,N_551);
nand U1332 (N_1332,N_566,N_959);
or U1333 (N_1333,N_584,N_585);
nand U1334 (N_1334,N_582,N_911);
or U1335 (N_1335,N_504,N_891);
nand U1336 (N_1336,N_976,N_632);
and U1337 (N_1337,N_858,N_595);
nand U1338 (N_1338,N_963,N_774);
nand U1339 (N_1339,N_835,N_770);
nand U1340 (N_1340,N_734,N_914);
and U1341 (N_1341,N_571,N_531);
nor U1342 (N_1342,N_787,N_956);
or U1343 (N_1343,N_533,N_847);
or U1344 (N_1344,N_750,N_795);
nand U1345 (N_1345,N_538,N_634);
nor U1346 (N_1346,N_996,N_820);
or U1347 (N_1347,N_850,N_867);
nand U1348 (N_1348,N_617,N_872);
nor U1349 (N_1349,N_957,N_866);
and U1350 (N_1350,N_750,N_606);
nand U1351 (N_1351,N_500,N_961);
nand U1352 (N_1352,N_863,N_868);
and U1353 (N_1353,N_573,N_944);
nand U1354 (N_1354,N_766,N_907);
nor U1355 (N_1355,N_953,N_776);
and U1356 (N_1356,N_656,N_809);
or U1357 (N_1357,N_857,N_704);
nand U1358 (N_1358,N_655,N_672);
nor U1359 (N_1359,N_844,N_863);
nand U1360 (N_1360,N_733,N_668);
nor U1361 (N_1361,N_579,N_620);
nand U1362 (N_1362,N_539,N_503);
nand U1363 (N_1363,N_788,N_950);
and U1364 (N_1364,N_903,N_650);
nand U1365 (N_1365,N_817,N_828);
nor U1366 (N_1366,N_681,N_996);
nand U1367 (N_1367,N_666,N_811);
xor U1368 (N_1368,N_666,N_577);
nor U1369 (N_1369,N_562,N_720);
or U1370 (N_1370,N_821,N_654);
or U1371 (N_1371,N_568,N_620);
or U1372 (N_1372,N_946,N_709);
or U1373 (N_1373,N_993,N_587);
nand U1374 (N_1374,N_895,N_842);
or U1375 (N_1375,N_922,N_535);
or U1376 (N_1376,N_583,N_735);
nand U1377 (N_1377,N_650,N_622);
nand U1378 (N_1378,N_987,N_707);
nor U1379 (N_1379,N_778,N_944);
nor U1380 (N_1380,N_831,N_785);
and U1381 (N_1381,N_535,N_929);
nand U1382 (N_1382,N_641,N_740);
nand U1383 (N_1383,N_860,N_663);
and U1384 (N_1384,N_654,N_572);
or U1385 (N_1385,N_991,N_773);
nand U1386 (N_1386,N_512,N_637);
and U1387 (N_1387,N_679,N_602);
nand U1388 (N_1388,N_524,N_810);
nor U1389 (N_1389,N_785,N_547);
and U1390 (N_1390,N_708,N_935);
and U1391 (N_1391,N_992,N_761);
nand U1392 (N_1392,N_841,N_687);
nand U1393 (N_1393,N_768,N_787);
nor U1394 (N_1394,N_919,N_903);
or U1395 (N_1395,N_514,N_918);
nor U1396 (N_1396,N_960,N_787);
or U1397 (N_1397,N_628,N_972);
nor U1398 (N_1398,N_770,N_951);
nor U1399 (N_1399,N_535,N_689);
nor U1400 (N_1400,N_987,N_889);
and U1401 (N_1401,N_951,N_810);
and U1402 (N_1402,N_532,N_568);
nor U1403 (N_1403,N_673,N_745);
or U1404 (N_1404,N_999,N_640);
nor U1405 (N_1405,N_731,N_677);
nand U1406 (N_1406,N_817,N_835);
nor U1407 (N_1407,N_994,N_659);
and U1408 (N_1408,N_695,N_890);
nor U1409 (N_1409,N_808,N_910);
nor U1410 (N_1410,N_564,N_849);
nor U1411 (N_1411,N_655,N_698);
and U1412 (N_1412,N_561,N_540);
and U1413 (N_1413,N_755,N_894);
nand U1414 (N_1414,N_577,N_764);
and U1415 (N_1415,N_745,N_792);
nor U1416 (N_1416,N_920,N_912);
or U1417 (N_1417,N_626,N_621);
or U1418 (N_1418,N_572,N_820);
nand U1419 (N_1419,N_701,N_824);
nor U1420 (N_1420,N_669,N_777);
and U1421 (N_1421,N_872,N_948);
and U1422 (N_1422,N_505,N_796);
or U1423 (N_1423,N_915,N_680);
or U1424 (N_1424,N_800,N_738);
and U1425 (N_1425,N_858,N_870);
or U1426 (N_1426,N_979,N_917);
and U1427 (N_1427,N_825,N_787);
and U1428 (N_1428,N_989,N_603);
and U1429 (N_1429,N_705,N_605);
or U1430 (N_1430,N_760,N_709);
and U1431 (N_1431,N_884,N_787);
or U1432 (N_1432,N_970,N_566);
nand U1433 (N_1433,N_893,N_782);
nand U1434 (N_1434,N_723,N_607);
and U1435 (N_1435,N_694,N_679);
nand U1436 (N_1436,N_919,N_984);
and U1437 (N_1437,N_718,N_720);
nand U1438 (N_1438,N_752,N_652);
or U1439 (N_1439,N_919,N_752);
nand U1440 (N_1440,N_913,N_622);
or U1441 (N_1441,N_546,N_600);
nor U1442 (N_1442,N_951,N_878);
nand U1443 (N_1443,N_773,N_849);
nand U1444 (N_1444,N_800,N_589);
nor U1445 (N_1445,N_754,N_681);
or U1446 (N_1446,N_796,N_777);
and U1447 (N_1447,N_809,N_985);
nor U1448 (N_1448,N_887,N_652);
nand U1449 (N_1449,N_753,N_601);
or U1450 (N_1450,N_842,N_833);
or U1451 (N_1451,N_891,N_769);
and U1452 (N_1452,N_663,N_856);
nand U1453 (N_1453,N_578,N_543);
nor U1454 (N_1454,N_931,N_590);
nand U1455 (N_1455,N_808,N_659);
or U1456 (N_1456,N_696,N_673);
or U1457 (N_1457,N_746,N_899);
xor U1458 (N_1458,N_850,N_892);
and U1459 (N_1459,N_892,N_934);
nand U1460 (N_1460,N_798,N_845);
nand U1461 (N_1461,N_673,N_560);
or U1462 (N_1462,N_928,N_899);
or U1463 (N_1463,N_918,N_756);
nand U1464 (N_1464,N_819,N_622);
nor U1465 (N_1465,N_614,N_594);
or U1466 (N_1466,N_707,N_730);
or U1467 (N_1467,N_971,N_682);
and U1468 (N_1468,N_870,N_799);
nand U1469 (N_1469,N_761,N_544);
or U1470 (N_1470,N_900,N_506);
or U1471 (N_1471,N_705,N_699);
nor U1472 (N_1472,N_869,N_688);
nor U1473 (N_1473,N_833,N_552);
nand U1474 (N_1474,N_930,N_651);
nor U1475 (N_1475,N_882,N_657);
nand U1476 (N_1476,N_816,N_516);
and U1477 (N_1477,N_652,N_699);
or U1478 (N_1478,N_713,N_686);
xnor U1479 (N_1479,N_751,N_915);
nand U1480 (N_1480,N_686,N_880);
nor U1481 (N_1481,N_903,N_982);
and U1482 (N_1482,N_752,N_533);
nor U1483 (N_1483,N_886,N_855);
nand U1484 (N_1484,N_762,N_516);
nor U1485 (N_1485,N_710,N_558);
or U1486 (N_1486,N_921,N_888);
or U1487 (N_1487,N_748,N_963);
nor U1488 (N_1488,N_831,N_733);
or U1489 (N_1489,N_581,N_874);
nor U1490 (N_1490,N_678,N_522);
nand U1491 (N_1491,N_532,N_853);
or U1492 (N_1492,N_706,N_622);
or U1493 (N_1493,N_504,N_918);
nor U1494 (N_1494,N_781,N_508);
and U1495 (N_1495,N_912,N_726);
nor U1496 (N_1496,N_867,N_815);
nor U1497 (N_1497,N_744,N_722);
nor U1498 (N_1498,N_706,N_969);
or U1499 (N_1499,N_888,N_802);
and U1500 (N_1500,N_1151,N_1112);
or U1501 (N_1501,N_1127,N_1173);
nand U1502 (N_1502,N_1291,N_1322);
or U1503 (N_1503,N_1286,N_1194);
nand U1504 (N_1504,N_1013,N_1165);
or U1505 (N_1505,N_1202,N_1155);
and U1506 (N_1506,N_1206,N_1083);
or U1507 (N_1507,N_1279,N_1265);
and U1508 (N_1508,N_1087,N_1189);
nand U1509 (N_1509,N_1191,N_1253);
or U1510 (N_1510,N_1409,N_1049);
nand U1511 (N_1511,N_1116,N_1019);
nor U1512 (N_1512,N_1042,N_1388);
and U1513 (N_1513,N_1306,N_1426);
and U1514 (N_1514,N_1115,N_1425);
nand U1515 (N_1515,N_1093,N_1382);
nand U1516 (N_1516,N_1031,N_1335);
and U1517 (N_1517,N_1256,N_1104);
or U1518 (N_1518,N_1328,N_1102);
nor U1519 (N_1519,N_1287,N_1456);
nor U1520 (N_1520,N_1177,N_1479);
nand U1521 (N_1521,N_1150,N_1313);
nor U1522 (N_1522,N_1169,N_1493);
nor U1523 (N_1523,N_1403,N_1252);
nand U1524 (N_1524,N_1167,N_1468);
xor U1525 (N_1525,N_1098,N_1489);
nor U1526 (N_1526,N_1117,N_1412);
nor U1527 (N_1527,N_1298,N_1204);
nand U1528 (N_1528,N_1354,N_1084);
and U1529 (N_1529,N_1273,N_1038);
nand U1530 (N_1530,N_1436,N_1028);
and U1531 (N_1531,N_1453,N_1339);
nand U1532 (N_1532,N_1334,N_1366);
and U1533 (N_1533,N_1471,N_1132);
nor U1534 (N_1534,N_1367,N_1076);
or U1535 (N_1535,N_1289,N_1159);
nand U1536 (N_1536,N_1103,N_1091);
nand U1537 (N_1537,N_1037,N_1090);
nand U1538 (N_1538,N_1374,N_1386);
nor U1539 (N_1539,N_1362,N_1119);
nor U1540 (N_1540,N_1363,N_1148);
nand U1541 (N_1541,N_1373,N_1276);
or U1542 (N_1542,N_1293,N_1187);
nor U1543 (N_1543,N_1008,N_1250);
or U1544 (N_1544,N_1251,N_1432);
nand U1545 (N_1545,N_1075,N_1133);
and U1546 (N_1546,N_1050,N_1303);
nor U1547 (N_1547,N_1405,N_1211);
and U1548 (N_1548,N_1469,N_1442);
and U1549 (N_1549,N_1413,N_1480);
and U1550 (N_1550,N_1094,N_1497);
nand U1551 (N_1551,N_1059,N_1141);
and U1552 (N_1552,N_1264,N_1437);
nor U1553 (N_1553,N_1427,N_1027);
and U1554 (N_1554,N_1284,N_1066);
nor U1555 (N_1555,N_1327,N_1079);
nor U1556 (N_1556,N_1240,N_1099);
and U1557 (N_1557,N_1229,N_1188);
and U1558 (N_1558,N_1353,N_1072);
or U1559 (N_1559,N_1356,N_1183);
and U1560 (N_1560,N_1496,N_1402);
nand U1561 (N_1561,N_1491,N_1419);
nor U1562 (N_1562,N_1452,N_1054);
nand U1563 (N_1563,N_1011,N_1325);
or U1564 (N_1564,N_1417,N_1305);
or U1565 (N_1565,N_1010,N_1434);
xnor U1566 (N_1566,N_1137,N_1156);
nand U1567 (N_1567,N_1473,N_1035);
nor U1568 (N_1568,N_1036,N_1213);
and U1569 (N_1569,N_1394,N_1120);
nand U1570 (N_1570,N_1359,N_1002);
xor U1571 (N_1571,N_1044,N_1218);
or U1572 (N_1572,N_1121,N_1448);
nor U1573 (N_1573,N_1166,N_1351);
or U1574 (N_1574,N_1267,N_1431);
or U1575 (N_1575,N_1312,N_1435);
nand U1576 (N_1576,N_1455,N_1336);
and U1577 (N_1577,N_1361,N_1107);
and U1578 (N_1578,N_1263,N_1170);
nor U1579 (N_1579,N_1332,N_1345);
and U1580 (N_1580,N_1193,N_1288);
or U1581 (N_1581,N_1467,N_1309);
and U1582 (N_1582,N_1350,N_1421);
or U1583 (N_1583,N_1294,N_1228);
nor U1584 (N_1584,N_1317,N_1182);
nor U1585 (N_1585,N_1341,N_1062);
nand U1586 (N_1586,N_1022,N_1108);
nor U1587 (N_1587,N_1389,N_1122);
nand U1588 (N_1588,N_1061,N_1329);
or U1589 (N_1589,N_1067,N_1360);
nand U1590 (N_1590,N_1478,N_1352);
nand U1591 (N_1591,N_1430,N_1343);
nor U1592 (N_1592,N_1198,N_1201);
nand U1593 (N_1593,N_1068,N_1423);
or U1594 (N_1594,N_1477,N_1315);
or U1595 (N_1595,N_1375,N_1368);
or U1596 (N_1596,N_1138,N_1307);
or U1597 (N_1597,N_1385,N_1499);
nand U1598 (N_1598,N_1472,N_1239);
and U1599 (N_1599,N_1406,N_1451);
nor U1600 (N_1600,N_1438,N_1227);
nor U1601 (N_1601,N_1040,N_1454);
or U1602 (N_1602,N_1106,N_1268);
and U1603 (N_1603,N_1494,N_1407);
and U1604 (N_1604,N_1290,N_1255);
and U1605 (N_1605,N_1249,N_1172);
and U1606 (N_1606,N_1383,N_1270);
nor U1607 (N_1607,N_1021,N_1408);
and U1608 (N_1608,N_1134,N_1297);
nand U1609 (N_1609,N_1258,N_1462);
nand U1610 (N_1610,N_1377,N_1179);
nand U1611 (N_1611,N_1387,N_1016);
nor U1612 (N_1612,N_1285,N_1178);
nand U1613 (N_1613,N_1358,N_1143);
nand U1614 (N_1614,N_1124,N_1277);
or U1615 (N_1615,N_1214,N_1278);
nand U1616 (N_1616,N_1039,N_1445);
nand U1617 (N_1617,N_1126,N_1081);
nand U1618 (N_1618,N_1295,N_1308);
nor U1619 (N_1619,N_1200,N_1244);
nor U1620 (N_1620,N_1418,N_1129);
or U1621 (N_1621,N_1230,N_1197);
and U1622 (N_1622,N_1057,N_1144);
nand U1623 (N_1623,N_1007,N_1488);
or U1624 (N_1624,N_1260,N_1242);
or U1625 (N_1625,N_1147,N_1004);
or U1626 (N_1626,N_1071,N_1415);
or U1627 (N_1627,N_1280,N_1225);
or U1628 (N_1628,N_1433,N_1272);
and U1629 (N_1629,N_1410,N_1347);
or U1630 (N_1630,N_1089,N_1158);
nor U1631 (N_1631,N_1444,N_1145);
nand U1632 (N_1632,N_1236,N_1365);
nand U1633 (N_1633,N_1020,N_1181);
and U1634 (N_1634,N_1396,N_1034);
or U1635 (N_1635,N_1461,N_1458);
or U1636 (N_1636,N_1047,N_1123);
or U1637 (N_1637,N_1370,N_1301);
xor U1638 (N_1638,N_1033,N_1395);
nand U1639 (N_1639,N_1208,N_1215);
or U1640 (N_1640,N_1248,N_1196);
nor U1641 (N_1641,N_1259,N_1243);
nand U1642 (N_1642,N_1466,N_1205);
nand U1643 (N_1643,N_1391,N_1069);
nand U1644 (N_1644,N_1238,N_1065);
or U1645 (N_1645,N_1078,N_1321);
and U1646 (N_1646,N_1490,N_1207);
nand U1647 (N_1647,N_1416,N_1160);
and U1648 (N_1648,N_1209,N_1046);
or U1649 (N_1649,N_1299,N_1338);
nand U1650 (N_1650,N_1149,N_1055);
or U1651 (N_1651,N_1131,N_1185);
nand U1652 (N_1652,N_1355,N_1443);
xnor U1653 (N_1653,N_1223,N_1018);
nor U1654 (N_1654,N_1222,N_1136);
nand U1655 (N_1655,N_1097,N_1369);
or U1656 (N_1656,N_1045,N_1146);
and U1657 (N_1657,N_1485,N_1446);
nand U1658 (N_1658,N_1135,N_1326);
or U1659 (N_1659,N_1224,N_1399);
nor U1660 (N_1660,N_1269,N_1281);
nand U1661 (N_1661,N_1379,N_1171);
or U1662 (N_1662,N_1457,N_1153);
and U1663 (N_1663,N_1095,N_1157);
nor U1664 (N_1664,N_1051,N_1475);
or U1665 (N_1665,N_1371,N_1195);
nor U1666 (N_1666,N_1470,N_1492);
and U1667 (N_1667,N_1261,N_1245);
and U1668 (N_1668,N_1113,N_1364);
nor U1669 (N_1669,N_1237,N_1476);
or U1670 (N_1670,N_1012,N_1246);
and U1671 (N_1671,N_1184,N_1221);
and U1672 (N_1672,N_1232,N_1411);
nand U1673 (N_1673,N_1052,N_1310);
and U1674 (N_1674,N_1398,N_1003);
nor U1675 (N_1675,N_1422,N_1486);
and U1676 (N_1676,N_1319,N_1381);
nor U1677 (N_1677,N_1210,N_1026);
nor U1678 (N_1678,N_1392,N_1043);
nor U1679 (N_1679,N_1015,N_1447);
nand U1680 (N_1680,N_1053,N_1266);
and U1681 (N_1681,N_1233,N_1304);
nor U1682 (N_1682,N_1041,N_1283);
or U1683 (N_1683,N_1154,N_1254);
nand U1684 (N_1684,N_1125,N_1346);
nand U1685 (N_1685,N_1064,N_1247);
nand U1686 (N_1686,N_1302,N_1024);
and U1687 (N_1687,N_1096,N_1176);
nand U1688 (N_1688,N_1384,N_1088);
nand U1689 (N_1689,N_1174,N_1393);
nor U1690 (N_1690,N_1161,N_1058);
nor U1691 (N_1691,N_1017,N_1186);
and U1692 (N_1692,N_1009,N_1073);
or U1693 (N_1693,N_1048,N_1463);
or U1694 (N_1694,N_1348,N_1140);
nor U1695 (N_1695,N_1400,N_1077);
or U1696 (N_1696,N_1282,N_1219);
and U1697 (N_1697,N_1152,N_1085);
and U1698 (N_1698,N_1275,N_1163);
nor U1699 (N_1699,N_1056,N_1231);
nand U1700 (N_1700,N_1001,N_1128);
and U1701 (N_1701,N_1111,N_1320);
nor U1702 (N_1702,N_1440,N_1380);
nor U1703 (N_1703,N_1226,N_1404);
or U1704 (N_1704,N_1234,N_1235);
nand U1705 (N_1705,N_1450,N_1005);
and U1706 (N_1706,N_1192,N_1428);
nor U1707 (N_1707,N_1372,N_1401);
nor U1708 (N_1708,N_1217,N_1331);
and U1709 (N_1709,N_1439,N_1316);
nor U1710 (N_1710,N_1481,N_1324);
nand U1711 (N_1711,N_1357,N_1271);
nor U1712 (N_1712,N_1474,N_1130);
or U1713 (N_1713,N_1063,N_1030);
nand U1714 (N_1714,N_1212,N_1257);
nand U1715 (N_1715,N_1484,N_1029);
or U1716 (N_1716,N_1070,N_1318);
nor U1717 (N_1717,N_1216,N_1142);
nand U1718 (N_1718,N_1241,N_1168);
nor U1719 (N_1719,N_1220,N_1086);
nand U1720 (N_1720,N_1376,N_1390);
nor U1721 (N_1721,N_1300,N_1465);
and U1722 (N_1722,N_1109,N_1420);
and U1723 (N_1723,N_1100,N_1495);
and U1724 (N_1724,N_1162,N_1311);
nor U1725 (N_1725,N_1092,N_1203);
nor U1726 (N_1726,N_1274,N_1424);
nand U1727 (N_1727,N_1342,N_1429);
nor U1728 (N_1728,N_1118,N_1482);
nand U1729 (N_1729,N_1340,N_1314);
or U1730 (N_1730,N_1397,N_1082);
and U1731 (N_1731,N_1139,N_1014);
nand U1732 (N_1732,N_1378,N_1074);
xnor U1733 (N_1733,N_1344,N_1483);
or U1734 (N_1734,N_1449,N_1414);
nor U1735 (N_1735,N_1349,N_1023);
or U1736 (N_1736,N_1296,N_1180);
and U1737 (N_1737,N_1498,N_1441);
nand U1738 (N_1738,N_1460,N_1000);
and U1739 (N_1739,N_1292,N_1105);
nand U1740 (N_1740,N_1101,N_1164);
or U1741 (N_1741,N_1330,N_1175);
nor U1742 (N_1742,N_1110,N_1262);
or U1743 (N_1743,N_1060,N_1114);
or U1744 (N_1744,N_1032,N_1199);
nor U1745 (N_1745,N_1337,N_1190);
nand U1746 (N_1746,N_1006,N_1464);
and U1747 (N_1747,N_1025,N_1459);
nor U1748 (N_1748,N_1333,N_1487);
or U1749 (N_1749,N_1080,N_1323);
or U1750 (N_1750,N_1215,N_1105);
nor U1751 (N_1751,N_1197,N_1425);
or U1752 (N_1752,N_1229,N_1386);
and U1753 (N_1753,N_1212,N_1431);
and U1754 (N_1754,N_1290,N_1090);
or U1755 (N_1755,N_1355,N_1136);
nand U1756 (N_1756,N_1253,N_1089);
and U1757 (N_1757,N_1301,N_1226);
or U1758 (N_1758,N_1101,N_1383);
and U1759 (N_1759,N_1061,N_1195);
nand U1760 (N_1760,N_1121,N_1262);
nor U1761 (N_1761,N_1316,N_1485);
or U1762 (N_1762,N_1101,N_1232);
nor U1763 (N_1763,N_1223,N_1100);
and U1764 (N_1764,N_1140,N_1178);
nor U1765 (N_1765,N_1393,N_1242);
nor U1766 (N_1766,N_1024,N_1159);
and U1767 (N_1767,N_1123,N_1187);
xnor U1768 (N_1768,N_1045,N_1399);
nand U1769 (N_1769,N_1412,N_1002);
and U1770 (N_1770,N_1480,N_1463);
xor U1771 (N_1771,N_1367,N_1040);
or U1772 (N_1772,N_1051,N_1153);
or U1773 (N_1773,N_1164,N_1044);
nand U1774 (N_1774,N_1239,N_1036);
nand U1775 (N_1775,N_1096,N_1373);
nor U1776 (N_1776,N_1296,N_1343);
nor U1777 (N_1777,N_1273,N_1229);
nand U1778 (N_1778,N_1465,N_1091);
and U1779 (N_1779,N_1463,N_1136);
or U1780 (N_1780,N_1181,N_1372);
nand U1781 (N_1781,N_1493,N_1217);
and U1782 (N_1782,N_1455,N_1429);
and U1783 (N_1783,N_1003,N_1334);
and U1784 (N_1784,N_1490,N_1031);
or U1785 (N_1785,N_1272,N_1392);
and U1786 (N_1786,N_1339,N_1361);
xor U1787 (N_1787,N_1465,N_1138);
nand U1788 (N_1788,N_1324,N_1143);
nand U1789 (N_1789,N_1387,N_1078);
nand U1790 (N_1790,N_1180,N_1492);
nand U1791 (N_1791,N_1041,N_1236);
and U1792 (N_1792,N_1177,N_1317);
nor U1793 (N_1793,N_1083,N_1241);
nor U1794 (N_1794,N_1038,N_1179);
or U1795 (N_1795,N_1340,N_1172);
or U1796 (N_1796,N_1044,N_1075);
nor U1797 (N_1797,N_1021,N_1298);
nor U1798 (N_1798,N_1478,N_1350);
nor U1799 (N_1799,N_1282,N_1036);
and U1800 (N_1800,N_1275,N_1412);
nand U1801 (N_1801,N_1285,N_1139);
nand U1802 (N_1802,N_1490,N_1323);
nand U1803 (N_1803,N_1103,N_1304);
or U1804 (N_1804,N_1221,N_1078);
and U1805 (N_1805,N_1078,N_1237);
and U1806 (N_1806,N_1380,N_1026);
nand U1807 (N_1807,N_1410,N_1108);
and U1808 (N_1808,N_1274,N_1013);
nand U1809 (N_1809,N_1082,N_1317);
or U1810 (N_1810,N_1424,N_1081);
nand U1811 (N_1811,N_1139,N_1422);
nand U1812 (N_1812,N_1219,N_1052);
and U1813 (N_1813,N_1399,N_1109);
nand U1814 (N_1814,N_1189,N_1187);
nand U1815 (N_1815,N_1463,N_1188);
and U1816 (N_1816,N_1413,N_1460);
or U1817 (N_1817,N_1373,N_1278);
nor U1818 (N_1818,N_1047,N_1133);
nand U1819 (N_1819,N_1448,N_1253);
or U1820 (N_1820,N_1281,N_1378);
nand U1821 (N_1821,N_1068,N_1241);
or U1822 (N_1822,N_1002,N_1365);
nor U1823 (N_1823,N_1146,N_1455);
nand U1824 (N_1824,N_1055,N_1218);
nand U1825 (N_1825,N_1308,N_1129);
and U1826 (N_1826,N_1305,N_1034);
and U1827 (N_1827,N_1218,N_1402);
nand U1828 (N_1828,N_1152,N_1145);
or U1829 (N_1829,N_1074,N_1293);
and U1830 (N_1830,N_1019,N_1409);
nor U1831 (N_1831,N_1097,N_1126);
and U1832 (N_1832,N_1135,N_1136);
nand U1833 (N_1833,N_1285,N_1397);
or U1834 (N_1834,N_1124,N_1123);
or U1835 (N_1835,N_1328,N_1106);
or U1836 (N_1836,N_1290,N_1286);
or U1837 (N_1837,N_1258,N_1224);
and U1838 (N_1838,N_1401,N_1034);
nor U1839 (N_1839,N_1480,N_1179);
nand U1840 (N_1840,N_1228,N_1072);
nor U1841 (N_1841,N_1295,N_1337);
nor U1842 (N_1842,N_1322,N_1268);
or U1843 (N_1843,N_1269,N_1307);
and U1844 (N_1844,N_1479,N_1387);
nor U1845 (N_1845,N_1365,N_1216);
nor U1846 (N_1846,N_1150,N_1328);
xor U1847 (N_1847,N_1140,N_1043);
nand U1848 (N_1848,N_1098,N_1476);
or U1849 (N_1849,N_1425,N_1160);
nor U1850 (N_1850,N_1378,N_1235);
and U1851 (N_1851,N_1034,N_1130);
and U1852 (N_1852,N_1181,N_1461);
and U1853 (N_1853,N_1440,N_1491);
xnor U1854 (N_1854,N_1034,N_1432);
nor U1855 (N_1855,N_1073,N_1016);
nand U1856 (N_1856,N_1228,N_1459);
or U1857 (N_1857,N_1278,N_1138);
or U1858 (N_1858,N_1296,N_1431);
nand U1859 (N_1859,N_1218,N_1098);
nor U1860 (N_1860,N_1275,N_1055);
nand U1861 (N_1861,N_1188,N_1314);
nor U1862 (N_1862,N_1258,N_1467);
or U1863 (N_1863,N_1072,N_1427);
and U1864 (N_1864,N_1401,N_1115);
and U1865 (N_1865,N_1424,N_1242);
nand U1866 (N_1866,N_1372,N_1036);
nor U1867 (N_1867,N_1029,N_1302);
or U1868 (N_1868,N_1072,N_1089);
nand U1869 (N_1869,N_1204,N_1040);
nor U1870 (N_1870,N_1308,N_1111);
nand U1871 (N_1871,N_1201,N_1120);
or U1872 (N_1872,N_1174,N_1372);
nor U1873 (N_1873,N_1030,N_1406);
nand U1874 (N_1874,N_1429,N_1272);
and U1875 (N_1875,N_1081,N_1456);
nand U1876 (N_1876,N_1316,N_1317);
nor U1877 (N_1877,N_1459,N_1468);
or U1878 (N_1878,N_1113,N_1289);
and U1879 (N_1879,N_1482,N_1018);
nor U1880 (N_1880,N_1230,N_1150);
nor U1881 (N_1881,N_1183,N_1412);
and U1882 (N_1882,N_1313,N_1289);
and U1883 (N_1883,N_1018,N_1015);
nor U1884 (N_1884,N_1285,N_1028);
nor U1885 (N_1885,N_1182,N_1152);
xnor U1886 (N_1886,N_1304,N_1203);
and U1887 (N_1887,N_1444,N_1296);
and U1888 (N_1888,N_1301,N_1211);
nand U1889 (N_1889,N_1463,N_1225);
nand U1890 (N_1890,N_1108,N_1221);
or U1891 (N_1891,N_1429,N_1215);
nand U1892 (N_1892,N_1406,N_1469);
nand U1893 (N_1893,N_1209,N_1179);
and U1894 (N_1894,N_1195,N_1425);
nor U1895 (N_1895,N_1245,N_1277);
nand U1896 (N_1896,N_1353,N_1306);
nand U1897 (N_1897,N_1434,N_1166);
nor U1898 (N_1898,N_1284,N_1125);
or U1899 (N_1899,N_1430,N_1301);
xnor U1900 (N_1900,N_1280,N_1350);
and U1901 (N_1901,N_1452,N_1294);
nor U1902 (N_1902,N_1457,N_1002);
nor U1903 (N_1903,N_1367,N_1056);
nor U1904 (N_1904,N_1016,N_1393);
or U1905 (N_1905,N_1121,N_1068);
or U1906 (N_1906,N_1052,N_1140);
or U1907 (N_1907,N_1282,N_1486);
and U1908 (N_1908,N_1016,N_1414);
nand U1909 (N_1909,N_1105,N_1107);
nor U1910 (N_1910,N_1161,N_1302);
nor U1911 (N_1911,N_1122,N_1339);
and U1912 (N_1912,N_1047,N_1300);
or U1913 (N_1913,N_1306,N_1472);
nor U1914 (N_1914,N_1205,N_1048);
and U1915 (N_1915,N_1331,N_1397);
and U1916 (N_1916,N_1408,N_1437);
nor U1917 (N_1917,N_1346,N_1271);
and U1918 (N_1918,N_1483,N_1463);
nand U1919 (N_1919,N_1342,N_1337);
nand U1920 (N_1920,N_1058,N_1000);
nor U1921 (N_1921,N_1241,N_1336);
or U1922 (N_1922,N_1145,N_1151);
and U1923 (N_1923,N_1245,N_1279);
and U1924 (N_1924,N_1158,N_1353);
nor U1925 (N_1925,N_1484,N_1482);
or U1926 (N_1926,N_1497,N_1147);
and U1927 (N_1927,N_1011,N_1164);
or U1928 (N_1928,N_1463,N_1441);
or U1929 (N_1929,N_1004,N_1312);
nand U1930 (N_1930,N_1319,N_1018);
and U1931 (N_1931,N_1341,N_1079);
xnor U1932 (N_1932,N_1062,N_1414);
or U1933 (N_1933,N_1012,N_1301);
or U1934 (N_1934,N_1498,N_1300);
and U1935 (N_1935,N_1334,N_1456);
nand U1936 (N_1936,N_1489,N_1202);
nor U1937 (N_1937,N_1066,N_1359);
or U1938 (N_1938,N_1476,N_1354);
nor U1939 (N_1939,N_1137,N_1030);
or U1940 (N_1940,N_1344,N_1046);
and U1941 (N_1941,N_1387,N_1258);
and U1942 (N_1942,N_1193,N_1083);
or U1943 (N_1943,N_1009,N_1318);
or U1944 (N_1944,N_1187,N_1473);
and U1945 (N_1945,N_1307,N_1135);
nor U1946 (N_1946,N_1460,N_1067);
or U1947 (N_1947,N_1009,N_1173);
or U1948 (N_1948,N_1128,N_1033);
nand U1949 (N_1949,N_1433,N_1353);
nand U1950 (N_1950,N_1494,N_1368);
nor U1951 (N_1951,N_1060,N_1135);
nor U1952 (N_1952,N_1462,N_1057);
and U1953 (N_1953,N_1459,N_1387);
nand U1954 (N_1954,N_1328,N_1257);
nand U1955 (N_1955,N_1473,N_1406);
nand U1956 (N_1956,N_1127,N_1243);
and U1957 (N_1957,N_1191,N_1446);
nand U1958 (N_1958,N_1417,N_1144);
and U1959 (N_1959,N_1186,N_1216);
nand U1960 (N_1960,N_1289,N_1205);
or U1961 (N_1961,N_1218,N_1296);
nand U1962 (N_1962,N_1417,N_1062);
or U1963 (N_1963,N_1071,N_1018);
and U1964 (N_1964,N_1347,N_1106);
or U1965 (N_1965,N_1160,N_1411);
nand U1966 (N_1966,N_1132,N_1441);
nand U1967 (N_1967,N_1175,N_1396);
and U1968 (N_1968,N_1038,N_1181);
nor U1969 (N_1969,N_1100,N_1190);
nor U1970 (N_1970,N_1429,N_1201);
nand U1971 (N_1971,N_1467,N_1192);
nand U1972 (N_1972,N_1476,N_1096);
nor U1973 (N_1973,N_1037,N_1353);
nor U1974 (N_1974,N_1245,N_1265);
nor U1975 (N_1975,N_1210,N_1045);
and U1976 (N_1976,N_1186,N_1389);
or U1977 (N_1977,N_1004,N_1131);
or U1978 (N_1978,N_1130,N_1107);
nand U1979 (N_1979,N_1079,N_1069);
nor U1980 (N_1980,N_1319,N_1353);
nand U1981 (N_1981,N_1361,N_1229);
nor U1982 (N_1982,N_1270,N_1384);
nor U1983 (N_1983,N_1485,N_1218);
and U1984 (N_1984,N_1484,N_1274);
nand U1985 (N_1985,N_1031,N_1340);
nor U1986 (N_1986,N_1099,N_1141);
or U1987 (N_1987,N_1229,N_1353);
and U1988 (N_1988,N_1133,N_1113);
or U1989 (N_1989,N_1136,N_1258);
nor U1990 (N_1990,N_1259,N_1205);
or U1991 (N_1991,N_1277,N_1169);
and U1992 (N_1992,N_1274,N_1283);
nand U1993 (N_1993,N_1437,N_1447);
nand U1994 (N_1994,N_1342,N_1062);
nor U1995 (N_1995,N_1322,N_1440);
nand U1996 (N_1996,N_1154,N_1435);
nor U1997 (N_1997,N_1399,N_1039);
nor U1998 (N_1998,N_1317,N_1184);
or U1999 (N_1999,N_1496,N_1203);
nand U2000 (N_2000,N_1964,N_1681);
or U2001 (N_2001,N_1564,N_1767);
and U2002 (N_2002,N_1870,N_1517);
and U2003 (N_2003,N_1757,N_1998);
nand U2004 (N_2004,N_1689,N_1558);
nor U2005 (N_2005,N_1541,N_1812);
nand U2006 (N_2006,N_1788,N_1738);
and U2007 (N_2007,N_1674,N_1945);
nor U2008 (N_2008,N_1616,N_1784);
and U2009 (N_2009,N_1652,N_1509);
nand U2010 (N_2010,N_1955,N_1817);
or U2011 (N_2011,N_1874,N_1553);
nand U2012 (N_2012,N_1831,N_1521);
or U2013 (N_2013,N_1792,N_1953);
and U2014 (N_2014,N_1718,N_1850);
and U2015 (N_2015,N_1502,N_1810);
and U2016 (N_2016,N_1914,N_1742);
or U2017 (N_2017,N_1770,N_1620);
xor U2018 (N_2018,N_1857,N_1847);
nor U2019 (N_2019,N_1546,N_1855);
nor U2020 (N_2020,N_1733,N_1697);
or U2021 (N_2021,N_1527,N_1725);
nor U2022 (N_2022,N_1882,N_1910);
and U2023 (N_2023,N_1677,N_1952);
and U2024 (N_2024,N_1904,N_1944);
nand U2025 (N_2025,N_1979,N_1795);
nand U2026 (N_2026,N_1853,N_1928);
or U2027 (N_2027,N_1606,N_1512);
and U2028 (N_2028,N_1591,N_1692);
nand U2029 (N_2029,N_1586,N_1961);
nor U2030 (N_2030,N_1838,N_1740);
xor U2031 (N_2031,N_1658,N_1634);
nor U2032 (N_2032,N_1637,N_1787);
nand U2033 (N_2033,N_1777,N_1960);
nor U2034 (N_2034,N_1806,N_1778);
nor U2035 (N_2035,N_1829,N_1837);
xor U2036 (N_2036,N_1891,N_1554);
or U2037 (N_2037,N_1585,N_1755);
and U2038 (N_2038,N_1747,N_1876);
nor U2039 (N_2039,N_1611,N_1514);
nand U2040 (N_2040,N_1576,N_1852);
xor U2041 (N_2041,N_1941,N_1511);
or U2042 (N_2042,N_1507,N_1522);
nor U2043 (N_2043,N_1743,N_1943);
or U2044 (N_2044,N_1972,N_1545);
or U2045 (N_2045,N_1594,N_1813);
or U2046 (N_2046,N_1655,N_1905);
or U2047 (N_2047,N_1645,N_1983);
and U2048 (N_2048,N_1846,N_1551);
and U2049 (N_2049,N_1722,N_1752);
or U2050 (N_2050,N_1986,N_1800);
nand U2051 (N_2051,N_1828,N_1704);
or U2052 (N_2052,N_1848,N_1937);
and U2053 (N_2053,N_1873,N_1956);
and U2054 (N_2054,N_1643,N_1917);
nor U2055 (N_2055,N_1613,N_1918);
or U2056 (N_2056,N_1950,N_1528);
or U2057 (N_2057,N_1995,N_1840);
and U2058 (N_2058,N_1574,N_1854);
nor U2059 (N_2059,N_1863,N_1627);
nand U2060 (N_2060,N_1808,N_1896);
and U2061 (N_2061,N_1650,N_1619);
nand U2062 (N_2062,N_1982,N_1825);
or U2063 (N_2063,N_1954,N_1844);
and U2064 (N_2064,N_1737,N_1851);
or U2065 (N_2065,N_1628,N_1782);
and U2066 (N_2066,N_1880,N_1642);
or U2067 (N_2067,N_1751,N_1878);
nor U2068 (N_2068,N_1572,N_1750);
nand U2069 (N_2069,N_1923,N_1590);
nor U2070 (N_2070,N_1993,N_1609);
or U2071 (N_2071,N_1839,N_1823);
and U2072 (N_2072,N_1543,N_1593);
and U2073 (N_2073,N_1670,N_1885);
or U2074 (N_2074,N_1868,N_1911);
nand U2075 (N_2075,N_1931,N_1799);
nor U2076 (N_2076,N_1781,N_1887);
nand U2077 (N_2077,N_1621,N_1809);
and U2078 (N_2078,N_1930,N_1673);
and U2079 (N_2079,N_1723,N_1513);
and U2080 (N_2080,N_1909,N_1780);
nand U2081 (N_2081,N_1536,N_1603);
and U2082 (N_2082,N_1833,N_1730);
or U2083 (N_2083,N_1649,N_1842);
nand U2084 (N_2084,N_1775,N_1765);
or U2085 (N_2085,N_1940,N_1819);
nand U2086 (N_2086,N_1990,N_1826);
nor U2087 (N_2087,N_1889,N_1530);
xor U2088 (N_2088,N_1818,N_1835);
nand U2089 (N_2089,N_1630,N_1776);
or U2090 (N_2090,N_1794,N_1562);
or U2091 (N_2091,N_1571,N_1753);
and U2092 (N_2092,N_1680,N_1699);
nand U2093 (N_2093,N_1890,N_1762);
or U2094 (N_2094,N_1821,N_1988);
or U2095 (N_2095,N_1602,N_1899);
or U2096 (N_2096,N_1734,N_1604);
nand U2097 (N_2097,N_1547,N_1695);
nor U2098 (N_2098,N_1802,N_1556);
and U2099 (N_2099,N_1764,N_1691);
nor U2100 (N_2100,N_1726,N_1610);
nor U2101 (N_2101,N_1938,N_1696);
nand U2102 (N_2102,N_1657,N_1612);
nand U2103 (N_2103,N_1688,N_1508);
and U2104 (N_2104,N_1834,N_1639);
nand U2105 (N_2105,N_1976,N_1744);
or U2106 (N_2106,N_1962,N_1540);
and U2107 (N_2107,N_1682,N_1915);
and U2108 (N_2108,N_1756,N_1721);
or U2109 (N_2109,N_1932,N_1820);
or U2110 (N_2110,N_1913,N_1779);
or U2111 (N_2111,N_1703,N_1686);
or U2112 (N_2112,N_1866,N_1500);
nor U2113 (N_2113,N_1647,N_1966);
or U2114 (N_2114,N_1600,N_1710);
or U2115 (N_2115,N_1713,N_1980);
nand U2116 (N_2116,N_1531,N_1897);
and U2117 (N_2117,N_1856,N_1958);
and U2118 (N_2118,N_1997,N_1774);
and U2119 (N_2119,N_1532,N_1676);
xor U2120 (N_2120,N_1969,N_1894);
nand U2121 (N_2121,N_1563,N_1957);
nand U2122 (N_2122,N_1929,N_1641);
nand U2123 (N_2123,N_1786,N_1661);
xor U2124 (N_2124,N_1903,N_1951);
xnor U2125 (N_2125,N_1525,N_1895);
nor U2126 (N_2126,N_1888,N_1783);
nand U2127 (N_2127,N_1559,N_1666);
and U2128 (N_2128,N_1769,N_1569);
xor U2129 (N_2129,N_1939,N_1701);
and U2130 (N_2130,N_1519,N_1790);
nand U2131 (N_2131,N_1815,N_1623);
and U2132 (N_2132,N_1675,N_1581);
and U2133 (N_2133,N_1595,N_1908);
or U2134 (N_2134,N_1996,N_1768);
and U2135 (N_2135,N_1567,N_1875);
and U2136 (N_2136,N_1663,N_1884);
nor U2137 (N_2137,N_1719,N_1754);
nand U2138 (N_2138,N_1845,N_1542);
nand U2139 (N_2139,N_1843,N_1566);
and U2140 (N_2140,N_1626,N_1667);
nor U2141 (N_2141,N_1516,N_1830);
and U2142 (N_2142,N_1529,N_1748);
and U2143 (N_2143,N_1946,N_1707);
or U2144 (N_2144,N_1632,N_1598);
nor U2145 (N_2145,N_1592,N_1700);
nor U2146 (N_2146,N_1805,N_1763);
nand U2147 (N_2147,N_1872,N_1577);
and U2148 (N_2148,N_1849,N_1535);
nand U2149 (N_2149,N_1865,N_1796);
or U2150 (N_2150,N_1599,N_1646);
or U2151 (N_2151,N_1936,N_1570);
and U2152 (N_2152,N_1879,N_1539);
and U2153 (N_2153,N_1816,N_1644);
nand U2154 (N_2154,N_1664,N_1978);
xor U2155 (N_2155,N_1948,N_1684);
and U2156 (N_2156,N_1503,N_1678);
and U2157 (N_2157,N_1501,N_1557);
nand U2158 (N_2158,N_1963,N_1862);
and U2159 (N_2159,N_1916,N_1860);
or U2160 (N_2160,N_1758,N_1971);
and U2161 (N_2161,N_1537,N_1968);
and U2162 (N_2162,N_1653,N_1702);
nor U2163 (N_2163,N_1538,N_1974);
nand U2164 (N_2164,N_1771,N_1807);
or U2165 (N_2165,N_1679,N_1708);
nor U2166 (N_2166,N_1714,N_1900);
or U2167 (N_2167,N_1892,N_1668);
nand U2168 (N_2168,N_1615,N_1662);
nor U2169 (N_2169,N_1902,N_1659);
nand U2170 (N_2170,N_1728,N_1669);
nor U2171 (N_2171,N_1793,N_1745);
nand U2172 (N_2172,N_1759,N_1822);
nand U2173 (N_2173,N_1732,N_1523);
and U2174 (N_2174,N_1797,N_1920);
or U2175 (N_2175,N_1548,N_1589);
nand U2176 (N_2176,N_1985,N_1515);
nor U2177 (N_2177,N_1975,N_1544);
nor U2178 (N_2178,N_1869,N_1731);
or U2179 (N_2179,N_1994,N_1859);
nand U2180 (N_2180,N_1935,N_1685);
nor U2181 (N_2181,N_1984,N_1579);
nand U2182 (N_2182,N_1886,N_1729);
nand U2183 (N_2183,N_1614,N_1942);
or U2184 (N_2184,N_1761,N_1864);
nand U2185 (N_2185,N_1970,N_1739);
nor U2186 (N_2186,N_1504,N_1631);
nor U2187 (N_2187,N_1801,N_1568);
nor U2188 (N_2188,N_1981,N_1605);
nand U2189 (N_2189,N_1618,N_1803);
or U2190 (N_2190,N_1683,N_1967);
nor U2191 (N_2191,N_1587,N_1992);
and U2192 (N_2192,N_1877,N_1912);
and U2193 (N_2193,N_1841,N_1883);
nor U2194 (N_2194,N_1624,N_1640);
or U2195 (N_2195,N_1711,N_1625);
or U2196 (N_2196,N_1933,N_1716);
nor U2197 (N_2197,N_1861,N_1565);
nor U2198 (N_2198,N_1607,N_1881);
nand U2199 (N_2199,N_1584,N_1991);
and U2200 (N_2200,N_1583,N_1580);
or U2201 (N_2201,N_1549,N_1694);
nor U2202 (N_2202,N_1550,N_1773);
and U2203 (N_2203,N_1921,N_1648);
nand U2204 (N_2204,N_1926,N_1617);
or U2205 (N_2205,N_1638,N_1832);
nand U2206 (N_2206,N_1687,N_1636);
nand U2207 (N_2207,N_1506,N_1949);
nand U2208 (N_2208,N_1922,N_1717);
and U2209 (N_2209,N_1526,N_1804);
or U2210 (N_2210,N_1578,N_1772);
and U2211 (N_2211,N_1660,N_1999);
or U2212 (N_2212,N_1907,N_1724);
and U2213 (N_2213,N_1520,N_1919);
or U2214 (N_2214,N_1505,N_1712);
nand U2215 (N_2215,N_1693,N_1977);
nand U2216 (N_2216,N_1601,N_1555);
or U2217 (N_2217,N_1629,N_1789);
nand U2218 (N_2218,N_1947,N_1760);
nand U2219 (N_2219,N_1824,N_1965);
nand U2220 (N_2220,N_1749,N_1582);
nor U2221 (N_2221,N_1706,N_1560);
and U2222 (N_2222,N_1552,N_1561);
nor U2223 (N_2223,N_1672,N_1720);
nand U2224 (N_2224,N_1898,N_1656);
or U2225 (N_2225,N_1934,N_1741);
and U2226 (N_2226,N_1871,N_1575);
and U2227 (N_2227,N_1901,N_1573);
nand U2228 (N_2228,N_1633,N_1973);
nor U2229 (N_2229,N_1814,N_1927);
nor U2230 (N_2230,N_1596,N_1533);
nor U2231 (N_2231,N_1518,N_1746);
nor U2232 (N_2232,N_1635,N_1867);
nor U2233 (N_2233,N_1798,N_1811);
and U2234 (N_2234,N_1827,N_1893);
nand U2235 (N_2235,N_1858,N_1608);
or U2236 (N_2236,N_1836,N_1987);
or U2237 (N_2237,N_1715,N_1735);
or U2238 (N_2238,N_1705,N_1989);
and U2239 (N_2239,N_1654,N_1709);
nor U2240 (N_2240,N_1510,N_1727);
and U2241 (N_2241,N_1766,N_1736);
and U2242 (N_2242,N_1651,N_1906);
or U2243 (N_2243,N_1671,N_1690);
and U2244 (N_2244,N_1698,N_1622);
and U2245 (N_2245,N_1791,N_1924);
nor U2246 (N_2246,N_1588,N_1959);
and U2247 (N_2247,N_1524,N_1785);
nor U2248 (N_2248,N_1665,N_1597);
or U2249 (N_2249,N_1925,N_1534);
nor U2250 (N_2250,N_1907,N_1623);
nand U2251 (N_2251,N_1934,N_1975);
or U2252 (N_2252,N_1848,N_1639);
nor U2253 (N_2253,N_1524,N_1502);
nand U2254 (N_2254,N_1689,N_1629);
nor U2255 (N_2255,N_1742,N_1863);
or U2256 (N_2256,N_1713,N_1885);
and U2257 (N_2257,N_1560,N_1806);
nand U2258 (N_2258,N_1647,N_1778);
and U2259 (N_2259,N_1571,N_1665);
and U2260 (N_2260,N_1899,N_1526);
or U2261 (N_2261,N_1654,N_1516);
nor U2262 (N_2262,N_1509,N_1899);
and U2263 (N_2263,N_1639,N_1904);
nor U2264 (N_2264,N_1871,N_1745);
and U2265 (N_2265,N_1981,N_1564);
nand U2266 (N_2266,N_1775,N_1734);
and U2267 (N_2267,N_1806,N_1698);
or U2268 (N_2268,N_1885,N_1596);
and U2269 (N_2269,N_1655,N_1964);
and U2270 (N_2270,N_1714,N_1993);
nand U2271 (N_2271,N_1679,N_1706);
and U2272 (N_2272,N_1717,N_1646);
or U2273 (N_2273,N_1671,N_1935);
or U2274 (N_2274,N_1883,N_1678);
nand U2275 (N_2275,N_1693,N_1596);
and U2276 (N_2276,N_1826,N_1923);
and U2277 (N_2277,N_1779,N_1724);
or U2278 (N_2278,N_1578,N_1803);
nor U2279 (N_2279,N_1581,N_1666);
and U2280 (N_2280,N_1731,N_1535);
nor U2281 (N_2281,N_1709,N_1689);
or U2282 (N_2282,N_1685,N_1977);
or U2283 (N_2283,N_1924,N_1931);
or U2284 (N_2284,N_1566,N_1575);
nand U2285 (N_2285,N_1691,N_1841);
nand U2286 (N_2286,N_1808,N_1820);
or U2287 (N_2287,N_1952,N_1827);
or U2288 (N_2288,N_1551,N_1630);
and U2289 (N_2289,N_1759,N_1887);
or U2290 (N_2290,N_1950,N_1981);
and U2291 (N_2291,N_1939,N_1532);
or U2292 (N_2292,N_1995,N_1955);
and U2293 (N_2293,N_1796,N_1813);
or U2294 (N_2294,N_1570,N_1818);
nand U2295 (N_2295,N_1940,N_1623);
and U2296 (N_2296,N_1931,N_1721);
or U2297 (N_2297,N_1722,N_1535);
nand U2298 (N_2298,N_1876,N_1914);
nor U2299 (N_2299,N_1918,N_1717);
or U2300 (N_2300,N_1618,N_1648);
nand U2301 (N_2301,N_1908,N_1589);
nor U2302 (N_2302,N_1983,N_1971);
nor U2303 (N_2303,N_1892,N_1713);
or U2304 (N_2304,N_1899,N_1923);
or U2305 (N_2305,N_1655,N_1854);
or U2306 (N_2306,N_1588,N_1507);
and U2307 (N_2307,N_1973,N_1907);
or U2308 (N_2308,N_1816,N_1737);
and U2309 (N_2309,N_1879,N_1905);
and U2310 (N_2310,N_1519,N_1651);
and U2311 (N_2311,N_1746,N_1733);
or U2312 (N_2312,N_1968,N_1933);
and U2313 (N_2313,N_1967,N_1665);
nand U2314 (N_2314,N_1587,N_1624);
or U2315 (N_2315,N_1926,N_1957);
nor U2316 (N_2316,N_1757,N_1666);
and U2317 (N_2317,N_1928,N_1740);
nand U2318 (N_2318,N_1698,N_1726);
or U2319 (N_2319,N_1829,N_1992);
nor U2320 (N_2320,N_1846,N_1882);
and U2321 (N_2321,N_1941,N_1958);
or U2322 (N_2322,N_1561,N_1857);
or U2323 (N_2323,N_1823,N_1551);
and U2324 (N_2324,N_1620,N_1950);
nor U2325 (N_2325,N_1885,N_1857);
or U2326 (N_2326,N_1928,N_1806);
or U2327 (N_2327,N_1616,N_1633);
or U2328 (N_2328,N_1977,N_1929);
nor U2329 (N_2329,N_1661,N_1622);
and U2330 (N_2330,N_1611,N_1641);
and U2331 (N_2331,N_1750,N_1954);
or U2332 (N_2332,N_1630,N_1683);
or U2333 (N_2333,N_1751,N_1735);
nand U2334 (N_2334,N_1765,N_1916);
nor U2335 (N_2335,N_1649,N_1958);
and U2336 (N_2336,N_1829,N_1788);
xnor U2337 (N_2337,N_1764,N_1743);
nor U2338 (N_2338,N_1663,N_1820);
nor U2339 (N_2339,N_1705,N_1621);
and U2340 (N_2340,N_1512,N_1665);
nand U2341 (N_2341,N_1609,N_1877);
and U2342 (N_2342,N_1878,N_1827);
nor U2343 (N_2343,N_1809,N_1679);
nand U2344 (N_2344,N_1732,N_1822);
nor U2345 (N_2345,N_1635,N_1610);
nand U2346 (N_2346,N_1556,N_1554);
or U2347 (N_2347,N_1890,N_1522);
and U2348 (N_2348,N_1520,N_1828);
and U2349 (N_2349,N_1511,N_1708);
or U2350 (N_2350,N_1808,N_1811);
or U2351 (N_2351,N_1601,N_1901);
and U2352 (N_2352,N_1594,N_1579);
and U2353 (N_2353,N_1944,N_1630);
nand U2354 (N_2354,N_1605,N_1767);
or U2355 (N_2355,N_1515,N_1509);
and U2356 (N_2356,N_1698,N_1658);
and U2357 (N_2357,N_1894,N_1594);
nor U2358 (N_2358,N_1847,N_1718);
or U2359 (N_2359,N_1711,N_1736);
nor U2360 (N_2360,N_1799,N_1828);
nand U2361 (N_2361,N_1738,N_1796);
and U2362 (N_2362,N_1652,N_1637);
nand U2363 (N_2363,N_1837,N_1525);
and U2364 (N_2364,N_1604,N_1664);
nand U2365 (N_2365,N_1703,N_1887);
or U2366 (N_2366,N_1681,N_1761);
or U2367 (N_2367,N_1941,N_1934);
nand U2368 (N_2368,N_1860,N_1850);
or U2369 (N_2369,N_1886,N_1853);
nand U2370 (N_2370,N_1845,N_1887);
nand U2371 (N_2371,N_1977,N_1696);
nor U2372 (N_2372,N_1639,N_1603);
and U2373 (N_2373,N_1555,N_1857);
nand U2374 (N_2374,N_1527,N_1865);
and U2375 (N_2375,N_1853,N_1840);
nand U2376 (N_2376,N_1694,N_1500);
or U2377 (N_2377,N_1709,N_1667);
nand U2378 (N_2378,N_1580,N_1941);
and U2379 (N_2379,N_1549,N_1792);
or U2380 (N_2380,N_1516,N_1858);
or U2381 (N_2381,N_1658,N_1740);
and U2382 (N_2382,N_1577,N_1580);
nor U2383 (N_2383,N_1524,N_1915);
nor U2384 (N_2384,N_1983,N_1942);
or U2385 (N_2385,N_1691,N_1569);
nor U2386 (N_2386,N_1747,N_1780);
nand U2387 (N_2387,N_1799,N_1652);
or U2388 (N_2388,N_1919,N_1958);
or U2389 (N_2389,N_1886,N_1658);
nor U2390 (N_2390,N_1628,N_1995);
nand U2391 (N_2391,N_1655,N_1679);
nor U2392 (N_2392,N_1896,N_1714);
nor U2393 (N_2393,N_1643,N_1943);
nor U2394 (N_2394,N_1600,N_1967);
and U2395 (N_2395,N_1935,N_1959);
nand U2396 (N_2396,N_1682,N_1564);
nand U2397 (N_2397,N_1701,N_1857);
or U2398 (N_2398,N_1584,N_1960);
xor U2399 (N_2399,N_1913,N_1553);
nand U2400 (N_2400,N_1900,N_1832);
and U2401 (N_2401,N_1979,N_1691);
nand U2402 (N_2402,N_1616,N_1765);
or U2403 (N_2403,N_1955,N_1691);
and U2404 (N_2404,N_1889,N_1509);
nand U2405 (N_2405,N_1661,N_1771);
and U2406 (N_2406,N_1763,N_1885);
and U2407 (N_2407,N_1614,N_1868);
nor U2408 (N_2408,N_1985,N_1927);
and U2409 (N_2409,N_1993,N_1912);
nor U2410 (N_2410,N_1939,N_1712);
and U2411 (N_2411,N_1753,N_1743);
or U2412 (N_2412,N_1609,N_1645);
nand U2413 (N_2413,N_1679,N_1658);
nor U2414 (N_2414,N_1969,N_1700);
nand U2415 (N_2415,N_1857,N_1683);
and U2416 (N_2416,N_1771,N_1800);
xor U2417 (N_2417,N_1711,N_1664);
or U2418 (N_2418,N_1736,N_1758);
nand U2419 (N_2419,N_1663,N_1971);
or U2420 (N_2420,N_1704,N_1813);
nor U2421 (N_2421,N_1998,N_1916);
and U2422 (N_2422,N_1661,N_1951);
nand U2423 (N_2423,N_1742,N_1675);
and U2424 (N_2424,N_1992,N_1645);
nand U2425 (N_2425,N_1686,N_1760);
and U2426 (N_2426,N_1710,N_1988);
and U2427 (N_2427,N_1862,N_1812);
nand U2428 (N_2428,N_1816,N_1519);
and U2429 (N_2429,N_1597,N_1984);
and U2430 (N_2430,N_1553,N_1924);
and U2431 (N_2431,N_1663,N_1928);
or U2432 (N_2432,N_1605,N_1881);
nand U2433 (N_2433,N_1980,N_1723);
and U2434 (N_2434,N_1861,N_1883);
nor U2435 (N_2435,N_1991,N_1520);
nor U2436 (N_2436,N_1762,N_1575);
and U2437 (N_2437,N_1859,N_1728);
nand U2438 (N_2438,N_1949,N_1944);
nand U2439 (N_2439,N_1911,N_1549);
nand U2440 (N_2440,N_1585,N_1608);
or U2441 (N_2441,N_1771,N_1684);
or U2442 (N_2442,N_1847,N_1769);
nand U2443 (N_2443,N_1602,N_1982);
nand U2444 (N_2444,N_1745,N_1744);
and U2445 (N_2445,N_1652,N_1985);
and U2446 (N_2446,N_1988,N_1550);
or U2447 (N_2447,N_1765,N_1901);
or U2448 (N_2448,N_1802,N_1986);
and U2449 (N_2449,N_1643,N_1863);
nand U2450 (N_2450,N_1948,N_1519);
nor U2451 (N_2451,N_1662,N_1970);
xor U2452 (N_2452,N_1826,N_1557);
or U2453 (N_2453,N_1984,N_1514);
nor U2454 (N_2454,N_1815,N_1848);
or U2455 (N_2455,N_1560,N_1982);
nor U2456 (N_2456,N_1901,N_1696);
and U2457 (N_2457,N_1676,N_1973);
or U2458 (N_2458,N_1872,N_1779);
nand U2459 (N_2459,N_1683,N_1677);
nand U2460 (N_2460,N_1640,N_1729);
nor U2461 (N_2461,N_1598,N_1735);
nor U2462 (N_2462,N_1864,N_1951);
nor U2463 (N_2463,N_1534,N_1715);
or U2464 (N_2464,N_1559,N_1934);
nand U2465 (N_2465,N_1669,N_1717);
and U2466 (N_2466,N_1891,N_1861);
or U2467 (N_2467,N_1502,N_1563);
nand U2468 (N_2468,N_1714,N_1999);
and U2469 (N_2469,N_1588,N_1548);
and U2470 (N_2470,N_1859,N_1794);
or U2471 (N_2471,N_1757,N_1873);
nor U2472 (N_2472,N_1505,N_1971);
or U2473 (N_2473,N_1780,N_1802);
or U2474 (N_2474,N_1948,N_1819);
or U2475 (N_2475,N_1767,N_1560);
nand U2476 (N_2476,N_1956,N_1929);
or U2477 (N_2477,N_1857,N_1998);
nor U2478 (N_2478,N_1567,N_1631);
nor U2479 (N_2479,N_1705,N_1993);
and U2480 (N_2480,N_1541,N_1595);
nand U2481 (N_2481,N_1653,N_1646);
nand U2482 (N_2482,N_1724,N_1813);
nand U2483 (N_2483,N_1887,N_1939);
and U2484 (N_2484,N_1791,N_1700);
or U2485 (N_2485,N_1571,N_1953);
nor U2486 (N_2486,N_1560,N_1536);
or U2487 (N_2487,N_1783,N_1772);
or U2488 (N_2488,N_1621,N_1823);
nand U2489 (N_2489,N_1741,N_1595);
nor U2490 (N_2490,N_1643,N_1971);
and U2491 (N_2491,N_1877,N_1812);
or U2492 (N_2492,N_1746,N_1868);
and U2493 (N_2493,N_1989,N_1992);
and U2494 (N_2494,N_1665,N_1518);
or U2495 (N_2495,N_1966,N_1902);
nand U2496 (N_2496,N_1694,N_1737);
nor U2497 (N_2497,N_1753,N_1805);
nor U2498 (N_2498,N_1681,N_1554);
nand U2499 (N_2499,N_1600,N_1535);
nor U2500 (N_2500,N_2405,N_2323);
nor U2501 (N_2501,N_2360,N_2358);
nand U2502 (N_2502,N_2257,N_2096);
nand U2503 (N_2503,N_2078,N_2347);
and U2504 (N_2504,N_2192,N_2178);
or U2505 (N_2505,N_2162,N_2349);
or U2506 (N_2506,N_2235,N_2007);
nand U2507 (N_2507,N_2270,N_2336);
or U2508 (N_2508,N_2116,N_2397);
nor U2509 (N_2509,N_2473,N_2390);
nand U2510 (N_2510,N_2008,N_2327);
nor U2511 (N_2511,N_2357,N_2155);
xor U2512 (N_2512,N_2317,N_2064);
nand U2513 (N_2513,N_2234,N_2062);
nand U2514 (N_2514,N_2383,N_2256);
nand U2515 (N_2515,N_2296,N_2493);
and U2516 (N_2516,N_2053,N_2458);
nor U2517 (N_2517,N_2247,N_2449);
or U2518 (N_2518,N_2117,N_2016);
nor U2519 (N_2519,N_2472,N_2034);
or U2520 (N_2520,N_2344,N_2470);
or U2521 (N_2521,N_2082,N_2128);
and U2522 (N_2522,N_2321,N_2393);
or U2523 (N_2523,N_2379,N_2381);
nor U2524 (N_2524,N_2319,N_2017);
or U2525 (N_2525,N_2076,N_2230);
nand U2526 (N_2526,N_2352,N_2005);
nand U2527 (N_2527,N_2119,N_2367);
nor U2528 (N_2528,N_2300,N_2399);
nor U2529 (N_2529,N_2228,N_2071);
nand U2530 (N_2530,N_2410,N_2464);
nor U2531 (N_2531,N_2063,N_2365);
nand U2532 (N_2532,N_2277,N_2196);
or U2533 (N_2533,N_2029,N_2477);
nand U2534 (N_2534,N_2129,N_2419);
or U2535 (N_2535,N_2471,N_2355);
nand U2536 (N_2536,N_2144,N_2406);
nand U2537 (N_2537,N_2214,N_2260);
or U2538 (N_2538,N_2147,N_2446);
nand U2539 (N_2539,N_2201,N_2246);
or U2540 (N_2540,N_2398,N_2299);
and U2541 (N_2541,N_2055,N_2261);
nand U2542 (N_2542,N_2320,N_2203);
nor U2543 (N_2543,N_2089,N_2309);
or U2544 (N_2544,N_2191,N_2272);
and U2545 (N_2545,N_2417,N_2429);
or U2546 (N_2546,N_2075,N_2036);
and U2547 (N_2547,N_2161,N_2452);
and U2548 (N_2548,N_2376,N_2179);
xnor U2549 (N_2549,N_2457,N_2254);
or U2550 (N_2550,N_2208,N_2242);
or U2551 (N_2551,N_2112,N_2118);
and U2552 (N_2552,N_2010,N_2157);
nor U2553 (N_2553,N_2488,N_2408);
or U2554 (N_2554,N_2154,N_2310);
nor U2555 (N_2555,N_2418,N_2197);
nor U2556 (N_2556,N_2202,N_2215);
nand U2557 (N_2557,N_2120,N_2479);
xnor U2558 (N_2558,N_2021,N_2106);
nand U2559 (N_2559,N_2187,N_2395);
nand U2560 (N_2560,N_2334,N_2314);
nor U2561 (N_2561,N_2145,N_2223);
and U2562 (N_2562,N_2474,N_2188);
nand U2563 (N_2563,N_2318,N_2003);
nand U2564 (N_2564,N_2439,N_2332);
and U2565 (N_2565,N_2394,N_2266);
nand U2566 (N_2566,N_2364,N_2366);
or U2567 (N_2567,N_2212,N_2158);
nand U2568 (N_2568,N_2194,N_2440);
and U2569 (N_2569,N_2425,N_2072);
nand U2570 (N_2570,N_2095,N_2380);
nor U2571 (N_2571,N_2404,N_2495);
and U2572 (N_2572,N_2416,N_2136);
nand U2573 (N_2573,N_2163,N_2295);
nand U2574 (N_2574,N_2020,N_2073);
or U2575 (N_2575,N_2285,N_2011);
nor U2576 (N_2576,N_2056,N_2373);
nand U2577 (N_2577,N_2359,N_2074);
xnor U2578 (N_2578,N_2281,N_2035);
and U2579 (N_2579,N_2308,N_2391);
nand U2580 (N_2580,N_2420,N_2258);
nor U2581 (N_2581,N_2123,N_2335);
or U2582 (N_2582,N_2177,N_2460);
nand U2583 (N_2583,N_2169,N_2040);
and U2584 (N_2584,N_2140,N_2100);
nor U2585 (N_2585,N_2019,N_2353);
nand U2586 (N_2586,N_2052,N_2450);
nand U2587 (N_2587,N_2108,N_2087);
nand U2588 (N_2588,N_2160,N_2047);
nand U2589 (N_2589,N_2138,N_2368);
or U2590 (N_2590,N_2276,N_2341);
and U2591 (N_2591,N_2243,N_2279);
nor U2592 (N_2592,N_2028,N_2233);
or U2593 (N_2593,N_2044,N_2356);
or U2594 (N_2594,N_2092,N_2079);
nand U2595 (N_2595,N_2122,N_2133);
nand U2596 (N_2596,N_2496,N_2485);
nand U2597 (N_2597,N_2486,N_2290);
or U2598 (N_2598,N_2181,N_2275);
nand U2599 (N_2599,N_2468,N_2442);
nor U2600 (N_2600,N_2375,N_2189);
nand U2601 (N_2601,N_2218,N_2291);
or U2602 (N_2602,N_2489,N_2057);
and U2603 (N_2603,N_2051,N_2232);
or U2604 (N_2604,N_2114,N_2283);
and U2605 (N_2605,N_2409,N_2292);
nand U2606 (N_2606,N_2432,N_2330);
and U2607 (N_2607,N_2451,N_2298);
nand U2608 (N_2608,N_2414,N_2022);
or U2609 (N_2609,N_2241,N_2059);
or U2610 (N_2610,N_2173,N_2012);
and U2611 (N_2611,N_2287,N_2206);
nor U2612 (N_2612,N_2186,N_2026);
nor U2613 (N_2613,N_2103,N_2067);
or U2614 (N_2614,N_2141,N_2264);
nor U2615 (N_2615,N_2494,N_2217);
or U2616 (N_2616,N_2475,N_2226);
nand U2617 (N_2617,N_2001,N_2263);
nand U2618 (N_2618,N_2094,N_2345);
nor U2619 (N_2619,N_2443,N_2433);
nor U2620 (N_2620,N_2156,N_2403);
nor U2621 (N_2621,N_2371,N_2412);
nor U2622 (N_2622,N_2113,N_2396);
or U2623 (N_2623,N_2061,N_2430);
xor U2624 (N_2624,N_2307,N_2483);
nor U2625 (N_2625,N_2484,N_2111);
nand U2626 (N_2626,N_2102,N_2027);
or U2627 (N_2627,N_2411,N_2286);
nand U2628 (N_2628,N_2236,N_2083);
or U2629 (N_2629,N_2467,N_2221);
nand U2630 (N_2630,N_2213,N_2343);
nand U2631 (N_2631,N_2250,N_2077);
and U2632 (N_2632,N_2374,N_2152);
or U2633 (N_2633,N_2448,N_2149);
or U2634 (N_2634,N_2305,N_2042);
nand U2635 (N_2635,N_2311,N_2342);
or U2636 (N_2636,N_2313,N_2240);
nand U2637 (N_2637,N_2024,N_2227);
nand U2638 (N_2638,N_2441,N_2269);
or U2639 (N_2639,N_2143,N_2065);
nand U2640 (N_2640,N_2015,N_2329);
nor U2641 (N_2641,N_2389,N_2306);
nor U2642 (N_2642,N_2031,N_2090);
and U2643 (N_2643,N_2370,N_2050);
or U2644 (N_2644,N_2339,N_2244);
xnor U2645 (N_2645,N_2265,N_2455);
nand U2646 (N_2646,N_2229,N_2351);
or U2647 (N_2647,N_2492,N_2006);
and U2648 (N_2648,N_2337,N_2205);
and U2649 (N_2649,N_2431,N_2248);
nor U2650 (N_2650,N_2293,N_2386);
nand U2651 (N_2651,N_2415,N_2025);
or U2652 (N_2652,N_2132,N_2436);
nand U2653 (N_2653,N_2098,N_2252);
nor U2654 (N_2654,N_2135,N_2032);
and U2655 (N_2655,N_2251,N_2190);
or U2656 (N_2656,N_2463,N_2107);
nor U2657 (N_2657,N_2387,N_2427);
nand U2658 (N_2658,N_2193,N_2469);
nor U2659 (N_2659,N_2456,N_2170);
or U2660 (N_2660,N_2382,N_2018);
or U2661 (N_2661,N_2153,N_2384);
or U2662 (N_2662,N_2361,N_2127);
or U2663 (N_2663,N_2126,N_2037);
and U2664 (N_2664,N_2426,N_2014);
nand U2665 (N_2665,N_2407,N_2400);
or U2666 (N_2666,N_2038,N_2326);
nor U2667 (N_2667,N_2224,N_2150);
nor U2668 (N_2668,N_2130,N_2183);
nor U2669 (N_2669,N_2346,N_2253);
and U2670 (N_2670,N_2487,N_2268);
or U2671 (N_2671,N_2238,N_2000);
nand U2672 (N_2672,N_2175,N_2207);
nand U2673 (N_2673,N_2099,N_2301);
nor U2674 (N_2674,N_2369,N_2091);
and U2675 (N_2675,N_2274,N_2434);
or U2676 (N_2676,N_2134,N_2041);
and U2677 (N_2677,N_2231,N_2304);
and U2678 (N_2678,N_2174,N_2462);
nand U2679 (N_2679,N_2478,N_2093);
and U2680 (N_2680,N_2362,N_2176);
and U2681 (N_2681,N_2294,N_2303);
or U2682 (N_2682,N_2033,N_2115);
and U2683 (N_2683,N_2198,N_2097);
and U2684 (N_2684,N_2385,N_2009);
and U2685 (N_2685,N_2168,N_2278);
or U2686 (N_2686,N_2363,N_2164);
or U2687 (N_2687,N_2348,N_2402);
or U2688 (N_2688,N_2219,N_2070);
nor U2689 (N_2689,N_2282,N_2039);
nor U2690 (N_2690,N_2328,N_2482);
nand U2691 (N_2691,N_2222,N_2185);
nand U2692 (N_2692,N_2491,N_2060);
nand U2693 (N_2693,N_2284,N_2139);
nand U2694 (N_2694,N_2171,N_2043);
nor U2695 (N_2695,N_2151,N_2104);
or U2696 (N_2696,N_2069,N_2437);
nand U2697 (N_2697,N_2372,N_2259);
or U2698 (N_2698,N_2216,N_2081);
nand U2699 (N_2699,N_2447,N_2288);
and U2700 (N_2700,N_2401,N_2239);
nand U2701 (N_2701,N_2030,N_2481);
nand U2702 (N_2702,N_2271,N_2220);
nor U2703 (N_2703,N_2167,N_2262);
and U2704 (N_2704,N_2422,N_2172);
and U2705 (N_2705,N_2124,N_2499);
nor U2706 (N_2706,N_2453,N_2454);
nor U2707 (N_2707,N_2249,N_2392);
nand U2708 (N_2708,N_2199,N_2424);
and U2709 (N_2709,N_2204,N_2497);
or U2710 (N_2710,N_2480,N_2200);
or U2711 (N_2711,N_2105,N_2125);
nor U2712 (N_2712,N_2109,N_2490);
nor U2713 (N_2713,N_2080,N_2068);
and U2714 (N_2714,N_2331,N_2476);
and U2715 (N_2715,N_2459,N_2498);
and U2716 (N_2716,N_2013,N_2350);
nor U2717 (N_2717,N_2273,N_2086);
nor U2718 (N_2718,N_2413,N_2209);
nand U2719 (N_2719,N_2101,N_2210);
and U2720 (N_2720,N_2049,N_2084);
nand U2721 (N_2721,N_2045,N_2166);
nor U2722 (N_2722,N_2023,N_2444);
nor U2723 (N_2723,N_2280,N_2388);
nand U2724 (N_2724,N_2002,N_2445);
and U2725 (N_2725,N_2137,N_2142);
or U2726 (N_2726,N_2333,N_2267);
nand U2727 (N_2727,N_2465,N_2322);
nand U2728 (N_2728,N_2354,N_2182);
and U2729 (N_2729,N_2004,N_2088);
and U2730 (N_2730,N_2435,N_2245);
or U2731 (N_2731,N_2131,N_2421);
nor U2732 (N_2732,N_2315,N_2110);
or U2733 (N_2733,N_2085,N_2195);
nand U2734 (N_2734,N_2461,N_2146);
or U2735 (N_2735,N_2340,N_2159);
and U2736 (N_2736,N_2165,N_2312);
or U2737 (N_2737,N_2316,N_2302);
nand U2738 (N_2738,N_2423,N_2211);
nand U2739 (N_2739,N_2324,N_2466);
or U2740 (N_2740,N_2184,N_2048);
nor U2741 (N_2741,N_2255,N_2054);
nand U2742 (N_2742,N_2148,N_2377);
or U2743 (N_2743,N_2046,N_2066);
and U2744 (N_2744,N_2428,N_2058);
nand U2745 (N_2745,N_2297,N_2289);
or U2746 (N_2746,N_2180,N_2121);
nor U2747 (N_2747,N_2438,N_2225);
or U2748 (N_2748,N_2325,N_2237);
nor U2749 (N_2749,N_2378,N_2338);
and U2750 (N_2750,N_2100,N_2480);
nand U2751 (N_2751,N_2226,N_2128);
nand U2752 (N_2752,N_2221,N_2360);
or U2753 (N_2753,N_2339,N_2211);
or U2754 (N_2754,N_2047,N_2345);
or U2755 (N_2755,N_2004,N_2141);
nand U2756 (N_2756,N_2078,N_2360);
and U2757 (N_2757,N_2367,N_2393);
nor U2758 (N_2758,N_2482,N_2316);
and U2759 (N_2759,N_2373,N_2020);
nor U2760 (N_2760,N_2140,N_2220);
or U2761 (N_2761,N_2446,N_2000);
or U2762 (N_2762,N_2410,N_2327);
nor U2763 (N_2763,N_2259,N_2215);
or U2764 (N_2764,N_2223,N_2243);
and U2765 (N_2765,N_2339,N_2250);
nand U2766 (N_2766,N_2427,N_2434);
xor U2767 (N_2767,N_2445,N_2151);
nor U2768 (N_2768,N_2435,N_2186);
xnor U2769 (N_2769,N_2047,N_2223);
nand U2770 (N_2770,N_2282,N_2029);
and U2771 (N_2771,N_2169,N_2495);
or U2772 (N_2772,N_2360,N_2015);
or U2773 (N_2773,N_2012,N_2367);
and U2774 (N_2774,N_2484,N_2425);
or U2775 (N_2775,N_2309,N_2020);
and U2776 (N_2776,N_2009,N_2104);
nor U2777 (N_2777,N_2353,N_2161);
or U2778 (N_2778,N_2182,N_2216);
or U2779 (N_2779,N_2243,N_2156);
or U2780 (N_2780,N_2384,N_2122);
nand U2781 (N_2781,N_2471,N_2209);
nand U2782 (N_2782,N_2087,N_2493);
xnor U2783 (N_2783,N_2176,N_2368);
or U2784 (N_2784,N_2372,N_2442);
and U2785 (N_2785,N_2144,N_2022);
nor U2786 (N_2786,N_2094,N_2410);
and U2787 (N_2787,N_2444,N_2384);
nand U2788 (N_2788,N_2390,N_2030);
nor U2789 (N_2789,N_2007,N_2434);
nor U2790 (N_2790,N_2427,N_2040);
and U2791 (N_2791,N_2097,N_2309);
nor U2792 (N_2792,N_2409,N_2079);
nor U2793 (N_2793,N_2351,N_2224);
nand U2794 (N_2794,N_2039,N_2318);
nor U2795 (N_2795,N_2248,N_2316);
nand U2796 (N_2796,N_2041,N_2127);
nor U2797 (N_2797,N_2106,N_2418);
and U2798 (N_2798,N_2337,N_2129);
or U2799 (N_2799,N_2336,N_2089);
nand U2800 (N_2800,N_2326,N_2033);
and U2801 (N_2801,N_2250,N_2166);
nand U2802 (N_2802,N_2498,N_2206);
nand U2803 (N_2803,N_2370,N_2194);
or U2804 (N_2804,N_2000,N_2443);
and U2805 (N_2805,N_2149,N_2397);
nand U2806 (N_2806,N_2392,N_2190);
nand U2807 (N_2807,N_2406,N_2254);
nand U2808 (N_2808,N_2214,N_2209);
nand U2809 (N_2809,N_2480,N_2376);
or U2810 (N_2810,N_2364,N_2136);
and U2811 (N_2811,N_2161,N_2463);
and U2812 (N_2812,N_2046,N_2100);
nand U2813 (N_2813,N_2056,N_2432);
and U2814 (N_2814,N_2428,N_2067);
and U2815 (N_2815,N_2243,N_2066);
or U2816 (N_2816,N_2325,N_2352);
nand U2817 (N_2817,N_2364,N_2350);
or U2818 (N_2818,N_2089,N_2067);
nor U2819 (N_2819,N_2295,N_2155);
nor U2820 (N_2820,N_2482,N_2314);
or U2821 (N_2821,N_2312,N_2322);
nand U2822 (N_2822,N_2457,N_2031);
nor U2823 (N_2823,N_2439,N_2418);
nand U2824 (N_2824,N_2117,N_2165);
nand U2825 (N_2825,N_2271,N_2132);
or U2826 (N_2826,N_2053,N_2238);
nand U2827 (N_2827,N_2234,N_2440);
nor U2828 (N_2828,N_2336,N_2111);
nand U2829 (N_2829,N_2144,N_2484);
or U2830 (N_2830,N_2148,N_2386);
or U2831 (N_2831,N_2490,N_2108);
nand U2832 (N_2832,N_2386,N_2164);
or U2833 (N_2833,N_2271,N_2111);
and U2834 (N_2834,N_2151,N_2212);
nor U2835 (N_2835,N_2328,N_2218);
xor U2836 (N_2836,N_2245,N_2261);
and U2837 (N_2837,N_2268,N_2259);
nor U2838 (N_2838,N_2242,N_2114);
and U2839 (N_2839,N_2334,N_2377);
nand U2840 (N_2840,N_2096,N_2054);
or U2841 (N_2841,N_2168,N_2326);
nand U2842 (N_2842,N_2074,N_2151);
or U2843 (N_2843,N_2232,N_2352);
nand U2844 (N_2844,N_2260,N_2164);
nand U2845 (N_2845,N_2335,N_2029);
nor U2846 (N_2846,N_2433,N_2188);
xor U2847 (N_2847,N_2224,N_2297);
or U2848 (N_2848,N_2371,N_2393);
nor U2849 (N_2849,N_2237,N_2414);
and U2850 (N_2850,N_2452,N_2193);
and U2851 (N_2851,N_2068,N_2424);
nand U2852 (N_2852,N_2110,N_2056);
nand U2853 (N_2853,N_2487,N_2218);
or U2854 (N_2854,N_2136,N_2375);
and U2855 (N_2855,N_2242,N_2256);
nand U2856 (N_2856,N_2359,N_2239);
nor U2857 (N_2857,N_2145,N_2052);
nand U2858 (N_2858,N_2069,N_2181);
nor U2859 (N_2859,N_2038,N_2223);
nor U2860 (N_2860,N_2355,N_2477);
and U2861 (N_2861,N_2041,N_2412);
and U2862 (N_2862,N_2058,N_2160);
and U2863 (N_2863,N_2417,N_2390);
or U2864 (N_2864,N_2479,N_2104);
or U2865 (N_2865,N_2190,N_2029);
and U2866 (N_2866,N_2170,N_2104);
and U2867 (N_2867,N_2295,N_2424);
and U2868 (N_2868,N_2497,N_2090);
and U2869 (N_2869,N_2170,N_2315);
and U2870 (N_2870,N_2020,N_2222);
nor U2871 (N_2871,N_2190,N_2482);
and U2872 (N_2872,N_2029,N_2489);
or U2873 (N_2873,N_2178,N_2119);
xnor U2874 (N_2874,N_2398,N_2189);
or U2875 (N_2875,N_2462,N_2256);
nor U2876 (N_2876,N_2023,N_2360);
nand U2877 (N_2877,N_2256,N_2085);
xor U2878 (N_2878,N_2294,N_2180);
or U2879 (N_2879,N_2128,N_2291);
nand U2880 (N_2880,N_2071,N_2062);
and U2881 (N_2881,N_2490,N_2205);
and U2882 (N_2882,N_2009,N_2456);
nand U2883 (N_2883,N_2010,N_2018);
nor U2884 (N_2884,N_2386,N_2439);
and U2885 (N_2885,N_2344,N_2380);
and U2886 (N_2886,N_2294,N_2462);
nor U2887 (N_2887,N_2268,N_2232);
nand U2888 (N_2888,N_2094,N_2259);
nand U2889 (N_2889,N_2022,N_2373);
or U2890 (N_2890,N_2458,N_2174);
nand U2891 (N_2891,N_2473,N_2134);
and U2892 (N_2892,N_2294,N_2093);
nand U2893 (N_2893,N_2077,N_2105);
or U2894 (N_2894,N_2196,N_2309);
nor U2895 (N_2895,N_2174,N_2265);
nor U2896 (N_2896,N_2382,N_2404);
nand U2897 (N_2897,N_2029,N_2308);
nor U2898 (N_2898,N_2139,N_2403);
nand U2899 (N_2899,N_2134,N_2191);
nand U2900 (N_2900,N_2323,N_2036);
nand U2901 (N_2901,N_2443,N_2462);
nand U2902 (N_2902,N_2455,N_2491);
and U2903 (N_2903,N_2243,N_2316);
xnor U2904 (N_2904,N_2283,N_2445);
nand U2905 (N_2905,N_2248,N_2353);
or U2906 (N_2906,N_2007,N_2263);
and U2907 (N_2907,N_2022,N_2093);
nand U2908 (N_2908,N_2356,N_2489);
nand U2909 (N_2909,N_2306,N_2353);
nand U2910 (N_2910,N_2374,N_2443);
or U2911 (N_2911,N_2219,N_2480);
nor U2912 (N_2912,N_2499,N_2161);
nor U2913 (N_2913,N_2483,N_2166);
and U2914 (N_2914,N_2149,N_2261);
nand U2915 (N_2915,N_2335,N_2042);
nand U2916 (N_2916,N_2313,N_2158);
nor U2917 (N_2917,N_2378,N_2389);
nand U2918 (N_2918,N_2005,N_2473);
or U2919 (N_2919,N_2140,N_2249);
nor U2920 (N_2920,N_2227,N_2133);
nor U2921 (N_2921,N_2067,N_2223);
nor U2922 (N_2922,N_2077,N_2364);
or U2923 (N_2923,N_2386,N_2192);
nor U2924 (N_2924,N_2083,N_2177);
or U2925 (N_2925,N_2071,N_2078);
nand U2926 (N_2926,N_2244,N_2180);
and U2927 (N_2927,N_2239,N_2079);
and U2928 (N_2928,N_2016,N_2452);
nand U2929 (N_2929,N_2030,N_2495);
or U2930 (N_2930,N_2477,N_2297);
nor U2931 (N_2931,N_2495,N_2172);
nor U2932 (N_2932,N_2342,N_2015);
or U2933 (N_2933,N_2327,N_2018);
nand U2934 (N_2934,N_2448,N_2039);
nand U2935 (N_2935,N_2440,N_2023);
nand U2936 (N_2936,N_2099,N_2446);
or U2937 (N_2937,N_2037,N_2270);
nor U2938 (N_2938,N_2064,N_2244);
or U2939 (N_2939,N_2144,N_2312);
and U2940 (N_2940,N_2492,N_2391);
or U2941 (N_2941,N_2356,N_2162);
nor U2942 (N_2942,N_2420,N_2210);
nand U2943 (N_2943,N_2240,N_2057);
nor U2944 (N_2944,N_2354,N_2378);
or U2945 (N_2945,N_2389,N_2298);
nor U2946 (N_2946,N_2132,N_2165);
nand U2947 (N_2947,N_2069,N_2220);
nor U2948 (N_2948,N_2398,N_2410);
and U2949 (N_2949,N_2349,N_2149);
xor U2950 (N_2950,N_2183,N_2395);
and U2951 (N_2951,N_2479,N_2099);
nor U2952 (N_2952,N_2431,N_2258);
nand U2953 (N_2953,N_2191,N_2014);
nor U2954 (N_2954,N_2067,N_2335);
nand U2955 (N_2955,N_2350,N_2119);
nand U2956 (N_2956,N_2202,N_2250);
nor U2957 (N_2957,N_2254,N_2325);
nand U2958 (N_2958,N_2466,N_2443);
nand U2959 (N_2959,N_2428,N_2391);
nand U2960 (N_2960,N_2064,N_2071);
or U2961 (N_2961,N_2242,N_2282);
xnor U2962 (N_2962,N_2259,N_2322);
or U2963 (N_2963,N_2431,N_2276);
nand U2964 (N_2964,N_2419,N_2391);
or U2965 (N_2965,N_2181,N_2312);
nor U2966 (N_2966,N_2404,N_2344);
or U2967 (N_2967,N_2424,N_2465);
nor U2968 (N_2968,N_2344,N_2322);
and U2969 (N_2969,N_2441,N_2308);
and U2970 (N_2970,N_2002,N_2023);
and U2971 (N_2971,N_2332,N_2441);
nand U2972 (N_2972,N_2248,N_2004);
nor U2973 (N_2973,N_2155,N_2491);
nor U2974 (N_2974,N_2144,N_2320);
nor U2975 (N_2975,N_2027,N_2489);
nor U2976 (N_2976,N_2050,N_2388);
nor U2977 (N_2977,N_2329,N_2012);
and U2978 (N_2978,N_2187,N_2453);
and U2979 (N_2979,N_2233,N_2115);
nand U2980 (N_2980,N_2273,N_2011);
and U2981 (N_2981,N_2055,N_2493);
nor U2982 (N_2982,N_2189,N_2200);
nand U2983 (N_2983,N_2450,N_2382);
nor U2984 (N_2984,N_2210,N_2009);
xor U2985 (N_2985,N_2460,N_2375);
xnor U2986 (N_2986,N_2056,N_2484);
and U2987 (N_2987,N_2474,N_2307);
nor U2988 (N_2988,N_2283,N_2221);
and U2989 (N_2989,N_2185,N_2394);
or U2990 (N_2990,N_2331,N_2394);
or U2991 (N_2991,N_2051,N_2029);
or U2992 (N_2992,N_2105,N_2009);
and U2993 (N_2993,N_2329,N_2040);
nand U2994 (N_2994,N_2405,N_2487);
nand U2995 (N_2995,N_2000,N_2416);
nor U2996 (N_2996,N_2240,N_2223);
and U2997 (N_2997,N_2323,N_2073);
nor U2998 (N_2998,N_2433,N_2463);
xnor U2999 (N_2999,N_2057,N_2261);
or UO_0 (O_0,N_2578,N_2708);
or UO_1 (O_1,N_2920,N_2635);
nand UO_2 (O_2,N_2768,N_2711);
nand UO_3 (O_3,N_2580,N_2511);
or UO_4 (O_4,N_2901,N_2770);
nand UO_5 (O_5,N_2588,N_2602);
or UO_6 (O_6,N_2935,N_2915);
nor UO_7 (O_7,N_2671,N_2828);
and UO_8 (O_8,N_2613,N_2722);
nand UO_9 (O_9,N_2514,N_2591);
and UO_10 (O_10,N_2834,N_2846);
nand UO_11 (O_11,N_2746,N_2579);
nand UO_12 (O_12,N_2535,N_2847);
xnor UO_13 (O_13,N_2844,N_2638);
and UO_14 (O_14,N_2748,N_2601);
nand UO_15 (O_15,N_2732,N_2887);
or UO_16 (O_16,N_2964,N_2769);
nor UO_17 (O_17,N_2968,N_2663);
or UO_18 (O_18,N_2909,N_2596);
nand UO_19 (O_19,N_2720,N_2633);
and UO_20 (O_20,N_2632,N_2636);
or UO_21 (O_21,N_2709,N_2500);
nand UO_22 (O_22,N_2698,N_2573);
nand UO_23 (O_23,N_2687,N_2541);
and UO_24 (O_24,N_2958,N_2657);
and UO_25 (O_25,N_2877,N_2517);
and UO_26 (O_26,N_2505,N_2614);
and UO_27 (O_27,N_2861,N_2704);
nor UO_28 (O_28,N_2533,N_2685);
nand UO_29 (O_29,N_2696,N_2705);
or UO_30 (O_30,N_2540,N_2907);
nand UO_31 (O_31,N_2959,N_2526);
or UO_32 (O_32,N_2554,N_2730);
or UO_33 (O_33,N_2830,N_2998);
nor UO_34 (O_34,N_2853,N_2572);
nand UO_35 (O_35,N_2949,N_2697);
nand UO_36 (O_36,N_2759,N_2950);
and UO_37 (O_37,N_2529,N_2912);
or UO_38 (O_38,N_2760,N_2512);
nand UO_39 (O_39,N_2963,N_2520);
nand UO_40 (O_40,N_2710,N_2878);
and UO_41 (O_41,N_2739,N_2783);
nand UO_42 (O_42,N_2800,N_2896);
or UO_43 (O_43,N_2557,N_2885);
and UO_44 (O_44,N_2568,N_2902);
xnor UO_45 (O_45,N_2795,N_2819);
and UO_46 (O_46,N_2599,N_2762);
or UO_47 (O_47,N_2651,N_2953);
and UO_48 (O_48,N_2808,N_2648);
and UO_49 (O_49,N_2680,N_2530);
nor UO_50 (O_50,N_2982,N_2818);
nand UO_51 (O_51,N_2618,N_2822);
and UO_52 (O_52,N_2753,N_2942);
nand UO_53 (O_53,N_2656,N_2791);
xor UO_54 (O_54,N_2700,N_2786);
nor UO_55 (O_55,N_2873,N_2874);
and UO_56 (O_56,N_2731,N_2924);
nor UO_57 (O_57,N_2794,N_2510);
nand UO_58 (O_58,N_2584,N_2867);
and UO_59 (O_59,N_2764,N_2987);
or UO_60 (O_60,N_2645,N_2930);
and UO_61 (O_61,N_2884,N_2779);
and UO_62 (O_62,N_2539,N_2501);
nand UO_63 (O_63,N_2558,N_2676);
and UO_64 (O_64,N_2978,N_2666);
nand UO_65 (O_65,N_2725,N_2889);
nand UO_66 (O_66,N_2669,N_2567);
nand UO_67 (O_67,N_2983,N_2823);
or UO_68 (O_68,N_2716,N_2681);
or UO_69 (O_69,N_2537,N_2985);
or UO_70 (O_70,N_2993,N_2544);
nand UO_71 (O_71,N_2707,N_2615);
or UO_72 (O_72,N_2560,N_2547);
or UO_73 (O_73,N_2804,N_2617);
nor UO_74 (O_74,N_2576,N_2522);
or UO_75 (O_75,N_2639,N_2532);
nand UO_76 (O_76,N_2937,N_2747);
nand UO_77 (O_77,N_2702,N_2542);
xor UO_78 (O_78,N_2852,N_2972);
and UO_79 (O_79,N_2839,N_2654);
nor UO_80 (O_80,N_2603,N_2631);
and UO_81 (O_81,N_2695,N_2995);
and UO_82 (O_82,N_2957,N_2548);
and UO_83 (O_83,N_2780,N_2506);
and UO_84 (O_84,N_2848,N_2620);
nand UO_85 (O_85,N_2655,N_2564);
and UO_86 (O_86,N_2575,N_2766);
nor UO_87 (O_87,N_2989,N_2590);
and UO_88 (O_88,N_2807,N_2918);
nor UO_89 (O_89,N_2742,N_2728);
or UO_90 (O_90,N_2965,N_2686);
nand UO_91 (O_91,N_2761,N_2970);
and UO_92 (O_92,N_2859,N_2771);
nor UO_93 (O_93,N_2967,N_2908);
nand UO_94 (O_94,N_2609,N_2851);
nand UO_95 (O_95,N_2876,N_2745);
nand UO_96 (O_96,N_2699,N_2677);
and UO_97 (O_97,N_2624,N_2837);
nand UO_98 (O_98,N_2717,N_2956);
and UO_99 (O_99,N_2842,N_2737);
nand UO_100 (O_100,N_2820,N_2879);
xor UO_101 (O_101,N_2977,N_2929);
and UO_102 (O_102,N_2821,N_2556);
and UO_103 (O_103,N_2606,N_2831);
and UO_104 (O_104,N_2527,N_2845);
and UO_105 (O_105,N_2589,N_2604);
nor UO_106 (O_106,N_2751,N_2583);
nor UO_107 (O_107,N_2736,N_2534);
nor UO_108 (O_108,N_2660,N_2503);
nand UO_109 (O_109,N_2598,N_2524);
nor UO_110 (O_110,N_2777,N_2775);
xor UO_111 (O_111,N_2653,N_2597);
nand UO_112 (O_112,N_2693,N_2750);
and UO_113 (O_113,N_2673,N_2713);
nor UO_114 (O_114,N_2741,N_2981);
and UO_115 (O_115,N_2927,N_2712);
nor UO_116 (O_116,N_2940,N_2814);
and UO_117 (O_117,N_2893,N_2797);
nor UO_118 (O_118,N_2835,N_2802);
nor UO_119 (O_119,N_2649,N_2860);
or UO_120 (O_120,N_2565,N_2857);
or UO_121 (O_121,N_2891,N_2974);
nand UO_122 (O_122,N_2793,N_2897);
and UO_123 (O_123,N_2763,N_2559);
nand UO_124 (O_124,N_2587,N_2829);
nor UO_125 (O_125,N_2774,N_2627);
nor UO_126 (O_126,N_2809,N_2605);
or UO_127 (O_127,N_2996,N_2933);
nand UO_128 (O_128,N_2850,N_2593);
or UO_129 (O_129,N_2553,N_2913);
nand UO_130 (O_130,N_2805,N_2812);
or UO_131 (O_131,N_2508,N_2919);
nand UO_132 (O_132,N_2898,N_2841);
xnor UO_133 (O_133,N_2836,N_2735);
nor UO_134 (O_134,N_2798,N_2744);
or UO_135 (O_135,N_2643,N_2815);
nor UO_136 (O_136,N_2675,N_2827);
or UO_137 (O_137,N_2543,N_2960);
nor UO_138 (O_138,N_2997,N_2755);
or UO_139 (O_139,N_2825,N_2999);
or UO_140 (O_140,N_2824,N_2625);
and UO_141 (O_141,N_2969,N_2734);
nand UO_142 (O_142,N_2525,N_2574);
nand UO_143 (O_143,N_2971,N_2951);
nand UO_144 (O_144,N_2917,N_2921);
nor UO_145 (O_145,N_2796,N_2743);
or UO_146 (O_146,N_2571,N_2718);
and UO_147 (O_147,N_2906,N_2550);
xor UO_148 (O_148,N_2621,N_2611);
xnor UO_149 (O_149,N_2900,N_2561);
nor UO_150 (O_150,N_2518,N_2934);
or UO_151 (O_151,N_2870,N_2899);
nor UO_152 (O_152,N_2507,N_2701);
or UO_153 (O_153,N_2922,N_2536);
nand UO_154 (O_154,N_2690,N_2646);
nand UO_155 (O_155,N_2756,N_2952);
nand UO_156 (O_156,N_2628,N_2630);
nand UO_157 (O_157,N_2608,N_2817);
nand UO_158 (O_158,N_2703,N_2577);
nor UO_159 (O_159,N_2883,N_2528);
nor UO_160 (O_160,N_2882,N_2941);
and UO_161 (O_161,N_2555,N_2816);
nand UO_162 (O_162,N_2833,N_2715);
nand UO_163 (O_163,N_2979,N_2838);
nor UO_164 (O_164,N_2694,N_2894);
nor UO_165 (O_165,N_2504,N_2749);
or UO_166 (O_166,N_2931,N_2832);
and UO_167 (O_167,N_2975,N_2661);
nand UO_168 (O_168,N_2781,N_2662);
nor UO_169 (O_169,N_2595,N_2665);
and UO_170 (O_170,N_2667,N_2678);
nor UO_171 (O_171,N_2672,N_2509);
and UO_172 (O_172,N_2622,N_2521);
nand UO_173 (O_173,N_2612,N_2757);
nand UO_174 (O_174,N_2943,N_2772);
nand UO_175 (O_175,N_2945,N_2585);
nor UO_176 (O_176,N_2637,N_2871);
nand UO_177 (O_177,N_2569,N_2910);
or UO_178 (O_178,N_2881,N_2776);
or UO_179 (O_179,N_2619,N_2855);
and UO_180 (O_180,N_2562,N_2914);
nor UO_181 (O_181,N_2936,N_2903);
or UO_182 (O_182,N_2724,N_2610);
nand UO_183 (O_183,N_2765,N_2890);
nand UO_184 (O_184,N_2858,N_2670);
and UO_185 (O_185,N_2523,N_2785);
nand UO_186 (O_186,N_2727,N_2990);
and UO_187 (O_187,N_2758,N_2880);
nand UO_188 (O_188,N_2674,N_2806);
and UO_189 (O_189,N_2515,N_2991);
and UO_190 (O_190,N_2992,N_2926);
nor UO_191 (O_191,N_2856,N_2546);
and UO_192 (O_192,N_2866,N_2811);
or UO_193 (O_193,N_2826,N_2519);
nand UO_194 (O_194,N_2586,N_2738);
nand UO_195 (O_195,N_2954,N_2966);
or UO_196 (O_196,N_2773,N_2531);
nor UO_197 (O_197,N_2911,N_2923);
nand UO_198 (O_198,N_2849,N_2551);
nor UO_199 (O_199,N_2642,N_2538);
and UO_200 (O_200,N_2594,N_2600);
and UO_201 (O_201,N_2947,N_2944);
nand UO_202 (O_202,N_2582,N_2644);
nand UO_203 (O_203,N_2986,N_2784);
or UO_204 (O_204,N_2723,N_2752);
and UO_205 (O_205,N_2650,N_2973);
nand UO_206 (O_206,N_2683,N_2962);
and UO_207 (O_207,N_2946,N_2801);
and UO_208 (O_208,N_2566,N_2719);
or UO_209 (O_209,N_2864,N_2668);
nor UO_210 (O_210,N_2925,N_2895);
nand UO_211 (O_211,N_2706,N_2616);
and UO_212 (O_212,N_2721,N_2563);
nor UO_213 (O_213,N_2754,N_2647);
nand UO_214 (O_214,N_2629,N_2869);
and UO_215 (O_215,N_2714,N_2810);
and UO_216 (O_216,N_2552,N_2976);
nor UO_217 (O_217,N_2581,N_2787);
or UO_218 (O_218,N_2840,N_2905);
nor UO_219 (O_219,N_2984,N_2658);
and UO_220 (O_220,N_2789,N_2607);
nor UO_221 (O_221,N_2872,N_2792);
or UO_222 (O_222,N_2843,N_2691);
or UO_223 (O_223,N_2961,N_2854);
or UO_224 (O_224,N_2513,N_2782);
or UO_225 (O_225,N_2641,N_2545);
and UO_226 (O_226,N_2892,N_2888);
nor UO_227 (O_227,N_2939,N_2733);
or UO_228 (O_228,N_2679,N_2626);
nor UO_229 (O_229,N_2788,N_2955);
and UO_230 (O_230,N_2904,N_2688);
or UO_231 (O_231,N_2592,N_2948);
and UO_232 (O_232,N_2868,N_2988);
nor UO_233 (O_233,N_2634,N_2729);
or UO_234 (O_234,N_2994,N_2684);
or UO_235 (O_235,N_2916,N_2928);
nor UO_236 (O_236,N_2682,N_2664);
and UO_237 (O_237,N_2813,N_2862);
or UO_238 (O_238,N_2863,N_2740);
and UO_239 (O_239,N_2549,N_2767);
nand UO_240 (O_240,N_2726,N_2875);
nor UO_241 (O_241,N_2790,N_2980);
or UO_242 (O_242,N_2516,N_2652);
or UO_243 (O_243,N_2799,N_2502);
nand UO_244 (O_244,N_2803,N_2778);
and UO_245 (O_245,N_2570,N_2692);
or UO_246 (O_246,N_2886,N_2640);
nor UO_247 (O_247,N_2623,N_2865);
nand UO_248 (O_248,N_2659,N_2938);
nand UO_249 (O_249,N_2932,N_2689);
and UO_250 (O_250,N_2791,N_2828);
or UO_251 (O_251,N_2989,N_2669);
and UO_252 (O_252,N_2948,N_2841);
and UO_253 (O_253,N_2584,N_2843);
nand UO_254 (O_254,N_2712,N_2730);
or UO_255 (O_255,N_2927,N_2525);
nand UO_256 (O_256,N_2888,N_2776);
nand UO_257 (O_257,N_2522,N_2912);
nand UO_258 (O_258,N_2519,N_2882);
nor UO_259 (O_259,N_2629,N_2842);
nor UO_260 (O_260,N_2899,N_2587);
or UO_261 (O_261,N_2736,N_2996);
nor UO_262 (O_262,N_2856,N_2538);
and UO_263 (O_263,N_2521,N_2774);
or UO_264 (O_264,N_2937,N_2789);
nor UO_265 (O_265,N_2638,N_2874);
nand UO_266 (O_266,N_2756,N_2613);
and UO_267 (O_267,N_2611,N_2944);
nand UO_268 (O_268,N_2599,N_2847);
nor UO_269 (O_269,N_2804,N_2509);
or UO_270 (O_270,N_2680,N_2763);
or UO_271 (O_271,N_2670,N_2750);
nand UO_272 (O_272,N_2881,N_2634);
nand UO_273 (O_273,N_2615,N_2560);
nand UO_274 (O_274,N_2888,N_2629);
nor UO_275 (O_275,N_2685,N_2562);
nor UO_276 (O_276,N_2679,N_2711);
nand UO_277 (O_277,N_2865,N_2915);
nand UO_278 (O_278,N_2996,N_2513);
or UO_279 (O_279,N_2673,N_2720);
nand UO_280 (O_280,N_2638,N_2972);
nor UO_281 (O_281,N_2588,N_2825);
nor UO_282 (O_282,N_2830,N_2983);
nor UO_283 (O_283,N_2954,N_2647);
nand UO_284 (O_284,N_2702,N_2635);
or UO_285 (O_285,N_2854,N_2759);
or UO_286 (O_286,N_2635,N_2528);
or UO_287 (O_287,N_2649,N_2982);
and UO_288 (O_288,N_2569,N_2802);
nor UO_289 (O_289,N_2731,N_2953);
nand UO_290 (O_290,N_2857,N_2829);
nand UO_291 (O_291,N_2659,N_2952);
nand UO_292 (O_292,N_2594,N_2557);
and UO_293 (O_293,N_2796,N_2870);
nor UO_294 (O_294,N_2666,N_2669);
or UO_295 (O_295,N_2599,N_2745);
nor UO_296 (O_296,N_2653,N_2759);
or UO_297 (O_297,N_2723,N_2826);
nor UO_298 (O_298,N_2990,N_2847);
and UO_299 (O_299,N_2836,N_2896);
and UO_300 (O_300,N_2840,N_2900);
and UO_301 (O_301,N_2893,N_2549);
nand UO_302 (O_302,N_2851,N_2763);
nor UO_303 (O_303,N_2983,N_2982);
nor UO_304 (O_304,N_2504,N_2763);
or UO_305 (O_305,N_2938,N_2787);
nand UO_306 (O_306,N_2768,N_2595);
xor UO_307 (O_307,N_2934,N_2999);
and UO_308 (O_308,N_2537,N_2857);
or UO_309 (O_309,N_2788,N_2669);
and UO_310 (O_310,N_2598,N_2789);
nand UO_311 (O_311,N_2656,N_2770);
and UO_312 (O_312,N_2894,N_2883);
nand UO_313 (O_313,N_2799,N_2537);
nor UO_314 (O_314,N_2585,N_2636);
nor UO_315 (O_315,N_2632,N_2817);
nor UO_316 (O_316,N_2546,N_2805);
nand UO_317 (O_317,N_2542,N_2619);
nor UO_318 (O_318,N_2972,N_2843);
nor UO_319 (O_319,N_2509,N_2875);
nand UO_320 (O_320,N_2928,N_2506);
nand UO_321 (O_321,N_2627,N_2865);
nor UO_322 (O_322,N_2748,N_2888);
or UO_323 (O_323,N_2982,N_2757);
or UO_324 (O_324,N_2673,N_2549);
nand UO_325 (O_325,N_2853,N_2791);
or UO_326 (O_326,N_2593,N_2883);
and UO_327 (O_327,N_2877,N_2976);
and UO_328 (O_328,N_2813,N_2518);
nor UO_329 (O_329,N_2564,N_2602);
nand UO_330 (O_330,N_2752,N_2575);
nor UO_331 (O_331,N_2805,N_2517);
and UO_332 (O_332,N_2865,N_2546);
and UO_333 (O_333,N_2527,N_2793);
nor UO_334 (O_334,N_2786,N_2732);
nand UO_335 (O_335,N_2853,N_2854);
or UO_336 (O_336,N_2912,N_2569);
and UO_337 (O_337,N_2597,N_2954);
nand UO_338 (O_338,N_2604,N_2742);
or UO_339 (O_339,N_2640,N_2677);
and UO_340 (O_340,N_2978,N_2536);
and UO_341 (O_341,N_2854,N_2833);
nand UO_342 (O_342,N_2717,N_2562);
or UO_343 (O_343,N_2514,N_2541);
or UO_344 (O_344,N_2630,N_2832);
or UO_345 (O_345,N_2985,N_2632);
and UO_346 (O_346,N_2838,N_2613);
and UO_347 (O_347,N_2919,N_2700);
nor UO_348 (O_348,N_2740,N_2640);
and UO_349 (O_349,N_2581,N_2922);
nand UO_350 (O_350,N_2892,N_2951);
or UO_351 (O_351,N_2641,N_2943);
or UO_352 (O_352,N_2889,N_2892);
or UO_353 (O_353,N_2825,N_2751);
nor UO_354 (O_354,N_2785,N_2783);
and UO_355 (O_355,N_2965,N_2697);
nand UO_356 (O_356,N_2779,N_2568);
nor UO_357 (O_357,N_2646,N_2655);
nor UO_358 (O_358,N_2618,N_2502);
nor UO_359 (O_359,N_2613,N_2842);
nand UO_360 (O_360,N_2858,N_2837);
nor UO_361 (O_361,N_2731,N_2597);
and UO_362 (O_362,N_2919,N_2707);
and UO_363 (O_363,N_2580,N_2609);
and UO_364 (O_364,N_2670,N_2957);
and UO_365 (O_365,N_2664,N_2736);
nand UO_366 (O_366,N_2730,N_2529);
or UO_367 (O_367,N_2577,N_2506);
or UO_368 (O_368,N_2819,N_2665);
nor UO_369 (O_369,N_2829,N_2657);
and UO_370 (O_370,N_2799,N_2528);
or UO_371 (O_371,N_2621,N_2674);
nand UO_372 (O_372,N_2946,N_2794);
and UO_373 (O_373,N_2588,N_2551);
and UO_374 (O_374,N_2954,N_2515);
and UO_375 (O_375,N_2760,N_2671);
or UO_376 (O_376,N_2913,N_2586);
nand UO_377 (O_377,N_2657,N_2879);
nand UO_378 (O_378,N_2898,N_2803);
nand UO_379 (O_379,N_2866,N_2865);
or UO_380 (O_380,N_2993,N_2880);
and UO_381 (O_381,N_2734,N_2996);
nor UO_382 (O_382,N_2869,N_2998);
nor UO_383 (O_383,N_2809,N_2894);
or UO_384 (O_384,N_2554,N_2632);
and UO_385 (O_385,N_2788,N_2711);
nand UO_386 (O_386,N_2518,N_2506);
and UO_387 (O_387,N_2575,N_2845);
or UO_388 (O_388,N_2973,N_2633);
xnor UO_389 (O_389,N_2628,N_2713);
or UO_390 (O_390,N_2681,N_2843);
and UO_391 (O_391,N_2646,N_2566);
or UO_392 (O_392,N_2547,N_2567);
and UO_393 (O_393,N_2914,N_2837);
or UO_394 (O_394,N_2680,N_2750);
nor UO_395 (O_395,N_2513,N_2592);
or UO_396 (O_396,N_2955,N_2606);
nor UO_397 (O_397,N_2870,N_2842);
nor UO_398 (O_398,N_2551,N_2637);
and UO_399 (O_399,N_2517,N_2959);
or UO_400 (O_400,N_2596,N_2523);
nand UO_401 (O_401,N_2781,N_2724);
nand UO_402 (O_402,N_2509,N_2905);
and UO_403 (O_403,N_2920,N_2779);
nand UO_404 (O_404,N_2779,N_2923);
and UO_405 (O_405,N_2714,N_2528);
or UO_406 (O_406,N_2918,N_2980);
nand UO_407 (O_407,N_2806,N_2631);
or UO_408 (O_408,N_2500,N_2802);
or UO_409 (O_409,N_2786,N_2724);
nor UO_410 (O_410,N_2924,N_2543);
and UO_411 (O_411,N_2804,N_2727);
and UO_412 (O_412,N_2750,N_2520);
or UO_413 (O_413,N_2855,N_2777);
and UO_414 (O_414,N_2661,N_2738);
nor UO_415 (O_415,N_2575,N_2542);
or UO_416 (O_416,N_2760,N_2809);
and UO_417 (O_417,N_2561,N_2564);
and UO_418 (O_418,N_2987,N_2616);
and UO_419 (O_419,N_2911,N_2710);
nor UO_420 (O_420,N_2736,N_2521);
and UO_421 (O_421,N_2717,N_2977);
or UO_422 (O_422,N_2786,N_2605);
nand UO_423 (O_423,N_2938,N_2841);
and UO_424 (O_424,N_2657,N_2765);
nor UO_425 (O_425,N_2680,N_2656);
and UO_426 (O_426,N_2808,N_2996);
nor UO_427 (O_427,N_2608,N_2582);
nor UO_428 (O_428,N_2910,N_2795);
or UO_429 (O_429,N_2535,N_2819);
or UO_430 (O_430,N_2764,N_2779);
xor UO_431 (O_431,N_2672,N_2514);
or UO_432 (O_432,N_2929,N_2837);
and UO_433 (O_433,N_2934,N_2504);
or UO_434 (O_434,N_2550,N_2647);
or UO_435 (O_435,N_2619,N_2810);
nor UO_436 (O_436,N_2932,N_2959);
and UO_437 (O_437,N_2796,N_2653);
and UO_438 (O_438,N_2688,N_2529);
nand UO_439 (O_439,N_2736,N_2539);
nor UO_440 (O_440,N_2874,N_2674);
nor UO_441 (O_441,N_2719,N_2822);
and UO_442 (O_442,N_2527,N_2720);
and UO_443 (O_443,N_2667,N_2664);
or UO_444 (O_444,N_2627,N_2788);
and UO_445 (O_445,N_2635,N_2994);
nor UO_446 (O_446,N_2758,N_2607);
and UO_447 (O_447,N_2984,N_2720);
or UO_448 (O_448,N_2501,N_2605);
nand UO_449 (O_449,N_2745,N_2998);
or UO_450 (O_450,N_2868,N_2916);
nand UO_451 (O_451,N_2589,N_2868);
nor UO_452 (O_452,N_2938,N_2531);
nand UO_453 (O_453,N_2881,N_2563);
nand UO_454 (O_454,N_2534,N_2847);
or UO_455 (O_455,N_2630,N_2899);
and UO_456 (O_456,N_2621,N_2992);
nor UO_457 (O_457,N_2641,N_2742);
or UO_458 (O_458,N_2619,N_2841);
and UO_459 (O_459,N_2525,N_2833);
nor UO_460 (O_460,N_2770,N_2698);
nor UO_461 (O_461,N_2863,N_2690);
and UO_462 (O_462,N_2986,N_2899);
nand UO_463 (O_463,N_2802,N_2870);
nor UO_464 (O_464,N_2655,N_2716);
nor UO_465 (O_465,N_2829,N_2914);
nand UO_466 (O_466,N_2528,N_2622);
or UO_467 (O_467,N_2790,N_2605);
nor UO_468 (O_468,N_2787,N_2606);
nand UO_469 (O_469,N_2839,N_2517);
nor UO_470 (O_470,N_2637,N_2902);
nand UO_471 (O_471,N_2682,N_2877);
nor UO_472 (O_472,N_2890,N_2881);
nor UO_473 (O_473,N_2771,N_2853);
nor UO_474 (O_474,N_2840,N_2793);
nor UO_475 (O_475,N_2988,N_2705);
nand UO_476 (O_476,N_2604,N_2632);
and UO_477 (O_477,N_2764,N_2952);
and UO_478 (O_478,N_2769,N_2628);
nor UO_479 (O_479,N_2570,N_2896);
and UO_480 (O_480,N_2714,N_2584);
or UO_481 (O_481,N_2690,N_2883);
xor UO_482 (O_482,N_2904,N_2748);
nor UO_483 (O_483,N_2539,N_2748);
nand UO_484 (O_484,N_2812,N_2582);
and UO_485 (O_485,N_2672,N_2601);
or UO_486 (O_486,N_2926,N_2775);
or UO_487 (O_487,N_2817,N_2931);
nor UO_488 (O_488,N_2815,N_2864);
or UO_489 (O_489,N_2645,N_2719);
nand UO_490 (O_490,N_2537,N_2767);
or UO_491 (O_491,N_2954,N_2937);
nor UO_492 (O_492,N_2899,N_2872);
nor UO_493 (O_493,N_2539,N_2788);
nand UO_494 (O_494,N_2540,N_2778);
and UO_495 (O_495,N_2868,N_2775);
nor UO_496 (O_496,N_2982,N_2870);
and UO_497 (O_497,N_2600,N_2927);
nand UO_498 (O_498,N_2848,N_2899);
and UO_499 (O_499,N_2646,N_2782);
endmodule