module basic_2500_25000_3000_25_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
or U0 (N_0,In_1339,In_1857);
nand U1 (N_1,In_2268,In_2077);
nand U2 (N_2,In_436,In_400);
nor U3 (N_3,In_1254,In_2270);
nor U4 (N_4,In_2421,In_1234);
nor U5 (N_5,In_188,In_2351);
and U6 (N_6,In_2279,In_1594);
xnor U7 (N_7,In_344,In_1534);
nor U8 (N_8,In_870,In_633);
nand U9 (N_9,In_169,In_2127);
nor U10 (N_10,In_1579,In_1576);
nor U11 (N_11,In_1068,In_449);
nand U12 (N_12,In_1568,In_2125);
xnor U13 (N_13,In_1349,In_234);
and U14 (N_14,In_542,In_375);
xnor U15 (N_15,In_2018,In_259);
xnor U16 (N_16,In_108,In_2199);
nor U17 (N_17,In_2340,In_1500);
nand U18 (N_18,In_686,In_2083);
and U19 (N_19,In_226,In_2286);
nand U20 (N_20,In_256,In_1885);
xnor U21 (N_21,In_1750,In_693);
xnor U22 (N_22,In_648,In_2094);
or U23 (N_23,In_14,In_1716);
nor U24 (N_24,In_255,In_660);
and U25 (N_25,In_1914,In_2240);
or U26 (N_26,In_1869,In_1962);
xnor U27 (N_27,In_1940,In_1346);
nand U28 (N_28,In_273,In_293);
xor U29 (N_29,In_2449,In_1042);
xnor U30 (N_30,In_837,In_1693);
and U31 (N_31,In_1620,In_658);
or U32 (N_32,In_523,In_1676);
nand U33 (N_33,In_1867,In_1243);
nor U34 (N_34,In_219,In_2046);
xor U35 (N_35,In_1744,In_1470);
nor U36 (N_36,In_2092,In_865);
or U37 (N_37,In_1499,In_1416);
xor U38 (N_38,In_676,In_311);
nand U39 (N_39,In_284,In_906);
or U40 (N_40,In_1749,In_1069);
and U41 (N_41,In_1368,In_2005);
nand U42 (N_42,In_2350,In_2411);
xnor U43 (N_43,In_856,In_190);
or U44 (N_44,In_2362,In_2168);
or U45 (N_45,In_1810,In_401);
or U46 (N_46,In_1851,In_1226);
nor U47 (N_47,In_151,In_1561);
and U48 (N_48,In_1988,In_599);
nor U49 (N_49,In_2023,In_2395);
and U50 (N_50,In_1514,In_1753);
nor U51 (N_51,In_172,In_1722);
and U52 (N_52,In_2236,In_1235);
or U53 (N_53,In_1077,In_1502);
and U54 (N_54,In_777,In_1574);
and U55 (N_55,In_1972,In_930);
or U56 (N_56,In_2149,In_1682);
xnor U57 (N_57,In_1495,In_1560);
xnor U58 (N_58,In_174,In_965);
and U59 (N_59,In_427,In_1858);
or U60 (N_60,In_721,In_1327);
xnor U61 (N_61,In_520,In_350);
nor U62 (N_62,In_1591,In_141);
nand U63 (N_63,In_2133,In_1652);
xnor U64 (N_64,In_1442,In_943);
nor U65 (N_65,In_407,In_1218);
nor U66 (N_66,In_73,In_2123);
and U67 (N_67,In_1369,In_2266);
xor U68 (N_68,In_666,In_2310);
or U69 (N_69,In_211,In_1925);
xnor U70 (N_70,In_2100,In_46);
xnor U71 (N_71,In_1870,In_708);
and U72 (N_72,In_1755,In_602);
or U73 (N_73,In_388,In_1151);
or U74 (N_74,In_221,In_815);
xnor U75 (N_75,In_593,In_1609);
xnor U76 (N_76,In_2379,In_2304);
and U77 (N_77,In_307,In_963);
nor U78 (N_78,In_1191,In_1479);
or U79 (N_79,In_1100,In_244);
nand U80 (N_80,In_2162,In_2180);
nor U81 (N_81,In_208,In_765);
or U82 (N_82,In_331,In_1832);
xor U83 (N_83,In_371,In_2106);
or U84 (N_84,In_1912,In_497);
and U85 (N_85,In_2384,In_209);
or U86 (N_86,In_1712,In_1187);
xnor U87 (N_87,In_571,In_812);
and U88 (N_88,In_1643,In_555);
or U89 (N_89,In_966,In_1038);
or U90 (N_90,In_1548,In_1689);
or U91 (N_91,In_1381,In_161);
or U92 (N_92,In_1786,In_1094);
nand U93 (N_93,In_2035,In_2399);
and U94 (N_94,In_1505,In_196);
nor U95 (N_95,In_2434,In_2032);
xor U96 (N_96,In_1679,In_2397);
or U97 (N_97,In_61,In_128);
nand U98 (N_98,In_160,In_1586);
and U99 (N_99,In_1539,In_365);
xnor U100 (N_100,In_1792,In_1315);
nor U101 (N_101,In_1703,In_873);
xor U102 (N_102,In_897,In_839);
or U103 (N_103,In_1250,In_2488);
nor U104 (N_104,In_1565,In_90);
nor U105 (N_105,In_1549,In_10);
nand U106 (N_106,In_1907,In_451);
nand U107 (N_107,In_1185,In_31);
nand U108 (N_108,In_1660,In_2405);
or U109 (N_109,In_985,In_2481);
or U110 (N_110,In_1666,In_125);
nand U111 (N_111,In_1598,In_1093);
or U112 (N_112,In_127,In_1376);
nand U113 (N_113,In_1850,In_1312);
or U114 (N_114,In_1075,In_29);
xor U115 (N_115,In_265,In_247);
nand U116 (N_116,In_1326,In_788);
or U117 (N_117,In_1303,In_466);
xnor U118 (N_118,In_598,In_1039);
nand U119 (N_119,In_2110,In_2118);
nand U120 (N_120,In_2060,In_691);
and U121 (N_121,In_422,In_460);
or U122 (N_122,In_2099,In_5);
nand U123 (N_123,In_737,In_2442);
and U124 (N_124,In_1866,In_2418);
or U125 (N_125,In_581,In_179);
nand U126 (N_126,In_527,In_1685);
and U127 (N_127,In_69,In_2489);
nand U128 (N_128,In_956,In_821);
nand U129 (N_129,In_1550,In_1302);
nand U130 (N_130,In_869,In_2081);
or U131 (N_131,In_463,In_1948);
or U132 (N_132,In_509,In_2020);
xor U133 (N_133,In_286,In_1415);
xor U134 (N_134,In_2355,In_2280);
nor U135 (N_135,In_175,In_356);
xnor U136 (N_136,In_1375,In_758);
or U137 (N_137,In_1709,In_1025);
nor U138 (N_138,In_1738,In_2471);
and U139 (N_139,In_1848,In_1783);
xnor U140 (N_140,In_780,In_1887);
and U141 (N_141,In_155,In_878);
or U142 (N_142,In_1814,In_2008);
nand U143 (N_143,In_855,In_1708);
or U144 (N_144,In_2055,In_516);
nand U145 (N_145,In_1966,In_1330);
or U146 (N_146,In_1820,In_1542);
or U147 (N_147,In_2239,In_102);
and U148 (N_148,In_752,In_1111);
nand U149 (N_149,In_409,In_1821);
xor U150 (N_150,In_1280,In_2329);
nand U151 (N_151,In_561,In_534);
nor U152 (N_152,In_884,In_1487);
or U153 (N_153,In_1868,In_2331);
and U154 (N_154,In_2215,In_1656);
and U155 (N_155,In_1190,In_1048);
and U156 (N_156,In_2370,In_2158);
xnor U157 (N_157,In_329,In_511);
and U158 (N_158,In_1941,In_40);
nand U159 (N_159,In_101,In_54);
or U160 (N_160,In_1872,In_352);
nor U161 (N_161,In_2145,In_1714);
nand U162 (N_162,In_2,In_149);
nand U163 (N_163,In_1704,In_305);
xnor U164 (N_164,In_601,In_2116);
and U165 (N_165,In_1454,In_280);
or U166 (N_166,In_1404,In_2166);
and U167 (N_167,In_2416,In_1189);
and U168 (N_168,In_672,In_1121);
and U169 (N_169,In_1472,In_1227);
or U170 (N_170,In_1232,In_1746);
xnor U171 (N_171,In_587,In_2157);
nand U172 (N_172,In_1958,In_2175);
and U173 (N_173,In_1041,In_1142);
and U174 (N_174,In_764,In_811);
or U175 (N_175,In_576,In_851);
xor U176 (N_176,In_1195,In_2438);
or U177 (N_177,In_146,In_1157);
or U178 (N_178,In_503,In_1913);
nor U179 (N_179,In_1634,In_1864);
or U180 (N_180,In_35,In_1604);
nor U181 (N_181,In_1959,In_2387);
xor U182 (N_182,In_1401,In_2378);
nand U183 (N_183,In_1840,In_917);
nor U184 (N_184,In_1691,In_1698);
or U185 (N_185,In_494,In_932);
xor U186 (N_186,In_899,In_2216);
xnor U187 (N_187,In_301,In_1555);
nor U188 (N_188,In_2204,In_421);
and U189 (N_189,In_2377,In_2021);
nor U190 (N_190,In_1469,In_1787);
and U191 (N_191,In_2206,In_382);
or U192 (N_192,In_1754,In_1137);
or U193 (N_193,In_1417,In_1603);
nor U194 (N_194,In_989,In_616);
nor U195 (N_195,In_15,In_584);
and U196 (N_196,In_281,In_349);
and U197 (N_197,In_2320,In_1937);
nor U198 (N_198,In_1646,In_1182);
and U199 (N_199,In_1970,In_1992);
nor U200 (N_200,In_113,In_1950);
nand U201 (N_201,In_1338,In_1461);
or U202 (N_202,In_292,In_982);
nand U203 (N_203,In_448,In_639);
xnor U204 (N_204,In_607,In_2235);
nor U205 (N_205,In_1529,In_354);
nor U206 (N_206,In_1455,In_2051);
xor U207 (N_207,In_786,In_701);
nand U208 (N_208,In_1447,In_1117);
nor U209 (N_209,In_1481,In_1888);
xnor U210 (N_210,In_1440,In_1730);
xor U211 (N_211,In_2446,In_66);
nand U212 (N_212,In_2171,In_718);
xor U213 (N_213,In_597,In_1158);
xnor U214 (N_214,In_1425,In_557);
xnor U215 (N_215,In_1406,In_37);
xor U216 (N_216,In_1238,In_1518);
and U217 (N_217,In_1874,In_1700);
or U218 (N_218,In_6,In_1762);
and U219 (N_219,In_590,In_620);
or U220 (N_220,In_1740,In_2097);
nor U221 (N_221,In_694,In_1806);
xnor U222 (N_222,In_1103,In_1323);
or U223 (N_223,In_166,In_1990);
xor U224 (N_224,In_1997,In_2181);
nor U225 (N_225,In_501,In_302);
xor U226 (N_226,In_1952,In_1337);
xnor U227 (N_227,In_1927,In_975);
nor U228 (N_228,In_696,In_2187);
xor U229 (N_229,In_774,In_670);
or U230 (N_230,In_204,In_1268);
xnor U231 (N_231,In_960,In_359);
nor U232 (N_232,In_1489,In_2102);
or U233 (N_233,In_1732,In_2154);
and U234 (N_234,In_617,In_1181);
or U235 (N_235,In_2385,In_2332);
or U236 (N_236,In_1116,In_1996);
xor U237 (N_237,In_419,In_1004);
nand U238 (N_238,In_2152,In_197);
xnor U239 (N_239,In_1233,In_1272);
xor U240 (N_240,In_1544,In_106);
nor U241 (N_241,In_1702,In_1706);
xor U242 (N_242,In_2334,In_2381);
nor U243 (N_243,In_1654,In_791);
and U244 (N_244,In_1681,In_714);
nor U245 (N_245,In_1955,In_1162);
xnor U246 (N_246,In_2009,In_236);
nor U247 (N_247,In_1031,In_689);
nor U248 (N_248,In_182,In_2183);
and U249 (N_249,In_1199,In_339);
and U250 (N_250,In_1605,In_1006);
nor U251 (N_251,In_1715,In_1322);
or U252 (N_252,In_1519,In_2232);
nand U253 (N_253,In_486,In_4);
xor U254 (N_254,In_1793,In_114);
xnor U255 (N_255,In_353,In_1072);
nor U256 (N_256,In_430,In_778);
xor U257 (N_257,In_546,In_261);
and U258 (N_258,In_944,In_628);
or U259 (N_259,In_1379,In_673);
xor U260 (N_260,In_988,In_1699);
and U261 (N_261,In_541,In_1552);
and U262 (N_262,In_1017,In_1623);
xor U263 (N_263,In_684,In_1733);
nor U264 (N_264,In_1405,In_2321);
and U265 (N_265,In_755,In_2044);
nand U266 (N_266,In_336,In_1220);
nor U267 (N_267,In_1289,In_2228);
and U268 (N_268,In_2307,In_475);
nand U269 (N_269,In_25,In_1908);
xnor U270 (N_270,In_540,In_1192);
xor U271 (N_271,In_1729,In_1266);
and U272 (N_272,In_1432,In_251);
and U273 (N_273,In_1766,In_1611);
nand U274 (N_274,In_2347,In_1240);
nor U275 (N_275,In_2289,In_818);
xor U276 (N_276,In_1491,In_665);
or U277 (N_277,In_1541,In_589);
or U278 (N_278,In_194,In_2042);
nor U279 (N_279,In_195,In_168);
xor U280 (N_280,In_435,In_1822);
or U281 (N_281,In_1807,In_1998);
xor U282 (N_282,In_332,In_2432);
xnor U283 (N_283,In_799,In_1843);
or U284 (N_284,In_1528,In_173);
xnor U285 (N_285,In_220,In_2074);
or U286 (N_286,In_913,In_2207);
and U287 (N_287,In_1933,In_1587);
xor U288 (N_288,In_785,In_1758);
nand U289 (N_289,In_1828,In_1597);
nor U290 (N_290,In_2062,In_641);
nor U291 (N_291,In_1517,In_386);
nor U292 (N_292,In_2041,In_861);
nand U293 (N_293,In_1278,In_1569);
xnor U294 (N_294,In_1893,In_1370);
and U295 (N_295,In_2262,In_2463);
or U296 (N_296,In_1015,In_751);
nor U297 (N_297,In_1136,In_2372);
xor U298 (N_298,In_1148,In_1956);
and U299 (N_299,In_1483,In_2271);
xnor U300 (N_300,In_1979,In_1304);
nand U301 (N_301,In_1924,In_834);
and U302 (N_302,In_1471,In_1207);
nand U303 (N_303,In_2079,In_447);
and U304 (N_304,In_2417,In_1677);
xor U305 (N_305,In_465,In_16);
nand U306 (N_306,In_1855,In_1882);
xnor U307 (N_307,In_804,In_2452);
xor U308 (N_308,In_1581,In_453);
and U309 (N_309,In_1779,In_1366);
nor U310 (N_310,In_2160,In_1036);
nor U311 (N_311,In_1836,In_2288);
xor U312 (N_312,In_1589,In_2223);
and U313 (N_313,In_502,In_2484);
and U314 (N_314,In_1089,In_133);
nor U315 (N_315,In_817,In_759);
nand U316 (N_316,In_1396,In_411);
xor U317 (N_317,In_176,In_1985);
and U318 (N_318,In_1949,In_2038);
nand U319 (N_319,In_846,In_2169);
nor U320 (N_320,In_748,In_1477);
xor U321 (N_321,In_1206,In_1824);
nor U322 (N_322,In_183,In_2324);
nand U323 (N_323,In_802,In_1661);
and U324 (N_324,In_213,In_827);
nor U325 (N_325,In_2193,In_1357);
and U326 (N_326,In_1551,In_950);
nand U327 (N_327,In_493,In_96);
xor U328 (N_328,In_1834,In_2210);
xor U329 (N_329,In_1902,In_2230);
nor U330 (N_330,In_1064,In_2265);
xor U331 (N_331,In_2052,In_585);
and U332 (N_332,In_1649,In_116);
nand U333 (N_333,In_715,In_2337);
xor U334 (N_334,In_309,In_1301);
nor U335 (N_335,In_872,In_374);
xor U336 (N_336,In_2076,In_1065);
and U337 (N_337,In_1389,In_1987);
or U338 (N_338,In_901,In_2058);
nand U339 (N_339,In_318,In_333);
and U340 (N_340,In_2354,In_1674);
nand U341 (N_341,In_1983,In_768);
or U342 (N_342,In_2172,In_1102);
and U343 (N_343,In_253,In_120);
xnor U344 (N_344,In_2170,In_1080);
or U345 (N_345,In_446,In_813);
or U346 (N_346,In_562,In_406);
nor U347 (N_347,In_2495,In_363);
xor U348 (N_348,In_568,In_51);
nor U349 (N_349,In_140,In_1718);
xor U350 (N_350,In_158,In_2349);
or U351 (N_351,In_287,In_2364);
nor U352 (N_352,In_1044,In_1827);
and U353 (N_353,In_1939,In_2292);
xor U354 (N_354,In_1147,In_2365);
or U355 (N_355,In_2333,In_822);
nand U356 (N_356,In_1745,In_1865);
and U357 (N_357,In_367,In_2469);
xnor U358 (N_358,In_1797,In_1001);
or U359 (N_359,In_1663,In_2080);
and U360 (N_360,In_2194,In_1600);
or U361 (N_361,In_1314,In_482);
or U362 (N_362,In_2410,In_863);
nor U363 (N_363,In_789,In_1149);
or U364 (N_364,In_1450,In_549);
nor U365 (N_365,In_2155,In_1653);
or U366 (N_366,In_1493,In_1256);
or U367 (N_367,In_2454,In_2264);
xor U368 (N_368,In_1028,In_854);
and U369 (N_369,In_836,In_1647);
nand U370 (N_370,In_800,In_653);
nand U371 (N_371,In_2071,In_1784);
nor U372 (N_372,In_484,In_784);
nor U373 (N_373,In_1642,In_2444);
xnor U374 (N_374,In_1335,In_437);
xnor U375 (N_375,In_1826,In_2474);
xor U376 (N_376,In_558,In_70);
xor U377 (N_377,In_410,In_1134);
xor U378 (N_378,In_844,In_625);
xnor U379 (N_379,In_1991,In_1021);
nor U380 (N_380,In_797,In_1225);
xnor U381 (N_381,In_1558,In_1705);
nor U382 (N_382,In_2404,In_1911);
nor U383 (N_383,In_2226,In_723);
nor U384 (N_384,In_2121,In_986);
nor U385 (N_385,In_1763,In_747);
nor U386 (N_386,In_1119,In_875);
or U387 (N_387,In_1767,In_376);
nand U388 (N_388,In_2108,In_24);
xor U389 (N_389,In_608,In_99);
xor U390 (N_390,In_2208,In_1593);
nor U391 (N_391,In_728,In_680);
nand U392 (N_392,In_2390,In_1537);
nor U393 (N_393,In_1607,In_1683);
nand U394 (N_394,In_1967,In_1723);
and U395 (N_395,In_766,In_299);
xnor U396 (N_396,In_583,In_1270);
or U397 (N_397,In_2394,In_726);
nand U398 (N_398,In_1411,In_842);
nor U399 (N_399,In_1115,In_1971);
nor U400 (N_400,In_1473,In_2140);
nor U401 (N_401,In_7,In_2001);
nand U402 (N_402,In_1362,In_122);
or U403 (N_403,In_79,In_2316);
nor U404 (N_404,In_184,In_252);
nand U405 (N_405,In_959,In_1391);
nor U406 (N_406,In_1894,In_1960);
and U407 (N_407,In_1143,In_277);
xnor U408 (N_408,In_1348,In_2440);
nor U409 (N_409,In_2217,In_115);
nor U410 (N_410,In_880,In_1486);
nand U411 (N_411,In_1079,In_1965);
nor U412 (N_412,In_1774,In_958);
xor U413 (N_413,In_574,In_1359);
nor U414 (N_414,In_519,In_1878);
and U415 (N_415,In_2222,In_1221);
nor U416 (N_416,In_1394,In_1790);
xnor U417 (N_417,In_1575,In_1980);
and U418 (N_418,In_2408,In_150);
nand U419 (N_419,In_488,In_738);
or U420 (N_420,In_849,In_560);
xor U421 (N_421,In_548,In_2195);
xnor U422 (N_422,In_937,In_1515);
nor U423 (N_423,In_2298,In_9);
nand U424 (N_424,In_2209,In_631);
and U425 (N_425,In_951,In_2451);
nand U426 (N_426,In_682,In_808);
nand U427 (N_427,In_330,In_2027);
nor U428 (N_428,In_2253,In_2415);
or U429 (N_429,In_2276,In_1946);
xor U430 (N_430,In_566,In_1687);
xor U431 (N_431,In_304,In_2016);
nand U432 (N_432,In_278,In_983);
or U433 (N_433,In_471,In_327);
nor U434 (N_434,In_1099,In_1764);
or U435 (N_435,In_1193,In_1005);
and U436 (N_436,In_1186,In_603);
nor U437 (N_437,In_2082,In_713);
nand U438 (N_438,In_1367,In_423);
nand U439 (N_439,In_912,In_1881);
or U440 (N_440,In_806,In_142);
nand U441 (N_441,In_2352,In_1167);
nor U442 (N_442,In_2414,In_993);
nand U443 (N_443,In_328,In_769);
and U444 (N_444,In_1222,In_1854);
nand U445 (N_445,In_1944,In_954);
xnor U446 (N_446,In_227,In_1049);
or U447 (N_447,In_2095,In_1352);
or U448 (N_448,In_1659,In_762);
xnor U449 (N_449,In_2360,In_415);
or U450 (N_450,In_1808,In_1695);
and U451 (N_451,In_1897,In_1782);
nor U452 (N_452,In_2000,In_105);
or U453 (N_453,In_1385,In_925);
nor U454 (N_454,In_1583,In_1769);
and U455 (N_455,In_319,In_2497);
xnor U456 (N_456,In_734,In_1059);
or U457 (N_457,In_1686,In_644);
or U458 (N_458,In_2087,In_425);
nand U459 (N_459,In_144,In_2294);
and U460 (N_460,In_823,In_746);
xor U461 (N_461,In_1994,In_1978);
or U462 (N_462,In_1619,In_725);
nand U463 (N_463,In_2382,In_1295);
or U464 (N_464,In_403,In_1976);
or U465 (N_465,In_1169,In_2202);
nor U466 (N_466,In_1131,In_1785);
and U467 (N_467,In_32,In_654);
xnor U468 (N_468,In_271,In_2141);
and U469 (N_469,In_835,In_1070);
and U470 (N_470,In_586,In_2012);
nand U471 (N_471,In_2243,In_1928);
xnor U472 (N_472,In_62,In_205);
nand U473 (N_473,In_829,In_1743);
xnor U474 (N_474,In_1237,In_1636);
nor U475 (N_475,In_1125,In_121);
nand U476 (N_476,In_1443,In_968);
nor U477 (N_477,In_1175,In_941);
nand U478 (N_478,In_2067,In_1331);
nand U479 (N_479,In_634,In_392);
xor U480 (N_480,In_1756,In_1298);
xnor U481 (N_481,In_1128,In_20);
or U482 (N_482,In_17,In_2260);
nand U483 (N_483,In_2031,In_266);
nor U484 (N_484,In_904,In_544);
nor U485 (N_485,In_2425,In_347);
nand U486 (N_486,In_185,In_888);
and U487 (N_487,In_798,In_889);
or U488 (N_488,In_2356,In_1176);
nand U489 (N_489,In_1420,In_338);
xnor U490 (N_490,In_651,In_1215);
nor U491 (N_491,In_1951,In_1239);
nand U492 (N_492,In_1961,In_2098);
xor U493 (N_493,In_903,In_698);
nand U494 (N_494,In_82,In_1291);
and U495 (N_495,In_2348,In_1061);
xnor U496 (N_496,In_826,In_454);
xnor U497 (N_497,In_891,In_1906);
xnor U498 (N_498,In_1856,In_1501);
xnor U499 (N_499,In_1513,In_2156);
nand U500 (N_500,In_543,In_1274);
nor U501 (N_501,In_2251,In_979);
nor U502 (N_502,In_383,In_1805);
and U503 (N_503,In_75,In_1617);
and U504 (N_504,In_615,In_577);
and U505 (N_505,In_1585,In_1794);
nor U506 (N_506,In_348,In_595);
nor U507 (N_507,In_2419,In_2103);
or U508 (N_508,In_189,In_1113);
nand U509 (N_509,In_907,In_820);
or U510 (N_510,In_2259,In_514);
nand U511 (N_511,In_1612,In_559);
xor U512 (N_512,In_2091,In_635);
nand U513 (N_513,In_1648,In_1353);
nand U514 (N_514,In_1088,In_588);
nand U515 (N_515,In_1651,In_874);
nand U516 (N_516,In_877,In_629);
or U517 (N_517,In_1920,In_1325);
nor U518 (N_518,In_2174,In_2011);
nand U519 (N_519,In_1484,In_775);
and U520 (N_520,In_2290,In_72);
nor U521 (N_521,In_1150,In_2420);
nor U522 (N_522,In_1091,In_2441);
or U523 (N_523,In_2109,In_2492);
or U524 (N_524,In_1839,In_2433);
nor U525 (N_525,In_1252,In_722);
and U526 (N_526,In_1588,In_377);
or U527 (N_527,In_742,In_59);
or U528 (N_528,In_398,In_1871);
nand U529 (N_529,In_1286,In_345);
xnor U530 (N_530,In_1178,In_2003);
and U531 (N_531,In_1285,In_1123);
nand U532 (N_532,In_1403,In_1726);
nor U533 (N_533,In_76,In_717);
nor U534 (N_534,In_2478,In_624);
xor U535 (N_535,In_908,In_1707);
xor U536 (N_536,In_312,In_36);
xnor U537 (N_537,In_1347,In_2330);
nand U538 (N_538,In_22,In_2479);
xor U539 (N_539,In_893,In_1577);
nand U540 (N_540,In_1290,In_91);
nand U541 (N_541,In_1875,In_469);
nand U542 (N_542,In_268,In_1110);
and U543 (N_543,In_729,In_687);
or U544 (N_544,In_2255,In_380);
nor U545 (N_545,In_563,In_942);
nor U546 (N_546,In_1640,In_2112);
or U547 (N_547,In_2148,In_1737);
or U548 (N_548,In_712,In_1208);
or U549 (N_549,In_413,In_927);
and U550 (N_550,In_1204,In_1511);
nor U551 (N_551,In_663,In_11);
or U552 (N_552,In_228,In_1196);
nand U553 (N_553,In_47,In_805);
nor U554 (N_554,In_1374,In_1400);
nand U555 (N_555,In_250,In_1632);
nand U556 (N_556,In_1900,In_1294);
nand U557 (N_557,In_496,In_522);
xor U558 (N_558,In_2338,In_1361);
nor U559 (N_559,In_887,In_2299);
xor U560 (N_560,In_2246,In_1921);
nand U561 (N_561,In_193,In_1496);
nor U562 (N_562,In_1557,In_935);
and U563 (N_563,In_1371,In_2269);
and U564 (N_564,In_1863,In_372);
or U565 (N_565,In_2325,In_1267);
nor U566 (N_566,In_2128,In_67);
xnor U567 (N_567,In_355,In_1022);
or U568 (N_568,In_860,In_2460);
or U569 (N_569,In_1441,In_604);
xnor U570 (N_570,In_2482,In_2291);
xnor U571 (N_571,In_433,In_1333);
or U572 (N_572,In_929,In_63);
xor U573 (N_573,In_1761,In_2458);
nor U574 (N_574,In_1624,In_1719);
or U575 (N_575,In_1156,In_2115);
nand U576 (N_576,In_655,In_1580);
or U577 (N_577,In_1465,In_2254);
nand U578 (N_578,In_2165,In_2173);
nor U579 (N_579,In_1212,In_978);
nand U580 (N_580,In_1141,In_2412);
nor U581 (N_581,In_491,In_1424);
xnor U582 (N_582,In_2105,In_2138);
or U583 (N_583,In_500,In_1884);
and U584 (N_584,In_248,In_235);
nand U585 (N_585,In_1688,In_2499);
or U586 (N_586,In_848,In_1019);
and U587 (N_587,In_360,In_2459);
and U588 (N_588,In_109,In_163);
xnor U589 (N_589,In_1492,In_346);
nor U590 (N_590,In_2007,In_2326);
nor U591 (N_591,In_2462,In_2258);
nand U592 (N_592,In_2429,In_1669);
xor U593 (N_593,In_760,In_1122);
or U594 (N_594,In_987,In_325);
or U595 (N_595,In_1462,In_528);
nand U596 (N_596,In_1800,In_532);
and U597 (N_597,In_1553,In_80);
nor U598 (N_598,In_882,In_241);
nand U599 (N_599,In_1510,In_1236);
and U600 (N_600,In_2143,In_1608);
or U601 (N_601,In_2150,In_1916);
xor U602 (N_602,In_2498,In_89);
xor U603 (N_603,In_1444,In_2006);
or U604 (N_604,In_2197,In_618);
nand U605 (N_605,In_810,In_1108);
and U606 (N_606,In_1482,In_1823);
nor U607 (N_607,In_1350,In_896);
xor U608 (N_608,In_1410,In_1963);
and U609 (N_609,In_1795,In_1328);
xnor U610 (N_610,In_2318,In_1018);
and U611 (N_611,In_2078,In_424);
and U612 (N_612,In_1090,In_1255);
and U613 (N_613,In_290,In_735);
or U614 (N_614,In_683,In_2319);
or U615 (N_615,In_1317,In_64);
xor U616 (N_616,In_1200,In_1000);
nand U617 (N_617,In_1095,In_740);
nor U618 (N_618,In_773,In_326);
and U619 (N_619,In_2263,In_1942);
xor U620 (N_620,In_1596,In_110);
and U621 (N_621,In_1650,In_2113);
xnor U622 (N_622,In_1747,In_341);
nor U623 (N_623,In_656,In_506);
or U624 (N_624,In_743,In_1426);
nand U625 (N_625,In_779,In_2391);
and U626 (N_626,In_432,In_892);
and U627 (N_627,In_2147,In_864);
xor U628 (N_628,In_2369,In_1098);
xor U629 (N_629,In_60,In_1701);
nor U630 (N_630,In_2376,In_643);
or U631 (N_631,In_1414,In_134);
xnor U632 (N_632,In_853,In_2037);
nand U633 (N_633,In_1096,In_1527);
xnor U634 (N_634,In_2424,In_2201);
and U635 (N_635,In_1035,In_218);
and U636 (N_636,In_704,In_1936);
or U637 (N_637,In_947,In_1164);
nand U638 (N_638,In_1056,In_117);
nor U639 (N_639,In_294,In_711);
xnor U640 (N_640,In_313,In_1665);
nand U641 (N_641,In_2443,In_1710);
nand U642 (N_642,In_1087,In_269);
xor U643 (N_643,In_1265,In_1393);
xor U644 (N_644,In_1264,In_2392);
and U645 (N_645,In_2069,In_709);
nand U646 (N_646,In_2466,In_1690);
nand U647 (N_647,In_1336,In_498);
nor U648 (N_648,In_551,In_1584);
nor U649 (N_649,In_2026,In_2303);
nand U650 (N_650,In_1757,In_1803);
nand U651 (N_651,In_1083,In_1132);
nor U652 (N_652,In_1862,In_2114);
and U653 (N_653,In_1435,In_1407);
or U654 (N_654,In_801,In_2457);
xor U655 (N_655,In_171,In_443);
xnor U656 (N_656,In_404,In_2389);
nor U657 (N_657,In_1316,In_2363);
nand U658 (N_658,In_2167,In_1421);
nor U659 (N_659,In_230,In_1572);
xor U660 (N_660,In_1051,In_1271);
and U661 (N_661,In_1344,In_1439);
and U662 (N_662,In_55,In_1107);
nor U663 (N_663,In_2407,In_611);
and U664 (N_664,In_1343,In_2019);
nor U665 (N_665,In_2196,In_749);
nand U666 (N_666,In_2437,In_610);
xor U667 (N_667,In_2144,In_1667);
xnor U668 (N_668,In_1340,In_1935);
nor U669 (N_669,In_914,In_1898);
nand U670 (N_670,In_202,In_198);
nand U671 (N_671,In_1139,In_1436);
and U672 (N_672,In_1082,In_2053);
or U673 (N_673,In_613,In_369);
nor U674 (N_674,In_1380,In_736);
or U675 (N_675,In_547,In_531);
or U676 (N_676,In_1024,In_156);
or U677 (N_677,In_1023,In_1860);
xnor U678 (N_678,In_1802,In_859);
xor U679 (N_679,In_2252,In_2430);
nand U680 (N_680,In_391,In_707);
nor U681 (N_681,In_2485,In_1886);
or U682 (N_682,In_2233,In_154);
nand U683 (N_683,In_1242,In_262);
xnor U684 (N_684,In_1045,In_2423);
and U685 (N_685,In_1168,In_254);
and U686 (N_686,In_2122,In_481);
xnor U687 (N_687,In_65,In_902);
nor U688 (N_688,In_1974,In_187);
xor U689 (N_689,In_1890,In_476);
xor U690 (N_690,In_1345,In_456);
xnor U691 (N_691,In_1844,In_1727);
and U692 (N_692,In_1109,In_2072);
nand U693 (N_693,In_2335,In_885);
nor U694 (N_694,In_129,In_678);
xnor U695 (N_695,In_894,In_342);
and U696 (N_696,In_1533,In_1466);
and U697 (N_697,In_890,In_1030);
xnor U698 (N_698,In_145,In_793);
nand U699 (N_699,In_373,In_1480);
xor U700 (N_700,In_487,In_621);
nor U701 (N_701,In_45,In_2059);
nor U702 (N_702,In_1320,In_2297);
and U703 (N_703,In_2132,In_1458);
nand U704 (N_704,In_1248,In_1504);
or U705 (N_705,In_485,In_1986);
nand U706 (N_706,In_480,In_868);
nor U707 (N_707,In_2361,In_229);
xor U708 (N_708,In_1358,In_2342);
xor U709 (N_709,In_1982,In_632);
nand U710 (N_710,In_961,In_135);
and U711 (N_711,In_1259,In_2277);
xnor U712 (N_712,In_1262,In_2311);
xor U713 (N_713,In_1684,In_1644);
nor U714 (N_714,In_792,In_1214);
and U715 (N_715,In_1402,In_2422);
nand U716 (N_716,In_1635,In_1060);
nor U717 (N_717,In_2244,In_852);
and U718 (N_718,In_1364,In_282);
nand U719 (N_719,In_402,In_1163);
xor U720 (N_720,In_879,In_776);
nor U721 (N_721,In_1880,In_973);
and U722 (N_722,In_1621,In_2135);
nor U723 (N_723,In_1748,In_1696);
xor U724 (N_724,In_2388,In_468);
and U725 (N_725,In_1395,In_1664);
xor U726 (N_726,In_1478,In_1628);
nand U727 (N_727,In_2309,In_1434);
and U728 (N_728,In_2427,In_1717);
or U729 (N_729,In_838,In_1382);
nand U730 (N_730,In_1662,In_1126);
xnor U731 (N_731,In_981,In_2475);
nor U732 (N_732,In_2163,In_2192);
xnor U733 (N_733,In_667,In_2017);
xnor U734 (N_734,In_1788,In_596);
and U735 (N_735,In_1188,In_2101);
nor U736 (N_736,In_1120,In_1734);
and U737 (N_737,In_841,In_553);
nand U738 (N_738,In_630,In_124);
nor U739 (N_739,In_1523,In_2345);
and U740 (N_740,In_317,In_662);
xor U741 (N_741,In_136,In_969);
and U742 (N_742,In_1773,In_1475);
nor U743 (N_743,In_900,In_1130);
or U744 (N_744,In_450,In_2313);
xor U745 (N_745,In_905,In_1852);
nor U746 (N_746,In_1768,In_1171);
and U747 (N_747,In_1697,In_77);
xnor U748 (N_748,In_2054,In_782);
xor U749 (N_749,In_1845,In_2257);
xnor U750 (N_750,In_384,In_472);
or U751 (N_751,In_1463,In_323);
or U752 (N_752,In_2346,In_957);
xor U753 (N_753,In_2045,In_28);
or U754 (N_754,In_700,In_1520);
or U755 (N_755,In_1431,In_2130);
nor U756 (N_756,In_831,In_393);
xnor U757 (N_757,In_41,In_1356);
or U758 (N_758,In_2028,In_924);
nor U759 (N_759,In_107,In_1058);
or U760 (N_760,In_232,In_1297);
and U761 (N_761,In_1672,In_970);
xnor U762 (N_762,In_1287,In_1835);
nand U763 (N_763,In_2131,In_1307);
nor U764 (N_764,In_119,In_1390);
nand U765 (N_765,In_362,In_1599);
xor U766 (N_766,In_1341,In_1751);
nor U767 (N_767,In_2341,In_535);
nand U768 (N_768,In_920,In_685);
nand U769 (N_769,In_803,In_1841);
or U770 (N_770,In_1926,In_1525);
xor U771 (N_771,In_408,In_690);
nor U772 (N_772,In_513,In_761);
xnor U773 (N_773,In_2242,In_2464);
or U774 (N_774,In_1046,In_1071);
or U775 (N_775,In_1507,In_216);
and U776 (N_776,In_847,In_1273);
nor U777 (N_777,In_669,In_1546);
nor U778 (N_778,In_1556,In_1033);
nor U779 (N_779,In_2490,In_1245);
or U780 (N_780,In_2476,In_1209);
and U781 (N_781,In_949,In_1645);
nor U782 (N_782,In_972,In_1321);
nand U783 (N_783,In_2056,In_1180);
xnor U784 (N_784,In_572,In_138);
or U785 (N_785,In_1896,In_2402);
nand U786 (N_786,In_1947,In_2050);
nand U787 (N_787,In_2426,In_1261);
nand U788 (N_788,In_1713,In_1050);
or U789 (N_789,In_2075,In_1127);
and U790 (N_790,In_1571,In_1815);
or U791 (N_791,In_300,In_224);
or U792 (N_792,In_2164,In_2400);
nor U793 (N_793,In_640,In_2119);
nor U794 (N_794,In_18,In_1968);
nand U795 (N_795,In_898,In_1459);
or U796 (N_796,In_1318,In_470);
nand U797 (N_797,In_272,In_1076);
nor U798 (N_798,In_1825,In_2487);
and U799 (N_799,In_971,In_2090);
xnor U800 (N_800,In_570,In_1067);
nor U801 (N_801,In_98,In_1283);
nor U802 (N_802,In_675,In_308);
nor U803 (N_803,In_275,In_2126);
and U804 (N_804,In_763,In_2151);
and U805 (N_805,In_1306,In_1741);
nand U806 (N_806,In_34,In_1263);
nor U807 (N_807,In_214,In_1363);
nand U808 (N_808,In_2491,In_2322);
nand U809 (N_809,In_1053,In_614);
xor U810 (N_810,In_2344,In_922);
xor U811 (N_811,In_26,In_1711);
and U812 (N_812,In_1485,In_2049);
nand U813 (N_813,In_1354,In_744);
nand U814 (N_814,In_1509,In_147);
xor U815 (N_815,In_2179,In_1910);
xor U816 (N_816,In_412,In_1626);
or U817 (N_817,In_1288,In_1154);
nand U818 (N_818,In_337,In_1251);
or U819 (N_819,In_1673,In_455);
and U820 (N_820,In_1428,In_533);
and U821 (N_821,In_1010,In_1837);
and U822 (N_822,In_637,In_2285);
or U823 (N_823,In_233,In_2225);
nor U824 (N_824,In_2153,In_1230);
and U825 (N_825,In_385,In_71);
or U826 (N_826,In_1721,In_237);
and U827 (N_827,In_668,In_2436);
nand U828 (N_828,In_1918,In_1977);
nand U829 (N_829,In_1995,In_754);
or U830 (N_830,In_191,In_1203);
and U831 (N_831,In_39,In_2409);
nor U832 (N_832,In_212,In_258);
nand U833 (N_833,In_681,In_442);
or U834 (N_834,In_716,In_1299);
xnor U835 (N_835,In_1922,In_94);
xnor U836 (N_836,In_2136,In_967);
and U837 (N_837,In_2403,In_1813);
and U838 (N_838,In_515,In_2191);
and U839 (N_839,In_1276,In_2010);
or U840 (N_840,In_2312,In_2205);
nand U841 (N_841,In_926,In_953);
xor U842 (N_842,In_461,In_980);
and U843 (N_843,In_592,In_1413);
nand U844 (N_844,In_1638,In_2029);
xor U845 (N_845,In_1931,In_0);
or U846 (N_846,In_948,In_2189);
xor U847 (N_847,In_833,In_322);
or U848 (N_848,In_2431,In_490);
xor U849 (N_849,In_1819,In_170);
or U850 (N_850,In_270,In_1037);
or U851 (N_851,In_1742,In_1559);
and U852 (N_852,In_2358,In_2439);
xnor U853 (N_853,In_2480,In_1817);
or U854 (N_854,In_2456,In_1838);
nor U855 (N_855,In_118,In_1543);
nor U856 (N_856,In_368,In_940);
xor U857 (N_857,In_606,In_1789);
nor U858 (N_858,In_1905,In_2025);
and U859 (N_859,In_2040,In_2366);
nor U860 (N_860,In_517,In_510);
or U861 (N_861,In_2357,In_569);
and U862 (N_862,In_1097,In_1989);
xor U863 (N_863,In_1903,In_1675);
nor U864 (N_864,In_38,In_867);
or U865 (N_865,In_19,In_1174);
nand U866 (N_866,In_1488,In_659);
or U867 (N_867,In_215,In_30);
nand U868 (N_868,In_1818,In_1144);
or U869 (N_869,In_2287,In_438);
or U870 (N_870,In_444,In_1724);
and U871 (N_871,In_1231,In_13);
xnor U872 (N_872,In_2182,In_1249);
and U873 (N_873,In_2039,In_911);
nor U874 (N_874,In_492,In_504);
nand U875 (N_875,In_207,In_1213);
xor U876 (N_876,In_2301,In_1430);
nor U877 (N_877,In_824,In_1975);
and U878 (N_878,In_1772,In_1614);
and U879 (N_879,In_321,In_964);
nand U880 (N_880,In_387,In_1224);
nand U881 (N_881,In_231,In_1412);
nor U882 (N_882,In_1873,In_2227);
and U883 (N_883,In_1508,In_1876);
or U884 (N_884,In_1476,In_795);
nand U885 (N_885,In_103,In_999);
or U886 (N_886,In_2470,In_1388);
nand U887 (N_887,In_1160,In_809);
nand U888 (N_888,In_249,In_1999);
nor U889 (N_889,In_2142,In_2124);
and U890 (N_890,In_157,In_2129);
or U891 (N_891,In_671,In_1879);
nand U892 (N_892,In_111,In_159);
nand U893 (N_893,In_396,In_1165);
and U894 (N_894,In_1601,In_1198);
nor U895 (N_895,In_830,In_2486);
nor U896 (N_896,In_623,In_816);
and U897 (N_897,In_2111,In_2296);
nand U898 (N_898,In_545,In_767);
and U899 (N_899,In_1205,In_2184);
and U900 (N_900,In_1247,In_2117);
or U901 (N_901,In_938,In_439);
and U902 (N_902,In_2406,In_1329);
xor U903 (N_903,In_1833,In_753);
nor U904 (N_904,In_324,In_85);
and U905 (N_905,In_131,In_1631);
xnor U906 (N_906,In_1981,In_2314);
and U907 (N_907,In_2096,In_1678);
and U908 (N_908,In_2448,In_1383);
xnor U909 (N_909,In_1637,In_1812);
or U910 (N_910,In_1625,In_1152);
or U911 (N_911,In_1279,In_334);
and U912 (N_912,In_274,In_1012);
or U913 (N_913,In_1610,In_206);
nor U914 (N_914,In_1360,In_390);
or U915 (N_915,In_962,In_2014);
or U916 (N_916,In_2461,In_536);
xnor U917 (N_917,In_2219,In_1521);
xnor U918 (N_918,In_361,In_2241);
nand U919 (N_919,In_936,In_2413);
and U920 (N_920,In_567,In_1114);
and U921 (N_921,In_1047,In_858);
nand U922 (N_922,In_1324,In_756);
nor U923 (N_923,In_739,In_1081);
nor U924 (N_924,In_167,In_2146);
nand U925 (N_925,In_524,In_931);
and U926 (N_926,In_1002,In_1013);
nor U927 (N_927,In_2468,In_130);
xor U928 (N_928,In_1210,In_222);
xnor U929 (N_929,In_242,In_378);
xnor U930 (N_930,In_794,In_2339);
nand U931 (N_931,In_1201,In_741);
nand U932 (N_932,In_2066,In_2493);
and U933 (N_933,In_474,In_1145);
xor U934 (N_934,In_955,In_2359);
nor U935 (N_935,In_1217,In_825);
nand U936 (N_936,In_2089,In_289);
and U937 (N_937,In_479,In_1101);
nor U938 (N_938,In_2004,In_1798);
xor U939 (N_939,In_165,In_2057);
and U940 (N_940,In_2278,In_674);
nand U941 (N_941,In_638,In_994);
nor U942 (N_942,In_1427,In_526);
nor U943 (N_943,In_695,In_1602);
or U944 (N_944,In_649,In_1526);
nand U945 (N_945,In_1258,In_2161);
or U946 (N_946,In_2328,In_1451);
xor U947 (N_947,In_467,In_1630);
or U948 (N_948,In_2343,In_2336);
or U949 (N_949,In_2084,In_1847);
and U950 (N_950,In_1140,In_279);
nand U951 (N_951,In_612,In_458);
or U952 (N_952,In_1135,In_2247);
nor U953 (N_953,In_1244,In_370);
and U954 (N_954,In_2002,In_389);
nand U955 (N_955,In_1849,In_622);
or U956 (N_956,In_1883,In_1173);
nor U957 (N_957,In_1310,In_2295);
or U958 (N_958,In_591,In_554);
and U959 (N_959,In_2398,In_923);
nand U960 (N_960,In_609,In_181);
xnor U961 (N_961,In_358,In_720);
or U962 (N_962,In_1530,In_1536);
or U963 (N_963,In_2088,In_1177);
and U964 (N_964,In_225,In_291);
xor U965 (N_965,In_910,In_100);
nand U966 (N_966,In_462,In_2317);
nor U967 (N_967,In_1892,In_1468);
and U968 (N_968,In_819,In_1564);
nand U969 (N_969,In_2267,In_1153);
or U970 (N_970,In_733,In_1464);
xor U971 (N_971,In_1448,In_1969);
or U972 (N_972,In_1112,In_850);
nand U973 (N_973,In_2465,In_1457);
and U974 (N_974,In_1964,In_137);
or U975 (N_975,In_2190,In_1026);
or U976 (N_976,In_2159,In_58);
or U977 (N_977,In_2323,In_518);
or U978 (N_978,In_990,In_1895);
or U979 (N_979,In_445,In_335);
or U980 (N_980,In_394,In_692);
and U981 (N_981,In_217,In_1277);
xor U982 (N_982,In_2300,In_48);
nor U983 (N_983,In_731,In_783);
nand U984 (N_984,In_1437,In_2275);
nor U985 (N_985,In_1538,In_508);
nor U986 (N_986,In_2450,In_647);
xnor U987 (N_987,In_1146,In_1032);
and U988 (N_988,In_2047,In_977);
nand U989 (N_989,In_1029,In_2186);
nor U990 (N_990,In_2386,In_2211);
and U991 (N_991,In_1954,In_1535);
nand U992 (N_992,In_74,In_1055);
or U993 (N_993,In_2022,In_52);
and U994 (N_994,In_1408,In_1775);
nand U995 (N_995,In_87,In_578);
nor U996 (N_996,In_1453,In_2435);
nor U997 (N_997,In_1211,In_1904);
nor U998 (N_998,In_1429,In_1460);
and U999 (N_999,In_2048,In_2063);
nor U1000 (N_1000,In_2229,N_659);
nor U1001 (N_1001,In_50,N_962);
and U1002 (N_1002,N_423,N_984);
or U1003 (N_1003,N_167,N_360);
nor U1004 (N_1004,In_1796,N_637);
nor U1005 (N_1005,In_727,In_95);
or U1006 (N_1006,N_623,N_965);
nor U1007 (N_1007,N_925,N_671);
and U1008 (N_1008,N_81,In_1319);
or U1009 (N_1009,N_933,N_688);
nor U1010 (N_1010,In_2375,N_705);
and U1011 (N_1011,N_924,N_567);
xnor U1012 (N_1012,N_38,N_416);
and U1013 (N_1013,In_529,N_900);
xor U1014 (N_1014,In_1801,N_472);
nor U1015 (N_1015,In_1957,N_452);
nand U1016 (N_1016,N_8,N_55);
and U1017 (N_1017,N_583,In_1229);
xnor U1018 (N_1018,N_304,N_836);
or U1019 (N_1019,N_752,In_895);
nand U1020 (N_1020,In_2218,In_770);
nor U1021 (N_1021,N_996,In_582);
xor U1022 (N_1022,N_830,N_297);
xnor U1023 (N_1023,In_2185,In_457);
xnor U1024 (N_1024,In_1066,N_676);
nand U1025 (N_1025,N_331,In_645);
nor U1026 (N_1026,N_200,N_683);
xnor U1027 (N_1027,N_34,In_1973);
nand U1028 (N_1028,N_308,In_1446);
xnor U1029 (N_1029,N_600,N_832);
and U1030 (N_1030,N_231,In_556);
or U1031 (N_1031,N_458,In_2371);
nor U1032 (N_1032,In_2188,In_871);
and U1033 (N_1033,N_440,N_233);
and U1034 (N_1034,In_303,N_376);
and U1035 (N_1035,N_222,In_1494);
nand U1036 (N_1036,In_1084,In_1334);
nand U1037 (N_1037,N_929,N_873);
xor U1038 (N_1038,N_427,In_1313);
xnor U1039 (N_1039,N_298,N_74);
nand U1040 (N_1040,In_790,N_151);
xor U1041 (N_1041,N_382,N_554);
or U1042 (N_1042,In_1804,N_442);
xnor U1043 (N_1043,N_299,N_886);
and U1044 (N_1044,N_588,N_111);
nor U1045 (N_1045,N_837,In_1104);
and U1046 (N_1046,N_301,N_461);
and U1047 (N_1047,N_257,In_405);
nand U1048 (N_1048,N_727,In_2401);
xor U1049 (N_1049,N_692,In_126);
and U1050 (N_1050,In_1452,N_644);
xnor U1051 (N_1051,N_765,N_205);
or U1052 (N_1052,N_168,N_796);
nand U1053 (N_1053,N_214,N_669);
or U1054 (N_1054,In_418,In_2107);
and U1055 (N_1055,In_730,N_920);
or U1056 (N_1056,In_706,N_101);
and U1057 (N_1057,N_485,N_280);
nand U1058 (N_1058,In_2373,In_1027);
xnor U1059 (N_1059,N_718,N_244);
or U1060 (N_1060,N_123,N_621);
nor U1061 (N_1061,N_534,N_916);
and U1062 (N_1062,N_690,In_2198);
and U1063 (N_1063,In_2065,N_358);
and U1064 (N_1064,In_605,N_456);
nand U1065 (N_1065,N_310,In_2380);
nand U1066 (N_1066,N_820,N_327);
xor U1067 (N_1067,In_512,In_652);
and U1068 (N_1068,N_682,N_763);
or U1069 (N_1069,N_236,N_569);
xnor U1070 (N_1070,In_1811,N_707);
or U1071 (N_1071,In_240,In_1655);
or U1072 (N_1072,N_26,N_894);
or U1073 (N_1073,N_895,N_29);
nand U1074 (N_1074,N_322,N_164);
and U1075 (N_1075,N_856,In_2467);
and U1076 (N_1076,In_2374,N_328);
nor U1077 (N_1077,In_2237,N_468);
nor U1078 (N_1078,In_2302,N_253);
or U1079 (N_1079,N_291,In_1889);
or U1080 (N_1080,N_50,N_961);
or U1081 (N_1081,N_861,N_343);
nor U1082 (N_1082,N_383,N_444);
xor U1083 (N_1083,N_911,In_1909);
nand U1084 (N_1084,N_77,In_1627);
and U1085 (N_1085,N_872,N_59);
nand U1086 (N_1086,N_899,N_636);
or U1087 (N_1087,N_364,N_309);
and U1088 (N_1088,In_2221,N_585);
xor U1089 (N_1089,In_1671,N_119);
nor U1090 (N_1090,N_125,In_340);
nor U1091 (N_1091,N_704,In_246);
xnor U1092 (N_1092,In_796,N_724);
nand U1093 (N_1093,N_448,N_450);
and U1094 (N_1094,In_1342,N_457);
or U1095 (N_1095,In_1670,In_1384);
xnor U1096 (N_1096,N_212,N_580);
and U1097 (N_1097,In_1456,N_991);
and U1098 (N_1098,In_186,In_192);
nand U1099 (N_1099,N_194,N_238);
nor U1100 (N_1100,In_697,N_481);
xnor U1101 (N_1101,In_43,N_968);
xor U1102 (N_1102,N_699,N_654);
nor U1103 (N_1103,In_1919,In_139);
nand U1104 (N_1104,N_694,N_435);
and U1105 (N_1105,In_781,N_797);
or U1106 (N_1106,In_1816,N_766);
xor U1107 (N_1107,In_507,N_201);
nand U1108 (N_1108,N_777,N_875);
nand U1109 (N_1109,In_1993,In_1293);
nand U1110 (N_1110,N_728,N_935);
nand U1111 (N_1111,N_32,N_169);
nand U1112 (N_1112,N_436,N_957);
and U1113 (N_1113,N_180,N_323);
nand U1114 (N_1114,N_192,N_104);
nor U1115 (N_1115,In_1074,N_197);
xor U1116 (N_1116,N_650,N_843);
or U1117 (N_1117,N_878,N_264);
xnor U1118 (N_1118,N_187,In_1197);
nor U1119 (N_1119,N_283,N_143);
or U1120 (N_1120,N_88,N_473);
and U1121 (N_1121,N_234,N_869);
nand U1122 (N_1122,In_565,In_1275);
or U1123 (N_1123,N_272,N_782);
nor U1124 (N_1124,N_801,N_702);
xnor U1125 (N_1125,In_1641,N_78);
xor U1126 (N_1126,In_1365,N_912);
or U1127 (N_1127,N_954,N_311);
and U1128 (N_1128,N_885,In_995);
and U1129 (N_1129,N_628,N_176);
nand U1130 (N_1130,N_386,In_946);
nor U1131 (N_1131,N_599,N_134);
nor U1132 (N_1132,N_446,In_1161);
nor U1133 (N_1133,N_516,N_206);
nand U1134 (N_1134,N_928,N_998);
and U1135 (N_1135,N_373,N_589);
nand U1136 (N_1136,N_3,In_1891);
or U1137 (N_1137,N_488,N_773);
and U1138 (N_1138,N_23,N_141);
nor U1139 (N_1139,N_983,N_825);
nor U1140 (N_1140,In_580,N_260);
or U1141 (N_1141,N_959,N_513);
nor U1142 (N_1142,In_2238,N_353);
or U1143 (N_1143,In_1281,N_161);
nand U1144 (N_1144,N_495,N_285);
nand U1145 (N_1145,N_767,N_384);
nor U1146 (N_1146,N_684,In_732);
and U1147 (N_1147,In_2383,In_399);
nor U1148 (N_1148,In_1054,N_73);
or U1149 (N_1149,In_2212,In_1945);
and U1150 (N_1150,N_235,N_1);
xnor U1151 (N_1151,In_1532,In_1092);
nand U1152 (N_1152,N_638,In_1377);
and U1153 (N_1153,In_379,N_131);
nand U1154 (N_1154,N_815,In_757);
or U1155 (N_1155,N_647,N_640);
and U1156 (N_1156,In_57,N_246);
and U1157 (N_1157,N_438,In_1567);
or U1158 (N_1158,N_145,N_336);
and U1159 (N_1159,In_1409,In_996);
nand U1160 (N_1160,N_598,In_357);
nand U1161 (N_1161,In_2033,In_2250);
xor U1162 (N_1162,In_2134,N_846);
nand U1163 (N_1163,In_164,N_806);
xor U1164 (N_1164,N_25,N_470);
or U1165 (N_1165,In_573,N_172);
nand U1166 (N_1166,N_30,N_421);
or U1167 (N_1167,N_956,N_918);
and U1168 (N_1168,N_594,In_661);
xor U1169 (N_1169,N_541,N_502);
or U1170 (N_1170,In_1522,In_2306);
nand U1171 (N_1171,In_1246,In_1765);
nor U1172 (N_1172,N_163,N_971);
and U1173 (N_1173,N_217,N_809);
and U1174 (N_1174,In_417,N_425);
or U1175 (N_1175,In_538,N_634);
or U1176 (N_1176,In_1570,In_1759);
or U1177 (N_1177,N_823,In_429);
and U1178 (N_1178,N_148,N_375);
nor U1179 (N_1179,N_678,N_276);
nand U1180 (N_1180,In_1923,In_1622);
and U1181 (N_1181,N_409,N_731);
xnor U1182 (N_1182,N_133,N_223);
nor U1183 (N_1183,N_91,N_35);
nand U1184 (N_1184,N_658,N_320);
xnor U1185 (N_1185,In_239,N_635);
nor U1186 (N_1186,N_279,N_687);
or U1187 (N_1187,In_1399,N_715);
nor U1188 (N_1188,In_1257,In_295);
nor U1189 (N_1189,N_615,In_2061);
or U1190 (N_1190,In_1387,N_219);
nand U1191 (N_1191,N_735,N_651);
xnor U1192 (N_1192,N_275,N_854);
nand U1193 (N_1193,In_260,N_207);
or U1194 (N_1194,N_760,N_330);
nand U1195 (N_1195,N_430,N_712);
or U1196 (N_1196,In_1842,N_14);
nor U1197 (N_1197,N_958,N_818);
nand U1198 (N_1198,In_364,N_392);
xor U1199 (N_1199,In_984,N_410);
and U1200 (N_1200,N_547,N_190);
xnor U1201 (N_1201,N_969,In_2305);
nor U1202 (N_1202,N_144,N_904);
xnor U1203 (N_1203,N_431,N_946);
and U1204 (N_1204,N_708,N_839);
nand U1205 (N_1205,In_1770,N_695);
xor U1206 (N_1206,In_945,N_936);
and U1207 (N_1207,N_986,In_1490);
nand U1208 (N_1208,In_86,N_942);
xor U1209 (N_1209,N_483,In_416);
nand U1210 (N_1210,N_879,In_2293);
and U1211 (N_1211,N_188,N_494);
and U1212 (N_1212,N_56,In_921);
nor U1213 (N_1213,N_261,N_390);
xor U1214 (N_1214,N_706,N_910);
nand U1215 (N_1215,N_867,In_223);
nor U1216 (N_1216,In_1932,N_371);
and U1217 (N_1217,N_582,N_913);
nor U1218 (N_1218,In_1085,N_573);
and U1219 (N_1219,In_245,In_1498);
and U1220 (N_1220,N_95,N_892);
or U1221 (N_1221,N_967,N_793);
xnor U1222 (N_1222,N_509,N_124);
nand U1223 (N_1223,N_697,In_203);
and U1224 (N_1224,In_162,N_814);
or U1225 (N_1225,N_155,N_855);
and U1226 (N_1226,N_531,N_645);
or U1227 (N_1227,N_514,In_2393);
and U1228 (N_1228,N_833,N_787);
and U1229 (N_1229,In_366,N_403);
nand U1230 (N_1230,In_2093,In_1859);
nor U1231 (N_1231,N_528,N_98);
nor U1232 (N_1232,In_2030,N_114);
xor U1233 (N_1233,N_496,N_432);
or U1234 (N_1234,N_117,In_1595);
xor U1235 (N_1235,N_917,In_123);
nor U1236 (N_1236,N_11,N_173);
or U1237 (N_1237,N_587,N_147);
or U1238 (N_1238,N_213,N_366);
nor U1239 (N_1239,N_783,In_267);
nor U1240 (N_1240,N_94,N_351);
nand U1241 (N_1241,N_893,In_1592);
and U1242 (N_1242,N_730,N_964);
xnor U1243 (N_1243,N_762,N_824);
nand U1244 (N_1244,N_443,N_550);
nand U1245 (N_1245,N_49,N_788);
or U1246 (N_1246,N_884,N_398);
nor U1247 (N_1247,In_1445,N_471);
xor U1248 (N_1248,N_743,In_1063);
nor U1249 (N_1249,In_1915,In_143);
nand U1250 (N_1250,In_1809,N_315);
and U1251 (N_1251,N_316,In_210);
and U1252 (N_1252,In_699,In_1618);
and U1253 (N_1253,In_3,In_1397);
xor U1254 (N_1254,N_252,In_594);
nor U1255 (N_1255,N_10,N_466);
nor U1256 (N_1256,N_868,In_1269);
xnor U1257 (N_1257,N_601,In_2231);
and U1258 (N_1258,In_2120,In_2137);
nand U1259 (N_1259,N_770,N_850);
xor U1260 (N_1260,N_510,N_520);
xor U1261 (N_1261,In_2496,N_953);
nand U1262 (N_1262,N_397,In_2445);
nand U1263 (N_1263,In_452,N_794);
nor U1264 (N_1264,N_296,N_539);
xor U1265 (N_1265,N_224,N_394);
or U1266 (N_1266,N_487,In_257);
nand U1267 (N_1267,N_838,N_237);
or U1268 (N_1268,N_858,N_527);
nor U1269 (N_1269,In_1613,In_657);
nand U1270 (N_1270,In_1953,N_877);
nor U1271 (N_1271,N_939,In_1778);
or U1272 (N_1272,In_1657,In_53);
xor U1273 (N_1273,N_726,N_52);
nand U1274 (N_1274,In_2024,N_198);
nand U1275 (N_1275,N_732,In_177);
nand U1276 (N_1276,N_862,In_288);
xnor U1277 (N_1277,In_1735,In_2064);
and U1278 (N_1278,N_250,N_37);
or U1279 (N_1279,In_1658,N_511);
nand U1280 (N_1280,N_307,In_1433);
and U1281 (N_1281,In_1129,In_539);
nor U1282 (N_1282,N_680,In_1007);
or U1283 (N_1283,N_860,N_691);
xnor U1284 (N_1284,N_980,N_749);
xor U1285 (N_1285,In_56,N_239);
and U1286 (N_1286,In_1355,In_2034);
or U1287 (N_1287,N_284,N_100);
and U1288 (N_1288,In_2013,N_191);
xor U1289 (N_1289,In_285,In_997);
nor U1290 (N_1290,In_8,N_734);
or U1291 (N_1291,N_548,N_2);
nor U1292 (N_1292,N_64,N_492);
nand U1293 (N_1293,N_372,N_48);
xor U1294 (N_1294,N_349,N_326);
nor U1295 (N_1295,N_247,N_245);
nor U1296 (N_1296,In_1917,N_632);
or U1297 (N_1297,N_553,In_886);
nand U1298 (N_1298,N_555,In_1194);
or U1299 (N_1299,N_666,In_1133);
or U1300 (N_1300,In_1791,N_278);
and U1301 (N_1301,N_480,N_719);
nor U1302 (N_1302,In_719,In_919);
nor U1303 (N_1303,In_1467,N_86);
or U1304 (N_1304,N_498,N_115);
nand U1305 (N_1305,N_993,N_604);
xnor U1306 (N_1306,N_748,N_350);
nor U1307 (N_1307,In_2224,N_211);
nor U1308 (N_1308,N_338,N_629);
xnor U1309 (N_1309,N_300,In_600);
nand U1310 (N_1310,In_1419,In_1003);
xnor U1311 (N_1311,N_887,N_419);
nor U1312 (N_1312,In_1,N_771);
nand U1313 (N_1313,N_69,In_473);
nand U1314 (N_1314,N_67,In_2213);
xnor U1315 (N_1315,N_464,In_1418);
or U1316 (N_1316,In_1138,In_104);
and U1317 (N_1317,In_1172,In_2473);
xor U1318 (N_1318,In_2281,N_288);
and U1319 (N_1319,N_515,In_1062);
xor U1320 (N_1320,N_947,N_714);
nor U1321 (N_1321,N_274,In_2139);
xnor U1322 (N_1322,In_710,In_1846);
nor U1323 (N_1323,In_1680,N_242);
nand U1324 (N_1324,N_324,N_677);
and U1325 (N_1325,N_158,N_761);
or U1326 (N_1326,N_68,In_42);
or U1327 (N_1327,N_60,N_13);
or U1328 (N_1328,N_630,N_566);
nor U1329 (N_1329,N_614,In_2353);
and U1330 (N_1330,N_340,N_344);
nor U1331 (N_1331,N_195,In_1547);
and U1332 (N_1332,N_926,N_533);
or U1333 (N_1333,N_411,N_227);
nand U1334 (N_1334,N_602,N_142);
nor U1335 (N_1335,In_495,In_2273);
and U1336 (N_1336,N_798,In_1516);
or U1337 (N_1337,In_1086,N_811);
and U1338 (N_1338,N_612,N_828);
xnor U1339 (N_1339,N_370,N_689);
or U1340 (N_1340,In_1578,N_179);
or U1341 (N_1341,N_290,In_1292);
nand U1342 (N_1342,In_1052,In_2447);
and U1343 (N_1343,N_551,In_1901);
and U1344 (N_1344,N_203,N_754);
nor U1345 (N_1345,N_150,N_624);
nand U1346 (N_1346,N_273,In_97);
or U1347 (N_1347,N_988,In_1183);
xnor U1348 (N_1348,N_778,N_292);
or U1349 (N_1349,In_1540,N_591);
or U1350 (N_1350,N_62,In_276);
nor U1351 (N_1351,N_329,N_717);
or U1352 (N_1352,N_518,In_1305);
xor U1353 (N_1353,N_166,In_397);
or U1354 (N_1354,In_1725,N_693);
nor U1355 (N_1355,N_22,In_1692);
xor U1356 (N_1356,In_2472,In_81);
or U1357 (N_1357,N_590,N_791);
or U1358 (N_1358,N_348,N_586);
nor U1359 (N_1359,N_16,N_361);
and U1360 (N_1360,N_345,N_903);
and U1361 (N_1361,N_625,N_199);
nor U1362 (N_1362,In_316,N_76);
or U1363 (N_1363,N_271,N_776);
nor U1364 (N_1364,N_93,N_422);
nand U1365 (N_1365,N_401,N_575);
nor U1366 (N_1366,In_428,N_96);
and U1367 (N_1367,N_467,In_2177);
xor U1368 (N_1368,N_122,N_816);
nand U1369 (N_1369,In_320,N_538);
nor U1370 (N_1370,N_126,N_407);
xnor U1371 (N_1371,N_129,N_226);
xor U1372 (N_1372,N_802,In_148);
or U1373 (N_1373,N_656,N_826);
nand U1374 (N_1374,N_611,In_1202);
and U1375 (N_1375,N_21,N_558);
or U1376 (N_1376,In_772,In_952);
or U1377 (N_1377,In_1398,N_426);
nor U1378 (N_1378,In_1831,N_46);
xor U1379 (N_1379,N_512,N_620);
or U1380 (N_1380,N_454,N_479);
and U1381 (N_1381,N_230,In_1554);
and U1382 (N_1382,N_396,In_1780);
xnor U1383 (N_1383,N_657,In_1506);
nor U1384 (N_1384,N_842,N_561);
or U1385 (N_1385,N_259,N_821);
nor U1386 (N_1386,N_453,N_500);
nor U1387 (N_1387,In_1720,N_503);
nor U1388 (N_1388,N_667,N_696);
and U1389 (N_1389,In_2245,N_646);
or U1390 (N_1390,N_408,N_840);
nor U1391 (N_1391,In_564,In_974);
nand U1392 (N_1392,N_429,In_992);
nand U1393 (N_1393,N_139,N_679);
and U1394 (N_1394,In_1590,In_2176);
xor U1395 (N_1395,N_412,N_757);
and U1396 (N_1396,In_1776,N_985);
nand U1397 (N_1397,N_342,In_1739);
nor U1398 (N_1398,N_741,N_943);
nand U1399 (N_1399,In_579,N_914);
nand U1400 (N_1400,N_149,N_932);
xnor U1401 (N_1401,In_489,N_922);
nor U1402 (N_1402,In_298,N_525);
or U1403 (N_1403,N_355,N_951);
or U1404 (N_1404,N_132,In_843);
nor U1405 (N_1405,In_1040,N_262);
nand U1406 (N_1406,N_156,N_759);
xnor U1407 (N_1407,N_42,In_1694);
xor U1408 (N_1408,In_750,N_889);
and U1409 (N_1409,N_152,In_12);
xnor U1410 (N_1410,In_499,N_622);
xor U1411 (N_1411,N_303,N_399);
xnor U1412 (N_1412,N_489,In_1545);
or U1413 (N_1413,N_507,N_109);
xnor U1414 (N_1414,N_774,In_976);
or U1415 (N_1415,N_75,N_803);
nand U1416 (N_1416,In_441,In_1777);
and U1417 (N_1417,N_750,N_381);
nor U1418 (N_1418,N_19,In_537);
nor U1419 (N_1419,N_389,N_966);
and U1420 (N_1420,N_451,N_817);
and U1421 (N_1421,N_701,N_822);
and U1422 (N_1422,N_15,N_536);
and U1423 (N_1423,In_283,N_995);
nand U1424 (N_1424,In_477,N_265);
xor U1425 (N_1425,N_805,N_930);
xnor U1426 (N_1426,N_359,N_116);
nor U1427 (N_1427,N_883,N_978);
nor U1428 (N_1428,N_529,N_295);
and U1429 (N_1429,N_848,N_263);
xnor U1430 (N_1430,In_866,N_356);
or U1431 (N_1431,In_2368,N_643);
and U1432 (N_1432,N_521,N_433);
and U1433 (N_1433,N_532,N_737);
nand U1434 (N_1434,N_989,N_576);
or U1435 (N_1435,In_201,N_474);
or U1436 (N_1436,N_661,N_919);
xor U1437 (N_1437,N_54,In_414);
nor U1438 (N_1438,N_110,N_792);
nor U1439 (N_1439,N_459,N_663);
xnor U1440 (N_1440,In_88,In_1300);
nor U1441 (N_1441,N_469,N_113);
xnor U1442 (N_1442,In_677,In_2282);
or U1443 (N_1443,N_901,N_41);
xnor U1444 (N_1444,In_459,N_321);
nand U1445 (N_1445,N_841,In_27);
nor U1446 (N_1446,In_1943,In_297);
xnor U1447 (N_1447,In_1166,N_834);
or U1448 (N_1448,N_723,N_546);
nor U1449 (N_1449,N_768,N_108);
nand U1450 (N_1450,N_58,N_225);
or U1451 (N_1451,In_2453,In_1309);
or U1452 (N_1452,N_53,In_2178);
nand U1453 (N_1453,N_347,N_670);
xnor U1454 (N_1454,In_1253,In_2086);
nor U1455 (N_1455,N_542,N_314);
nor U1456 (N_1456,In_1830,N_970);
nand U1457 (N_1457,In_2327,N_255);
or U1458 (N_1458,N_672,N_121);
xor U1459 (N_1459,N_790,N_388);
xnor U1460 (N_1460,N_595,In_1184);
xnor U1461 (N_1461,In_2284,N_103);
xor U1462 (N_1462,N_859,In_1582);
nand U1463 (N_1463,N_57,N_434);
and U1464 (N_1464,N_501,N_975);
nand U1465 (N_1465,N_387,N_477);
or U1466 (N_1466,In_343,In_1930);
nand U1467 (N_1467,N_758,N_949);
xnor U1468 (N_1468,N_313,N_18);
xnor U1469 (N_1469,N_6,N_9);
nor U1470 (N_1470,In_1562,In_2220);
xnor U1471 (N_1471,N_248,N_847);
and U1472 (N_1472,N_577,N_405);
nand U1473 (N_1473,N_317,N_333);
nor U1474 (N_1474,N_543,N_486);
or U1475 (N_1475,N_112,N_963);
nor U1476 (N_1476,N_346,In_1282);
nand U1477 (N_1477,In_1179,N_24);
nor U1478 (N_1478,In_1639,N_36);
xor U1479 (N_1479,N_92,In_1372);
nor U1480 (N_1480,In_2249,In_310);
or U1481 (N_1481,N_746,N_795);
nor U1482 (N_1482,N_153,In_1011);
nor U1483 (N_1483,N_574,N_742);
nand U1484 (N_1484,N_85,In_881);
xnor U1485 (N_1485,In_1159,N_530);
nand U1486 (N_1486,N_844,In_1118);
nor U1487 (N_1487,In_1829,N_537);
and U1488 (N_1488,N_559,In_1934);
xnor U1489 (N_1489,N_812,N_413);
nor U1490 (N_1490,N_999,N_228);
xnor U1491 (N_1491,N_979,N_385);
nor U1492 (N_1492,N_293,N_681);
nand U1493 (N_1493,N_404,N_269);
xor U1494 (N_1494,N_584,In_575);
xnor U1495 (N_1495,N_65,In_1563);
xnor U1496 (N_1496,N_47,N_138);
nor U1497 (N_1497,N_703,N_556);
nor U1498 (N_1498,N_420,N_713);
nand U1499 (N_1499,N_71,N_258);
or U1500 (N_1500,In_2261,N_987);
or U1501 (N_1501,N_437,N_720);
and U1502 (N_1502,N_931,In_702);
nor U1503 (N_1503,In_2428,N_655);
xor U1504 (N_1504,In_264,N_977);
nor U1505 (N_1505,N_921,In_44);
or U1506 (N_1506,In_1781,N_549);
and U1507 (N_1507,N_685,N_424);
or U1508 (N_1508,N_193,N_849);
or U1509 (N_1509,N_578,N_973);
nand U1510 (N_1510,N_908,In_1668);
and U1511 (N_1511,N_334,N_249);
nor U1512 (N_1512,N_365,N_606);
xnor U1513 (N_1513,N_552,N_981);
or U1514 (N_1514,In_152,In_296);
or U1515 (N_1515,In_2396,In_420);
xor U1516 (N_1516,N_952,N_415);
nand U1517 (N_1517,N_305,N_229);
nand U1518 (N_1518,N_170,In_1073);
or U1519 (N_1519,In_915,N_618);
or U1520 (N_1520,N_974,In_1008);
and U1521 (N_1521,N_475,N_445);
nor U1522 (N_1522,In_21,In_1106);
or U1523 (N_1523,N_905,N_617);
xnor U1524 (N_1524,N_597,In_1170);
xnor U1525 (N_1525,N_747,N_175);
or U1526 (N_1526,N_572,In_1861);
xor U1527 (N_1527,N_764,N_368);
xnor U1528 (N_1528,N_455,In_2477);
xnor U1529 (N_1529,In_153,N_874);
and U1530 (N_1530,In_1877,In_1078);
xnor U1531 (N_1531,In_646,N_851);
nand U1532 (N_1532,N_40,N_897);
or U1533 (N_1533,N_891,N_813);
xor U1534 (N_1534,N_186,In_78);
nand U1535 (N_1535,In_1853,N_950);
and U1536 (N_1536,In_1043,N_80);
xnor U1537 (N_1537,N_325,N_740);
nand U1538 (N_1538,N_162,N_819);
or U1539 (N_1539,N_352,In_2256);
nand U1540 (N_1540,N_845,N_232);
xor U1541 (N_1541,N_84,N_540);
nand U1542 (N_1542,N_902,N_898);
and U1543 (N_1543,N_357,In_688);
or U1544 (N_1544,N_120,In_1423);
and U1545 (N_1545,In_1016,N_626);
nor U1546 (N_1546,N_560,In_840);
nor U1547 (N_1547,N_711,N_302);
xnor U1548 (N_1548,N_571,N_105);
and U1549 (N_1549,In_2203,In_934);
and U1550 (N_1550,In_132,In_84);
xnor U1551 (N_1551,N_220,N_652);
xor U1552 (N_1552,N_240,N_277);
nor U1553 (N_1553,N_140,N_136);
nor U1554 (N_1554,N_99,In_440);
and U1555 (N_1555,N_7,In_1752);
nand U1556 (N_1556,In_83,N_639);
and U1557 (N_1557,In_505,N_948);
and U1558 (N_1558,N_130,In_178);
or U1559 (N_1559,N_33,N_738);
nor U1560 (N_1560,N_208,In_2214);
or U1561 (N_1561,N_772,N_960);
xor U1562 (N_1562,N_866,N_880);
nand U1563 (N_1563,In_426,N_870);
nand U1564 (N_1564,In_1615,N_535);
nor U1565 (N_1565,N_135,In_2073);
nand U1566 (N_1566,In_909,In_1629);
or U1567 (N_1567,In_1124,N_428);
nor U1568 (N_1568,N_853,N_596);
and U1569 (N_1569,N_20,In_626);
xor U1570 (N_1570,N_159,N_87);
xnor U1571 (N_1571,In_1573,N_890);
and U1572 (N_1572,In_49,N_829);
xnor U1573 (N_1573,N_994,N_465);
xnor U1574 (N_1574,N_522,N_675);
nor U1575 (N_1575,In_619,In_483);
nand U1576 (N_1576,N_736,In_1512);
nor U1577 (N_1577,In_464,N_506);
and U1578 (N_1578,N_775,N_395);
xor U1579 (N_1579,N_863,N_254);
nand U1580 (N_1580,N_784,N_256);
nor U1581 (N_1581,N_739,N_379);
or U1582 (N_1582,N_896,N_827);
or U1583 (N_1583,N_380,In_991);
xnor U1584 (N_1584,N_722,N_941);
xor U1585 (N_1585,In_180,N_579);
nor U1586 (N_1586,N_729,In_1606);
and U1587 (N_1587,N_484,In_550);
xnor U1588 (N_1588,N_45,In_1731);
and U1589 (N_1589,N_478,In_68);
and U1590 (N_1590,N_785,N_733);
nor U1591 (N_1591,N_955,N_716);
or U1592 (N_1592,N_27,N_852);
nor U1593 (N_1593,In_1219,N_0);
nor U1594 (N_1594,In_1284,In_2315);
nor U1595 (N_1595,N_882,N_865);
and U1596 (N_1596,N_641,In_1105);
xor U1597 (N_1597,In_351,N_810);
or U1598 (N_1598,N_165,N_944);
nor U1599 (N_1599,N_562,N_725);
nand U1600 (N_1600,N_171,In_478);
nand U1601 (N_1601,In_679,N_441);
or U1602 (N_1602,N_146,In_2068);
xor U1603 (N_1603,N_306,N_721);
or U1604 (N_1604,In_1311,In_724);
nand U1605 (N_1605,N_66,N_267);
and U1606 (N_1606,N_341,N_519);
nor U1607 (N_1607,In_1378,N_786);
nand U1608 (N_1608,In_998,In_263);
nand U1609 (N_1609,N_505,In_1616);
nand U1610 (N_1610,N_5,N_476);
nand U1611 (N_1611,In_862,N_43);
and U1612 (N_1612,N_660,N_648);
nand U1613 (N_1613,N_44,N_493);
nand U1614 (N_1614,N_369,N_154);
nor U1615 (N_1615,In_1332,In_1984);
nand U1616 (N_1616,In_1531,In_1386);
and U1617 (N_1617,In_1524,N_215);
nor U1618 (N_1618,In_1392,N_745);
or U1619 (N_1619,N_831,N_439);
nor U1620 (N_1620,In_33,N_178);
nand U1621 (N_1621,In_1449,N_934);
or U1622 (N_1622,In_705,N_418);
nand U1623 (N_1623,N_835,N_700);
nand U1624 (N_1624,In_2200,N_565);
nor U1625 (N_1625,In_2248,N_282);
or U1626 (N_1626,N_270,In_933);
nand U1627 (N_1627,N_613,In_2367);
xnor U1628 (N_1628,In_1014,N_61);
nand U1629 (N_1629,N_976,N_940);
or U1630 (N_1630,N_294,In_918);
xor U1631 (N_1631,In_703,N_605);
nor U1632 (N_1632,N_482,N_593);
and U1633 (N_1633,N_881,In_2455);
xnor U1634 (N_1634,N_524,N_490);
nand U1635 (N_1635,In_93,N_102);
and U1636 (N_1636,N_992,In_1216);
or U1637 (N_1637,N_997,In_315);
nor U1638 (N_1638,N_603,N_243);
xnor U1639 (N_1639,In_636,In_1241);
nand U1640 (N_1640,N_289,In_521);
nor U1641 (N_1641,N_354,N_12);
or U1642 (N_1642,In_876,N_607);
or U1643 (N_1643,In_650,N_990);
xor U1644 (N_1644,N_698,N_497);
or U1645 (N_1645,In_1728,N_377);
nand U1646 (N_1646,N_800,N_804);
or U1647 (N_1647,N_367,In_1799);
nor U1648 (N_1648,N_751,N_491);
or U1649 (N_1649,N_756,In_530);
or U1650 (N_1650,N_189,N_972);
xor U1651 (N_1651,In_381,In_1771);
nand U1652 (N_1652,In_1503,N_633);
and U1653 (N_1653,N_927,N_523);
and U1654 (N_1654,N_923,N_241);
or U1655 (N_1655,In_1228,N_417);
xnor U1656 (N_1656,N_363,N_799);
nor U1657 (N_1657,In_1034,N_51);
xnor U1658 (N_1658,In_1566,In_2283);
nand U1659 (N_1659,In_2494,N_70);
xor U1660 (N_1660,N_216,N_339);
and U1661 (N_1661,N_204,N_137);
or U1662 (N_1662,N_710,N_499);
nor U1663 (N_1663,N_378,In_2274);
and U1664 (N_1664,N_177,N_202);
or U1665 (N_1665,N_755,N_608);
and U1666 (N_1666,N_221,N_196);
nand U1667 (N_1667,N_185,In_395);
nand U1668 (N_1668,N_335,In_1308);
nand U1669 (N_1669,N_907,In_199);
xnor U1670 (N_1670,N_789,N_665);
nor U1671 (N_1671,In_1422,N_266);
and U1672 (N_1672,N_406,In_112);
xor U1673 (N_1673,N_753,N_463);
nor U1674 (N_1674,N_545,In_857);
or U1675 (N_1675,N_218,N_544);
or U1676 (N_1676,N_393,In_434);
and U1677 (N_1677,In_939,N_668);
xor U1678 (N_1678,In_928,N_807);
nand U1679 (N_1679,N_709,N_945);
or U1680 (N_1680,In_828,In_2015);
and U1681 (N_1681,In_2308,N_281);
or U1682 (N_1682,N_182,In_771);
and U1683 (N_1683,In_1474,In_627);
and U1684 (N_1684,N_251,N_808);
xor U1685 (N_1685,In_92,In_1155);
xnor U1686 (N_1686,N_653,N_17);
nor U1687 (N_1687,In_1351,In_200);
and U1688 (N_1688,N_63,N_4);
nor U1689 (N_1689,N_319,N_857);
xnor U1690 (N_1690,In_642,In_845);
nor U1691 (N_1691,N_90,In_787);
nor U1692 (N_1692,N_312,N_449);
xor U1693 (N_1693,N_557,N_286);
nor U1694 (N_1694,N_619,N_674);
or U1695 (N_1695,N_128,N_627);
nor U1696 (N_1696,In_23,N_107);
nor U1697 (N_1697,N_982,In_1497);
nand U1698 (N_1698,N_318,N_82);
and U1699 (N_1699,N_157,N_184);
and U1700 (N_1700,N_888,In_1736);
or U1701 (N_1701,N_673,In_238);
and U1702 (N_1702,In_745,N_72);
and U1703 (N_1703,N_616,N_89);
nor U1704 (N_1704,N_402,In_2036);
and U1705 (N_1705,N_871,N_609);
or U1706 (N_1706,In_664,N_210);
nand U1707 (N_1707,In_1760,N_183);
or U1708 (N_1708,N_460,N_39);
or U1709 (N_1709,N_209,N_779);
nor U1710 (N_1710,N_31,N_28);
and U1711 (N_1711,N_780,In_1057);
nor U1712 (N_1712,N_568,N_337);
nand U1713 (N_1713,N_938,N_631);
or U1714 (N_1714,In_1373,In_2104);
nor U1715 (N_1715,N_937,N_462);
and U1716 (N_1716,In_431,N_517);
xnor U1717 (N_1717,N_610,In_2272);
or U1718 (N_1718,N_563,N_118);
and U1719 (N_1719,N_268,In_916);
nand U1720 (N_1720,In_2043,In_883);
xnor U1721 (N_1721,N_864,N_526);
xor U1722 (N_1722,N_414,In_306);
nand U1723 (N_1723,N_769,N_97);
and U1724 (N_1724,In_2234,N_909);
and U1725 (N_1725,In_1296,N_686);
nand U1726 (N_1726,N_508,N_106);
nor U1727 (N_1727,N_642,N_400);
nand U1728 (N_1728,N_915,In_832);
nor U1729 (N_1729,In_525,In_1633);
nand U1730 (N_1730,N_564,N_127);
xnor U1731 (N_1731,In_1899,In_1938);
nand U1732 (N_1732,N_664,N_374);
xor U1733 (N_1733,N_83,In_552);
and U1734 (N_1734,In_1929,In_1020);
xor U1735 (N_1735,N_181,In_1223);
or U1736 (N_1736,N_174,N_362);
xnor U1737 (N_1737,N_391,N_332);
or U1738 (N_1738,In_2483,In_1260);
nand U1739 (N_1739,N_662,N_744);
and U1740 (N_1740,N_649,In_2085);
and U1741 (N_1741,In_1009,In_807);
nand U1742 (N_1742,In_2070,N_160);
and U1743 (N_1743,N_287,N_876);
or U1744 (N_1744,N_570,N_581);
and U1745 (N_1745,N_781,N_79);
or U1746 (N_1746,In_1438,In_243);
nor U1747 (N_1747,In_814,N_504);
nor U1748 (N_1748,N_592,N_906);
nor U1749 (N_1749,N_447,In_314);
nand U1750 (N_1750,In_1054,N_816);
nor U1751 (N_1751,N_872,In_1861);
nor U1752 (N_1752,N_737,N_466);
and U1753 (N_1753,In_1282,N_873);
xnor U1754 (N_1754,N_654,In_552);
or U1755 (N_1755,N_847,N_425);
xor U1756 (N_1756,In_1063,N_272);
xor U1757 (N_1757,In_267,N_993);
xnor U1758 (N_1758,N_132,In_2220);
nor U1759 (N_1759,N_815,N_371);
nor U1760 (N_1760,N_396,N_40);
nand U1761 (N_1761,N_997,In_1595);
and U1762 (N_1762,In_1313,N_939);
xor U1763 (N_1763,N_815,In_263);
and U1764 (N_1764,In_2070,N_400);
and U1765 (N_1765,N_919,N_175);
or U1766 (N_1766,N_479,In_2212);
and U1767 (N_1767,N_904,In_27);
or U1768 (N_1768,In_703,N_986);
and U1769 (N_1769,N_244,N_356);
or U1770 (N_1770,N_346,N_532);
nand U1771 (N_1771,N_523,In_1830);
and U1772 (N_1772,N_415,N_668);
or U1773 (N_1773,N_295,In_1799);
nand U1774 (N_1774,N_451,In_310);
xor U1775 (N_1775,N_464,N_657);
or U1776 (N_1776,In_1859,N_213);
and U1777 (N_1777,In_1009,In_314);
nor U1778 (N_1778,In_1269,N_142);
and U1779 (N_1779,In_2068,In_1172);
or U1780 (N_1780,N_811,In_1984);
nand U1781 (N_1781,In_1934,N_909);
nand U1782 (N_1782,N_757,N_964);
or U1783 (N_1783,N_701,N_765);
nand U1784 (N_1784,In_477,N_298);
and U1785 (N_1785,N_640,N_570);
nand U1786 (N_1786,N_23,N_311);
or U1787 (N_1787,In_1901,N_952);
nand U1788 (N_1788,In_1084,In_2137);
xnor U1789 (N_1789,N_429,N_773);
nand U1790 (N_1790,N_188,In_996);
and U1791 (N_1791,N_882,N_873);
nand U1792 (N_1792,In_688,N_507);
nor U1793 (N_1793,N_933,N_451);
or U1794 (N_1794,In_1627,N_190);
nand U1795 (N_1795,N_306,N_161);
and U1796 (N_1796,N_365,N_370);
xor U1797 (N_1797,In_2220,In_1197);
nand U1798 (N_1798,In_1633,N_106);
xor U1799 (N_1799,In_550,In_1777);
and U1800 (N_1800,N_600,N_607);
or U1801 (N_1801,N_529,N_579);
or U1802 (N_1802,In_201,N_920);
nand U1803 (N_1803,In_1334,In_2139);
and U1804 (N_1804,N_510,In_405);
or U1805 (N_1805,N_142,In_441);
nor U1806 (N_1806,N_897,N_583);
xnor U1807 (N_1807,In_1054,N_751);
nor U1808 (N_1808,N_857,In_1658);
and U1809 (N_1809,N_517,In_178);
nand U1810 (N_1810,N_398,In_1804);
nor U1811 (N_1811,In_1179,In_727);
xor U1812 (N_1812,N_195,N_56);
nor U1813 (N_1813,N_59,In_688);
and U1814 (N_1814,N_27,N_988);
and U1815 (N_1815,N_984,N_105);
nor U1816 (N_1816,N_946,In_1418);
xnor U1817 (N_1817,N_304,N_328);
nor U1818 (N_1818,In_984,In_727);
xor U1819 (N_1819,N_812,N_595);
nor U1820 (N_1820,N_412,N_466);
nor U1821 (N_1821,N_238,N_744);
and U1822 (N_1822,In_1007,In_699);
nand U1823 (N_1823,N_331,N_621);
and U1824 (N_1824,N_438,N_414);
xor U1825 (N_1825,N_40,N_659);
nor U1826 (N_1826,N_448,N_290);
or U1827 (N_1827,N_267,In_97);
nor U1828 (N_1828,N_456,N_404);
nor U1829 (N_1829,N_846,N_46);
and U1830 (N_1830,N_151,N_71);
or U1831 (N_1831,N_2,In_1622);
and U1832 (N_1832,N_473,N_710);
nand U1833 (N_1833,In_921,N_204);
nand U1834 (N_1834,In_53,N_6);
xor U1835 (N_1835,In_1578,N_352);
xnor U1836 (N_1836,In_645,N_500);
or U1837 (N_1837,N_62,In_1008);
nand U1838 (N_1838,In_316,In_1540);
nor U1839 (N_1839,N_820,N_79);
xnor U1840 (N_1840,N_836,N_878);
nand U1841 (N_1841,N_899,N_878);
or U1842 (N_1842,In_2120,N_139);
nand U1843 (N_1843,N_408,In_288);
xor U1844 (N_1844,In_1296,N_777);
or U1845 (N_1845,N_539,In_1246);
nand U1846 (N_1846,N_790,N_734);
xnor U1847 (N_1847,N_450,N_651);
nand U1848 (N_1848,In_1932,In_1387);
and U1849 (N_1849,N_358,N_837);
xnor U1850 (N_1850,N_847,N_496);
nand U1851 (N_1851,In_267,In_1311);
nand U1852 (N_1852,N_408,N_726);
nor U1853 (N_1853,N_224,N_241);
nand U1854 (N_1854,In_1657,In_2293);
xnor U1855 (N_1855,N_873,In_1780);
xnor U1856 (N_1856,N_851,N_473);
or U1857 (N_1857,N_946,N_707);
and U1858 (N_1858,N_231,N_498);
xnor U1859 (N_1859,In_1957,N_9);
nor U1860 (N_1860,N_362,In_1106);
xor U1861 (N_1861,N_835,N_681);
nand U1862 (N_1862,In_1859,N_899);
xor U1863 (N_1863,N_997,In_1078);
or U1864 (N_1864,N_834,N_213);
nand U1865 (N_1865,In_1309,N_401);
xor U1866 (N_1866,N_730,N_721);
nand U1867 (N_1867,In_1799,N_741);
nor U1868 (N_1868,In_1293,N_661);
and U1869 (N_1869,N_874,In_573);
xor U1870 (N_1870,N_126,N_215);
and U1871 (N_1871,N_428,N_778);
nor U1872 (N_1872,In_126,N_151);
or U1873 (N_1873,In_732,N_432);
xnor U1874 (N_1874,N_405,In_946);
xnor U1875 (N_1875,In_1104,N_491);
xnor U1876 (N_1876,N_614,N_343);
xor U1877 (N_1877,N_650,N_234);
or U1878 (N_1878,In_92,N_327);
xor U1879 (N_1879,N_575,In_1615);
nand U1880 (N_1880,In_199,N_279);
nand U1881 (N_1881,In_441,N_333);
nor U1882 (N_1882,In_314,N_535);
and U1883 (N_1883,N_68,N_657);
or U1884 (N_1884,N_16,N_455);
or U1885 (N_1885,In_1,N_78);
nand U1886 (N_1886,N_851,N_396);
nand U1887 (N_1887,N_212,In_1409);
and U1888 (N_1888,In_1877,N_207);
or U1889 (N_1889,N_710,In_1720);
nand U1890 (N_1890,N_46,N_4);
and U1891 (N_1891,N_620,N_316);
nand U1892 (N_1892,N_579,N_718);
or U1893 (N_1893,N_944,N_947);
xor U1894 (N_1894,N_860,N_698);
or U1895 (N_1895,In_2013,N_229);
nand U1896 (N_1896,N_757,In_2308);
nand U1897 (N_1897,N_821,In_2374);
or U1898 (N_1898,N_76,In_1770);
xnor U1899 (N_1899,In_457,In_2368);
and U1900 (N_1900,N_825,In_1984);
nand U1901 (N_1901,In_507,N_173);
xnor U1902 (N_1902,N_70,N_229);
xor U1903 (N_1903,N_679,N_873);
and U1904 (N_1904,N_110,In_1578);
and U1905 (N_1905,In_1305,In_2383);
or U1906 (N_1906,N_199,N_813);
xor U1907 (N_1907,In_1531,N_329);
xor U1908 (N_1908,N_912,N_34);
and U1909 (N_1909,In_996,N_981);
nand U1910 (N_1910,N_841,N_696);
and U1911 (N_1911,N_416,In_2274);
nand U1912 (N_1912,N_85,In_636);
nor U1913 (N_1913,N_857,In_2306);
nand U1914 (N_1914,N_672,In_257);
nor U1915 (N_1915,In_2428,N_673);
nand U1916 (N_1916,In_974,In_246);
xor U1917 (N_1917,In_1062,In_164);
xnor U1918 (N_1918,In_1613,N_338);
and U1919 (N_1919,N_740,In_1062);
xnor U1920 (N_1920,In_84,N_699);
or U1921 (N_1921,N_149,N_432);
nand U1922 (N_1922,In_2086,In_2178);
xnor U1923 (N_1923,N_738,In_2368);
nand U1924 (N_1924,In_1378,N_419);
xor U1925 (N_1925,N_93,N_49);
nand U1926 (N_1926,N_952,N_653);
xor U1927 (N_1927,In_357,N_443);
xor U1928 (N_1928,N_387,N_89);
nor U1929 (N_1929,N_609,In_710);
or U1930 (N_1930,In_200,N_757);
or U1931 (N_1931,N_590,In_1057);
nor U1932 (N_1932,In_939,N_271);
or U1933 (N_1933,In_441,N_279);
nor U1934 (N_1934,N_941,N_308);
xnor U1935 (N_1935,N_162,N_658);
and U1936 (N_1936,N_968,In_697);
or U1937 (N_1937,N_581,N_612);
or U1938 (N_1938,N_514,N_594);
and U1939 (N_1939,N_165,N_226);
xor U1940 (N_1940,N_989,N_713);
and U1941 (N_1941,N_500,N_830);
xor U1942 (N_1942,N_234,N_275);
nor U1943 (N_1943,N_511,N_251);
nand U1944 (N_1944,N_854,N_790);
or U1945 (N_1945,N_327,N_330);
xnor U1946 (N_1946,N_599,N_972);
or U1947 (N_1947,N_392,N_961);
xnor U1948 (N_1948,N_788,In_414);
and U1949 (N_1949,In_1735,N_533);
nor U1950 (N_1950,N_295,N_486);
nand U1951 (N_1951,N_449,N_544);
xnor U1952 (N_1952,N_550,N_345);
nand U1953 (N_1953,In_1566,N_199);
nor U1954 (N_1954,N_109,In_1085);
nand U1955 (N_1955,In_478,In_1639);
nand U1956 (N_1956,N_416,N_431);
nand U1957 (N_1957,N_141,N_67);
and U1958 (N_1958,N_551,N_445);
xnor U1959 (N_1959,N_292,N_65);
xnor U1960 (N_1960,N_756,N_250);
or U1961 (N_1961,N_362,N_360);
nand U1962 (N_1962,N_587,N_873);
xnor U1963 (N_1963,In_1392,N_582);
and U1964 (N_1964,N_310,N_994);
nor U1965 (N_1965,In_1945,N_584);
or U1966 (N_1966,In_1074,N_962);
xor U1967 (N_1967,N_508,N_425);
and U1968 (N_1968,N_748,N_962);
nor U1969 (N_1969,In_397,In_1842);
or U1970 (N_1970,In_1085,N_594);
nand U1971 (N_1971,N_801,In_395);
nor U1972 (N_1972,N_738,In_1891);
xnor U1973 (N_1973,N_275,In_1562);
and U1974 (N_1974,In_1194,N_694);
nand U1975 (N_1975,N_702,N_896);
nand U1976 (N_1976,N_220,N_699);
nand U1977 (N_1977,In_2383,In_1512);
and U1978 (N_1978,N_68,N_163);
and U1979 (N_1979,N_164,In_2327);
xnor U1980 (N_1980,N_853,In_162);
and U1981 (N_1981,N_949,N_339);
and U1982 (N_1982,N_417,In_507);
nand U1983 (N_1983,N_830,In_81);
nor U1984 (N_1984,N_918,N_649);
or U1985 (N_1985,In_2234,In_992);
or U1986 (N_1986,N_191,N_837);
xnor U1987 (N_1987,In_1516,N_93);
and U1988 (N_1988,In_2013,N_754);
and U1989 (N_1989,In_1351,In_883);
or U1990 (N_1990,N_964,N_208);
nand U1991 (N_1991,In_790,N_679);
xor U1992 (N_1992,N_420,In_1161);
nand U1993 (N_1993,In_1595,N_242);
or U1994 (N_1994,N_806,N_918);
and U1995 (N_1995,N_82,N_358);
or U1996 (N_1996,N_710,In_1801);
or U1997 (N_1997,In_379,N_341);
nand U1998 (N_1998,N_456,In_1494);
nand U1999 (N_1999,In_1973,N_298);
and U2000 (N_2000,N_1706,N_1703);
and U2001 (N_2001,N_1521,N_1998);
and U2002 (N_2002,N_1982,N_1532);
or U2003 (N_2003,N_1987,N_1062);
nor U2004 (N_2004,N_1383,N_1822);
nor U2005 (N_2005,N_1684,N_1835);
xor U2006 (N_2006,N_1573,N_1032);
or U2007 (N_2007,N_1675,N_1237);
xor U2008 (N_2008,N_1325,N_1587);
nand U2009 (N_2009,N_1764,N_1869);
nor U2010 (N_2010,N_1460,N_1780);
xor U2011 (N_2011,N_1480,N_1507);
xor U2012 (N_2012,N_1911,N_1468);
nand U2013 (N_2013,N_1541,N_1864);
nor U2014 (N_2014,N_1090,N_1920);
and U2015 (N_2015,N_1022,N_1348);
xor U2016 (N_2016,N_1264,N_1786);
xnor U2017 (N_2017,N_1417,N_1568);
or U2018 (N_2018,N_1669,N_1029);
or U2019 (N_2019,N_1825,N_1650);
or U2020 (N_2020,N_1380,N_1902);
or U2021 (N_2021,N_1394,N_1601);
nor U2022 (N_2022,N_1451,N_1308);
and U2023 (N_2023,N_1853,N_1761);
nand U2024 (N_2024,N_1148,N_1574);
xor U2025 (N_2025,N_1852,N_1104);
and U2026 (N_2026,N_1859,N_1083);
or U2027 (N_2027,N_1595,N_1628);
nand U2028 (N_2028,N_1929,N_1923);
or U2029 (N_2029,N_1198,N_1978);
or U2030 (N_2030,N_1774,N_1158);
nor U2031 (N_2031,N_1539,N_1155);
nor U2032 (N_2032,N_1166,N_1046);
nor U2033 (N_2033,N_1826,N_1252);
and U2034 (N_2034,N_1326,N_1959);
nor U2035 (N_2035,N_1291,N_1003);
or U2036 (N_2036,N_1951,N_1938);
nand U2037 (N_2037,N_1755,N_1243);
nor U2038 (N_2038,N_1097,N_1447);
nand U2039 (N_2039,N_1932,N_1333);
xnor U2040 (N_2040,N_1000,N_1748);
xnor U2041 (N_2041,N_1047,N_1346);
xnor U2042 (N_2042,N_1194,N_1176);
nand U2043 (N_2043,N_1278,N_1948);
xnor U2044 (N_2044,N_1096,N_1505);
nand U2045 (N_2045,N_1736,N_1411);
or U2046 (N_2046,N_1379,N_1906);
nor U2047 (N_2047,N_1810,N_1921);
nor U2048 (N_2048,N_1156,N_1110);
or U2049 (N_2049,N_1449,N_1455);
xor U2050 (N_2050,N_1214,N_1304);
nor U2051 (N_2051,N_1154,N_1162);
and U2052 (N_2052,N_1433,N_1694);
or U2053 (N_2053,N_1847,N_1591);
nand U2054 (N_2054,N_1809,N_1497);
and U2055 (N_2055,N_1882,N_1458);
xor U2056 (N_2056,N_1772,N_1121);
xor U2057 (N_2057,N_1749,N_1477);
xor U2058 (N_2058,N_1345,N_1973);
nor U2059 (N_2059,N_1049,N_1353);
xnor U2060 (N_2060,N_1210,N_1089);
or U2061 (N_2061,N_1909,N_1999);
nor U2062 (N_2062,N_1995,N_1860);
xor U2063 (N_2063,N_1400,N_1406);
or U2064 (N_2064,N_1217,N_1500);
and U2065 (N_2065,N_1160,N_1710);
xor U2066 (N_2066,N_1656,N_1147);
or U2067 (N_2067,N_1294,N_1692);
nand U2068 (N_2068,N_1887,N_1054);
xnor U2069 (N_2069,N_1506,N_1716);
and U2070 (N_2070,N_1880,N_1623);
nor U2071 (N_2071,N_1401,N_1438);
nor U2072 (N_2072,N_1408,N_1550);
nor U2073 (N_2073,N_1721,N_1750);
or U2074 (N_2074,N_1907,N_1363);
or U2075 (N_2075,N_1361,N_1958);
and U2076 (N_2076,N_1385,N_1720);
and U2077 (N_2077,N_1905,N_1708);
xnor U2078 (N_2078,N_1330,N_1114);
and U2079 (N_2079,N_1366,N_1510);
or U2080 (N_2080,N_1578,N_1640);
nand U2081 (N_2081,N_1785,N_1233);
or U2082 (N_2082,N_1084,N_1286);
and U2083 (N_2083,N_1391,N_1903);
xnor U2084 (N_2084,N_1130,N_1473);
nand U2085 (N_2085,N_1280,N_1877);
xor U2086 (N_2086,N_1292,N_1102);
xor U2087 (N_2087,N_1612,N_1966);
nor U2088 (N_2088,N_1465,N_1374);
nand U2089 (N_2089,N_1878,N_1949);
and U2090 (N_2090,N_1056,N_1830);
or U2091 (N_2091,N_1901,N_1562);
xor U2092 (N_2092,N_1001,N_1413);
xor U2093 (N_2093,N_1791,N_1662);
and U2094 (N_2094,N_1360,N_1037);
nand U2095 (N_2095,N_1174,N_1834);
and U2096 (N_2096,N_1050,N_1884);
or U2097 (N_2097,N_1087,N_1251);
or U2098 (N_2098,N_1793,N_1602);
and U2099 (N_2099,N_1017,N_1422);
nor U2100 (N_2100,N_1953,N_1627);
nand U2101 (N_2101,N_1129,N_1118);
nor U2102 (N_2102,N_1020,N_1435);
or U2103 (N_2103,N_1013,N_1688);
or U2104 (N_2104,N_1946,N_1040);
xnor U2105 (N_2105,N_1546,N_1059);
nor U2106 (N_2106,N_1896,N_1072);
nor U2107 (N_2107,N_1192,N_1801);
nor U2108 (N_2108,N_1425,N_1461);
xnor U2109 (N_2109,N_1495,N_1913);
or U2110 (N_2110,N_1520,N_1754);
xor U2111 (N_2111,N_1857,N_1557);
xor U2112 (N_2112,N_1289,N_1693);
nor U2113 (N_2113,N_1808,N_1952);
xnor U2114 (N_2114,N_1329,N_1305);
xnor U2115 (N_2115,N_1874,N_1523);
nand U2116 (N_2116,N_1077,N_1225);
and U2117 (N_2117,N_1041,N_1430);
or U2118 (N_2118,N_1841,N_1301);
and U2119 (N_2119,N_1027,N_1547);
or U2120 (N_2120,N_1424,N_1961);
and U2121 (N_2121,N_1078,N_1220);
nor U2122 (N_2122,N_1842,N_1616);
or U2123 (N_2123,N_1789,N_1898);
and U2124 (N_2124,N_1554,N_1454);
or U2125 (N_2125,N_1594,N_1356);
and U2126 (N_2126,N_1799,N_1827);
nor U2127 (N_2127,N_1262,N_1651);
nor U2128 (N_2128,N_1629,N_1180);
nand U2129 (N_2129,N_1881,N_1957);
or U2130 (N_2130,N_1545,N_1051);
nand U2131 (N_2131,N_1516,N_1767);
nand U2132 (N_2132,N_1831,N_1939);
nor U2133 (N_2133,N_1357,N_1188);
nand U2134 (N_2134,N_1642,N_1377);
and U2135 (N_2135,N_1914,N_1531);
xnor U2136 (N_2136,N_1610,N_1711);
nand U2137 (N_2137,N_1781,N_1010);
xnor U2138 (N_2138,N_1218,N_1025);
or U2139 (N_2139,N_1904,N_1343);
or U2140 (N_2140,N_1804,N_1770);
xor U2141 (N_2141,N_1567,N_1570);
and U2142 (N_2142,N_1542,N_1211);
xnor U2143 (N_2143,N_1034,N_1502);
xnor U2144 (N_2144,N_1015,N_1974);
nor U2145 (N_2145,N_1828,N_1762);
nor U2146 (N_2146,N_1073,N_1604);
or U2147 (N_2147,N_1419,N_1576);
xnor U2148 (N_2148,N_1886,N_1437);
nand U2149 (N_2149,N_1249,N_1971);
nand U2150 (N_2150,N_1475,N_1596);
or U2151 (N_2151,N_1668,N_1418);
or U2152 (N_2152,N_1002,N_1742);
nand U2153 (N_2153,N_1729,N_1765);
nor U2154 (N_2154,N_1759,N_1312);
or U2155 (N_2155,N_1151,N_1099);
nand U2156 (N_2156,N_1396,N_1227);
xnor U2157 (N_2157,N_1508,N_1075);
and U2158 (N_2158,N_1402,N_1016);
or U2159 (N_2159,N_1168,N_1712);
and U2160 (N_2160,N_1849,N_1565);
and U2161 (N_2161,N_1979,N_1434);
xnor U2162 (N_2162,N_1970,N_1645);
and U2163 (N_2163,N_1744,N_1984);
xor U2164 (N_2164,N_1322,N_1861);
and U2165 (N_2165,N_1031,N_1942);
xor U2166 (N_2166,N_1779,N_1496);
nor U2167 (N_2167,N_1341,N_1815);
nand U2168 (N_2168,N_1023,N_1518);
or U2169 (N_2169,N_1368,N_1392);
nor U2170 (N_2170,N_1572,N_1782);
xnor U2171 (N_2171,N_1637,N_1199);
nand U2172 (N_2172,N_1163,N_1846);
nand U2173 (N_2173,N_1275,N_1229);
and U2174 (N_2174,N_1281,N_1661);
nor U2175 (N_2175,N_1235,N_1763);
or U2176 (N_2176,N_1985,N_1664);
xor U2177 (N_2177,N_1014,N_1239);
nor U2178 (N_2178,N_1036,N_1479);
nand U2179 (N_2179,N_1445,N_1224);
nand U2180 (N_2180,N_1582,N_1279);
xnor U2181 (N_2181,N_1723,N_1108);
and U2182 (N_2182,N_1064,N_1871);
nor U2183 (N_2183,N_1190,N_1035);
or U2184 (N_2184,N_1687,N_1757);
xnor U2185 (N_2185,N_1685,N_1365);
and U2186 (N_2186,N_1686,N_1498);
or U2187 (N_2187,N_1823,N_1443);
or U2188 (N_2188,N_1098,N_1030);
nor U2189 (N_2189,N_1676,N_1634);
xnor U2190 (N_2190,N_1100,N_1695);
and U2191 (N_2191,N_1665,N_1577);
or U2192 (N_2192,N_1283,N_1559);
nand U2193 (N_2193,N_1248,N_1583);
or U2194 (N_2194,N_1875,N_1756);
nand U2195 (N_2195,N_1528,N_1691);
xor U2196 (N_2196,N_1739,N_1592);
xor U2197 (N_2197,N_1812,N_1055);
nand U2198 (N_2198,N_1331,N_1488);
nor U2199 (N_2199,N_1579,N_1021);
or U2200 (N_2200,N_1071,N_1316);
or U2201 (N_2201,N_1486,N_1843);
xor U2202 (N_2202,N_1420,N_1328);
xnor U2203 (N_2203,N_1947,N_1483);
nand U2204 (N_2204,N_1513,N_1463);
or U2205 (N_2205,N_1126,N_1910);
nand U2206 (N_2206,N_1673,N_1773);
nor U2207 (N_2207,N_1306,N_1127);
and U2208 (N_2208,N_1590,N_1297);
or U2209 (N_2209,N_1800,N_1336);
xnor U2210 (N_2210,N_1992,N_1766);
or U2211 (N_2211,N_1260,N_1821);
nand U2212 (N_2212,N_1060,N_1204);
xor U2213 (N_2213,N_1698,N_1494);
nand U2214 (N_2214,N_1735,N_1120);
nor U2215 (N_2215,N_1146,N_1648);
nand U2216 (N_2216,N_1922,N_1165);
nand U2217 (N_2217,N_1816,N_1323);
nand U2218 (N_2218,N_1339,N_1805);
and U2219 (N_2219,N_1028,N_1890);
nand U2220 (N_2220,N_1792,N_1274);
nand U2221 (N_2221,N_1092,N_1196);
nand U2222 (N_2222,N_1824,N_1209);
nor U2223 (N_2223,N_1441,N_1106);
or U2224 (N_2224,N_1512,N_1813);
nand U2225 (N_2225,N_1265,N_1139);
nor U2226 (N_2226,N_1674,N_1080);
or U2227 (N_2227,N_1314,N_1501);
nor U2228 (N_2228,N_1088,N_1484);
nand U2229 (N_2229,N_1608,N_1515);
xnor U2230 (N_2230,N_1646,N_1918);
and U2231 (N_2231,N_1536,N_1912);
xnor U2232 (N_2232,N_1241,N_1647);
nand U2233 (N_2233,N_1159,N_1276);
and U2234 (N_2234,N_1128,N_1599);
nor U2235 (N_2235,N_1777,N_1614);
nor U2236 (N_2236,N_1429,N_1795);
nor U2237 (N_2237,N_1436,N_1266);
nor U2238 (N_2238,N_1369,N_1644);
nor U2239 (N_2239,N_1927,N_1273);
nor U2240 (N_2240,N_1802,N_1862);
or U2241 (N_2241,N_1743,N_1149);
nand U2242 (N_2242,N_1045,N_1839);
nand U2243 (N_2243,N_1285,N_1868);
and U2244 (N_2244,N_1103,N_1421);
nand U2245 (N_2245,N_1186,N_1972);
nor U2246 (N_2246,N_1169,N_1619);
xnor U2247 (N_2247,N_1143,N_1788);
and U2248 (N_2248,N_1888,N_1983);
or U2249 (N_2249,N_1925,N_1267);
or U2250 (N_2250,N_1033,N_1960);
nand U2251 (N_2251,N_1538,N_1311);
nand U2252 (N_2252,N_1867,N_1179);
nor U2253 (N_2253,N_1244,N_1734);
and U2254 (N_2254,N_1471,N_1704);
and U2255 (N_2255,N_1551,N_1928);
xnor U2256 (N_2256,N_1145,N_1746);
xor U2257 (N_2257,N_1485,N_1845);
nor U2258 (N_2258,N_1751,N_1172);
nor U2259 (N_2259,N_1019,N_1112);
nand U2260 (N_2260,N_1269,N_1334);
and U2261 (N_2261,N_1702,N_1446);
nor U2262 (N_2262,N_1005,N_1141);
nor U2263 (N_2263,N_1250,N_1175);
nand U2264 (N_2264,N_1137,N_1295);
or U2265 (N_2265,N_1919,N_1585);
or U2266 (N_2266,N_1620,N_1533);
nor U2267 (N_2267,N_1259,N_1431);
and U2268 (N_2268,N_1635,N_1490);
and U2269 (N_2269,N_1261,N_1643);
and U2270 (N_2270,N_1870,N_1397);
nor U2271 (N_2271,N_1018,N_1197);
nand U2272 (N_2272,N_1563,N_1462);
and U2273 (N_2273,N_1895,N_1737);
nor U2274 (N_2274,N_1234,N_1061);
or U2275 (N_2275,N_1069,N_1797);
nand U2276 (N_2276,N_1600,N_1456);
and U2277 (N_2277,N_1277,N_1296);
nor U2278 (N_2278,N_1844,N_1833);
xnor U2279 (N_2279,N_1606,N_1509);
xnor U2280 (N_2280,N_1879,N_1641);
and U2281 (N_2281,N_1611,N_1941);
xnor U2282 (N_2282,N_1967,N_1355);
or U2283 (N_2283,N_1367,N_1517);
and U2284 (N_2284,N_1935,N_1553);
xor U2285 (N_2285,N_1581,N_1375);
and U2286 (N_2286,N_1226,N_1588);
nor U2287 (N_2287,N_1228,N_1707);
or U2288 (N_2288,N_1571,N_1299);
nand U2289 (N_2289,N_1549,N_1965);
xor U2290 (N_2290,N_1784,N_1364);
nor U2291 (N_2291,N_1633,N_1666);
xor U2292 (N_2292,N_1556,N_1519);
nor U2293 (N_2293,N_1962,N_1371);
nor U2294 (N_2294,N_1290,N_1012);
nor U2295 (N_2295,N_1850,N_1254);
nor U2296 (N_2296,N_1378,N_1714);
and U2297 (N_2297,N_1745,N_1448);
xor U2298 (N_2298,N_1621,N_1205);
nand U2299 (N_2299,N_1405,N_1416);
nand U2300 (N_2300,N_1564,N_1063);
nor U2301 (N_2301,N_1232,N_1851);
and U2302 (N_2302,N_1924,N_1133);
and U2303 (N_2303,N_1111,N_1955);
nor U2304 (N_2304,N_1373,N_1086);
xor U2305 (N_2305,N_1344,N_1082);
and U2306 (N_2306,N_1426,N_1107);
xor U2307 (N_2307,N_1185,N_1393);
xor U2308 (N_2308,N_1885,N_1769);
nor U2309 (N_2309,N_1395,N_1410);
xor U2310 (N_2310,N_1883,N_1511);
nand U2311 (N_2311,N_1231,N_1522);
xnor U2312 (N_2312,N_1771,N_1135);
or U2313 (N_2313,N_1598,N_1288);
and U2314 (N_2314,N_1652,N_1407);
nand U2315 (N_2315,N_1964,N_1618);
or U2316 (N_2316,N_1136,N_1153);
nand U2317 (N_2317,N_1124,N_1819);
nor U2318 (N_2318,N_1164,N_1575);
or U2319 (N_2319,N_1740,N_1926);
and U2320 (N_2320,N_1854,N_1349);
nor U2321 (N_2321,N_1183,N_1963);
xnor U2322 (N_2322,N_1132,N_1215);
and U2323 (N_2323,N_1258,N_1543);
nor U2324 (N_2324,N_1131,N_1432);
and U2325 (N_2325,N_1206,N_1991);
xor U2326 (N_2326,N_1491,N_1358);
or U2327 (N_2327,N_1863,N_1866);
xnor U2328 (N_2328,N_1981,N_1384);
xnor U2329 (N_2329,N_1741,N_1727);
nor U2330 (N_2330,N_1760,N_1790);
nand U2331 (N_2331,N_1362,N_1113);
and U2332 (N_2332,N_1659,N_1310);
and U2333 (N_2333,N_1453,N_1409);
or U2334 (N_2334,N_1658,N_1622);
nor U2335 (N_2335,N_1725,N_1263);
xor U2336 (N_2336,N_1677,N_1238);
and U2337 (N_2337,N_1412,N_1271);
nand U2338 (N_2338,N_1937,N_1332);
or U2339 (N_2339,N_1615,N_1829);
nor U2340 (N_2340,N_1667,N_1242);
or U2341 (N_2341,N_1101,N_1931);
nand U2342 (N_2342,N_1457,N_1440);
and U2343 (N_2343,N_1255,N_1048);
nor U2344 (N_2344,N_1404,N_1530);
nor U2345 (N_2345,N_1855,N_1184);
or U2346 (N_2346,N_1655,N_1387);
xor U2347 (N_2347,N_1681,N_1605);
nand U2348 (N_2348,N_1302,N_1134);
and U2349 (N_2349,N_1024,N_1631);
xor U2350 (N_2350,N_1117,N_1894);
nor U2351 (N_2351,N_1680,N_1338);
nand U2352 (N_2352,N_1607,N_1452);
xor U2353 (N_2353,N_1679,N_1728);
nand U2354 (N_2354,N_1470,N_1219);
nand U2355 (N_2355,N_1376,N_1649);
or U2356 (N_2356,N_1945,N_1977);
and U2357 (N_2357,N_1713,N_1527);
and U2358 (N_2358,N_1058,N_1068);
nor U2359 (N_2359,N_1207,N_1672);
or U2360 (N_2360,N_1584,N_1682);
and U2361 (N_2361,N_1638,N_1427);
and U2362 (N_2362,N_1144,N_1492);
xor U2363 (N_2363,N_1700,N_1915);
xnor U2364 (N_2364,N_1318,N_1444);
nor U2365 (N_2365,N_1351,N_1811);
or U2366 (N_2366,N_1347,N_1317);
nor U2367 (N_2367,N_1690,N_1337);
xor U2368 (N_2368,N_1370,N_1042);
nand U2369 (N_2369,N_1776,N_1459);
or U2370 (N_2370,N_1954,N_1988);
or U2371 (N_2371,N_1287,N_1996);
nor U2372 (N_2372,N_1423,N_1093);
nand U2373 (N_2373,N_1152,N_1203);
or U2374 (N_2374,N_1319,N_1548);
or U2375 (N_2375,N_1832,N_1566);
xor U2376 (N_2376,N_1593,N_1738);
nand U2377 (N_2377,N_1715,N_1555);
and U2378 (N_2378,N_1388,N_1315);
nand U2379 (N_2379,N_1382,N_1892);
nor U2380 (N_2380,N_1936,N_1624);
and U2381 (N_2381,N_1472,N_1719);
xnor U2382 (N_2382,N_1008,N_1980);
nor U2383 (N_2383,N_1876,N_1889);
or U2384 (N_2384,N_1817,N_1683);
nor U2385 (N_2385,N_1300,N_1007);
or U2386 (N_2386,N_1803,N_1775);
and U2387 (N_2387,N_1167,N_1178);
or U2388 (N_2388,N_1514,N_1481);
nand U2389 (N_2389,N_1115,N_1415);
xor U2390 (N_2390,N_1758,N_1768);
nor U2391 (N_2391,N_1350,N_1940);
or U2392 (N_2392,N_1524,N_1718);
or U2393 (N_2393,N_1678,N_1181);
nor U2394 (N_2394,N_1428,N_1730);
nand U2395 (N_2395,N_1717,N_1726);
or U2396 (N_2396,N_1105,N_1968);
nand U2397 (N_2397,N_1335,N_1990);
and U2398 (N_2398,N_1943,N_1222);
xor U2399 (N_2399,N_1157,N_1930);
xnor U2400 (N_2400,N_1893,N_1150);
and U2401 (N_2401,N_1245,N_1246);
nor U2402 (N_2402,N_1840,N_1293);
or U2403 (N_2403,N_1856,N_1173);
or U2404 (N_2404,N_1389,N_1609);
and U2405 (N_2405,N_1381,N_1223);
or U2406 (N_2406,N_1873,N_1848);
xor U2407 (N_2407,N_1778,N_1796);
nor U2408 (N_2408,N_1950,N_1006);
or U2409 (N_2409,N_1212,N_1140);
nor U2410 (N_2410,N_1561,N_1065);
or U2411 (N_2411,N_1309,N_1247);
nor U2412 (N_2412,N_1464,N_1125);
and U2413 (N_2413,N_1067,N_1256);
xnor U2414 (N_2414,N_1352,N_1625);
nand U2415 (N_2415,N_1586,N_1724);
and U2416 (N_2416,N_1891,N_1091);
and U2417 (N_2417,N_1701,N_1221);
nor U2418 (N_2418,N_1070,N_1200);
or U2419 (N_2419,N_1403,N_1558);
nor U2420 (N_2420,N_1138,N_1414);
nand U2421 (N_2421,N_1944,N_1177);
nor U2422 (N_2422,N_1123,N_1899);
or U2423 (N_2423,N_1537,N_1170);
nor U2424 (N_2424,N_1663,N_1504);
nand U2425 (N_2425,N_1066,N_1202);
and U2426 (N_2426,N_1753,N_1193);
or U2427 (N_2427,N_1696,N_1529);
nor U2428 (N_2428,N_1076,N_1321);
or U2429 (N_2429,N_1597,N_1390);
nand U2430 (N_2430,N_1109,N_1195);
nand U2431 (N_2431,N_1818,N_1630);
or U2432 (N_2432,N_1858,N_1201);
nand U2433 (N_2433,N_1705,N_1613);
nor U2434 (N_2434,N_1011,N_1085);
nor U2435 (N_2435,N_1026,N_1916);
nor U2436 (N_2436,N_1359,N_1732);
or U2437 (N_2437,N_1569,N_1142);
nor U2438 (N_2438,N_1997,N_1989);
or U2439 (N_2439,N_1044,N_1654);
and U2440 (N_2440,N_1208,N_1467);
or U2441 (N_2441,N_1240,N_1969);
nand U2442 (N_2442,N_1257,N_1639);
nor U2443 (N_2443,N_1731,N_1603);
nor U2444 (N_2444,N_1324,N_1489);
and U2445 (N_2445,N_1079,N_1493);
nor U2446 (N_2446,N_1439,N_1787);
or U2447 (N_2447,N_1094,N_1552);
nand U2448 (N_2448,N_1993,N_1399);
or U2449 (N_2449,N_1191,N_1442);
and U2450 (N_2450,N_1908,N_1540);
and U2451 (N_2451,N_1386,N_1053);
nand U2452 (N_2452,N_1722,N_1794);
and U2453 (N_2453,N_1956,N_1009);
and U2454 (N_2454,N_1689,N_1189);
nor U2455 (N_2455,N_1660,N_1526);
nand U2456 (N_2456,N_1872,N_1670);
nor U2457 (N_2457,N_1372,N_1733);
xor U2458 (N_2458,N_1268,N_1216);
and U2459 (N_2459,N_1476,N_1095);
or U2460 (N_2460,N_1122,N_1340);
nand U2461 (N_2461,N_1986,N_1282);
nand U2462 (N_2462,N_1626,N_1272);
or U2463 (N_2463,N_1298,N_1580);
nor U2464 (N_2464,N_1820,N_1976);
and U2465 (N_2465,N_1284,N_1709);
and U2466 (N_2466,N_1213,N_1354);
or U2467 (N_2467,N_1398,N_1466);
xnor U2468 (N_2468,N_1236,N_1653);
and U2469 (N_2469,N_1900,N_1535);
and U2470 (N_2470,N_1934,N_1342);
and U2471 (N_2471,N_1450,N_1161);
nand U2472 (N_2472,N_1182,N_1836);
xor U2473 (N_2473,N_1897,N_1838);
xor U2474 (N_2474,N_1171,N_1270);
or U2475 (N_2475,N_1783,N_1469);
xor U2476 (N_2476,N_1052,N_1752);
nand U2477 (N_2477,N_1657,N_1837);
and U2478 (N_2478,N_1617,N_1589);
or U2479 (N_2479,N_1994,N_1043);
or U2480 (N_2480,N_1038,N_1307);
or U2481 (N_2481,N_1917,N_1327);
xnor U2482 (N_2482,N_1865,N_1975);
xnor U2483 (N_2483,N_1004,N_1499);
nand U2484 (N_2484,N_1807,N_1482);
nor U2485 (N_2485,N_1081,N_1697);
nor U2486 (N_2486,N_1487,N_1814);
xnor U2487 (N_2487,N_1253,N_1039);
nand U2488 (N_2488,N_1187,N_1747);
nand U2489 (N_2489,N_1636,N_1474);
nand U2490 (N_2490,N_1671,N_1632);
nor U2491 (N_2491,N_1230,N_1057);
xnor U2492 (N_2492,N_1933,N_1699);
nand U2493 (N_2493,N_1503,N_1798);
nand U2494 (N_2494,N_1116,N_1478);
or U2495 (N_2495,N_1806,N_1320);
xor U2496 (N_2496,N_1534,N_1119);
nor U2497 (N_2497,N_1303,N_1313);
nand U2498 (N_2498,N_1560,N_1544);
or U2499 (N_2499,N_1525,N_1074);
nand U2500 (N_2500,N_1477,N_1498);
nand U2501 (N_2501,N_1706,N_1730);
xor U2502 (N_2502,N_1920,N_1411);
and U2503 (N_2503,N_1436,N_1137);
or U2504 (N_2504,N_1771,N_1005);
and U2505 (N_2505,N_1743,N_1292);
and U2506 (N_2506,N_1740,N_1564);
and U2507 (N_2507,N_1451,N_1354);
nand U2508 (N_2508,N_1184,N_1254);
nand U2509 (N_2509,N_1164,N_1897);
xor U2510 (N_2510,N_1401,N_1360);
or U2511 (N_2511,N_1779,N_1301);
nor U2512 (N_2512,N_1219,N_1538);
or U2513 (N_2513,N_1607,N_1343);
or U2514 (N_2514,N_1906,N_1140);
and U2515 (N_2515,N_1702,N_1561);
nor U2516 (N_2516,N_1788,N_1357);
and U2517 (N_2517,N_1323,N_1447);
and U2518 (N_2518,N_1512,N_1541);
and U2519 (N_2519,N_1462,N_1457);
or U2520 (N_2520,N_1345,N_1643);
or U2521 (N_2521,N_1731,N_1703);
and U2522 (N_2522,N_1081,N_1486);
or U2523 (N_2523,N_1307,N_1428);
xnor U2524 (N_2524,N_1143,N_1710);
or U2525 (N_2525,N_1732,N_1004);
nor U2526 (N_2526,N_1683,N_1572);
or U2527 (N_2527,N_1281,N_1696);
xnor U2528 (N_2528,N_1942,N_1633);
and U2529 (N_2529,N_1373,N_1008);
xnor U2530 (N_2530,N_1738,N_1249);
xor U2531 (N_2531,N_1827,N_1213);
nor U2532 (N_2532,N_1037,N_1344);
or U2533 (N_2533,N_1534,N_1442);
and U2534 (N_2534,N_1872,N_1055);
nor U2535 (N_2535,N_1769,N_1508);
and U2536 (N_2536,N_1436,N_1931);
nor U2537 (N_2537,N_1720,N_1109);
nand U2538 (N_2538,N_1185,N_1335);
xnor U2539 (N_2539,N_1756,N_1535);
nand U2540 (N_2540,N_1710,N_1351);
and U2541 (N_2541,N_1208,N_1877);
or U2542 (N_2542,N_1128,N_1731);
and U2543 (N_2543,N_1722,N_1741);
xnor U2544 (N_2544,N_1716,N_1167);
and U2545 (N_2545,N_1642,N_1128);
and U2546 (N_2546,N_1618,N_1490);
nand U2547 (N_2547,N_1630,N_1324);
or U2548 (N_2548,N_1059,N_1414);
nor U2549 (N_2549,N_1733,N_1875);
nor U2550 (N_2550,N_1821,N_1091);
nor U2551 (N_2551,N_1256,N_1516);
nand U2552 (N_2552,N_1017,N_1494);
nor U2553 (N_2553,N_1238,N_1640);
and U2554 (N_2554,N_1566,N_1756);
and U2555 (N_2555,N_1414,N_1539);
xnor U2556 (N_2556,N_1473,N_1294);
nand U2557 (N_2557,N_1704,N_1885);
nor U2558 (N_2558,N_1592,N_1218);
nor U2559 (N_2559,N_1613,N_1611);
xor U2560 (N_2560,N_1223,N_1586);
nand U2561 (N_2561,N_1119,N_1234);
nand U2562 (N_2562,N_1379,N_1272);
or U2563 (N_2563,N_1898,N_1134);
and U2564 (N_2564,N_1813,N_1598);
and U2565 (N_2565,N_1426,N_1813);
nor U2566 (N_2566,N_1796,N_1912);
and U2567 (N_2567,N_1935,N_1581);
and U2568 (N_2568,N_1567,N_1623);
nand U2569 (N_2569,N_1598,N_1478);
xnor U2570 (N_2570,N_1867,N_1453);
nand U2571 (N_2571,N_1574,N_1076);
and U2572 (N_2572,N_1023,N_1596);
nand U2573 (N_2573,N_1043,N_1774);
nand U2574 (N_2574,N_1547,N_1546);
nor U2575 (N_2575,N_1995,N_1954);
nor U2576 (N_2576,N_1825,N_1363);
nor U2577 (N_2577,N_1691,N_1121);
nand U2578 (N_2578,N_1119,N_1447);
or U2579 (N_2579,N_1891,N_1418);
nor U2580 (N_2580,N_1406,N_1451);
nor U2581 (N_2581,N_1218,N_1427);
xor U2582 (N_2582,N_1874,N_1142);
and U2583 (N_2583,N_1552,N_1955);
and U2584 (N_2584,N_1126,N_1460);
nand U2585 (N_2585,N_1215,N_1650);
xnor U2586 (N_2586,N_1725,N_1904);
or U2587 (N_2587,N_1664,N_1607);
nor U2588 (N_2588,N_1065,N_1791);
or U2589 (N_2589,N_1850,N_1580);
and U2590 (N_2590,N_1493,N_1022);
nand U2591 (N_2591,N_1475,N_1632);
and U2592 (N_2592,N_1100,N_1362);
or U2593 (N_2593,N_1518,N_1512);
and U2594 (N_2594,N_1959,N_1025);
nor U2595 (N_2595,N_1128,N_1654);
nor U2596 (N_2596,N_1080,N_1501);
xor U2597 (N_2597,N_1290,N_1930);
xor U2598 (N_2598,N_1150,N_1475);
nand U2599 (N_2599,N_1975,N_1049);
xor U2600 (N_2600,N_1063,N_1264);
and U2601 (N_2601,N_1685,N_1283);
and U2602 (N_2602,N_1798,N_1858);
nor U2603 (N_2603,N_1961,N_1193);
or U2604 (N_2604,N_1373,N_1258);
or U2605 (N_2605,N_1813,N_1886);
and U2606 (N_2606,N_1376,N_1084);
and U2607 (N_2607,N_1360,N_1868);
xnor U2608 (N_2608,N_1157,N_1648);
nand U2609 (N_2609,N_1676,N_1836);
xor U2610 (N_2610,N_1036,N_1804);
nor U2611 (N_2611,N_1141,N_1339);
nand U2612 (N_2612,N_1258,N_1304);
nor U2613 (N_2613,N_1032,N_1012);
nor U2614 (N_2614,N_1271,N_1867);
nand U2615 (N_2615,N_1508,N_1242);
xor U2616 (N_2616,N_1493,N_1410);
nor U2617 (N_2617,N_1697,N_1108);
nand U2618 (N_2618,N_1867,N_1059);
nor U2619 (N_2619,N_1566,N_1408);
xnor U2620 (N_2620,N_1349,N_1657);
or U2621 (N_2621,N_1559,N_1435);
nand U2622 (N_2622,N_1906,N_1224);
nand U2623 (N_2623,N_1487,N_1191);
nand U2624 (N_2624,N_1590,N_1350);
or U2625 (N_2625,N_1700,N_1105);
xor U2626 (N_2626,N_1354,N_1832);
nor U2627 (N_2627,N_1671,N_1014);
and U2628 (N_2628,N_1336,N_1170);
xnor U2629 (N_2629,N_1543,N_1870);
xnor U2630 (N_2630,N_1506,N_1642);
nand U2631 (N_2631,N_1836,N_1192);
and U2632 (N_2632,N_1430,N_1447);
or U2633 (N_2633,N_1072,N_1367);
nor U2634 (N_2634,N_1959,N_1994);
nand U2635 (N_2635,N_1712,N_1317);
and U2636 (N_2636,N_1178,N_1454);
nand U2637 (N_2637,N_1574,N_1138);
nor U2638 (N_2638,N_1526,N_1728);
and U2639 (N_2639,N_1261,N_1210);
nor U2640 (N_2640,N_1467,N_1548);
xnor U2641 (N_2641,N_1354,N_1024);
nor U2642 (N_2642,N_1967,N_1328);
or U2643 (N_2643,N_1385,N_1445);
nor U2644 (N_2644,N_1069,N_1461);
xnor U2645 (N_2645,N_1354,N_1991);
xor U2646 (N_2646,N_1433,N_1624);
or U2647 (N_2647,N_1917,N_1507);
nor U2648 (N_2648,N_1833,N_1510);
xnor U2649 (N_2649,N_1713,N_1049);
or U2650 (N_2650,N_1268,N_1191);
or U2651 (N_2651,N_1980,N_1312);
and U2652 (N_2652,N_1732,N_1509);
nand U2653 (N_2653,N_1292,N_1883);
nand U2654 (N_2654,N_1976,N_1470);
xnor U2655 (N_2655,N_1441,N_1088);
and U2656 (N_2656,N_1676,N_1242);
and U2657 (N_2657,N_1586,N_1255);
nor U2658 (N_2658,N_1223,N_1525);
nand U2659 (N_2659,N_1774,N_1379);
or U2660 (N_2660,N_1932,N_1181);
nand U2661 (N_2661,N_1794,N_1088);
or U2662 (N_2662,N_1061,N_1686);
and U2663 (N_2663,N_1424,N_1890);
nor U2664 (N_2664,N_1279,N_1586);
xnor U2665 (N_2665,N_1248,N_1280);
or U2666 (N_2666,N_1291,N_1681);
nor U2667 (N_2667,N_1947,N_1022);
nand U2668 (N_2668,N_1410,N_1476);
xor U2669 (N_2669,N_1628,N_1960);
nand U2670 (N_2670,N_1636,N_1275);
nand U2671 (N_2671,N_1291,N_1869);
or U2672 (N_2672,N_1815,N_1617);
or U2673 (N_2673,N_1102,N_1809);
and U2674 (N_2674,N_1670,N_1218);
nand U2675 (N_2675,N_1395,N_1200);
or U2676 (N_2676,N_1624,N_1086);
or U2677 (N_2677,N_1149,N_1841);
and U2678 (N_2678,N_1236,N_1173);
xnor U2679 (N_2679,N_1881,N_1132);
and U2680 (N_2680,N_1361,N_1730);
nor U2681 (N_2681,N_1389,N_1460);
and U2682 (N_2682,N_1917,N_1368);
nand U2683 (N_2683,N_1326,N_1725);
nor U2684 (N_2684,N_1698,N_1292);
xnor U2685 (N_2685,N_1931,N_1416);
xor U2686 (N_2686,N_1132,N_1302);
and U2687 (N_2687,N_1546,N_1371);
or U2688 (N_2688,N_1760,N_1120);
xnor U2689 (N_2689,N_1951,N_1658);
nor U2690 (N_2690,N_1892,N_1284);
and U2691 (N_2691,N_1121,N_1210);
and U2692 (N_2692,N_1266,N_1680);
xor U2693 (N_2693,N_1078,N_1285);
nand U2694 (N_2694,N_1494,N_1325);
xnor U2695 (N_2695,N_1127,N_1208);
or U2696 (N_2696,N_1318,N_1876);
nor U2697 (N_2697,N_1431,N_1477);
and U2698 (N_2698,N_1135,N_1232);
nand U2699 (N_2699,N_1828,N_1364);
nand U2700 (N_2700,N_1245,N_1019);
or U2701 (N_2701,N_1299,N_1007);
nand U2702 (N_2702,N_1476,N_1856);
xor U2703 (N_2703,N_1580,N_1926);
and U2704 (N_2704,N_1090,N_1672);
nor U2705 (N_2705,N_1769,N_1491);
and U2706 (N_2706,N_1098,N_1597);
xor U2707 (N_2707,N_1588,N_1541);
or U2708 (N_2708,N_1906,N_1025);
nor U2709 (N_2709,N_1843,N_1833);
nor U2710 (N_2710,N_1150,N_1108);
nand U2711 (N_2711,N_1920,N_1783);
xnor U2712 (N_2712,N_1955,N_1912);
nand U2713 (N_2713,N_1386,N_1071);
nor U2714 (N_2714,N_1591,N_1012);
and U2715 (N_2715,N_1499,N_1515);
xnor U2716 (N_2716,N_1754,N_1214);
or U2717 (N_2717,N_1633,N_1901);
nand U2718 (N_2718,N_1451,N_1900);
xor U2719 (N_2719,N_1969,N_1899);
and U2720 (N_2720,N_1097,N_1502);
or U2721 (N_2721,N_1069,N_1779);
and U2722 (N_2722,N_1579,N_1495);
nand U2723 (N_2723,N_1950,N_1843);
or U2724 (N_2724,N_1384,N_1128);
and U2725 (N_2725,N_1290,N_1817);
nand U2726 (N_2726,N_1761,N_1062);
or U2727 (N_2727,N_1452,N_1422);
nor U2728 (N_2728,N_1900,N_1274);
nand U2729 (N_2729,N_1193,N_1217);
or U2730 (N_2730,N_1333,N_1464);
or U2731 (N_2731,N_1671,N_1158);
nand U2732 (N_2732,N_1985,N_1814);
nor U2733 (N_2733,N_1212,N_1850);
xnor U2734 (N_2734,N_1382,N_1017);
or U2735 (N_2735,N_1382,N_1798);
nor U2736 (N_2736,N_1513,N_1536);
and U2737 (N_2737,N_1253,N_1995);
xnor U2738 (N_2738,N_1510,N_1499);
xnor U2739 (N_2739,N_1075,N_1037);
nor U2740 (N_2740,N_1426,N_1858);
nor U2741 (N_2741,N_1346,N_1572);
nor U2742 (N_2742,N_1787,N_1386);
nor U2743 (N_2743,N_1388,N_1702);
and U2744 (N_2744,N_1471,N_1256);
and U2745 (N_2745,N_1810,N_1719);
nor U2746 (N_2746,N_1302,N_1140);
or U2747 (N_2747,N_1809,N_1932);
nor U2748 (N_2748,N_1929,N_1637);
nand U2749 (N_2749,N_1419,N_1313);
and U2750 (N_2750,N_1096,N_1155);
and U2751 (N_2751,N_1314,N_1662);
xnor U2752 (N_2752,N_1296,N_1518);
and U2753 (N_2753,N_1708,N_1260);
or U2754 (N_2754,N_1867,N_1124);
nor U2755 (N_2755,N_1747,N_1746);
xnor U2756 (N_2756,N_1782,N_1470);
and U2757 (N_2757,N_1859,N_1515);
nand U2758 (N_2758,N_1690,N_1480);
or U2759 (N_2759,N_1289,N_1690);
and U2760 (N_2760,N_1247,N_1397);
xnor U2761 (N_2761,N_1594,N_1593);
xnor U2762 (N_2762,N_1684,N_1238);
or U2763 (N_2763,N_1175,N_1926);
and U2764 (N_2764,N_1639,N_1632);
or U2765 (N_2765,N_1085,N_1766);
and U2766 (N_2766,N_1589,N_1107);
nor U2767 (N_2767,N_1301,N_1275);
xnor U2768 (N_2768,N_1281,N_1769);
or U2769 (N_2769,N_1303,N_1500);
or U2770 (N_2770,N_1187,N_1155);
xor U2771 (N_2771,N_1396,N_1063);
or U2772 (N_2772,N_1921,N_1964);
nand U2773 (N_2773,N_1146,N_1974);
nor U2774 (N_2774,N_1873,N_1832);
nor U2775 (N_2775,N_1811,N_1292);
nand U2776 (N_2776,N_1339,N_1342);
xor U2777 (N_2777,N_1782,N_1739);
nor U2778 (N_2778,N_1878,N_1722);
nor U2779 (N_2779,N_1489,N_1772);
and U2780 (N_2780,N_1846,N_1635);
nand U2781 (N_2781,N_1621,N_1603);
or U2782 (N_2782,N_1418,N_1789);
or U2783 (N_2783,N_1410,N_1996);
or U2784 (N_2784,N_1085,N_1442);
xor U2785 (N_2785,N_1191,N_1185);
or U2786 (N_2786,N_1699,N_1985);
xor U2787 (N_2787,N_1162,N_1770);
and U2788 (N_2788,N_1443,N_1861);
nand U2789 (N_2789,N_1585,N_1704);
or U2790 (N_2790,N_1550,N_1079);
nor U2791 (N_2791,N_1506,N_1295);
and U2792 (N_2792,N_1482,N_1655);
nor U2793 (N_2793,N_1235,N_1919);
or U2794 (N_2794,N_1085,N_1999);
nor U2795 (N_2795,N_1921,N_1358);
and U2796 (N_2796,N_1082,N_1054);
nand U2797 (N_2797,N_1689,N_1289);
nand U2798 (N_2798,N_1614,N_1294);
and U2799 (N_2799,N_1290,N_1166);
or U2800 (N_2800,N_1445,N_1223);
and U2801 (N_2801,N_1079,N_1899);
or U2802 (N_2802,N_1001,N_1941);
nor U2803 (N_2803,N_1398,N_1512);
nand U2804 (N_2804,N_1262,N_1171);
or U2805 (N_2805,N_1151,N_1800);
xnor U2806 (N_2806,N_1943,N_1972);
nor U2807 (N_2807,N_1280,N_1686);
and U2808 (N_2808,N_1103,N_1621);
nand U2809 (N_2809,N_1000,N_1407);
and U2810 (N_2810,N_1532,N_1087);
and U2811 (N_2811,N_1364,N_1217);
xnor U2812 (N_2812,N_1085,N_1327);
and U2813 (N_2813,N_1013,N_1051);
nor U2814 (N_2814,N_1392,N_1128);
xor U2815 (N_2815,N_1219,N_1375);
nor U2816 (N_2816,N_1725,N_1477);
xor U2817 (N_2817,N_1550,N_1303);
or U2818 (N_2818,N_1045,N_1489);
xnor U2819 (N_2819,N_1517,N_1040);
nor U2820 (N_2820,N_1920,N_1476);
and U2821 (N_2821,N_1007,N_1297);
nor U2822 (N_2822,N_1586,N_1628);
xor U2823 (N_2823,N_1573,N_1694);
and U2824 (N_2824,N_1054,N_1359);
and U2825 (N_2825,N_1035,N_1940);
and U2826 (N_2826,N_1796,N_1192);
xor U2827 (N_2827,N_1598,N_1059);
nand U2828 (N_2828,N_1039,N_1650);
or U2829 (N_2829,N_1524,N_1376);
xnor U2830 (N_2830,N_1028,N_1241);
xor U2831 (N_2831,N_1279,N_1680);
xor U2832 (N_2832,N_1371,N_1847);
or U2833 (N_2833,N_1884,N_1396);
nor U2834 (N_2834,N_1693,N_1260);
xor U2835 (N_2835,N_1535,N_1331);
nand U2836 (N_2836,N_1780,N_1956);
or U2837 (N_2837,N_1396,N_1782);
nand U2838 (N_2838,N_1675,N_1351);
or U2839 (N_2839,N_1093,N_1955);
or U2840 (N_2840,N_1574,N_1154);
and U2841 (N_2841,N_1485,N_1061);
xnor U2842 (N_2842,N_1174,N_1217);
nor U2843 (N_2843,N_1604,N_1029);
nand U2844 (N_2844,N_1676,N_1209);
and U2845 (N_2845,N_1041,N_1998);
and U2846 (N_2846,N_1139,N_1854);
xnor U2847 (N_2847,N_1560,N_1772);
nor U2848 (N_2848,N_1182,N_1657);
and U2849 (N_2849,N_1102,N_1516);
nand U2850 (N_2850,N_1120,N_1654);
and U2851 (N_2851,N_1555,N_1243);
and U2852 (N_2852,N_1985,N_1796);
nand U2853 (N_2853,N_1082,N_1138);
or U2854 (N_2854,N_1271,N_1786);
or U2855 (N_2855,N_1477,N_1246);
xor U2856 (N_2856,N_1641,N_1071);
xnor U2857 (N_2857,N_1212,N_1641);
nand U2858 (N_2858,N_1075,N_1540);
and U2859 (N_2859,N_1823,N_1857);
nor U2860 (N_2860,N_1136,N_1219);
and U2861 (N_2861,N_1365,N_1174);
nand U2862 (N_2862,N_1963,N_1983);
nor U2863 (N_2863,N_1660,N_1302);
and U2864 (N_2864,N_1353,N_1994);
nand U2865 (N_2865,N_1156,N_1625);
xnor U2866 (N_2866,N_1914,N_1623);
xor U2867 (N_2867,N_1716,N_1717);
and U2868 (N_2868,N_1588,N_1889);
xor U2869 (N_2869,N_1995,N_1184);
nor U2870 (N_2870,N_1599,N_1865);
nor U2871 (N_2871,N_1526,N_1822);
or U2872 (N_2872,N_1824,N_1496);
xor U2873 (N_2873,N_1948,N_1363);
or U2874 (N_2874,N_1330,N_1948);
xnor U2875 (N_2875,N_1637,N_1875);
and U2876 (N_2876,N_1428,N_1360);
or U2877 (N_2877,N_1981,N_1193);
and U2878 (N_2878,N_1850,N_1479);
xor U2879 (N_2879,N_1673,N_1790);
nand U2880 (N_2880,N_1795,N_1820);
xnor U2881 (N_2881,N_1389,N_1789);
nand U2882 (N_2882,N_1238,N_1069);
nand U2883 (N_2883,N_1215,N_1525);
xnor U2884 (N_2884,N_1023,N_1643);
nand U2885 (N_2885,N_1849,N_1746);
and U2886 (N_2886,N_1840,N_1365);
or U2887 (N_2887,N_1889,N_1978);
and U2888 (N_2888,N_1969,N_1606);
nor U2889 (N_2889,N_1481,N_1105);
or U2890 (N_2890,N_1282,N_1688);
nor U2891 (N_2891,N_1515,N_1336);
xor U2892 (N_2892,N_1940,N_1382);
nor U2893 (N_2893,N_1295,N_1926);
xnor U2894 (N_2894,N_1968,N_1257);
nor U2895 (N_2895,N_1285,N_1544);
nand U2896 (N_2896,N_1875,N_1494);
or U2897 (N_2897,N_1022,N_1651);
xor U2898 (N_2898,N_1246,N_1937);
xor U2899 (N_2899,N_1068,N_1672);
nor U2900 (N_2900,N_1737,N_1543);
nor U2901 (N_2901,N_1037,N_1280);
xnor U2902 (N_2902,N_1283,N_1947);
and U2903 (N_2903,N_1314,N_1221);
nand U2904 (N_2904,N_1472,N_1586);
nor U2905 (N_2905,N_1414,N_1194);
xnor U2906 (N_2906,N_1607,N_1187);
or U2907 (N_2907,N_1964,N_1055);
nor U2908 (N_2908,N_1477,N_1572);
xnor U2909 (N_2909,N_1799,N_1914);
or U2910 (N_2910,N_1545,N_1658);
and U2911 (N_2911,N_1977,N_1893);
and U2912 (N_2912,N_1521,N_1594);
nor U2913 (N_2913,N_1471,N_1842);
nor U2914 (N_2914,N_1920,N_1937);
nor U2915 (N_2915,N_1882,N_1792);
and U2916 (N_2916,N_1891,N_1893);
nor U2917 (N_2917,N_1896,N_1164);
or U2918 (N_2918,N_1926,N_1486);
and U2919 (N_2919,N_1610,N_1571);
or U2920 (N_2920,N_1946,N_1030);
nor U2921 (N_2921,N_1479,N_1328);
nand U2922 (N_2922,N_1082,N_1359);
and U2923 (N_2923,N_1434,N_1282);
and U2924 (N_2924,N_1284,N_1620);
xor U2925 (N_2925,N_1840,N_1670);
nor U2926 (N_2926,N_1093,N_1615);
nor U2927 (N_2927,N_1843,N_1697);
and U2928 (N_2928,N_1718,N_1248);
or U2929 (N_2929,N_1137,N_1441);
nand U2930 (N_2930,N_1171,N_1863);
and U2931 (N_2931,N_1879,N_1406);
nand U2932 (N_2932,N_1442,N_1682);
xnor U2933 (N_2933,N_1612,N_1469);
nor U2934 (N_2934,N_1764,N_1860);
xor U2935 (N_2935,N_1208,N_1634);
nor U2936 (N_2936,N_1585,N_1198);
and U2937 (N_2937,N_1426,N_1909);
and U2938 (N_2938,N_1167,N_1542);
nand U2939 (N_2939,N_1692,N_1540);
and U2940 (N_2940,N_1719,N_1274);
nand U2941 (N_2941,N_1171,N_1842);
or U2942 (N_2942,N_1003,N_1692);
xnor U2943 (N_2943,N_1470,N_1401);
or U2944 (N_2944,N_1337,N_1119);
nor U2945 (N_2945,N_1600,N_1166);
or U2946 (N_2946,N_1371,N_1031);
and U2947 (N_2947,N_1231,N_1161);
and U2948 (N_2948,N_1235,N_1003);
nand U2949 (N_2949,N_1269,N_1663);
xnor U2950 (N_2950,N_1193,N_1191);
xnor U2951 (N_2951,N_1578,N_1220);
nor U2952 (N_2952,N_1878,N_1743);
nor U2953 (N_2953,N_1112,N_1319);
nor U2954 (N_2954,N_1172,N_1256);
xor U2955 (N_2955,N_1718,N_1258);
nor U2956 (N_2956,N_1180,N_1166);
or U2957 (N_2957,N_1502,N_1057);
xor U2958 (N_2958,N_1171,N_1454);
and U2959 (N_2959,N_1209,N_1628);
nor U2960 (N_2960,N_1148,N_1664);
or U2961 (N_2961,N_1002,N_1706);
nand U2962 (N_2962,N_1130,N_1873);
nor U2963 (N_2963,N_1681,N_1944);
xor U2964 (N_2964,N_1896,N_1312);
xnor U2965 (N_2965,N_1464,N_1302);
or U2966 (N_2966,N_1500,N_1459);
and U2967 (N_2967,N_1304,N_1540);
and U2968 (N_2968,N_1261,N_1152);
nor U2969 (N_2969,N_1046,N_1485);
nand U2970 (N_2970,N_1367,N_1834);
and U2971 (N_2971,N_1186,N_1942);
nor U2972 (N_2972,N_1787,N_1055);
nor U2973 (N_2973,N_1205,N_1515);
and U2974 (N_2974,N_1785,N_1088);
nand U2975 (N_2975,N_1813,N_1319);
nor U2976 (N_2976,N_1399,N_1241);
or U2977 (N_2977,N_1688,N_1618);
xnor U2978 (N_2978,N_1802,N_1406);
xnor U2979 (N_2979,N_1763,N_1250);
nand U2980 (N_2980,N_1223,N_1501);
xnor U2981 (N_2981,N_1631,N_1513);
nor U2982 (N_2982,N_1324,N_1782);
xnor U2983 (N_2983,N_1397,N_1643);
nand U2984 (N_2984,N_1136,N_1516);
nand U2985 (N_2985,N_1561,N_1423);
nand U2986 (N_2986,N_1415,N_1295);
nand U2987 (N_2987,N_1427,N_1978);
and U2988 (N_2988,N_1142,N_1881);
xnor U2989 (N_2989,N_1361,N_1081);
or U2990 (N_2990,N_1065,N_1379);
xnor U2991 (N_2991,N_1652,N_1102);
xor U2992 (N_2992,N_1217,N_1568);
nor U2993 (N_2993,N_1562,N_1648);
xor U2994 (N_2994,N_1931,N_1913);
nor U2995 (N_2995,N_1652,N_1963);
xnor U2996 (N_2996,N_1010,N_1480);
nor U2997 (N_2997,N_1332,N_1023);
nor U2998 (N_2998,N_1330,N_1261);
xnor U2999 (N_2999,N_1511,N_1913);
and U3000 (N_3000,N_2697,N_2444);
or U3001 (N_3001,N_2391,N_2270);
nor U3002 (N_3002,N_2803,N_2913);
xnor U3003 (N_3003,N_2548,N_2583);
nor U3004 (N_3004,N_2810,N_2647);
or U3005 (N_3005,N_2685,N_2287);
and U3006 (N_3006,N_2946,N_2582);
xnor U3007 (N_3007,N_2961,N_2394);
nand U3008 (N_3008,N_2484,N_2944);
nand U3009 (N_3009,N_2112,N_2260);
nor U3010 (N_3010,N_2301,N_2235);
or U3011 (N_3011,N_2906,N_2641);
xor U3012 (N_3012,N_2355,N_2700);
and U3013 (N_3013,N_2242,N_2238);
and U3014 (N_3014,N_2711,N_2390);
nor U3015 (N_3015,N_2233,N_2471);
nor U3016 (N_3016,N_2150,N_2783);
xor U3017 (N_3017,N_2476,N_2300);
or U3018 (N_3018,N_2674,N_2488);
xor U3019 (N_3019,N_2194,N_2175);
xor U3020 (N_3020,N_2369,N_2097);
nor U3021 (N_3021,N_2283,N_2473);
and U3022 (N_3022,N_2225,N_2578);
or U3023 (N_3023,N_2011,N_2148);
and U3024 (N_3024,N_2110,N_2989);
or U3025 (N_3025,N_2635,N_2593);
nor U3026 (N_3026,N_2228,N_2629);
or U3027 (N_3027,N_2642,N_2190);
nor U3028 (N_3028,N_2559,N_2265);
nor U3029 (N_3029,N_2928,N_2604);
or U3030 (N_3030,N_2033,N_2269);
or U3031 (N_3031,N_2510,N_2663);
xnor U3032 (N_3032,N_2757,N_2790);
nor U3033 (N_3033,N_2761,N_2813);
nand U3034 (N_3034,N_2078,N_2506);
and U3035 (N_3035,N_2345,N_2249);
xnor U3036 (N_3036,N_2643,N_2977);
or U3037 (N_3037,N_2948,N_2198);
nand U3038 (N_3038,N_2061,N_2037);
and U3039 (N_3039,N_2512,N_2828);
nor U3040 (N_3040,N_2121,N_2808);
or U3041 (N_3041,N_2395,N_2323);
nor U3042 (N_3042,N_2104,N_2497);
xnor U3043 (N_3043,N_2503,N_2768);
nand U3044 (N_3044,N_2479,N_2539);
nor U3045 (N_3045,N_2555,N_2010);
and U3046 (N_3046,N_2428,N_2698);
nand U3047 (N_3047,N_2405,N_2897);
xnor U3048 (N_3048,N_2611,N_2001);
and U3049 (N_3049,N_2968,N_2086);
nor U3050 (N_3050,N_2205,N_2665);
nor U3051 (N_3051,N_2147,N_2831);
and U3052 (N_3052,N_2807,N_2220);
and U3053 (N_3053,N_2914,N_2204);
nand U3054 (N_3054,N_2754,N_2219);
xor U3055 (N_3055,N_2045,N_2915);
nor U3056 (N_3056,N_2883,N_2053);
nand U3057 (N_3057,N_2119,N_2972);
nor U3058 (N_3058,N_2015,N_2986);
and U3059 (N_3059,N_2494,N_2367);
xnor U3060 (N_3060,N_2307,N_2419);
and U3061 (N_3061,N_2836,N_2975);
xor U3062 (N_3062,N_2450,N_2858);
or U3063 (N_3063,N_2823,N_2157);
or U3064 (N_3064,N_2180,N_2921);
or U3065 (N_3065,N_2107,N_2358);
nand U3066 (N_3066,N_2266,N_2406);
or U3067 (N_3067,N_2255,N_2026);
nor U3068 (N_3068,N_2118,N_2480);
xor U3069 (N_3069,N_2692,N_2139);
nand U3070 (N_3070,N_2776,N_2438);
or U3071 (N_3071,N_2923,N_2126);
or U3072 (N_3072,N_2145,N_2085);
xnor U3073 (N_3073,N_2751,N_2889);
xor U3074 (N_3074,N_2268,N_2544);
and U3075 (N_3075,N_2842,N_2922);
and U3076 (N_3076,N_2368,N_2445);
nor U3077 (N_3077,N_2974,N_2523);
nand U3078 (N_3078,N_2123,N_2141);
and U3079 (N_3079,N_2749,N_2014);
nand U3080 (N_3080,N_2144,N_2540);
xor U3081 (N_3081,N_2688,N_2967);
xnor U3082 (N_3082,N_2645,N_2735);
nand U3083 (N_3083,N_2028,N_2091);
nor U3084 (N_3084,N_2414,N_2491);
nand U3085 (N_3085,N_2694,N_2873);
or U3086 (N_3086,N_2602,N_2365);
nand U3087 (N_3087,N_2134,N_2256);
and U3088 (N_3088,N_2092,N_2032);
xnor U3089 (N_3089,N_2214,N_2983);
nand U3090 (N_3090,N_2704,N_2039);
nor U3091 (N_3091,N_2328,N_2952);
or U3092 (N_3092,N_2447,N_2937);
nand U3093 (N_3093,N_2357,N_2174);
xor U3094 (N_3094,N_2284,N_2764);
xnor U3095 (N_3095,N_2377,N_2599);
nor U3096 (N_3096,N_2076,N_2400);
nand U3097 (N_3097,N_2586,N_2898);
xnor U3098 (N_3098,N_2770,N_2223);
and U3099 (N_3099,N_2077,N_2890);
xnor U3100 (N_3100,N_2335,N_2507);
xnor U3101 (N_3101,N_2155,N_2030);
xnor U3102 (N_3102,N_2362,N_2140);
nor U3103 (N_3103,N_2988,N_2666);
or U3104 (N_3104,N_2880,N_2664);
xnor U3105 (N_3105,N_2295,N_2064);
nor U3106 (N_3106,N_2797,N_2251);
or U3107 (N_3107,N_2384,N_2908);
nor U3108 (N_3108,N_2756,N_2442);
and U3109 (N_3109,N_2226,N_2837);
or U3110 (N_3110,N_2662,N_2392);
xor U3111 (N_3111,N_2505,N_2049);
and U3112 (N_3112,N_2459,N_2533);
and U3113 (N_3113,N_2575,N_2185);
nand U3114 (N_3114,N_2441,N_2859);
or U3115 (N_3115,N_2521,N_2597);
or U3116 (N_3116,N_2250,N_2321);
or U3117 (N_3117,N_2477,N_2197);
or U3118 (N_3118,N_2302,N_2954);
and U3119 (N_3119,N_2690,N_2035);
nor U3120 (N_3120,N_2970,N_2201);
nor U3121 (N_3121,N_2332,N_2278);
nand U3122 (N_3122,N_2087,N_2649);
nand U3123 (N_3123,N_2614,N_2127);
or U3124 (N_3124,N_2565,N_2741);
and U3125 (N_3125,N_2101,N_2845);
and U3126 (N_3126,N_2452,N_2370);
xor U3127 (N_3127,N_2239,N_2257);
xnor U3128 (N_3128,N_2387,N_2654);
and U3129 (N_3129,N_2360,N_2043);
xor U3130 (N_3130,N_2976,N_2341);
and U3131 (N_3131,N_2158,N_2153);
nor U3132 (N_3132,N_2486,N_2755);
nor U3133 (N_3133,N_2122,N_2364);
xnor U3134 (N_3134,N_2388,N_2788);
or U3135 (N_3135,N_2769,N_2574);
or U3136 (N_3136,N_2031,N_2534);
nor U3137 (N_3137,N_2580,N_2258);
nand U3138 (N_3138,N_2397,N_2463);
nor U3139 (N_3139,N_2267,N_2612);
or U3140 (N_3140,N_2562,N_2451);
nor U3141 (N_3141,N_2531,N_2561);
nor U3142 (N_3142,N_2294,N_2940);
nand U3143 (N_3143,N_2729,N_2276);
and U3144 (N_3144,N_2855,N_2798);
nor U3145 (N_3145,N_2708,N_2900);
nor U3146 (N_3146,N_2965,N_2615);
nor U3147 (N_3147,N_2209,N_2192);
or U3148 (N_3148,N_2835,N_2263);
nand U3149 (N_3149,N_2947,N_2609);
xor U3150 (N_3150,N_2423,N_2273);
and U3151 (N_3151,N_2746,N_2038);
nand U3152 (N_3152,N_2703,N_2762);
xor U3153 (N_3153,N_2417,N_2535);
or U3154 (N_3154,N_2082,N_2563);
nand U3155 (N_3155,N_2717,N_2796);
nor U3156 (N_3156,N_2920,N_2721);
nand U3157 (N_3157,N_2100,N_2689);
nor U3158 (N_3158,N_2289,N_2829);
nor U3159 (N_3159,N_2051,N_2820);
nand U3160 (N_3160,N_2546,N_2046);
nor U3161 (N_3161,N_2044,N_2894);
or U3162 (N_3162,N_2792,N_2824);
or U3163 (N_3163,N_2063,N_2142);
nor U3164 (N_3164,N_2125,N_2775);
and U3165 (N_3165,N_2380,N_2543);
xor U3166 (N_3166,N_2389,N_2128);
nand U3167 (N_3167,N_2728,N_2777);
nand U3168 (N_3168,N_2800,N_2115);
and U3169 (N_3169,N_2917,N_2517);
xnor U3170 (N_3170,N_2680,N_2293);
and U3171 (N_3171,N_2945,N_2591);
or U3172 (N_3172,N_2589,N_2522);
nor U3173 (N_3173,N_2427,N_2084);
and U3174 (N_3174,N_2464,N_2924);
xnor U3175 (N_3175,N_2090,N_2374);
or U3176 (N_3176,N_2131,N_2111);
nor U3177 (N_3177,N_2686,N_2933);
nor U3178 (N_3178,N_2785,N_2640);
xnor U3179 (N_3179,N_2839,N_2315);
and U3180 (N_3180,N_2072,N_2203);
xnor U3181 (N_3181,N_2786,N_2093);
nand U3182 (N_3182,N_2590,N_2661);
nand U3183 (N_3183,N_2843,N_2518);
nand U3184 (N_3184,N_2630,N_2288);
nand U3185 (N_3185,N_2443,N_2350);
nand U3186 (N_3186,N_2418,N_2271);
or U3187 (N_3187,N_2213,N_2252);
nand U3188 (N_3188,N_2648,N_2159);
and U3189 (N_3189,N_2245,N_2361);
or U3190 (N_3190,N_2679,N_2719);
nand U3191 (N_3191,N_2929,N_2655);
xnor U3192 (N_3192,N_2537,N_2573);
nand U3193 (N_3193,N_2433,N_2812);
and U3194 (N_3194,N_2339,N_2652);
and U3195 (N_3195,N_2519,N_2865);
and U3196 (N_3196,N_2079,N_2313);
xor U3197 (N_3197,N_2860,N_2726);
xnor U3198 (N_3198,N_2936,N_2000);
xnor U3199 (N_3199,N_2806,N_2195);
nor U3200 (N_3200,N_2230,N_2402);
nor U3201 (N_3201,N_2892,N_2376);
and U3202 (N_3202,N_2234,N_2605);
nand U3203 (N_3203,N_2018,N_2556);
and U3204 (N_3204,N_2996,N_2019);
xnor U3205 (N_3205,N_2366,N_2303);
nand U3206 (N_3206,N_2457,N_2191);
xnor U3207 (N_3207,N_2877,N_2876);
or U3208 (N_3208,N_2187,N_2541);
nand U3209 (N_3209,N_2639,N_2551);
and U3210 (N_3210,N_2472,N_2375);
nor U3211 (N_3211,N_2149,N_2896);
xnor U3212 (N_3212,N_2168,N_2567);
nor U3213 (N_3213,N_2993,N_2334);
nand U3214 (N_3214,N_2216,N_2706);
xor U3215 (N_3215,N_2596,N_2971);
nand U3216 (N_3216,N_2918,N_2025);
xnor U3217 (N_3217,N_2919,N_2595);
xnor U3218 (N_3218,N_2004,N_2272);
and U3219 (N_3219,N_2298,N_2964);
nand U3220 (N_3220,N_2088,N_2677);
xor U3221 (N_3221,N_2841,N_2143);
nor U3222 (N_3222,N_2902,N_2676);
and U3223 (N_3223,N_2616,N_2878);
nand U3224 (N_3224,N_2048,N_2290);
nor U3225 (N_3225,N_2424,N_2325);
xnor U3226 (N_3226,N_2055,N_2075);
nand U3227 (N_3227,N_2312,N_2930);
nand U3228 (N_3228,N_2748,N_2513);
xnor U3229 (N_3229,N_2598,N_2372);
or U3230 (N_3230,N_2236,N_2867);
nand U3231 (N_3231,N_2791,N_2520);
or U3232 (N_3232,N_2469,N_2330);
xnor U3233 (N_3233,N_2322,N_2868);
nand U3234 (N_3234,N_2215,N_2413);
or U3235 (N_3235,N_2910,N_2094);
nand U3236 (N_3236,N_2737,N_2040);
xor U3237 (N_3237,N_2132,N_2552);
and U3238 (N_3238,N_2421,N_2830);
or U3239 (N_3239,N_2453,N_2847);
nor U3240 (N_3240,N_2024,N_2712);
nor U3241 (N_3241,N_2102,N_2193);
nor U3242 (N_3242,N_2802,N_2886);
nand U3243 (N_3243,N_2722,N_2714);
nor U3244 (N_3244,N_2179,N_2297);
nand U3245 (N_3245,N_2545,N_2991);
nor U3246 (N_3246,N_2285,N_2327);
xor U3247 (N_3247,N_2724,N_2492);
or U3248 (N_3248,N_2718,N_2047);
nand U3249 (N_3249,N_2211,N_2863);
or U3250 (N_3250,N_2296,N_2470);
nand U3251 (N_3251,N_2960,N_2412);
nor U3252 (N_3252,N_2317,N_2166);
nand U3253 (N_3253,N_2584,N_2344);
nor U3254 (N_3254,N_2627,N_2529);
xnor U3255 (N_3255,N_2958,N_2637);
nand U3256 (N_3256,N_2628,N_2992);
and U3257 (N_3257,N_2753,N_2449);
nor U3258 (N_3258,N_2939,N_2740);
nand U3259 (N_3259,N_2959,N_2059);
and U3260 (N_3260,N_2437,N_2516);
nand U3261 (N_3261,N_2730,N_2695);
nand U3262 (N_3262,N_2408,N_2398);
nand U3263 (N_3263,N_2196,N_2727);
nor U3264 (N_3264,N_2742,N_2008);
xor U3265 (N_3265,N_2027,N_2834);
nor U3266 (N_3266,N_2985,N_2074);
and U3267 (N_3267,N_2953,N_2982);
xnor U3268 (N_3268,N_2626,N_2879);
nand U3269 (N_3269,N_2618,N_2036);
nand U3270 (N_3270,N_2467,N_2221);
nor U3271 (N_3271,N_2651,N_2261);
xnor U3272 (N_3272,N_2997,N_2435);
or U3273 (N_3273,N_2710,N_2969);
xnor U3274 (N_3274,N_2246,N_2096);
or U3275 (N_3275,N_2550,N_2911);
nor U3276 (N_3276,N_2851,N_2660);
nor U3277 (N_3277,N_2114,N_2675);
nor U3278 (N_3278,N_2904,N_2005);
nor U3279 (N_3279,N_2475,N_2081);
nand U3280 (N_3280,N_2188,N_2241);
nor U3281 (N_3281,N_2318,N_2041);
nor U3282 (N_3282,N_2154,N_2787);
or U3283 (N_3283,N_2671,N_2162);
nand U3284 (N_3284,N_2819,N_2884);
nor U3285 (N_3285,N_2862,N_2814);
or U3286 (N_3286,N_2934,N_2962);
nand U3287 (N_3287,N_2304,N_2262);
xor U3288 (N_3288,N_2231,N_2903);
nand U3289 (N_3289,N_2822,N_2254);
nand U3290 (N_3290,N_2186,N_2243);
or U3291 (N_3291,N_2581,N_2429);
and U3292 (N_3292,N_2178,N_2342);
nand U3293 (N_3293,N_2386,N_2483);
xor U3294 (N_3294,N_2793,N_2696);
nor U3295 (N_3295,N_2532,N_2594);
and U3296 (N_3296,N_2684,N_2699);
nor U3297 (N_3297,N_2515,N_2440);
nand U3298 (N_3298,N_2980,N_2073);
nand U3299 (N_3299,N_2347,N_2881);
and U3300 (N_3300,N_2171,N_2981);
xnor U3301 (N_3301,N_2489,N_2650);
nor U3302 (N_3302,N_2003,N_2393);
and U3303 (N_3303,N_2274,N_2653);
and U3304 (N_3304,N_2184,N_2071);
nand U3305 (N_3305,N_2106,N_2089);
nand U3306 (N_3306,N_2508,N_2481);
nor U3307 (N_3307,N_2485,N_2938);
nor U3308 (N_3308,N_2432,N_2326);
nand U3309 (N_3309,N_2425,N_2554);
and U3310 (N_3310,N_2264,N_2848);
nand U3311 (N_3311,N_2632,N_2657);
and U3312 (N_3312,N_2693,N_2524);
nor U3313 (N_3313,N_2382,N_2600);
or U3314 (N_3314,N_2856,N_2869);
nand U3315 (N_3315,N_2871,N_2407);
nand U3316 (N_3316,N_2176,N_2189);
and U3317 (N_3317,N_2702,N_2247);
or U3318 (N_3318,N_2199,N_2763);
nor U3319 (N_3319,N_2750,N_2579);
nor U3320 (N_3320,N_2129,N_2482);
nand U3321 (N_3321,N_2984,N_2337);
and U3322 (N_3322,N_2415,N_2277);
and U3323 (N_3323,N_2888,N_2052);
or U3324 (N_3324,N_2781,N_2882);
and U3325 (N_3325,N_2857,N_2673);
nand U3326 (N_3326,N_2109,N_2854);
or U3327 (N_3327,N_2784,N_2778);
and U3328 (N_3328,N_2866,N_2681);
nand U3329 (N_3329,N_2426,N_2133);
and U3330 (N_3330,N_2732,N_2745);
nand U3331 (N_3331,N_2638,N_2404);
and U3332 (N_3332,N_2499,N_2617);
or U3333 (N_3333,N_2009,N_2765);
or U3334 (N_3334,N_2504,N_2229);
xnor U3335 (N_3335,N_2259,N_2135);
or U3336 (N_3336,N_2430,N_2656);
xor U3337 (N_3337,N_2603,N_2891);
xnor U3338 (N_3338,N_2782,N_2156);
nor U3339 (N_3339,N_2420,N_2108);
nand U3340 (N_3340,N_2941,N_2352);
and U3341 (N_3341,N_2202,N_2013);
and U3342 (N_3342,N_2951,N_2774);
nand U3343 (N_3343,N_2151,N_2098);
nor U3344 (N_3344,N_2282,N_2012);
or U3345 (N_3345,N_2029,N_2530);
and U3346 (N_3346,N_2716,N_2576);
xnor U3347 (N_3347,N_2874,N_2978);
or U3348 (N_3348,N_2333,N_2987);
or U3349 (N_3349,N_2912,N_2678);
nor U3350 (N_3350,N_2496,N_2998);
and U3351 (N_3351,N_2138,N_2838);
xor U3352 (N_3352,N_2068,N_2170);
nor U3353 (N_3353,N_2146,N_2023);
xor U3354 (N_3354,N_2731,N_2343);
and U3355 (N_3355,N_2577,N_2130);
nor U3356 (N_3356,N_2210,N_2849);
and U3357 (N_3357,N_2329,N_2670);
or U3358 (N_3358,N_2493,N_2371);
nand U3359 (N_3359,N_2536,N_2124);
xor U3360 (N_3360,N_2163,N_2458);
xnor U3361 (N_3361,N_2455,N_2963);
or U3362 (N_3362,N_2624,N_2725);
nor U3363 (N_3363,N_2474,N_2621);
or U3364 (N_3364,N_2227,N_2709);
nor U3365 (N_3365,N_2502,N_2572);
or U3366 (N_3366,N_2066,N_2527);
xor U3367 (N_3367,N_2744,N_2083);
or U3368 (N_3368,N_2773,N_2446);
and U3369 (N_3369,N_2117,N_2557);
and U3370 (N_3370,N_2080,N_2821);
and U3371 (N_3371,N_2772,N_2291);
and U3372 (N_3372,N_2487,N_2613);
xor U3373 (N_3373,N_2916,N_2054);
and U3374 (N_3374,N_2990,N_2490);
and U3375 (N_3375,N_2634,N_2999);
nor U3376 (N_3376,N_2065,N_2275);
or U3377 (N_3377,N_2566,N_2720);
nor U3378 (N_3378,N_2631,N_2955);
nand U3379 (N_3379,N_2116,N_2422);
and U3380 (N_3380,N_2217,N_2336);
nand U3381 (N_3381,N_2509,N_2165);
or U3382 (N_3382,N_2587,N_2498);
xnor U3383 (N_3383,N_2495,N_2305);
and U3384 (N_3384,N_2253,N_2340);
and U3385 (N_3385,N_2771,N_2547);
and U3386 (N_3386,N_2468,N_2973);
or U3387 (N_3387,N_2713,N_2758);
nor U3388 (N_3388,N_2826,N_2050);
xor U3389 (N_3389,N_2832,N_2931);
xor U3390 (N_3390,N_2137,N_2411);
nor U3391 (N_3391,N_2478,N_2373);
or U3392 (N_3392,N_2120,N_2069);
nor U3393 (N_3393,N_2528,N_2571);
xor U3394 (N_3394,N_2899,N_2852);
nor U3395 (N_3395,N_2668,N_2017);
nand U3396 (N_3396,N_2281,N_2349);
and U3397 (N_3397,N_2016,N_2319);
or U3398 (N_3398,N_2942,N_2683);
nand U3399 (N_3399,N_2956,N_2378);
nor U3400 (N_3400,N_2058,N_2353);
and U3401 (N_3401,N_2570,N_2549);
and U3402 (N_3402,N_2060,N_2218);
nor U3403 (N_3403,N_2306,N_2811);
nor U3404 (N_3404,N_2794,N_2943);
xor U3405 (N_3405,N_2514,N_2324);
or U3406 (N_3406,N_2825,N_2299);
or U3407 (N_3407,N_2995,N_2316);
xnor U3408 (N_3408,N_2560,N_2850);
and U3409 (N_3409,N_2062,N_2542);
and U3410 (N_3410,N_2320,N_2606);
xor U3411 (N_3411,N_2887,N_2401);
xnor U3412 (N_3412,N_2431,N_2525);
xor U3413 (N_3413,N_2607,N_2846);
nor U3414 (N_3414,N_2585,N_2105);
xor U3415 (N_3415,N_2416,N_2363);
xnor U3416 (N_3416,N_2608,N_2927);
xnor U3417 (N_3417,N_2739,N_2002);
or U3418 (N_3418,N_2687,N_2331);
nand U3419 (N_3419,N_2399,N_2456);
or U3420 (N_3420,N_2095,N_2244);
or U3421 (N_3421,N_2760,N_2669);
xnor U3422 (N_3422,N_2006,N_2733);
nand U3423 (N_3423,N_2734,N_2682);
and U3424 (N_3424,N_2905,N_2844);
nand U3425 (N_3425,N_2644,N_2454);
xnor U3426 (N_3426,N_2893,N_2691);
nand U3427 (N_3427,N_2208,N_2620);
nand U3428 (N_3428,N_2780,N_2658);
and U3429 (N_3429,N_2462,N_2379);
and U3430 (N_3430,N_2280,N_2853);
and U3431 (N_3431,N_2907,N_2801);
nand U3432 (N_3432,N_2351,N_2789);
nor U3433 (N_3433,N_2466,N_2434);
nor U3434 (N_3434,N_2224,N_2248);
or U3435 (N_3435,N_2346,N_2177);
nand U3436 (N_3436,N_2672,N_2925);
xor U3437 (N_3437,N_2099,N_2292);
or U3438 (N_3438,N_2747,N_2827);
nor U3439 (N_3439,N_2359,N_2169);
nand U3440 (N_3440,N_2240,N_2526);
nand U3441 (N_3441,N_2385,N_2610);
nand U3442 (N_3442,N_2795,N_2701);
nand U3443 (N_3443,N_2056,N_2619);
xor U3444 (N_3444,N_2182,N_2805);
and U3445 (N_3445,N_2705,N_2707);
nor U3446 (N_3446,N_2659,N_2861);
and U3447 (N_3447,N_2436,N_2500);
nor U3448 (N_3448,N_2625,N_2381);
or U3449 (N_3449,N_2553,N_2173);
nand U3450 (N_3450,N_2237,N_2736);
or U3451 (N_3451,N_2310,N_2767);
nand U3452 (N_3452,N_2809,N_2864);
and U3453 (N_3453,N_2994,N_2592);
nand U3454 (N_3454,N_2875,N_2348);
xnor U3455 (N_3455,N_2160,N_2901);
or U3456 (N_3456,N_2979,N_2383);
nand U3457 (N_3457,N_2439,N_2738);
and U3458 (N_3458,N_2354,N_2932);
xnor U3459 (N_3459,N_2870,N_2715);
and U3460 (N_3460,N_2799,N_2152);
and U3461 (N_3461,N_2766,N_2164);
and U3462 (N_3462,N_2136,N_2314);
or U3463 (N_3463,N_2167,N_2034);
nor U3464 (N_3464,N_2396,N_2623);
and U3465 (N_3465,N_2511,N_2636);
nand U3466 (N_3466,N_2232,N_2410);
or U3467 (N_3467,N_2279,N_2667);
and U3468 (N_3468,N_2057,N_2222);
and U3469 (N_3469,N_2815,N_2804);
nor U3470 (N_3470,N_2161,N_2723);
xnor U3471 (N_3471,N_2935,N_2212);
nand U3472 (N_3472,N_2622,N_2538);
xnor U3473 (N_3473,N_2338,N_2183);
nor U3474 (N_3474,N_2356,N_2286);
xnor U3475 (N_3475,N_2103,N_2872);
nand U3476 (N_3476,N_2308,N_2949);
or U3477 (N_3477,N_2779,N_2588);
and U3478 (N_3478,N_2633,N_2403);
and U3479 (N_3479,N_2460,N_2817);
nand U3480 (N_3480,N_2752,N_2558);
nand U3481 (N_3481,N_2461,N_2020);
nor U3482 (N_3482,N_2465,N_2895);
and U3483 (N_3483,N_2601,N_2926);
and U3484 (N_3484,N_2957,N_2409);
or U3485 (N_3485,N_2070,N_2007);
or U3486 (N_3486,N_2743,N_2309);
xor U3487 (N_3487,N_2966,N_2909);
nand U3488 (N_3488,N_2022,N_2569);
nor U3489 (N_3489,N_2759,N_2818);
nor U3490 (N_3490,N_2840,N_2207);
nand U3491 (N_3491,N_2501,N_2885);
nand U3492 (N_3492,N_2816,N_2021);
and U3493 (N_3493,N_2311,N_2646);
nor U3494 (N_3494,N_2200,N_2206);
and U3495 (N_3495,N_2181,N_2448);
and U3496 (N_3496,N_2113,N_2067);
nor U3497 (N_3497,N_2568,N_2833);
and U3498 (N_3498,N_2042,N_2172);
and U3499 (N_3499,N_2564,N_2950);
and U3500 (N_3500,N_2048,N_2424);
or U3501 (N_3501,N_2079,N_2457);
xnor U3502 (N_3502,N_2959,N_2619);
xnor U3503 (N_3503,N_2442,N_2143);
nor U3504 (N_3504,N_2449,N_2976);
nand U3505 (N_3505,N_2092,N_2173);
xor U3506 (N_3506,N_2939,N_2149);
xor U3507 (N_3507,N_2411,N_2776);
nand U3508 (N_3508,N_2993,N_2623);
nand U3509 (N_3509,N_2837,N_2759);
or U3510 (N_3510,N_2755,N_2868);
nor U3511 (N_3511,N_2413,N_2788);
nand U3512 (N_3512,N_2022,N_2256);
or U3513 (N_3513,N_2197,N_2510);
or U3514 (N_3514,N_2344,N_2549);
nand U3515 (N_3515,N_2703,N_2563);
or U3516 (N_3516,N_2389,N_2298);
nor U3517 (N_3517,N_2858,N_2664);
nand U3518 (N_3518,N_2897,N_2860);
nor U3519 (N_3519,N_2465,N_2025);
nand U3520 (N_3520,N_2086,N_2003);
nand U3521 (N_3521,N_2766,N_2070);
and U3522 (N_3522,N_2860,N_2881);
xnor U3523 (N_3523,N_2551,N_2379);
nand U3524 (N_3524,N_2680,N_2517);
and U3525 (N_3525,N_2796,N_2674);
xor U3526 (N_3526,N_2318,N_2701);
xnor U3527 (N_3527,N_2894,N_2509);
and U3528 (N_3528,N_2706,N_2070);
and U3529 (N_3529,N_2963,N_2706);
or U3530 (N_3530,N_2915,N_2064);
or U3531 (N_3531,N_2992,N_2942);
and U3532 (N_3532,N_2765,N_2493);
and U3533 (N_3533,N_2946,N_2801);
nor U3534 (N_3534,N_2279,N_2778);
or U3535 (N_3535,N_2551,N_2195);
or U3536 (N_3536,N_2021,N_2398);
and U3537 (N_3537,N_2438,N_2687);
or U3538 (N_3538,N_2358,N_2543);
or U3539 (N_3539,N_2250,N_2978);
nor U3540 (N_3540,N_2290,N_2932);
or U3541 (N_3541,N_2394,N_2821);
nor U3542 (N_3542,N_2509,N_2575);
nand U3543 (N_3543,N_2722,N_2573);
and U3544 (N_3544,N_2443,N_2010);
nand U3545 (N_3545,N_2460,N_2867);
nor U3546 (N_3546,N_2668,N_2141);
nand U3547 (N_3547,N_2746,N_2724);
xnor U3548 (N_3548,N_2080,N_2138);
nand U3549 (N_3549,N_2237,N_2328);
nor U3550 (N_3550,N_2209,N_2353);
and U3551 (N_3551,N_2583,N_2587);
nand U3552 (N_3552,N_2445,N_2621);
xnor U3553 (N_3553,N_2337,N_2787);
or U3554 (N_3554,N_2015,N_2191);
and U3555 (N_3555,N_2607,N_2623);
xor U3556 (N_3556,N_2117,N_2066);
nor U3557 (N_3557,N_2049,N_2478);
and U3558 (N_3558,N_2763,N_2380);
and U3559 (N_3559,N_2244,N_2908);
nand U3560 (N_3560,N_2669,N_2158);
or U3561 (N_3561,N_2131,N_2385);
and U3562 (N_3562,N_2113,N_2281);
nand U3563 (N_3563,N_2620,N_2016);
nand U3564 (N_3564,N_2254,N_2350);
and U3565 (N_3565,N_2795,N_2743);
nand U3566 (N_3566,N_2965,N_2873);
xor U3567 (N_3567,N_2688,N_2788);
or U3568 (N_3568,N_2503,N_2314);
and U3569 (N_3569,N_2823,N_2204);
and U3570 (N_3570,N_2016,N_2840);
and U3571 (N_3571,N_2441,N_2668);
and U3572 (N_3572,N_2121,N_2308);
nand U3573 (N_3573,N_2175,N_2225);
or U3574 (N_3574,N_2110,N_2761);
nand U3575 (N_3575,N_2912,N_2334);
nor U3576 (N_3576,N_2150,N_2658);
xor U3577 (N_3577,N_2551,N_2481);
and U3578 (N_3578,N_2359,N_2600);
nor U3579 (N_3579,N_2156,N_2464);
or U3580 (N_3580,N_2259,N_2612);
nand U3581 (N_3581,N_2865,N_2326);
and U3582 (N_3582,N_2022,N_2348);
or U3583 (N_3583,N_2571,N_2629);
nand U3584 (N_3584,N_2953,N_2983);
xnor U3585 (N_3585,N_2526,N_2328);
and U3586 (N_3586,N_2160,N_2428);
or U3587 (N_3587,N_2827,N_2012);
xnor U3588 (N_3588,N_2049,N_2255);
or U3589 (N_3589,N_2256,N_2194);
and U3590 (N_3590,N_2275,N_2154);
and U3591 (N_3591,N_2002,N_2810);
or U3592 (N_3592,N_2116,N_2504);
nor U3593 (N_3593,N_2098,N_2874);
nand U3594 (N_3594,N_2338,N_2064);
or U3595 (N_3595,N_2741,N_2510);
xor U3596 (N_3596,N_2944,N_2027);
xor U3597 (N_3597,N_2468,N_2340);
nand U3598 (N_3598,N_2498,N_2099);
nand U3599 (N_3599,N_2291,N_2415);
or U3600 (N_3600,N_2714,N_2400);
nand U3601 (N_3601,N_2802,N_2879);
nand U3602 (N_3602,N_2898,N_2003);
or U3603 (N_3603,N_2641,N_2959);
or U3604 (N_3604,N_2494,N_2165);
or U3605 (N_3605,N_2666,N_2230);
or U3606 (N_3606,N_2880,N_2817);
and U3607 (N_3607,N_2805,N_2054);
nor U3608 (N_3608,N_2984,N_2167);
xnor U3609 (N_3609,N_2345,N_2889);
and U3610 (N_3610,N_2998,N_2973);
and U3611 (N_3611,N_2031,N_2030);
or U3612 (N_3612,N_2919,N_2287);
nor U3613 (N_3613,N_2677,N_2746);
nand U3614 (N_3614,N_2440,N_2671);
or U3615 (N_3615,N_2722,N_2314);
and U3616 (N_3616,N_2712,N_2240);
or U3617 (N_3617,N_2676,N_2830);
or U3618 (N_3618,N_2654,N_2619);
xnor U3619 (N_3619,N_2319,N_2700);
xor U3620 (N_3620,N_2251,N_2936);
xor U3621 (N_3621,N_2106,N_2643);
or U3622 (N_3622,N_2426,N_2671);
and U3623 (N_3623,N_2898,N_2170);
and U3624 (N_3624,N_2338,N_2030);
or U3625 (N_3625,N_2733,N_2554);
and U3626 (N_3626,N_2216,N_2542);
or U3627 (N_3627,N_2741,N_2190);
nor U3628 (N_3628,N_2044,N_2714);
nand U3629 (N_3629,N_2752,N_2074);
nor U3630 (N_3630,N_2864,N_2591);
xnor U3631 (N_3631,N_2144,N_2690);
nor U3632 (N_3632,N_2686,N_2406);
and U3633 (N_3633,N_2040,N_2155);
xor U3634 (N_3634,N_2325,N_2100);
nand U3635 (N_3635,N_2577,N_2239);
or U3636 (N_3636,N_2285,N_2659);
xnor U3637 (N_3637,N_2317,N_2650);
nor U3638 (N_3638,N_2195,N_2138);
nand U3639 (N_3639,N_2887,N_2460);
nand U3640 (N_3640,N_2308,N_2993);
nand U3641 (N_3641,N_2930,N_2732);
nand U3642 (N_3642,N_2054,N_2730);
and U3643 (N_3643,N_2053,N_2074);
and U3644 (N_3644,N_2176,N_2604);
xor U3645 (N_3645,N_2496,N_2140);
nand U3646 (N_3646,N_2426,N_2769);
nor U3647 (N_3647,N_2758,N_2217);
nor U3648 (N_3648,N_2424,N_2898);
or U3649 (N_3649,N_2070,N_2638);
nor U3650 (N_3650,N_2223,N_2057);
nand U3651 (N_3651,N_2378,N_2676);
or U3652 (N_3652,N_2337,N_2267);
nand U3653 (N_3653,N_2564,N_2732);
nor U3654 (N_3654,N_2298,N_2379);
nor U3655 (N_3655,N_2842,N_2696);
and U3656 (N_3656,N_2314,N_2148);
nor U3657 (N_3657,N_2862,N_2488);
nor U3658 (N_3658,N_2450,N_2079);
nor U3659 (N_3659,N_2755,N_2267);
and U3660 (N_3660,N_2061,N_2148);
xor U3661 (N_3661,N_2031,N_2944);
nand U3662 (N_3662,N_2072,N_2661);
and U3663 (N_3663,N_2053,N_2005);
or U3664 (N_3664,N_2481,N_2473);
xor U3665 (N_3665,N_2790,N_2104);
xor U3666 (N_3666,N_2425,N_2471);
nand U3667 (N_3667,N_2350,N_2834);
xor U3668 (N_3668,N_2865,N_2610);
xnor U3669 (N_3669,N_2121,N_2466);
and U3670 (N_3670,N_2833,N_2926);
or U3671 (N_3671,N_2554,N_2398);
or U3672 (N_3672,N_2464,N_2836);
nand U3673 (N_3673,N_2732,N_2512);
nand U3674 (N_3674,N_2130,N_2608);
xnor U3675 (N_3675,N_2200,N_2821);
or U3676 (N_3676,N_2674,N_2123);
xnor U3677 (N_3677,N_2979,N_2093);
nor U3678 (N_3678,N_2670,N_2205);
nor U3679 (N_3679,N_2918,N_2874);
nand U3680 (N_3680,N_2278,N_2705);
xnor U3681 (N_3681,N_2262,N_2429);
nor U3682 (N_3682,N_2376,N_2610);
and U3683 (N_3683,N_2622,N_2964);
nand U3684 (N_3684,N_2344,N_2693);
or U3685 (N_3685,N_2538,N_2407);
nand U3686 (N_3686,N_2695,N_2541);
nor U3687 (N_3687,N_2901,N_2033);
and U3688 (N_3688,N_2726,N_2471);
and U3689 (N_3689,N_2972,N_2041);
and U3690 (N_3690,N_2856,N_2470);
nor U3691 (N_3691,N_2776,N_2001);
nand U3692 (N_3692,N_2377,N_2634);
xor U3693 (N_3693,N_2175,N_2916);
nor U3694 (N_3694,N_2469,N_2325);
nand U3695 (N_3695,N_2732,N_2570);
nand U3696 (N_3696,N_2668,N_2372);
xor U3697 (N_3697,N_2052,N_2560);
or U3698 (N_3698,N_2894,N_2948);
nand U3699 (N_3699,N_2799,N_2422);
nor U3700 (N_3700,N_2473,N_2661);
nand U3701 (N_3701,N_2240,N_2414);
and U3702 (N_3702,N_2898,N_2732);
xnor U3703 (N_3703,N_2636,N_2204);
xnor U3704 (N_3704,N_2193,N_2296);
nand U3705 (N_3705,N_2847,N_2934);
nand U3706 (N_3706,N_2117,N_2903);
and U3707 (N_3707,N_2273,N_2082);
nand U3708 (N_3708,N_2091,N_2683);
and U3709 (N_3709,N_2743,N_2621);
or U3710 (N_3710,N_2149,N_2256);
nand U3711 (N_3711,N_2226,N_2819);
or U3712 (N_3712,N_2922,N_2488);
or U3713 (N_3713,N_2380,N_2756);
and U3714 (N_3714,N_2182,N_2253);
and U3715 (N_3715,N_2559,N_2412);
nor U3716 (N_3716,N_2097,N_2197);
and U3717 (N_3717,N_2718,N_2553);
nand U3718 (N_3718,N_2432,N_2581);
nor U3719 (N_3719,N_2710,N_2591);
nand U3720 (N_3720,N_2833,N_2945);
xor U3721 (N_3721,N_2994,N_2742);
and U3722 (N_3722,N_2145,N_2770);
and U3723 (N_3723,N_2971,N_2555);
nand U3724 (N_3724,N_2101,N_2202);
or U3725 (N_3725,N_2228,N_2967);
nand U3726 (N_3726,N_2520,N_2423);
nand U3727 (N_3727,N_2012,N_2472);
nand U3728 (N_3728,N_2922,N_2381);
and U3729 (N_3729,N_2106,N_2944);
xor U3730 (N_3730,N_2462,N_2566);
and U3731 (N_3731,N_2966,N_2443);
xor U3732 (N_3732,N_2340,N_2533);
xnor U3733 (N_3733,N_2483,N_2059);
nor U3734 (N_3734,N_2921,N_2466);
xnor U3735 (N_3735,N_2361,N_2206);
nor U3736 (N_3736,N_2132,N_2423);
and U3737 (N_3737,N_2104,N_2713);
or U3738 (N_3738,N_2687,N_2750);
or U3739 (N_3739,N_2447,N_2901);
nand U3740 (N_3740,N_2680,N_2248);
nand U3741 (N_3741,N_2629,N_2460);
or U3742 (N_3742,N_2875,N_2826);
xor U3743 (N_3743,N_2468,N_2736);
nand U3744 (N_3744,N_2610,N_2762);
nor U3745 (N_3745,N_2210,N_2546);
nor U3746 (N_3746,N_2346,N_2771);
and U3747 (N_3747,N_2950,N_2980);
nor U3748 (N_3748,N_2797,N_2091);
xnor U3749 (N_3749,N_2000,N_2933);
xor U3750 (N_3750,N_2897,N_2816);
xnor U3751 (N_3751,N_2377,N_2312);
or U3752 (N_3752,N_2660,N_2669);
nor U3753 (N_3753,N_2045,N_2831);
and U3754 (N_3754,N_2221,N_2653);
and U3755 (N_3755,N_2536,N_2687);
and U3756 (N_3756,N_2316,N_2986);
or U3757 (N_3757,N_2840,N_2724);
and U3758 (N_3758,N_2433,N_2470);
nor U3759 (N_3759,N_2735,N_2798);
nand U3760 (N_3760,N_2652,N_2901);
nand U3761 (N_3761,N_2849,N_2703);
nor U3762 (N_3762,N_2914,N_2501);
xor U3763 (N_3763,N_2784,N_2329);
nand U3764 (N_3764,N_2771,N_2667);
xnor U3765 (N_3765,N_2264,N_2999);
nor U3766 (N_3766,N_2640,N_2843);
or U3767 (N_3767,N_2231,N_2870);
nor U3768 (N_3768,N_2514,N_2060);
nor U3769 (N_3769,N_2454,N_2934);
nor U3770 (N_3770,N_2612,N_2060);
xnor U3771 (N_3771,N_2887,N_2716);
xor U3772 (N_3772,N_2155,N_2701);
and U3773 (N_3773,N_2405,N_2465);
xor U3774 (N_3774,N_2953,N_2391);
nand U3775 (N_3775,N_2739,N_2825);
nand U3776 (N_3776,N_2400,N_2207);
and U3777 (N_3777,N_2460,N_2270);
and U3778 (N_3778,N_2387,N_2520);
xnor U3779 (N_3779,N_2154,N_2040);
xor U3780 (N_3780,N_2085,N_2275);
and U3781 (N_3781,N_2689,N_2105);
nand U3782 (N_3782,N_2295,N_2583);
or U3783 (N_3783,N_2645,N_2504);
xor U3784 (N_3784,N_2547,N_2134);
nor U3785 (N_3785,N_2801,N_2777);
and U3786 (N_3786,N_2273,N_2256);
and U3787 (N_3787,N_2243,N_2386);
nand U3788 (N_3788,N_2596,N_2164);
nand U3789 (N_3789,N_2002,N_2808);
or U3790 (N_3790,N_2393,N_2688);
xnor U3791 (N_3791,N_2161,N_2577);
and U3792 (N_3792,N_2650,N_2284);
or U3793 (N_3793,N_2044,N_2329);
or U3794 (N_3794,N_2220,N_2977);
xnor U3795 (N_3795,N_2045,N_2914);
nand U3796 (N_3796,N_2217,N_2404);
and U3797 (N_3797,N_2786,N_2698);
and U3798 (N_3798,N_2043,N_2297);
and U3799 (N_3799,N_2553,N_2323);
nor U3800 (N_3800,N_2893,N_2019);
xnor U3801 (N_3801,N_2012,N_2387);
nor U3802 (N_3802,N_2322,N_2389);
nand U3803 (N_3803,N_2768,N_2499);
and U3804 (N_3804,N_2297,N_2321);
or U3805 (N_3805,N_2011,N_2535);
and U3806 (N_3806,N_2072,N_2697);
and U3807 (N_3807,N_2473,N_2355);
or U3808 (N_3808,N_2759,N_2118);
and U3809 (N_3809,N_2420,N_2153);
nor U3810 (N_3810,N_2546,N_2035);
or U3811 (N_3811,N_2041,N_2598);
nor U3812 (N_3812,N_2425,N_2502);
or U3813 (N_3813,N_2894,N_2802);
nor U3814 (N_3814,N_2638,N_2649);
nand U3815 (N_3815,N_2586,N_2119);
nor U3816 (N_3816,N_2168,N_2252);
or U3817 (N_3817,N_2890,N_2296);
or U3818 (N_3818,N_2840,N_2094);
and U3819 (N_3819,N_2443,N_2363);
xnor U3820 (N_3820,N_2581,N_2502);
or U3821 (N_3821,N_2955,N_2227);
nand U3822 (N_3822,N_2718,N_2900);
and U3823 (N_3823,N_2051,N_2770);
or U3824 (N_3824,N_2376,N_2751);
or U3825 (N_3825,N_2676,N_2588);
nor U3826 (N_3826,N_2103,N_2169);
nand U3827 (N_3827,N_2008,N_2823);
nor U3828 (N_3828,N_2735,N_2127);
or U3829 (N_3829,N_2552,N_2032);
xnor U3830 (N_3830,N_2038,N_2049);
and U3831 (N_3831,N_2128,N_2190);
xnor U3832 (N_3832,N_2868,N_2533);
and U3833 (N_3833,N_2083,N_2176);
nor U3834 (N_3834,N_2753,N_2397);
nand U3835 (N_3835,N_2694,N_2051);
xnor U3836 (N_3836,N_2097,N_2233);
or U3837 (N_3837,N_2836,N_2844);
nor U3838 (N_3838,N_2429,N_2874);
or U3839 (N_3839,N_2121,N_2778);
nand U3840 (N_3840,N_2701,N_2414);
nand U3841 (N_3841,N_2966,N_2939);
or U3842 (N_3842,N_2772,N_2047);
nor U3843 (N_3843,N_2116,N_2234);
xor U3844 (N_3844,N_2206,N_2782);
nand U3845 (N_3845,N_2985,N_2143);
xnor U3846 (N_3846,N_2352,N_2164);
nor U3847 (N_3847,N_2805,N_2368);
nor U3848 (N_3848,N_2330,N_2260);
nand U3849 (N_3849,N_2490,N_2127);
nor U3850 (N_3850,N_2054,N_2191);
or U3851 (N_3851,N_2308,N_2128);
xnor U3852 (N_3852,N_2843,N_2723);
nor U3853 (N_3853,N_2448,N_2968);
and U3854 (N_3854,N_2440,N_2582);
nand U3855 (N_3855,N_2989,N_2165);
and U3856 (N_3856,N_2854,N_2918);
and U3857 (N_3857,N_2913,N_2429);
or U3858 (N_3858,N_2238,N_2766);
and U3859 (N_3859,N_2145,N_2641);
nor U3860 (N_3860,N_2146,N_2596);
and U3861 (N_3861,N_2058,N_2413);
nor U3862 (N_3862,N_2747,N_2826);
and U3863 (N_3863,N_2698,N_2565);
xnor U3864 (N_3864,N_2323,N_2219);
nand U3865 (N_3865,N_2505,N_2318);
and U3866 (N_3866,N_2500,N_2886);
or U3867 (N_3867,N_2280,N_2332);
xor U3868 (N_3868,N_2097,N_2686);
or U3869 (N_3869,N_2081,N_2201);
or U3870 (N_3870,N_2948,N_2807);
or U3871 (N_3871,N_2534,N_2397);
nand U3872 (N_3872,N_2379,N_2123);
nand U3873 (N_3873,N_2371,N_2345);
xnor U3874 (N_3874,N_2197,N_2525);
nand U3875 (N_3875,N_2685,N_2402);
or U3876 (N_3876,N_2284,N_2507);
or U3877 (N_3877,N_2816,N_2937);
or U3878 (N_3878,N_2811,N_2217);
nor U3879 (N_3879,N_2042,N_2136);
nand U3880 (N_3880,N_2044,N_2219);
nand U3881 (N_3881,N_2373,N_2984);
nor U3882 (N_3882,N_2167,N_2993);
nor U3883 (N_3883,N_2259,N_2187);
xnor U3884 (N_3884,N_2063,N_2889);
and U3885 (N_3885,N_2820,N_2898);
xor U3886 (N_3886,N_2547,N_2881);
nand U3887 (N_3887,N_2615,N_2473);
or U3888 (N_3888,N_2570,N_2149);
nand U3889 (N_3889,N_2640,N_2442);
xor U3890 (N_3890,N_2517,N_2430);
and U3891 (N_3891,N_2315,N_2092);
nor U3892 (N_3892,N_2782,N_2343);
nor U3893 (N_3893,N_2381,N_2999);
nor U3894 (N_3894,N_2225,N_2600);
and U3895 (N_3895,N_2779,N_2431);
and U3896 (N_3896,N_2737,N_2022);
nand U3897 (N_3897,N_2556,N_2678);
and U3898 (N_3898,N_2568,N_2140);
nand U3899 (N_3899,N_2320,N_2857);
nand U3900 (N_3900,N_2869,N_2663);
and U3901 (N_3901,N_2655,N_2373);
nor U3902 (N_3902,N_2490,N_2846);
nand U3903 (N_3903,N_2104,N_2625);
or U3904 (N_3904,N_2193,N_2005);
and U3905 (N_3905,N_2819,N_2447);
nand U3906 (N_3906,N_2644,N_2136);
xnor U3907 (N_3907,N_2057,N_2935);
nor U3908 (N_3908,N_2679,N_2804);
and U3909 (N_3909,N_2916,N_2642);
and U3910 (N_3910,N_2353,N_2814);
xor U3911 (N_3911,N_2139,N_2855);
xnor U3912 (N_3912,N_2454,N_2384);
nand U3913 (N_3913,N_2994,N_2591);
nor U3914 (N_3914,N_2224,N_2371);
nand U3915 (N_3915,N_2579,N_2720);
and U3916 (N_3916,N_2184,N_2660);
xor U3917 (N_3917,N_2421,N_2963);
or U3918 (N_3918,N_2994,N_2396);
and U3919 (N_3919,N_2429,N_2303);
nand U3920 (N_3920,N_2249,N_2169);
and U3921 (N_3921,N_2936,N_2276);
nor U3922 (N_3922,N_2980,N_2767);
and U3923 (N_3923,N_2964,N_2642);
and U3924 (N_3924,N_2294,N_2911);
or U3925 (N_3925,N_2878,N_2985);
nor U3926 (N_3926,N_2806,N_2165);
nand U3927 (N_3927,N_2546,N_2323);
xor U3928 (N_3928,N_2287,N_2743);
nand U3929 (N_3929,N_2682,N_2579);
or U3930 (N_3930,N_2896,N_2137);
nand U3931 (N_3931,N_2219,N_2581);
nand U3932 (N_3932,N_2583,N_2960);
and U3933 (N_3933,N_2196,N_2108);
nor U3934 (N_3934,N_2940,N_2201);
or U3935 (N_3935,N_2014,N_2004);
xor U3936 (N_3936,N_2624,N_2328);
and U3937 (N_3937,N_2412,N_2273);
nand U3938 (N_3938,N_2489,N_2013);
xor U3939 (N_3939,N_2078,N_2432);
nor U3940 (N_3940,N_2641,N_2442);
nor U3941 (N_3941,N_2784,N_2382);
xor U3942 (N_3942,N_2958,N_2508);
and U3943 (N_3943,N_2755,N_2029);
and U3944 (N_3944,N_2559,N_2505);
and U3945 (N_3945,N_2134,N_2104);
or U3946 (N_3946,N_2909,N_2402);
xnor U3947 (N_3947,N_2755,N_2832);
or U3948 (N_3948,N_2821,N_2446);
nor U3949 (N_3949,N_2820,N_2344);
nor U3950 (N_3950,N_2802,N_2846);
nor U3951 (N_3951,N_2803,N_2215);
nor U3952 (N_3952,N_2977,N_2111);
and U3953 (N_3953,N_2262,N_2254);
nor U3954 (N_3954,N_2736,N_2326);
or U3955 (N_3955,N_2872,N_2372);
nand U3956 (N_3956,N_2944,N_2011);
nor U3957 (N_3957,N_2862,N_2366);
or U3958 (N_3958,N_2230,N_2705);
nand U3959 (N_3959,N_2646,N_2261);
nor U3960 (N_3960,N_2518,N_2776);
nor U3961 (N_3961,N_2407,N_2508);
or U3962 (N_3962,N_2534,N_2900);
and U3963 (N_3963,N_2275,N_2743);
nor U3964 (N_3964,N_2781,N_2334);
and U3965 (N_3965,N_2851,N_2448);
and U3966 (N_3966,N_2500,N_2374);
and U3967 (N_3967,N_2560,N_2357);
or U3968 (N_3968,N_2541,N_2206);
nor U3969 (N_3969,N_2930,N_2694);
nor U3970 (N_3970,N_2410,N_2717);
nor U3971 (N_3971,N_2955,N_2778);
nor U3972 (N_3972,N_2825,N_2997);
xnor U3973 (N_3973,N_2265,N_2009);
or U3974 (N_3974,N_2986,N_2950);
nand U3975 (N_3975,N_2565,N_2003);
nor U3976 (N_3976,N_2834,N_2750);
nor U3977 (N_3977,N_2650,N_2892);
and U3978 (N_3978,N_2937,N_2943);
or U3979 (N_3979,N_2990,N_2610);
and U3980 (N_3980,N_2069,N_2304);
nor U3981 (N_3981,N_2183,N_2924);
and U3982 (N_3982,N_2660,N_2083);
xor U3983 (N_3983,N_2548,N_2582);
xnor U3984 (N_3984,N_2973,N_2559);
and U3985 (N_3985,N_2351,N_2078);
nand U3986 (N_3986,N_2557,N_2308);
or U3987 (N_3987,N_2925,N_2335);
nand U3988 (N_3988,N_2625,N_2195);
and U3989 (N_3989,N_2672,N_2642);
and U3990 (N_3990,N_2046,N_2597);
or U3991 (N_3991,N_2813,N_2160);
nand U3992 (N_3992,N_2340,N_2930);
nand U3993 (N_3993,N_2370,N_2847);
and U3994 (N_3994,N_2504,N_2111);
nor U3995 (N_3995,N_2961,N_2053);
and U3996 (N_3996,N_2558,N_2805);
nor U3997 (N_3997,N_2264,N_2181);
nand U3998 (N_3998,N_2534,N_2550);
or U3999 (N_3999,N_2023,N_2861);
nor U4000 (N_4000,N_3065,N_3616);
nor U4001 (N_4001,N_3774,N_3486);
and U4002 (N_4002,N_3802,N_3717);
xnor U4003 (N_4003,N_3607,N_3861);
and U4004 (N_4004,N_3565,N_3702);
or U4005 (N_4005,N_3442,N_3892);
nand U4006 (N_4006,N_3675,N_3686);
nand U4007 (N_4007,N_3636,N_3356);
and U4008 (N_4008,N_3160,N_3258);
nor U4009 (N_4009,N_3757,N_3429);
or U4010 (N_4010,N_3804,N_3230);
or U4011 (N_4011,N_3974,N_3282);
xor U4012 (N_4012,N_3700,N_3495);
nor U4013 (N_4013,N_3621,N_3452);
and U4014 (N_4014,N_3790,N_3186);
or U4015 (N_4015,N_3481,N_3149);
nand U4016 (N_4016,N_3448,N_3959);
nor U4017 (N_4017,N_3826,N_3660);
and U4018 (N_4018,N_3887,N_3390);
or U4019 (N_4019,N_3900,N_3142);
nor U4020 (N_4020,N_3745,N_3658);
and U4021 (N_4021,N_3140,N_3270);
xor U4022 (N_4022,N_3935,N_3051);
nor U4023 (N_4023,N_3419,N_3195);
xnor U4024 (N_4024,N_3551,N_3680);
nand U4025 (N_4025,N_3013,N_3848);
nor U4026 (N_4026,N_3317,N_3432);
and U4027 (N_4027,N_3446,N_3285);
and U4028 (N_4028,N_3005,N_3685);
nand U4029 (N_4029,N_3350,N_3241);
and U4030 (N_4030,N_3523,N_3601);
xnor U4031 (N_4031,N_3605,N_3278);
nor U4032 (N_4032,N_3336,N_3237);
and U4033 (N_4033,N_3044,N_3889);
and U4034 (N_4034,N_3875,N_3595);
nor U4035 (N_4035,N_3520,N_3944);
nor U4036 (N_4036,N_3067,N_3096);
xnor U4037 (N_4037,N_3535,N_3733);
nor U4038 (N_4038,N_3943,N_3344);
xnor U4039 (N_4039,N_3379,N_3009);
or U4040 (N_4040,N_3076,N_3247);
nand U4041 (N_4041,N_3990,N_3644);
or U4042 (N_4042,N_3995,N_3633);
xnor U4043 (N_4043,N_3184,N_3425);
and U4044 (N_4044,N_3870,N_3951);
and U4045 (N_4045,N_3938,N_3279);
xnor U4046 (N_4046,N_3460,N_3928);
xnor U4047 (N_4047,N_3192,N_3805);
nand U4048 (N_4048,N_3271,N_3866);
nor U4049 (N_4049,N_3820,N_3054);
and U4050 (N_4050,N_3365,N_3347);
xor U4051 (N_4051,N_3631,N_3079);
nand U4052 (N_4052,N_3075,N_3619);
and U4053 (N_4053,N_3458,N_3896);
or U4054 (N_4054,N_3583,N_3464);
nor U4055 (N_4055,N_3272,N_3570);
nand U4056 (N_4056,N_3921,N_3123);
nand U4057 (N_4057,N_3868,N_3785);
nand U4058 (N_4058,N_3791,N_3806);
nand U4059 (N_4059,N_3440,N_3941);
nor U4060 (N_4060,N_3867,N_3321);
nor U4061 (N_4061,N_3634,N_3590);
nor U4062 (N_4062,N_3764,N_3420);
xor U4063 (N_4063,N_3954,N_3093);
nor U4064 (N_4064,N_3226,N_3871);
xnor U4065 (N_4065,N_3476,N_3880);
or U4066 (N_4066,N_3510,N_3152);
or U4067 (N_4067,N_3787,N_3980);
or U4068 (N_4068,N_3594,N_3087);
nand U4069 (N_4069,N_3933,N_3228);
xnor U4070 (N_4070,N_3988,N_3800);
nor U4071 (N_4071,N_3740,N_3626);
nand U4072 (N_4072,N_3857,N_3414);
and U4073 (N_4073,N_3275,N_3413);
or U4074 (N_4074,N_3337,N_3406);
nor U4075 (N_4075,N_3055,N_3630);
xnor U4076 (N_4076,N_3524,N_3796);
xor U4077 (N_4077,N_3654,N_3412);
xnor U4078 (N_4078,N_3860,N_3765);
and U4079 (N_4079,N_3451,N_3885);
nor U4080 (N_4080,N_3086,N_3238);
nand U4081 (N_4081,N_3224,N_3743);
nand U4082 (N_4082,N_3080,N_3391);
xnor U4083 (N_4083,N_3670,N_3372);
and U4084 (N_4084,N_3109,N_3457);
or U4085 (N_4085,N_3699,N_3308);
nand U4086 (N_4086,N_3752,N_3507);
and U4087 (N_4087,N_3261,N_3483);
or U4088 (N_4088,N_3937,N_3821);
and U4089 (N_4089,N_3137,N_3666);
or U4090 (N_4090,N_3903,N_3094);
nand U4091 (N_4091,N_3841,N_3695);
xor U4092 (N_4092,N_3479,N_3610);
nor U4093 (N_4093,N_3737,N_3383);
or U4094 (N_4094,N_3681,N_3894);
nand U4095 (N_4095,N_3297,N_3789);
nand U4096 (N_4096,N_3314,N_3557);
nand U4097 (N_4097,N_3244,N_3166);
or U4098 (N_4098,N_3588,N_3130);
nand U4099 (N_4099,N_3537,N_3053);
or U4100 (N_4100,N_3734,N_3940);
nor U4101 (N_4101,N_3639,N_3389);
or U4102 (N_4102,N_3615,N_3216);
and U4103 (N_4103,N_3746,N_3577);
and U4104 (N_4104,N_3924,N_3792);
xor U4105 (N_4105,N_3664,N_3795);
or U4106 (N_4106,N_3918,N_3319);
nor U4107 (N_4107,N_3533,N_3931);
xnor U4108 (N_4108,N_3978,N_3694);
or U4109 (N_4109,N_3649,N_3597);
nor U4110 (N_4110,N_3910,N_3772);
xor U4111 (N_4111,N_3380,N_3568);
nand U4112 (N_4112,N_3388,N_3326);
nor U4113 (N_4113,N_3946,N_3183);
nor U4114 (N_4114,N_3421,N_3330);
or U4115 (N_4115,N_3437,N_3274);
and U4116 (N_4116,N_3267,N_3089);
or U4117 (N_4117,N_3068,N_3444);
nand U4118 (N_4118,N_3538,N_3828);
or U4119 (N_4119,N_3602,N_3839);
xnor U4120 (N_4120,N_3180,N_3422);
nor U4121 (N_4121,N_3713,N_3083);
or U4122 (N_4122,N_3002,N_3541);
or U4123 (N_4123,N_3478,N_3163);
xor U4124 (N_4124,N_3655,N_3512);
xor U4125 (N_4125,N_3898,N_3961);
xnor U4126 (N_4126,N_3581,N_3480);
and U4127 (N_4127,N_3416,N_3555);
xnor U4128 (N_4128,N_3129,N_3084);
nor U4129 (N_4129,N_3807,N_3017);
xnor U4130 (N_4130,N_3584,N_3286);
and U4131 (N_4131,N_3307,N_3677);
and U4132 (N_4132,N_3987,N_3957);
xnor U4133 (N_4133,N_3148,N_3975);
nor U4134 (N_4134,N_3121,N_3563);
xor U4135 (N_4135,N_3641,N_3852);
and U4136 (N_4136,N_3225,N_3667);
and U4137 (N_4137,N_3811,N_3788);
nand U4138 (N_4138,N_3032,N_3052);
nand U4139 (N_4139,N_3450,N_3118);
xor U4140 (N_4140,N_3291,N_3172);
xor U4141 (N_4141,N_3834,N_3914);
or U4142 (N_4142,N_3998,N_3977);
xnor U4143 (N_4143,N_3742,N_3467);
nor U4144 (N_4144,N_3404,N_3612);
nor U4145 (N_4145,N_3108,N_3447);
and U4146 (N_4146,N_3780,N_3728);
nand U4147 (N_4147,N_3659,N_3808);
xor U4148 (N_4148,N_3441,N_3474);
or U4149 (N_4149,N_3313,N_3045);
nand U4150 (N_4150,N_3357,N_3124);
or U4151 (N_4151,N_3876,N_3643);
xnor U4152 (N_4152,N_3505,N_3428);
xor U4153 (N_4153,N_3882,N_3179);
or U4154 (N_4154,N_3922,N_3126);
and U4155 (N_4155,N_3628,N_3823);
xnor U4156 (N_4156,N_3374,N_3251);
or U4157 (N_4157,N_3037,N_3622);
or U4158 (N_4158,N_3212,N_3306);
or U4159 (N_4159,N_3682,N_3611);
xor U4160 (N_4160,N_3298,N_3345);
and U4161 (N_4161,N_3661,N_3689);
and U4162 (N_4162,N_3145,N_3955);
and U4163 (N_4163,N_3221,N_3909);
nand U4164 (N_4164,N_3007,N_3503);
nand U4165 (N_4165,N_3168,N_3092);
xnor U4166 (N_4166,N_3066,N_3198);
nand U4167 (N_4167,N_3691,N_3901);
nand U4168 (N_4168,N_3242,N_3606);
xor U4169 (N_4169,N_3574,N_3335);
nand U4170 (N_4170,N_3836,N_3239);
and U4171 (N_4171,N_3339,N_3672);
nand U4172 (N_4172,N_3328,N_3793);
xnor U4173 (N_4173,N_3292,N_3646);
and U4174 (N_4174,N_3283,N_3731);
nand U4175 (N_4175,N_3135,N_3603);
and U4176 (N_4176,N_3105,N_3814);
nand U4177 (N_4177,N_3354,N_3647);
nand U4178 (N_4178,N_3418,N_3926);
xor U4179 (N_4179,N_3508,N_3276);
or U4180 (N_4180,N_3469,N_3041);
or U4181 (N_4181,N_3942,N_3958);
and U4182 (N_4182,N_3090,N_3552);
or U4183 (N_4183,N_3254,N_3854);
or U4184 (N_4184,N_3167,N_3562);
or U4185 (N_4185,N_3531,N_3593);
and U4186 (N_4186,N_3240,N_3468);
xor U4187 (N_4187,N_3651,N_3770);
or U4188 (N_4188,N_3515,N_3705);
nor U4189 (N_4189,N_3436,N_3930);
xor U4190 (N_4190,N_3057,N_3015);
nor U4191 (N_4191,N_3579,N_3150);
xnor U4192 (N_4192,N_3561,N_3214);
nor U4193 (N_4193,N_3360,N_3599);
xor U4194 (N_4194,N_3022,N_3100);
nand U4195 (N_4195,N_3984,N_3618);
nand U4196 (N_4196,N_3801,N_3099);
nand U4197 (N_4197,N_3039,N_3426);
nand U4198 (N_4198,N_3608,N_3684);
or U4199 (N_4199,N_3560,N_3434);
xor U4200 (N_4200,N_3704,N_3494);
xnor U4201 (N_4201,N_3604,N_3056);
and U4202 (N_4202,N_3913,N_3676);
nor U4203 (N_4203,N_3683,N_3174);
nor U4204 (N_4204,N_3262,N_3578);
and U4205 (N_4205,N_3762,N_3164);
nand U4206 (N_4206,N_3915,N_3217);
nor U4207 (N_4207,N_3950,N_3582);
xor U4208 (N_4208,N_3830,N_3521);
nand U4209 (N_4209,N_3200,N_3732);
xnor U4210 (N_4210,N_3569,N_3662);
or U4211 (N_4211,N_3019,N_3753);
nor U4212 (N_4212,N_3956,N_3156);
nor U4213 (N_4213,N_3316,N_3250);
xor U4214 (N_4214,N_3288,N_3587);
nand U4215 (N_4215,N_3025,N_3653);
xor U4216 (N_4216,N_3818,N_3073);
nand U4217 (N_4217,N_3449,N_3960);
and U4218 (N_4218,N_3210,N_3257);
nand U4219 (N_4219,N_3373,N_3318);
xor U4220 (N_4220,N_3844,N_3119);
nor U4221 (N_4221,N_3349,N_3899);
or U4222 (N_4222,N_3750,N_3912);
nor U4223 (N_4223,N_3132,N_3969);
or U4224 (N_4224,N_3829,N_3033);
and U4225 (N_4225,N_3177,N_3331);
nand U4226 (N_4226,N_3222,N_3060);
and U4227 (N_4227,N_3359,N_3465);
and U4228 (N_4228,N_3632,N_3280);
xnor U4229 (N_4229,N_3169,N_3263);
nand U4230 (N_4230,N_3236,N_3847);
nor U4231 (N_4231,N_3338,N_3923);
or U4232 (N_4232,N_3652,N_3502);
or U4233 (N_4233,N_3727,N_3231);
and U4234 (N_4234,N_3273,N_3424);
xor U4235 (N_4235,N_3989,N_3971);
and U4236 (N_4236,N_3491,N_3352);
xor U4237 (N_4237,N_3966,N_3863);
nor U4238 (N_4238,N_3598,N_3264);
and U4239 (N_4239,N_3739,N_3062);
nor U4240 (N_4240,N_3548,N_3819);
nor U4241 (N_4241,N_3725,N_3289);
xnor U4242 (N_4242,N_3783,N_3884);
nand U4243 (N_4243,N_3229,N_3485);
or U4244 (N_4244,N_3377,N_3919);
and U4245 (N_4245,N_3382,N_3799);
or U4246 (N_4246,N_3706,N_3994);
xor U4247 (N_4247,N_3077,N_3114);
nor U4248 (N_4248,N_3435,N_3766);
and U4249 (N_4249,N_3620,N_3245);
or U4250 (N_4250,N_3845,N_3034);
nor U4251 (N_4251,N_3962,N_3206);
or U4252 (N_4252,N_3650,N_3014);
and U4253 (N_4253,N_3473,N_3856);
and U4254 (N_4254,N_3175,N_3157);
and U4255 (N_4255,N_3106,N_3453);
nand U4256 (N_4256,N_3749,N_3720);
nor U4257 (N_4257,N_3853,N_3088);
nor U4258 (N_4258,N_3572,N_3072);
nor U4259 (N_4259,N_3904,N_3061);
nand U4260 (N_4260,N_3098,N_3546);
and U4261 (N_4261,N_3952,N_3635);
nand U4262 (N_4262,N_3387,N_3897);
nand U4263 (N_4263,N_3190,N_3895);
and U4264 (N_4264,N_3532,N_3081);
nand U4265 (N_4265,N_3368,N_3456);
and U4266 (N_4266,N_3663,N_3050);
xor U4267 (N_4267,N_3063,N_3322);
nand U4268 (N_4268,N_3320,N_3542);
and U4269 (N_4269,N_3300,N_3202);
or U4270 (N_4270,N_3310,N_3775);
and U4271 (N_4271,N_3679,N_3196);
nand U4272 (N_4272,N_3295,N_3095);
or U4273 (N_4273,N_3996,N_3735);
and U4274 (N_4274,N_3837,N_3953);
and U4275 (N_4275,N_3835,N_3711);
nor U4276 (N_4276,N_3375,N_3128);
nor U4277 (N_4277,N_3623,N_3591);
or U4278 (N_4278,N_3397,N_3769);
nor U4279 (N_4279,N_3536,N_3511);
and U4280 (N_4280,N_3692,N_3656);
nand U4281 (N_4281,N_3405,N_3431);
and U4282 (N_4282,N_3115,N_3540);
xor U4283 (N_4283,N_3763,N_3873);
xor U4284 (N_4284,N_3116,N_3609);
nand U4285 (N_4285,N_3268,N_3751);
and U4286 (N_4286,N_3293,N_3147);
nor U4287 (N_4287,N_3155,N_3235);
nand U4288 (N_4288,N_3193,N_3248);
nor U4289 (N_4289,N_3776,N_3269);
nand U4290 (N_4290,N_3417,N_3462);
nand U4291 (N_4291,N_3755,N_3199);
and U4292 (N_4292,N_3514,N_3327);
or U4293 (N_4293,N_3883,N_3657);
nor U4294 (N_4294,N_3690,N_3991);
nor U4295 (N_4295,N_3864,N_3840);
nand U4296 (N_4296,N_3803,N_3454);
nand U4297 (N_4297,N_3171,N_3613);
and U4298 (N_4298,N_3187,N_3394);
xor U4299 (N_4299,N_3869,N_3550);
or U4300 (N_4300,N_3302,N_3754);
nand U4301 (N_4301,N_3078,N_3112);
nand U4302 (N_4302,N_3046,N_3916);
and U4303 (N_4303,N_3500,N_3558);
nor U4304 (N_4304,N_3211,N_3234);
and U4305 (N_4305,N_3920,N_3284);
and U4306 (N_4306,N_3255,N_3110);
and U4307 (N_4307,N_3744,N_3049);
and U4308 (N_4308,N_3246,N_3817);
nor U4309 (N_4309,N_3153,N_3010);
nor U4310 (N_4310,N_3091,N_3771);
nor U4311 (N_4311,N_3484,N_3809);
nor U4312 (N_4312,N_3340,N_3362);
nand U4313 (N_4313,N_3724,N_3648);
or U4314 (N_4314,N_3985,N_3929);
and U4315 (N_4315,N_3410,N_3567);
nor U4316 (N_4316,N_3812,N_3949);
or U4317 (N_4317,N_3008,N_3981);
nand U4318 (N_4318,N_3773,N_3201);
nor U4319 (N_4319,N_3035,N_3525);
xnor U4320 (N_4320,N_3838,N_3346);
or U4321 (N_4321,N_3369,N_3006);
xnor U4322 (N_4322,N_3312,N_3223);
or U4323 (N_4323,N_3718,N_3948);
or U4324 (N_4324,N_3461,N_3408);
nor U4325 (N_4325,N_3696,N_3997);
and U4326 (N_4326,N_3784,N_3207);
xnor U4327 (N_4327,N_3194,N_3471);
nor U4328 (N_4328,N_3526,N_3736);
or U4329 (N_4329,N_3498,N_3516);
nand U4330 (N_4330,N_3999,N_3294);
xor U4331 (N_4331,N_3085,N_3138);
nor U4332 (N_4332,N_3120,N_3760);
nand U4333 (N_4333,N_3965,N_3716);
nor U4334 (N_4334,N_3208,N_3188);
or U4335 (N_4335,N_3253,N_3544);
and U4336 (N_4336,N_3182,N_3439);
nand U4337 (N_4337,N_3392,N_3709);
and U4338 (N_4338,N_3290,N_3758);
and U4339 (N_4339,N_3497,N_3723);
nor U4340 (N_4340,N_3509,N_3842);
nand U4341 (N_4341,N_3355,N_3325);
xor U4342 (N_4342,N_3393,N_3069);
nand U4343 (N_4343,N_3596,N_3266);
or U4344 (N_4344,N_3058,N_3107);
and U4345 (N_4345,N_3968,N_3134);
and U4346 (N_4346,N_3693,N_3906);
nor U4347 (N_4347,N_3455,N_3122);
or U4348 (N_4348,N_3580,N_3554);
and U4349 (N_4349,N_3566,N_3833);
or U4350 (N_4350,N_3191,N_3043);
and U4351 (N_4351,N_3071,N_3499);
or U4352 (N_4352,N_3012,N_3674);
or U4353 (N_4353,N_3703,N_3824);
and U4354 (N_4354,N_3165,N_3233);
or U4355 (N_4355,N_3865,N_3024);
nand U4356 (N_4356,N_3136,N_3333);
or U4357 (N_4357,N_3721,N_3047);
xnor U4358 (N_4358,N_3779,N_3070);
nor U4359 (N_4359,N_3000,N_3260);
xor U4360 (N_4360,N_3399,N_3185);
or U4361 (N_4361,N_3026,N_3204);
nand U4362 (N_4362,N_3232,N_3983);
or U4363 (N_4363,N_3589,N_3178);
and U4364 (N_4364,N_3627,N_3992);
or U4365 (N_4365,N_3522,N_3296);
or U4366 (N_4366,N_3688,N_3850);
nor U4367 (N_4367,N_3517,N_3370);
nand U4368 (N_4368,N_3011,N_3879);
xor U4369 (N_4369,N_3712,N_3205);
and U4370 (N_4370,N_3342,N_3501);
xnor U4371 (N_4371,N_3074,N_3348);
nor U4372 (N_4372,N_3518,N_3381);
nand U4373 (N_4373,N_3872,N_3710);
xor U4374 (N_4374,N_3097,N_3181);
xor U4375 (N_4375,N_3637,N_3890);
nor U4376 (N_4376,N_3496,N_3741);
nor U4377 (N_4377,N_3549,N_3492);
xnor U4378 (N_4378,N_3001,N_3443);
xnor U4379 (N_4379,N_3963,N_3714);
or U4380 (N_4380,N_3893,N_3874);
and U4381 (N_4381,N_3016,N_3559);
nor U4382 (N_4382,N_3825,N_3385);
nor U4383 (N_4383,N_3030,N_3028);
nor U4384 (N_4384,N_3970,N_3299);
or U4385 (N_4385,N_3888,N_3701);
or U4386 (N_4386,N_3729,N_3665);
or U4387 (N_4387,N_3127,N_3220);
or U4388 (N_4388,N_3539,N_3301);
xnor U4389 (N_4389,N_3048,N_3982);
nand U4390 (N_4390,N_3738,N_3101);
nand U4391 (N_4391,N_3143,N_3475);
nand U4392 (N_4392,N_3151,N_3891);
or U4393 (N_4393,N_3378,N_3343);
and U4394 (N_4394,N_3719,N_3463);
and U4395 (N_4395,N_3427,N_3529);
xor U4396 (N_4396,N_3158,N_3846);
nand U4397 (N_4397,N_3423,N_3911);
or U4398 (N_4398,N_3020,N_3947);
nor U4399 (N_4399,N_3315,N_3925);
and U4400 (N_4400,N_3213,N_3161);
nor U4401 (N_4401,N_3722,N_3708);
and U4402 (N_4402,N_3575,N_3967);
and U4403 (N_4403,N_3881,N_3878);
and U4404 (N_4404,N_3341,N_3102);
xor U4405 (N_4405,N_3396,N_3945);
xnor U4406 (N_4406,N_3329,N_3671);
and U4407 (N_4407,N_3939,N_3530);
nor U4408 (N_4408,N_3778,N_3877);
nand U4409 (N_4409,N_3936,N_3173);
xnor U4410 (N_4410,N_3082,N_3459);
or U4411 (N_4411,N_3932,N_3614);
nor U4412 (N_4412,N_3794,N_3504);
nand U4413 (N_4413,N_3402,N_3029);
or U4414 (N_4414,N_3902,N_3576);
xor U4415 (N_4415,N_3858,N_3018);
and U4416 (N_4416,N_3843,N_3040);
nand U4417 (N_4417,N_3361,N_3748);
and U4418 (N_4418,N_3403,N_3400);
or U4419 (N_4419,N_3592,N_3332);
and U4420 (N_4420,N_3859,N_3125);
nand U4421 (N_4421,N_3642,N_3287);
or U4422 (N_4422,N_3543,N_3004);
nor U4423 (N_4423,N_3917,N_3358);
or U4424 (N_4424,N_3934,N_3993);
nor U4425 (N_4425,N_3488,N_3064);
nor U4426 (N_4426,N_3027,N_3144);
or U4427 (N_4427,N_3133,N_3218);
nor U4428 (N_4428,N_3305,N_3747);
or U4429 (N_4429,N_3798,N_3038);
nand U4430 (N_4430,N_3490,N_3023);
and U4431 (N_4431,N_3227,N_3986);
and U4432 (N_4432,N_3401,N_3810);
nand U4433 (N_4433,N_3827,N_3629);
or U4434 (N_4434,N_3862,N_3219);
or U4435 (N_4435,N_3031,N_3907);
xnor U4436 (N_4436,N_3493,N_3265);
xnor U4437 (N_4437,N_3489,N_3687);
or U4438 (N_4438,N_3281,N_3176);
nor U4439 (N_4439,N_3767,N_3252);
and U4440 (N_4440,N_3777,N_3527);
xor U4441 (N_4441,N_3438,N_3600);
or U4442 (N_4442,N_3756,N_3534);
nand U4443 (N_4443,N_3813,N_3303);
nor U4444 (N_4444,N_3506,N_3972);
nor U4445 (N_4445,N_3851,N_3249);
xnor U4446 (N_4446,N_3973,N_3976);
nand U4447 (N_4447,N_3886,N_3215);
xnor U4448 (N_4448,N_3832,N_3831);
and U4449 (N_4449,N_3964,N_3395);
nor U4450 (N_4450,N_3466,N_3624);
and U4451 (N_4451,N_3117,N_3409);
nand U4452 (N_4452,N_3376,N_3797);
and U4453 (N_4453,N_3131,N_3513);
or U4454 (N_4454,N_3849,N_3759);
or U4455 (N_4455,N_3154,N_3556);
nand U4456 (N_4456,N_3715,N_3927);
and U4457 (N_4457,N_3707,N_3189);
xnor U4458 (N_4458,N_3203,N_3324);
nor U4459 (N_4459,N_3645,N_3673);
xor U4460 (N_4460,N_3786,N_3141);
xnor U4461 (N_4461,N_3364,N_3617);
xnor U4462 (N_4462,N_3698,N_3761);
nand U4463 (N_4463,N_3640,N_3547);
or U4464 (N_4464,N_3519,N_3036);
nand U4465 (N_4465,N_3669,N_3482);
and U4466 (N_4466,N_3477,N_3528);
or U4467 (N_4467,N_3855,N_3256);
nand U4468 (N_4468,N_3781,N_3564);
nor U4469 (N_4469,N_3334,N_3545);
nor U4470 (N_4470,N_3304,N_3768);
or U4471 (N_4471,N_3170,N_3625);
nor U4472 (N_4472,N_3059,N_3553);
nor U4473 (N_4473,N_3470,N_3726);
xnor U4474 (N_4474,N_3209,N_3309);
xor U4475 (N_4475,N_3197,N_3351);
and U4476 (N_4476,N_3585,N_3908);
xor U4477 (N_4477,N_3678,N_3433);
nor U4478 (N_4478,N_3103,N_3146);
and U4479 (N_4479,N_3822,N_3311);
nand U4480 (N_4480,N_3586,N_3386);
or U4481 (N_4481,N_3415,N_3782);
nand U4482 (N_4482,N_3104,N_3363);
or U4483 (N_4483,N_3243,N_3139);
and U4484 (N_4484,N_3697,N_3366);
nand U4485 (N_4485,N_3571,N_3668);
nor U4486 (N_4486,N_3815,N_3353);
xor U4487 (N_4487,N_3638,N_3111);
nand U4488 (N_4488,N_3367,N_3472);
or U4489 (N_4489,N_3398,N_3979);
and U4490 (N_4490,N_3159,N_3277);
nor U4491 (N_4491,N_3573,N_3371);
nand U4492 (N_4492,N_3021,N_3430);
nor U4493 (N_4493,N_3003,N_3905);
nand U4494 (N_4494,N_3816,N_3487);
and U4495 (N_4495,N_3162,N_3411);
and U4496 (N_4496,N_3113,N_3323);
or U4497 (N_4497,N_3445,N_3259);
nor U4498 (N_4498,N_3407,N_3730);
nor U4499 (N_4499,N_3042,N_3384);
nand U4500 (N_4500,N_3169,N_3484);
and U4501 (N_4501,N_3887,N_3842);
nand U4502 (N_4502,N_3608,N_3622);
or U4503 (N_4503,N_3453,N_3591);
nand U4504 (N_4504,N_3540,N_3344);
and U4505 (N_4505,N_3196,N_3884);
xor U4506 (N_4506,N_3180,N_3687);
xnor U4507 (N_4507,N_3694,N_3237);
or U4508 (N_4508,N_3031,N_3819);
and U4509 (N_4509,N_3735,N_3874);
or U4510 (N_4510,N_3187,N_3014);
or U4511 (N_4511,N_3398,N_3104);
or U4512 (N_4512,N_3643,N_3582);
nand U4513 (N_4513,N_3829,N_3614);
or U4514 (N_4514,N_3024,N_3868);
xor U4515 (N_4515,N_3695,N_3572);
xor U4516 (N_4516,N_3697,N_3445);
and U4517 (N_4517,N_3038,N_3023);
and U4518 (N_4518,N_3217,N_3927);
xnor U4519 (N_4519,N_3300,N_3891);
and U4520 (N_4520,N_3324,N_3037);
and U4521 (N_4521,N_3625,N_3050);
nand U4522 (N_4522,N_3309,N_3836);
xnor U4523 (N_4523,N_3403,N_3739);
xor U4524 (N_4524,N_3686,N_3823);
xor U4525 (N_4525,N_3427,N_3511);
or U4526 (N_4526,N_3817,N_3807);
and U4527 (N_4527,N_3806,N_3845);
nor U4528 (N_4528,N_3315,N_3161);
nand U4529 (N_4529,N_3758,N_3157);
nor U4530 (N_4530,N_3407,N_3069);
nand U4531 (N_4531,N_3357,N_3189);
nand U4532 (N_4532,N_3617,N_3529);
nor U4533 (N_4533,N_3982,N_3209);
and U4534 (N_4534,N_3039,N_3301);
nand U4535 (N_4535,N_3375,N_3112);
nor U4536 (N_4536,N_3243,N_3921);
xor U4537 (N_4537,N_3971,N_3130);
nand U4538 (N_4538,N_3022,N_3718);
or U4539 (N_4539,N_3834,N_3125);
xnor U4540 (N_4540,N_3456,N_3880);
nor U4541 (N_4541,N_3058,N_3144);
and U4542 (N_4542,N_3056,N_3212);
nand U4543 (N_4543,N_3820,N_3847);
and U4544 (N_4544,N_3564,N_3466);
nand U4545 (N_4545,N_3245,N_3155);
or U4546 (N_4546,N_3175,N_3599);
xnor U4547 (N_4547,N_3191,N_3366);
or U4548 (N_4548,N_3235,N_3510);
or U4549 (N_4549,N_3983,N_3026);
xnor U4550 (N_4550,N_3979,N_3191);
xnor U4551 (N_4551,N_3974,N_3290);
nor U4552 (N_4552,N_3059,N_3411);
nor U4553 (N_4553,N_3703,N_3154);
and U4554 (N_4554,N_3895,N_3808);
or U4555 (N_4555,N_3106,N_3807);
or U4556 (N_4556,N_3149,N_3058);
and U4557 (N_4557,N_3295,N_3822);
nand U4558 (N_4558,N_3791,N_3365);
nand U4559 (N_4559,N_3983,N_3191);
nand U4560 (N_4560,N_3036,N_3740);
nor U4561 (N_4561,N_3475,N_3160);
or U4562 (N_4562,N_3200,N_3146);
xnor U4563 (N_4563,N_3568,N_3879);
and U4564 (N_4564,N_3982,N_3424);
nor U4565 (N_4565,N_3213,N_3122);
or U4566 (N_4566,N_3222,N_3128);
xnor U4567 (N_4567,N_3982,N_3217);
and U4568 (N_4568,N_3223,N_3453);
xor U4569 (N_4569,N_3091,N_3818);
or U4570 (N_4570,N_3484,N_3132);
and U4571 (N_4571,N_3270,N_3301);
and U4572 (N_4572,N_3251,N_3896);
and U4573 (N_4573,N_3339,N_3114);
and U4574 (N_4574,N_3828,N_3109);
nor U4575 (N_4575,N_3137,N_3922);
xor U4576 (N_4576,N_3311,N_3450);
nand U4577 (N_4577,N_3608,N_3686);
nand U4578 (N_4578,N_3629,N_3126);
nor U4579 (N_4579,N_3271,N_3903);
and U4580 (N_4580,N_3506,N_3059);
xnor U4581 (N_4581,N_3491,N_3661);
nand U4582 (N_4582,N_3975,N_3225);
and U4583 (N_4583,N_3987,N_3548);
and U4584 (N_4584,N_3607,N_3867);
nand U4585 (N_4585,N_3265,N_3477);
xnor U4586 (N_4586,N_3757,N_3371);
nor U4587 (N_4587,N_3436,N_3511);
and U4588 (N_4588,N_3874,N_3378);
and U4589 (N_4589,N_3917,N_3386);
nor U4590 (N_4590,N_3870,N_3545);
xor U4591 (N_4591,N_3320,N_3089);
nor U4592 (N_4592,N_3282,N_3020);
nand U4593 (N_4593,N_3012,N_3158);
or U4594 (N_4594,N_3138,N_3443);
nor U4595 (N_4595,N_3468,N_3428);
nand U4596 (N_4596,N_3567,N_3814);
or U4597 (N_4597,N_3494,N_3842);
and U4598 (N_4598,N_3414,N_3869);
and U4599 (N_4599,N_3227,N_3520);
xnor U4600 (N_4600,N_3063,N_3860);
nor U4601 (N_4601,N_3771,N_3529);
nand U4602 (N_4602,N_3451,N_3874);
nand U4603 (N_4603,N_3718,N_3912);
xnor U4604 (N_4604,N_3893,N_3328);
or U4605 (N_4605,N_3850,N_3184);
and U4606 (N_4606,N_3632,N_3970);
and U4607 (N_4607,N_3244,N_3934);
xor U4608 (N_4608,N_3774,N_3440);
or U4609 (N_4609,N_3325,N_3256);
xor U4610 (N_4610,N_3958,N_3244);
nor U4611 (N_4611,N_3265,N_3633);
nand U4612 (N_4612,N_3569,N_3217);
or U4613 (N_4613,N_3487,N_3056);
xor U4614 (N_4614,N_3351,N_3479);
xnor U4615 (N_4615,N_3175,N_3696);
xor U4616 (N_4616,N_3549,N_3576);
nand U4617 (N_4617,N_3390,N_3380);
xor U4618 (N_4618,N_3856,N_3366);
nand U4619 (N_4619,N_3179,N_3780);
and U4620 (N_4620,N_3545,N_3061);
nand U4621 (N_4621,N_3812,N_3638);
and U4622 (N_4622,N_3039,N_3908);
or U4623 (N_4623,N_3051,N_3802);
nand U4624 (N_4624,N_3503,N_3336);
nand U4625 (N_4625,N_3039,N_3262);
and U4626 (N_4626,N_3335,N_3189);
and U4627 (N_4627,N_3507,N_3006);
nand U4628 (N_4628,N_3432,N_3287);
and U4629 (N_4629,N_3678,N_3000);
nand U4630 (N_4630,N_3201,N_3722);
or U4631 (N_4631,N_3858,N_3178);
nor U4632 (N_4632,N_3092,N_3309);
nor U4633 (N_4633,N_3848,N_3536);
and U4634 (N_4634,N_3689,N_3747);
and U4635 (N_4635,N_3172,N_3730);
xor U4636 (N_4636,N_3486,N_3713);
or U4637 (N_4637,N_3465,N_3393);
and U4638 (N_4638,N_3148,N_3751);
or U4639 (N_4639,N_3103,N_3655);
nor U4640 (N_4640,N_3963,N_3685);
nor U4641 (N_4641,N_3765,N_3774);
xor U4642 (N_4642,N_3996,N_3583);
or U4643 (N_4643,N_3906,N_3372);
or U4644 (N_4644,N_3965,N_3572);
nor U4645 (N_4645,N_3849,N_3658);
and U4646 (N_4646,N_3079,N_3287);
xnor U4647 (N_4647,N_3940,N_3152);
or U4648 (N_4648,N_3076,N_3290);
nand U4649 (N_4649,N_3120,N_3991);
nor U4650 (N_4650,N_3206,N_3633);
xor U4651 (N_4651,N_3939,N_3028);
or U4652 (N_4652,N_3678,N_3953);
or U4653 (N_4653,N_3637,N_3931);
nor U4654 (N_4654,N_3547,N_3052);
nand U4655 (N_4655,N_3361,N_3768);
or U4656 (N_4656,N_3377,N_3415);
nand U4657 (N_4657,N_3899,N_3632);
and U4658 (N_4658,N_3549,N_3653);
xor U4659 (N_4659,N_3523,N_3435);
or U4660 (N_4660,N_3579,N_3958);
or U4661 (N_4661,N_3742,N_3937);
and U4662 (N_4662,N_3310,N_3453);
and U4663 (N_4663,N_3464,N_3557);
xor U4664 (N_4664,N_3441,N_3580);
and U4665 (N_4665,N_3551,N_3148);
nand U4666 (N_4666,N_3115,N_3358);
and U4667 (N_4667,N_3243,N_3215);
or U4668 (N_4668,N_3405,N_3170);
or U4669 (N_4669,N_3280,N_3053);
nand U4670 (N_4670,N_3684,N_3053);
nor U4671 (N_4671,N_3393,N_3962);
nor U4672 (N_4672,N_3606,N_3484);
nand U4673 (N_4673,N_3168,N_3152);
xor U4674 (N_4674,N_3608,N_3446);
xnor U4675 (N_4675,N_3234,N_3670);
and U4676 (N_4676,N_3501,N_3119);
or U4677 (N_4677,N_3258,N_3803);
xor U4678 (N_4678,N_3166,N_3797);
xor U4679 (N_4679,N_3961,N_3493);
or U4680 (N_4680,N_3782,N_3755);
nand U4681 (N_4681,N_3916,N_3326);
xor U4682 (N_4682,N_3200,N_3571);
and U4683 (N_4683,N_3760,N_3564);
nor U4684 (N_4684,N_3313,N_3630);
or U4685 (N_4685,N_3405,N_3496);
or U4686 (N_4686,N_3829,N_3275);
or U4687 (N_4687,N_3072,N_3741);
nor U4688 (N_4688,N_3896,N_3044);
nand U4689 (N_4689,N_3413,N_3210);
nor U4690 (N_4690,N_3792,N_3189);
or U4691 (N_4691,N_3541,N_3496);
and U4692 (N_4692,N_3697,N_3097);
nand U4693 (N_4693,N_3660,N_3083);
or U4694 (N_4694,N_3756,N_3957);
nand U4695 (N_4695,N_3961,N_3743);
and U4696 (N_4696,N_3385,N_3996);
or U4697 (N_4697,N_3216,N_3170);
xnor U4698 (N_4698,N_3287,N_3388);
nand U4699 (N_4699,N_3725,N_3027);
xor U4700 (N_4700,N_3280,N_3803);
nor U4701 (N_4701,N_3770,N_3986);
and U4702 (N_4702,N_3304,N_3152);
xnor U4703 (N_4703,N_3550,N_3263);
nand U4704 (N_4704,N_3161,N_3174);
nor U4705 (N_4705,N_3499,N_3402);
or U4706 (N_4706,N_3471,N_3787);
xor U4707 (N_4707,N_3367,N_3750);
and U4708 (N_4708,N_3113,N_3734);
xor U4709 (N_4709,N_3006,N_3096);
or U4710 (N_4710,N_3108,N_3681);
nor U4711 (N_4711,N_3391,N_3398);
nor U4712 (N_4712,N_3443,N_3266);
nor U4713 (N_4713,N_3246,N_3105);
nor U4714 (N_4714,N_3679,N_3122);
nor U4715 (N_4715,N_3576,N_3176);
and U4716 (N_4716,N_3419,N_3169);
and U4717 (N_4717,N_3698,N_3241);
and U4718 (N_4718,N_3411,N_3507);
nor U4719 (N_4719,N_3093,N_3258);
xor U4720 (N_4720,N_3604,N_3079);
or U4721 (N_4721,N_3022,N_3809);
and U4722 (N_4722,N_3471,N_3691);
nor U4723 (N_4723,N_3100,N_3894);
and U4724 (N_4724,N_3686,N_3267);
or U4725 (N_4725,N_3712,N_3240);
nand U4726 (N_4726,N_3501,N_3733);
xnor U4727 (N_4727,N_3163,N_3280);
and U4728 (N_4728,N_3135,N_3924);
xor U4729 (N_4729,N_3780,N_3700);
nand U4730 (N_4730,N_3585,N_3935);
nand U4731 (N_4731,N_3325,N_3794);
or U4732 (N_4732,N_3922,N_3458);
nand U4733 (N_4733,N_3630,N_3242);
nor U4734 (N_4734,N_3075,N_3349);
nand U4735 (N_4735,N_3009,N_3022);
or U4736 (N_4736,N_3727,N_3109);
nand U4737 (N_4737,N_3183,N_3987);
or U4738 (N_4738,N_3599,N_3570);
nor U4739 (N_4739,N_3872,N_3502);
nand U4740 (N_4740,N_3707,N_3092);
and U4741 (N_4741,N_3930,N_3419);
or U4742 (N_4742,N_3616,N_3711);
xor U4743 (N_4743,N_3727,N_3414);
or U4744 (N_4744,N_3713,N_3278);
or U4745 (N_4745,N_3976,N_3094);
and U4746 (N_4746,N_3774,N_3697);
nand U4747 (N_4747,N_3776,N_3497);
nor U4748 (N_4748,N_3436,N_3957);
nand U4749 (N_4749,N_3051,N_3284);
and U4750 (N_4750,N_3028,N_3050);
or U4751 (N_4751,N_3591,N_3671);
nor U4752 (N_4752,N_3716,N_3725);
or U4753 (N_4753,N_3808,N_3017);
and U4754 (N_4754,N_3472,N_3459);
nor U4755 (N_4755,N_3830,N_3638);
or U4756 (N_4756,N_3085,N_3180);
or U4757 (N_4757,N_3005,N_3881);
nand U4758 (N_4758,N_3664,N_3076);
and U4759 (N_4759,N_3036,N_3885);
nand U4760 (N_4760,N_3044,N_3627);
nor U4761 (N_4761,N_3936,N_3974);
xnor U4762 (N_4762,N_3687,N_3090);
xor U4763 (N_4763,N_3178,N_3280);
xor U4764 (N_4764,N_3828,N_3263);
xor U4765 (N_4765,N_3812,N_3477);
nor U4766 (N_4766,N_3400,N_3585);
and U4767 (N_4767,N_3465,N_3735);
xor U4768 (N_4768,N_3036,N_3484);
nor U4769 (N_4769,N_3516,N_3613);
xor U4770 (N_4770,N_3942,N_3256);
nand U4771 (N_4771,N_3017,N_3228);
nand U4772 (N_4772,N_3060,N_3016);
xnor U4773 (N_4773,N_3099,N_3522);
nand U4774 (N_4774,N_3603,N_3471);
nand U4775 (N_4775,N_3144,N_3987);
xnor U4776 (N_4776,N_3897,N_3702);
or U4777 (N_4777,N_3822,N_3464);
or U4778 (N_4778,N_3856,N_3111);
or U4779 (N_4779,N_3043,N_3347);
or U4780 (N_4780,N_3468,N_3483);
nand U4781 (N_4781,N_3162,N_3188);
xnor U4782 (N_4782,N_3538,N_3949);
xor U4783 (N_4783,N_3181,N_3926);
nand U4784 (N_4784,N_3643,N_3013);
or U4785 (N_4785,N_3931,N_3429);
nand U4786 (N_4786,N_3305,N_3822);
nor U4787 (N_4787,N_3886,N_3846);
or U4788 (N_4788,N_3807,N_3577);
nand U4789 (N_4789,N_3196,N_3369);
and U4790 (N_4790,N_3831,N_3184);
nor U4791 (N_4791,N_3846,N_3037);
and U4792 (N_4792,N_3243,N_3606);
and U4793 (N_4793,N_3367,N_3659);
nor U4794 (N_4794,N_3074,N_3554);
xor U4795 (N_4795,N_3519,N_3959);
xor U4796 (N_4796,N_3051,N_3437);
nand U4797 (N_4797,N_3742,N_3069);
and U4798 (N_4798,N_3660,N_3525);
nand U4799 (N_4799,N_3526,N_3197);
or U4800 (N_4800,N_3526,N_3182);
or U4801 (N_4801,N_3991,N_3371);
or U4802 (N_4802,N_3207,N_3586);
nand U4803 (N_4803,N_3149,N_3748);
xor U4804 (N_4804,N_3697,N_3742);
xor U4805 (N_4805,N_3491,N_3969);
nand U4806 (N_4806,N_3722,N_3719);
nand U4807 (N_4807,N_3848,N_3349);
or U4808 (N_4808,N_3899,N_3083);
nor U4809 (N_4809,N_3608,N_3896);
xnor U4810 (N_4810,N_3505,N_3482);
and U4811 (N_4811,N_3560,N_3190);
or U4812 (N_4812,N_3355,N_3330);
xnor U4813 (N_4813,N_3303,N_3583);
nor U4814 (N_4814,N_3809,N_3841);
xor U4815 (N_4815,N_3675,N_3540);
nand U4816 (N_4816,N_3624,N_3130);
nand U4817 (N_4817,N_3569,N_3410);
nor U4818 (N_4818,N_3134,N_3769);
xor U4819 (N_4819,N_3193,N_3473);
or U4820 (N_4820,N_3993,N_3783);
nand U4821 (N_4821,N_3142,N_3834);
nor U4822 (N_4822,N_3707,N_3473);
and U4823 (N_4823,N_3567,N_3612);
nand U4824 (N_4824,N_3103,N_3795);
or U4825 (N_4825,N_3906,N_3477);
xnor U4826 (N_4826,N_3189,N_3345);
nand U4827 (N_4827,N_3762,N_3692);
or U4828 (N_4828,N_3267,N_3184);
or U4829 (N_4829,N_3001,N_3088);
xnor U4830 (N_4830,N_3815,N_3678);
nand U4831 (N_4831,N_3958,N_3704);
and U4832 (N_4832,N_3422,N_3557);
and U4833 (N_4833,N_3005,N_3368);
or U4834 (N_4834,N_3568,N_3036);
and U4835 (N_4835,N_3850,N_3122);
xnor U4836 (N_4836,N_3176,N_3666);
nand U4837 (N_4837,N_3217,N_3133);
nor U4838 (N_4838,N_3104,N_3568);
nand U4839 (N_4839,N_3253,N_3026);
nor U4840 (N_4840,N_3564,N_3069);
nand U4841 (N_4841,N_3692,N_3608);
xor U4842 (N_4842,N_3340,N_3371);
nand U4843 (N_4843,N_3337,N_3934);
nand U4844 (N_4844,N_3975,N_3648);
nor U4845 (N_4845,N_3941,N_3747);
or U4846 (N_4846,N_3855,N_3635);
and U4847 (N_4847,N_3851,N_3351);
nor U4848 (N_4848,N_3846,N_3298);
nand U4849 (N_4849,N_3588,N_3963);
xnor U4850 (N_4850,N_3817,N_3717);
or U4851 (N_4851,N_3830,N_3141);
nor U4852 (N_4852,N_3569,N_3775);
nor U4853 (N_4853,N_3276,N_3297);
xnor U4854 (N_4854,N_3465,N_3567);
or U4855 (N_4855,N_3009,N_3790);
and U4856 (N_4856,N_3116,N_3038);
nand U4857 (N_4857,N_3445,N_3681);
and U4858 (N_4858,N_3852,N_3199);
nand U4859 (N_4859,N_3574,N_3893);
xnor U4860 (N_4860,N_3699,N_3258);
or U4861 (N_4861,N_3008,N_3676);
nand U4862 (N_4862,N_3572,N_3544);
or U4863 (N_4863,N_3617,N_3501);
nand U4864 (N_4864,N_3735,N_3498);
and U4865 (N_4865,N_3332,N_3920);
nor U4866 (N_4866,N_3587,N_3130);
nor U4867 (N_4867,N_3104,N_3595);
nand U4868 (N_4868,N_3796,N_3255);
or U4869 (N_4869,N_3140,N_3482);
and U4870 (N_4870,N_3757,N_3029);
nand U4871 (N_4871,N_3000,N_3776);
and U4872 (N_4872,N_3190,N_3708);
nor U4873 (N_4873,N_3436,N_3698);
nor U4874 (N_4874,N_3337,N_3837);
nor U4875 (N_4875,N_3641,N_3024);
and U4876 (N_4876,N_3075,N_3660);
and U4877 (N_4877,N_3825,N_3063);
or U4878 (N_4878,N_3648,N_3614);
nor U4879 (N_4879,N_3285,N_3011);
nor U4880 (N_4880,N_3759,N_3804);
or U4881 (N_4881,N_3919,N_3050);
or U4882 (N_4882,N_3757,N_3388);
or U4883 (N_4883,N_3589,N_3994);
nand U4884 (N_4884,N_3918,N_3650);
or U4885 (N_4885,N_3480,N_3367);
or U4886 (N_4886,N_3937,N_3227);
and U4887 (N_4887,N_3745,N_3480);
nand U4888 (N_4888,N_3794,N_3780);
nand U4889 (N_4889,N_3994,N_3811);
nand U4890 (N_4890,N_3291,N_3477);
nand U4891 (N_4891,N_3604,N_3941);
nand U4892 (N_4892,N_3825,N_3369);
nand U4893 (N_4893,N_3074,N_3957);
or U4894 (N_4894,N_3020,N_3747);
nand U4895 (N_4895,N_3693,N_3992);
xnor U4896 (N_4896,N_3711,N_3286);
xor U4897 (N_4897,N_3141,N_3160);
or U4898 (N_4898,N_3359,N_3838);
xor U4899 (N_4899,N_3059,N_3296);
nor U4900 (N_4900,N_3213,N_3290);
nor U4901 (N_4901,N_3592,N_3708);
nand U4902 (N_4902,N_3984,N_3800);
and U4903 (N_4903,N_3446,N_3002);
nor U4904 (N_4904,N_3867,N_3013);
xor U4905 (N_4905,N_3032,N_3115);
or U4906 (N_4906,N_3887,N_3259);
xor U4907 (N_4907,N_3637,N_3644);
nor U4908 (N_4908,N_3218,N_3769);
xor U4909 (N_4909,N_3427,N_3334);
or U4910 (N_4910,N_3197,N_3368);
or U4911 (N_4911,N_3830,N_3092);
xor U4912 (N_4912,N_3736,N_3804);
or U4913 (N_4913,N_3657,N_3997);
xor U4914 (N_4914,N_3912,N_3898);
and U4915 (N_4915,N_3077,N_3127);
or U4916 (N_4916,N_3782,N_3941);
and U4917 (N_4917,N_3715,N_3496);
and U4918 (N_4918,N_3102,N_3545);
xnor U4919 (N_4919,N_3363,N_3009);
nor U4920 (N_4920,N_3410,N_3446);
and U4921 (N_4921,N_3750,N_3010);
nand U4922 (N_4922,N_3112,N_3007);
xnor U4923 (N_4923,N_3318,N_3810);
nand U4924 (N_4924,N_3376,N_3642);
and U4925 (N_4925,N_3155,N_3562);
or U4926 (N_4926,N_3541,N_3088);
or U4927 (N_4927,N_3768,N_3450);
nor U4928 (N_4928,N_3174,N_3589);
nor U4929 (N_4929,N_3098,N_3184);
nand U4930 (N_4930,N_3001,N_3698);
xnor U4931 (N_4931,N_3507,N_3128);
nand U4932 (N_4932,N_3824,N_3627);
and U4933 (N_4933,N_3138,N_3155);
xnor U4934 (N_4934,N_3838,N_3678);
or U4935 (N_4935,N_3143,N_3034);
xnor U4936 (N_4936,N_3590,N_3311);
xnor U4937 (N_4937,N_3098,N_3725);
and U4938 (N_4938,N_3947,N_3622);
nand U4939 (N_4939,N_3207,N_3021);
or U4940 (N_4940,N_3431,N_3259);
xor U4941 (N_4941,N_3205,N_3648);
and U4942 (N_4942,N_3122,N_3714);
xor U4943 (N_4943,N_3977,N_3018);
nand U4944 (N_4944,N_3798,N_3749);
and U4945 (N_4945,N_3921,N_3811);
nand U4946 (N_4946,N_3752,N_3817);
xor U4947 (N_4947,N_3694,N_3385);
or U4948 (N_4948,N_3262,N_3631);
nor U4949 (N_4949,N_3775,N_3373);
xor U4950 (N_4950,N_3769,N_3266);
nand U4951 (N_4951,N_3240,N_3258);
nor U4952 (N_4952,N_3286,N_3911);
and U4953 (N_4953,N_3121,N_3128);
or U4954 (N_4954,N_3796,N_3745);
or U4955 (N_4955,N_3504,N_3812);
xor U4956 (N_4956,N_3576,N_3253);
nor U4957 (N_4957,N_3171,N_3819);
nor U4958 (N_4958,N_3477,N_3339);
or U4959 (N_4959,N_3136,N_3842);
and U4960 (N_4960,N_3469,N_3252);
nor U4961 (N_4961,N_3856,N_3511);
or U4962 (N_4962,N_3467,N_3602);
and U4963 (N_4963,N_3640,N_3430);
nor U4964 (N_4964,N_3159,N_3917);
nand U4965 (N_4965,N_3968,N_3949);
nor U4966 (N_4966,N_3348,N_3331);
xnor U4967 (N_4967,N_3356,N_3558);
xnor U4968 (N_4968,N_3824,N_3768);
nand U4969 (N_4969,N_3372,N_3227);
nand U4970 (N_4970,N_3248,N_3136);
and U4971 (N_4971,N_3447,N_3142);
and U4972 (N_4972,N_3149,N_3721);
and U4973 (N_4973,N_3665,N_3724);
or U4974 (N_4974,N_3097,N_3201);
or U4975 (N_4975,N_3502,N_3385);
nor U4976 (N_4976,N_3478,N_3484);
or U4977 (N_4977,N_3580,N_3596);
nand U4978 (N_4978,N_3668,N_3908);
or U4979 (N_4979,N_3167,N_3715);
or U4980 (N_4980,N_3725,N_3114);
nor U4981 (N_4981,N_3835,N_3808);
nand U4982 (N_4982,N_3320,N_3355);
and U4983 (N_4983,N_3525,N_3264);
nor U4984 (N_4984,N_3773,N_3502);
xor U4985 (N_4985,N_3904,N_3219);
nand U4986 (N_4986,N_3004,N_3190);
nor U4987 (N_4987,N_3883,N_3174);
nor U4988 (N_4988,N_3866,N_3433);
xnor U4989 (N_4989,N_3329,N_3586);
and U4990 (N_4990,N_3447,N_3143);
nor U4991 (N_4991,N_3607,N_3427);
xor U4992 (N_4992,N_3735,N_3485);
xor U4993 (N_4993,N_3202,N_3208);
or U4994 (N_4994,N_3219,N_3368);
xor U4995 (N_4995,N_3320,N_3874);
xnor U4996 (N_4996,N_3458,N_3938);
nand U4997 (N_4997,N_3235,N_3294);
xor U4998 (N_4998,N_3044,N_3619);
and U4999 (N_4999,N_3825,N_3387);
and U5000 (N_5000,N_4861,N_4667);
and U5001 (N_5001,N_4398,N_4289);
xor U5002 (N_5002,N_4178,N_4939);
nand U5003 (N_5003,N_4181,N_4032);
and U5004 (N_5004,N_4639,N_4144);
or U5005 (N_5005,N_4275,N_4095);
nor U5006 (N_5006,N_4969,N_4125);
xor U5007 (N_5007,N_4572,N_4294);
nand U5008 (N_5008,N_4299,N_4613);
nor U5009 (N_5009,N_4386,N_4431);
nor U5010 (N_5010,N_4111,N_4618);
nand U5011 (N_5011,N_4088,N_4955);
and U5012 (N_5012,N_4137,N_4217);
or U5013 (N_5013,N_4641,N_4376);
and U5014 (N_5014,N_4688,N_4664);
nor U5015 (N_5015,N_4026,N_4717);
or U5016 (N_5016,N_4744,N_4107);
and U5017 (N_5017,N_4435,N_4280);
xnor U5018 (N_5018,N_4771,N_4420);
nand U5019 (N_5019,N_4225,N_4127);
or U5020 (N_5020,N_4701,N_4138);
xor U5021 (N_5021,N_4951,N_4441);
or U5022 (N_5022,N_4516,N_4789);
nand U5023 (N_5023,N_4073,N_4965);
nor U5024 (N_5024,N_4953,N_4364);
xor U5025 (N_5025,N_4469,N_4240);
and U5026 (N_5026,N_4703,N_4592);
nor U5027 (N_5027,N_4086,N_4967);
and U5028 (N_5028,N_4675,N_4005);
nor U5029 (N_5029,N_4200,N_4436);
nand U5030 (N_5030,N_4952,N_4040);
nor U5031 (N_5031,N_4583,N_4543);
and U5032 (N_5032,N_4707,N_4503);
or U5033 (N_5033,N_4341,N_4253);
nor U5034 (N_5034,N_4860,N_4630);
nand U5035 (N_5035,N_4783,N_4266);
nor U5036 (N_5036,N_4896,N_4576);
or U5037 (N_5037,N_4083,N_4637);
or U5038 (N_5038,N_4120,N_4906);
xor U5039 (N_5039,N_4742,N_4692);
nand U5040 (N_5040,N_4291,N_4843);
nor U5041 (N_5041,N_4395,N_4957);
nand U5042 (N_5042,N_4207,N_4594);
nor U5043 (N_5043,N_4540,N_4242);
xnor U5044 (N_5044,N_4980,N_4855);
xor U5045 (N_5045,N_4549,N_4362);
and U5046 (N_5046,N_4907,N_4854);
and U5047 (N_5047,N_4923,N_4008);
nor U5048 (N_5048,N_4187,N_4356);
nand U5049 (N_5049,N_4748,N_4683);
xnor U5050 (N_5050,N_4129,N_4841);
nand U5051 (N_5051,N_4171,N_4239);
xnor U5052 (N_5052,N_4929,N_4329);
nor U5053 (N_5053,N_4821,N_4279);
xnor U5054 (N_5054,N_4625,N_4072);
nor U5055 (N_5055,N_4784,N_4098);
or U5056 (N_5056,N_4085,N_4350);
nor U5057 (N_5057,N_4782,N_4468);
xnor U5058 (N_5058,N_4193,N_4296);
or U5059 (N_5059,N_4943,N_4589);
nor U5060 (N_5060,N_4714,N_4614);
and U5061 (N_5061,N_4002,N_4657);
nand U5062 (N_5062,N_4882,N_4970);
and U5063 (N_5063,N_4756,N_4825);
or U5064 (N_5064,N_4726,N_4766);
nor U5065 (N_5065,N_4495,N_4197);
nand U5066 (N_5066,N_4258,N_4670);
xnor U5067 (N_5067,N_4814,N_4808);
or U5068 (N_5068,N_4824,N_4229);
and U5069 (N_5069,N_4968,N_4273);
nor U5070 (N_5070,N_4787,N_4303);
xor U5071 (N_5071,N_4373,N_4548);
xor U5072 (N_5072,N_4151,N_4711);
and U5073 (N_5073,N_4477,N_4852);
nand U5074 (N_5074,N_4284,N_4570);
nor U5075 (N_5075,N_4182,N_4772);
nand U5076 (N_5076,N_4868,N_4321);
or U5077 (N_5077,N_4505,N_4145);
and U5078 (N_5078,N_4326,N_4932);
xor U5079 (N_5079,N_4461,N_4451);
and U5080 (N_5080,N_4765,N_4716);
xnor U5081 (N_5081,N_4898,N_4050);
nor U5082 (N_5082,N_4631,N_4224);
nand U5083 (N_5083,N_4926,N_4562);
xor U5084 (N_5084,N_4757,N_4745);
and U5085 (N_5085,N_4316,N_4698);
nor U5086 (N_5086,N_4066,N_4177);
or U5087 (N_5087,N_4330,N_4908);
xor U5088 (N_5088,N_4723,N_4816);
nand U5089 (N_5089,N_4586,N_4312);
nand U5090 (N_5090,N_4881,N_4558);
and U5091 (N_5091,N_4663,N_4801);
nor U5092 (N_5092,N_4743,N_4672);
and U5093 (N_5093,N_4322,N_4930);
xnor U5094 (N_5094,N_4009,N_4813);
nor U5095 (N_5095,N_4013,N_4916);
xnor U5096 (N_5096,N_4874,N_4278);
or U5097 (N_5097,N_4449,N_4447);
nor U5098 (N_5098,N_4498,N_4180);
nor U5099 (N_5099,N_4654,N_4243);
nor U5100 (N_5100,N_4523,N_4949);
nor U5101 (N_5101,N_4262,N_4453);
xnor U5102 (N_5102,N_4118,N_4038);
nor U5103 (N_5103,N_4897,N_4946);
or U5104 (N_5104,N_4295,N_4646);
nor U5105 (N_5105,N_4252,N_4097);
nor U5106 (N_5106,N_4656,N_4371);
xnor U5107 (N_5107,N_4018,N_4638);
xnor U5108 (N_5108,N_4864,N_4610);
and U5109 (N_5109,N_4261,N_4049);
and U5110 (N_5110,N_4658,N_4560);
nor U5111 (N_5111,N_4859,N_4578);
and U5112 (N_5112,N_4135,N_4622);
and U5113 (N_5113,N_4042,N_4057);
nand U5114 (N_5114,N_4828,N_4101);
nor U5115 (N_5115,N_4623,N_4839);
nor U5116 (N_5116,N_4858,N_4994);
and U5117 (N_5117,N_4173,N_4478);
nor U5118 (N_5118,N_4154,N_4763);
or U5119 (N_5119,N_4747,N_4609);
nand U5120 (N_5120,N_4941,N_4835);
and U5121 (N_5121,N_4168,N_4331);
xnor U5122 (N_5122,N_4434,N_4297);
or U5123 (N_5123,N_4140,N_4323);
nand U5124 (N_5124,N_4082,N_4532);
nor U5125 (N_5125,N_4978,N_4515);
and U5126 (N_5126,N_4687,N_4408);
nand U5127 (N_5127,N_4818,N_4301);
xnor U5128 (N_5128,N_4444,N_4497);
or U5129 (N_5129,N_4029,N_4564);
nor U5130 (N_5130,N_4223,N_4734);
and U5131 (N_5131,N_4494,N_4931);
or U5132 (N_5132,N_4377,N_4267);
nor U5133 (N_5133,N_4944,N_4936);
and U5134 (N_5134,N_4000,N_4666);
nand U5135 (N_5135,N_4191,N_4851);
or U5136 (N_5136,N_4774,N_4448);
nand U5137 (N_5137,N_4838,N_4606);
and U5138 (N_5138,N_4693,N_4091);
and U5139 (N_5139,N_4110,N_4423);
xor U5140 (N_5140,N_4710,N_4319);
nand U5141 (N_5141,N_4739,N_4112);
or U5142 (N_5142,N_4749,N_4422);
nor U5143 (N_5143,N_4697,N_4651);
nand U5144 (N_5144,N_4529,N_4293);
nand U5145 (N_5145,N_4017,N_4192);
xnor U5146 (N_5146,N_4195,N_4090);
nand U5147 (N_5147,N_4327,N_4149);
nor U5148 (N_5148,N_4387,N_4343);
nand U5149 (N_5149,N_4361,N_4715);
and U5150 (N_5150,N_4642,N_4348);
nand U5151 (N_5151,N_4349,N_4254);
or U5152 (N_5152,N_4249,N_4102);
or U5153 (N_5153,N_4450,N_4521);
nor U5154 (N_5154,N_4643,N_4561);
or U5155 (N_5155,N_4012,N_4159);
nand U5156 (N_5156,N_4826,N_4781);
xnor U5157 (N_5157,N_4611,N_4413);
xor U5158 (N_5158,N_4831,N_4034);
xnor U5159 (N_5159,N_4372,N_4446);
xor U5160 (N_5160,N_4231,N_4893);
nor U5161 (N_5161,N_4652,N_4134);
or U5162 (N_5162,N_4769,N_4731);
nor U5163 (N_5163,N_4028,N_4593);
and U5164 (N_5164,N_4876,N_4704);
xnor U5165 (N_5165,N_4557,N_4313);
nor U5166 (N_5166,N_4466,N_4309);
xor U5167 (N_5167,N_4222,N_4728);
xor U5168 (N_5168,N_4496,N_4945);
xor U5169 (N_5169,N_4452,N_4023);
and U5170 (N_5170,N_4619,N_4481);
xor U5171 (N_5171,N_4136,N_4604);
nand U5172 (N_5172,N_4179,N_4513);
and U5173 (N_5173,N_4388,N_4210);
xor U5174 (N_5174,N_4298,N_4850);
xnor U5175 (N_5175,N_4036,N_4153);
and U5176 (N_5176,N_4918,N_4456);
nand U5177 (N_5177,N_4509,N_4369);
or U5178 (N_5178,N_4215,N_4119);
or U5179 (N_5179,N_4158,N_4359);
xnor U5180 (N_5180,N_4848,N_4829);
xor U5181 (N_5181,N_4352,N_4577);
nor U5182 (N_5182,N_4588,N_4964);
or U5183 (N_5183,N_4706,N_4832);
nand U5184 (N_5184,N_4199,N_4580);
nor U5185 (N_5185,N_4347,N_4411);
nand U5186 (N_5186,N_4753,N_4281);
or U5187 (N_5187,N_4519,N_4437);
xor U5188 (N_5188,N_4624,N_4574);
nor U5189 (N_5189,N_4919,N_4338);
nor U5190 (N_5190,N_4800,N_4694);
or U5191 (N_5191,N_4535,N_4581);
nand U5192 (N_5192,N_4194,N_4847);
and U5193 (N_5193,N_4659,N_4233);
xor U5194 (N_5194,N_4074,N_4522);
nor U5195 (N_5195,N_4476,N_4428);
nor U5196 (N_5196,N_4671,N_4457);
xnor U5197 (N_5197,N_4845,N_4232);
or U5198 (N_5198,N_4130,N_4269);
nor U5199 (N_5199,N_4092,N_4070);
or U5200 (N_5200,N_4184,N_4089);
or U5201 (N_5201,N_4003,N_4205);
nor U5202 (N_5202,N_4512,N_4069);
nand U5203 (N_5203,N_4628,N_4212);
or U5204 (N_5204,N_4811,N_4024);
or U5205 (N_5205,N_4492,N_4989);
nor U5206 (N_5206,N_4649,N_4152);
nand U5207 (N_5207,N_4573,N_4375);
nor U5208 (N_5208,N_4527,N_4320);
nand U5209 (N_5209,N_4702,N_4315);
nand U5210 (N_5210,N_4912,N_4162);
nand U5211 (N_5211,N_4966,N_4059);
nand U5212 (N_5212,N_4141,N_4484);
xnor U5213 (N_5213,N_4425,N_4133);
nand U5214 (N_5214,N_4963,N_4934);
or U5215 (N_5215,N_4567,N_4201);
and U5216 (N_5216,N_4385,N_4877);
xor U5217 (N_5217,N_4442,N_4645);
nand U5218 (N_5218,N_4406,N_4142);
nor U5219 (N_5219,N_4064,N_4004);
xor U5220 (N_5220,N_4598,N_4514);
xnor U5221 (N_5221,N_4462,N_4394);
or U5222 (N_5222,N_4555,N_4238);
nand U5223 (N_5223,N_4014,N_4595);
and U5224 (N_5224,N_4459,N_4307);
nor U5225 (N_5225,N_4950,N_4530);
nand U5226 (N_5226,N_4937,N_4900);
nand U5227 (N_5227,N_4685,N_4202);
or U5228 (N_5228,N_4292,N_4430);
nor U5229 (N_5229,N_4081,N_4791);
xor U5230 (N_5230,N_4536,N_4116);
nor U5231 (N_5231,N_4956,N_4695);
nor U5232 (N_5232,N_4650,N_4662);
nor U5233 (N_5233,N_4048,N_4684);
nor U5234 (N_5234,N_4977,N_4909);
and U5235 (N_5235,N_4396,N_4817);
or U5236 (N_5236,N_4888,N_4998);
nor U5237 (N_5237,N_4402,N_4500);
xor U5238 (N_5238,N_4105,N_4054);
xor U5239 (N_5239,N_4043,N_4827);
and U5240 (N_5240,N_4164,N_4020);
and U5241 (N_5241,N_4318,N_4972);
or U5242 (N_5242,N_4735,N_4354);
nor U5243 (N_5243,N_4910,N_4960);
or U5244 (N_5244,N_4464,N_4308);
nand U5245 (N_5245,N_4221,N_4542);
nand U5246 (N_5246,N_4366,N_4230);
and U5247 (N_5247,N_4661,N_4996);
and U5248 (N_5248,N_4482,N_4310);
and U5249 (N_5249,N_4099,N_4304);
xor U5250 (N_5250,N_4467,N_4914);
nand U5251 (N_5251,N_4443,N_4669);
xnor U5252 (N_5252,N_4220,N_4725);
and U5253 (N_5253,N_4336,N_4283);
nand U5254 (N_5254,N_4006,N_4021);
nand U5255 (N_5255,N_4235,N_4732);
xor U5256 (N_5256,N_4504,N_4682);
nand U5257 (N_5257,N_4999,N_4306);
and U5258 (N_5258,N_4520,N_4027);
or U5259 (N_5259,N_4156,N_4426);
nand U5260 (N_5260,N_4849,N_4344);
nor U5261 (N_5261,N_4087,N_4337);
xnor U5262 (N_5262,N_4227,N_4837);
xor U5263 (N_5263,N_4615,N_4078);
or U5264 (N_5264,N_4880,N_4668);
nand U5265 (N_5265,N_4730,N_4044);
and U5266 (N_5266,N_4871,N_4165);
nand U5267 (N_5267,N_4626,N_4899);
nor U5268 (N_5268,N_4046,N_4737);
and U5269 (N_5269,N_4062,N_4750);
nor U5270 (N_5270,N_4256,N_4475);
or U5271 (N_5271,N_4103,N_4597);
or U5272 (N_5272,N_4740,N_4196);
nand U5273 (N_5273,N_4792,N_4139);
or U5274 (N_5274,N_4804,N_4143);
nor U5275 (N_5275,N_4209,N_4264);
nand U5276 (N_5276,N_4265,N_4245);
xnor U5277 (N_5277,N_4257,N_4905);
nor U5278 (N_5278,N_4853,N_4131);
xnor U5279 (N_5279,N_4517,N_4775);
nor U5280 (N_5280,N_4241,N_4547);
or U5281 (N_5281,N_4384,N_4833);
nand U5282 (N_5282,N_4213,N_4403);
and U5283 (N_5283,N_4351,N_4401);
nor U5284 (N_5284,N_4857,N_4988);
xor U5285 (N_5285,N_4079,N_4001);
nand U5286 (N_5286,N_4015,N_4440);
nor U5287 (N_5287,N_4890,N_4166);
nor U5288 (N_5288,N_4114,N_4836);
nor U5289 (N_5289,N_4339,N_4188);
xor U5290 (N_5290,N_4115,N_4629);
nor U5291 (N_5291,N_4758,N_4128);
or U5292 (N_5292,N_4607,N_4155);
and U5293 (N_5293,N_4603,N_4633);
and U5294 (N_5294,N_4709,N_4991);
nor U5295 (N_5295,N_4493,N_4404);
and U5296 (N_5296,N_4342,N_4473);
xor U5297 (N_5297,N_4379,N_4620);
nor U5298 (N_5298,N_4236,N_4370);
nor U5299 (N_5299,N_4104,N_4391);
and U5300 (N_5300,N_4903,N_4096);
and U5301 (N_5301,N_4713,N_4802);
xnor U5302 (N_5302,N_4454,N_4681);
and U5303 (N_5303,N_4035,N_4077);
nor U5304 (N_5304,N_4997,N_4305);
and U5305 (N_5305,N_4634,N_4290);
or U5306 (N_5306,N_4708,N_4365);
nand U5307 (N_5307,N_4767,N_4485);
nand U5308 (N_5308,N_4429,N_4925);
nand U5309 (N_5309,N_4834,N_4084);
xnor U5310 (N_5310,N_4510,N_4263);
xor U5311 (N_5311,N_4334,N_4234);
and U5312 (N_5312,N_4992,N_4807);
and U5313 (N_5313,N_4830,N_4080);
or U5314 (N_5314,N_4106,N_4647);
or U5315 (N_5315,N_4754,N_4602);
and U5316 (N_5316,N_4762,N_4979);
nor U5317 (N_5317,N_4248,N_4314);
nor U5318 (N_5318,N_4959,N_4690);
and U5319 (N_5319,N_4472,N_4585);
and U5320 (N_5320,N_4559,N_4973);
and U5321 (N_5321,N_4729,N_4790);
xor U5322 (N_5322,N_4842,N_4333);
and U5323 (N_5323,N_4268,N_4427);
or U5324 (N_5324,N_4823,N_4058);
or U5325 (N_5325,N_4938,N_4544);
nor U5326 (N_5326,N_4806,N_4974);
or U5327 (N_5327,N_4617,N_4525);
nor U5328 (N_5328,N_4552,N_4653);
and U5329 (N_5329,N_4768,N_4325);
or U5330 (N_5330,N_4226,N_4550);
or U5331 (N_5331,N_4405,N_4590);
nor U5332 (N_5332,N_4219,N_4150);
and U5333 (N_5333,N_4380,N_4863);
nand U5334 (N_5334,N_4546,N_4174);
xor U5335 (N_5335,N_4389,N_4499);
nor U5336 (N_5336,N_4124,N_4990);
and U5337 (N_5337,N_4502,N_4534);
nand U5338 (N_5338,N_4636,N_4582);
nor U5339 (N_5339,N_4324,N_4100);
xnor U5340 (N_5340,N_4678,N_4797);
nor U5341 (N_5341,N_4700,N_4186);
or U5342 (N_5342,N_4019,N_4538);
nor U5343 (N_5343,N_4198,N_4374);
or U5344 (N_5344,N_4883,N_4755);
and U5345 (N_5345,N_4752,N_4302);
nor U5346 (N_5346,N_4873,N_4355);
xnor U5347 (N_5347,N_4568,N_4862);
or U5348 (N_5348,N_4031,N_4410);
nor U5349 (N_5349,N_4528,N_4600);
nand U5350 (N_5350,N_4785,N_4846);
and U5351 (N_5351,N_4720,N_4438);
and U5352 (N_5352,N_4724,N_4208);
or U5353 (N_5353,N_4524,N_4587);
xnor U5354 (N_5354,N_4840,N_4122);
and U5355 (N_5355,N_4689,N_4185);
nor U5356 (N_5356,N_4237,N_4067);
xor U5357 (N_5357,N_4927,N_4526);
xor U5358 (N_5358,N_4346,N_4676);
nor U5359 (N_5359,N_4093,N_4971);
nor U5360 (N_5360,N_4416,N_4820);
nand U5361 (N_5361,N_4803,N_4612);
nor U5362 (N_5362,N_4727,N_4433);
xor U5363 (N_5363,N_4541,N_4691);
and U5364 (N_5364,N_4211,N_4889);
nand U5365 (N_5365,N_4479,N_4866);
or U5366 (N_5366,N_4065,N_4465);
xor U5367 (N_5367,N_4363,N_4400);
nor U5368 (N_5368,N_4677,N_4798);
nand U5369 (N_5369,N_4983,N_4418);
xor U5370 (N_5370,N_4511,N_4928);
xor U5371 (N_5371,N_4640,N_4439);
nand U5372 (N_5372,N_4246,N_4037);
xor U5373 (N_5373,N_4063,N_4718);
xnor U5374 (N_5374,N_4381,N_4872);
xor U5375 (N_5375,N_4160,N_4022);
nor U5376 (N_5376,N_4986,N_4958);
xor U5377 (N_5377,N_4189,N_4169);
nand U5378 (N_5378,N_4533,N_4746);
nor U5379 (N_5379,N_4076,N_4601);
or U5380 (N_5380,N_4770,N_4660);
xor U5381 (N_5381,N_4865,N_4940);
nand U5382 (N_5382,N_4474,N_4214);
nand U5383 (N_5383,N_4608,N_4407);
or U5384 (N_5384,N_4271,N_4875);
and U5385 (N_5385,N_4961,N_4382);
xor U5386 (N_5386,N_4025,N_4556);
xnor U5387 (N_5387,N_4247,N_4760);
xnor U5388 (N_5388,N_4895,N_4679);
xor U5389 (N_5389,N_4490,N_4360);
nor U5390 (N_5390,N_4167,N_4170);
nand U5391 (N_5391,N_4007,N_4867);
nor U5392 (N_5392,N_4751,N_4869);
nand U5393 (N_5393,N_4415,N_4132);
xnor U5394 (N_5394,N_4810,N_4705);
or U5395 (N_5395,N_4335,N_4421);
and U5396 (N_5396,N_4984,N_4052);
nor U5397 (N_5397,N_4470,N_4795);
nand U5398 (N_5398,N_4982,N_4759);
xor U5399 (N_5399,N_4993,N_4489);
nor U5400 (N_5400,N_4913,N_4176);
nor U5401 (N_5401,N_4332,N_4041);
nand U5402 (N_5402,N_4733,N_4175);
nor U5403 (N_5403,N_4412,N_4796);
or U5404 (N_5404,N_4244,N_4856);
nor U5405 (N_5405,N_4537,N_4591);
nand U5406 (N_5406,N_4566,N_4885);
nor U5407 (N_5407,N_4056,N_4061);
xnor U5408 (N_5408,N_4203,N_4047);
xnor U5409 (N_5409,N_4995,N_4935);
nor U5410 (N_5410,N_4545,N_4892);
xnor U5411 (N_5411,N_4367,N_4471);
xor U5412 (N_5412,N_4571,N_4539);
xnor U5413 (N_5413,N_4575,N_4358);
nand U5414 (N_5414,N_4648,N_4117);
nand U5415 (N_5415,N_4030,N_4764);
and U5416 (N_5416,N_4353,N_4146);
nand U5417 (N_5417,N_4383,N_4644);
nand U5418 (N_5418,N_4901,N_4460);
nand U5419 (N_5419,N_4917,N_4445);
nand U5420 (N_5420,N_4799,N_4719);
and U5421 (N_5421,N_4458,N_4696);
or U5422 (N_5422,N_4419,N_4599);
xor U5423 (N_5423,N_4033,N_4920);
nand U5424 (N_5424,N_4933,N_4397);
and U5425 (N_5425,N_4819,N_4699);
and U5426 (N_5426,N_4844,N_4879);
xor U5427 (N_5427,N_4812,N_4393);
xor U5428 (N_5428,N_4870,N_4463);
xor U5429 (N_5429,N_4409,N_4531);
nand U5430 (N_5430,N_4894,N_4285);
or U5431 (N_5431,N_4776,N_4068);
nor U5432 (N_5432,N_4311,N_4922);
or U5433 (N_5433,N_4216,N_4147);
nand U5434 (N_5434,N_4317,N_4904);
and U5435 (N_5435,N_4204,N_4738);
xnor U5436 (N_5436,N_4328,N_4163);
and U5437 (N_5437,N_4911,N_4260);
and U5438 (N_5438,N_4786,N_4891);
nand U5439 (N_5439,N_4553,N_4399);
xor U5440 (N_5440,N_4282,N_4815);
and U5441 (N_5441,N_4686,N_4722);
or U5442 (N_5442,N_4286,N_4094);
or U5443 (N_5443,N_4596,N_4228);
nor U5444 (N_5444,N_4218,N_4761);
nand U5445 (N_5445,N_4778,N_4368);
nor U5446 (N_5446,N_4055,N_4113);
nor U5447 (N_5447,N_4390,N_4071);
nand U5448 (N_5448,N_4424,N_4975);
or U5449 (N_5449,N_4712,N_4345);
xnor U5450 (N_5450,N_4183,N_4010);
nor U5451 (N_5451,N_4157,N_4501);
nor U5452 (N_5452,N_4161,N_4277);
and U5453 (N_5453,N_4584,N_4655);
xnor U5454 (N_5454,N_4665,N_4518);
nand U5455 (N_5455,N_4491,N_4051);
and U5456 (N_5456,N_4190,N_4414);
and U5457 (N_5457,N_4884,N_4123);
or U5458 (N_5458,N_4616,N_4579);
and U5459 (N_5459,N_4886,N_4773);
nand U5460 (N_5460,N_4809,N_4109);
xor U5461 (N_5461,N_4680,N_4016);
or U5462 (N_5462,N_4270,N_4942);
xnor U5463 (N_5463,N_4822,N_4378);
nor U5464 (N_5464,N_4793,N_4075);
xnor U5465 (N_5465,N_4563,N_4508);
or U5466 (N_5466,N_4794,N_4487);
nor U5467 (N_5467,N_4011,N_4887);
nor U5468 (N_5468,N_4551,N_4621);
nand U5469 (N_5469,N_4987,N_4981);
nor U5470 (N_5470,N_4148,N_4172);
nand U5471 (N_5471,N_4741,N_4053);
xnor U5472 (N_5472,N_4921,N_4962);
and U5473 (N_5473,N_4483,N_4251);
and U5474 (N_5474,N_4288,N_4357);
or U5475 (N_5475,N_4736,N_4985);
nand U5476 (N_5476,N_4780,N_4569);
xnor U5477 (N_5477,N_4915,N_4250);
xnor U5478 (N_5478,N_4287,N_4506);
nor U5479 (N_5479,N_4272,N_4432);
nand U5480 (N_5480,N_4340,N_4627);
or U5481 (N_5481,N_4674,N_4948);
nor U5482 (N_5482,N_4635,N_4788);
nor U5483 (N_5483,N_4206,N_4417);
nor U5484 (N_5484,N_4060,N_4605);
and U5485 (N_5485,N_4976,N_4108);
nor U5486 (N_5486,N_4565,N_4480);
nor U5487 (N_5487,N_4039,N_4507);
or U5488 (N_5488,N_4274,N_4259);
nor U5489 (N_5489,N_4721,N_4779);
nand U5490 (N_5490,N_4126,N_4878);
nor U5491 (N_5491,N_4777,N_4632);
or U5492 (N_5492,N_4455,N_4805);
nand U5493 (N_5493,N_4300,N_4673);
nor U5494 (N_5494,N_4947,N_4392);
nor U5495 (N_5495,N_4554,N_4954);
nor U5496 (N_5496,N_4902,N_4924);
or U5497 (N_5497,N_4121,N_4486);
or U5498 (N_5498,N_4276,N_4255);
and U5499 (N_5499,N_4488,N_4045);
and U5500 (N_5500,N_4718,N_4311);
xnor U5501 (N_5501,N_4793,N_4812);
nand U5502 (N_5502,N_4697,N_4593);
or U5503 (N_5503,N_4156,N_4417);
or U5504 (N_5504,N_4159,N_4891);
or U5505 (N_5505,N_4411,N_4093);
or U5506 (N_5506,N_4146,N_4857);
xor U5507 (N_5507,N_4872,N_4888);
nand U5508 (N_5508,N_4098,N_4179);
xnor U5509 (N_5509,N_4608,N_4914);
and U5510 (N_5510,N_4195,N_4489);
and U5511 (N_5511,N_4337,N_4728);
nor U5512 (N_5512,N_4215,N_4434);
and U5513 (N_5513,N_4155,N_4114);
and U5514 (N_5514,N_4523,N_4027);
and U5515 (N_5515,N_4057,N_4562);
or U5516 (N_5516,N_4813,N_4149);
xor U5517 (N_5517,N_4131,N_4573);
nor U5518 (N_5518,N_4518,N_4970);
nand U5519 (N_5519,N_4417,N_4923);
and U5520 (N_5520,N_4439,N_4537);
nor U5521 (N_5521,N_4139,N_4842);
xnor U5522 (N_5522,N_4132,N_4109);
and U5523 (N_5523,N_4781,N_4570);
and U5524 (N_5524,N_4579,N_4452);
and U5525 (N_5525,N_4514,N_4495);
nor U5526 (N_5526,N_4688,N_4824);
xor U5527 (N_5527,N_4988,N_4682);
or U5528 (N_5528,N_4642,N_4458);
xnor U5529 (N_5529,N_4304,N_4014);
nor U5530 (N_5530,N_4501,N_4524);
nand U5531 (N_5531,N_4502,N_4988);
and U5532 (N_5532,N_4894,N_4123);
nor U5533 (N_5533,N_4088,N_4412);
nor U5534 (N_5534,N_4760,N_4552);
xnor U5535 (N_5535,N_4038,N_4732);
nand U5536 (N_5536,N_4048,N_4289);
or U5537 (N_5537,N_4267,N_4093);
xnor U5538 (N_5538,N_4528,N_4962);
or U5539 (N_5539,N_4267,N_4567);
nor U5540 (N_5540,N_4909,N_4040);
nand U5541 (N_5541,N_4291,N_4965);
xnor U5542 (N_5542,N_4327,N_4235);
or U5543 (N_5543,N_4012,N_4489);
or U5544 (N_5544,N_4695,N_4692);
and U5545 (N_5545,N_4679,N_4274);
or U5546 (N_5546,N_4803,N_4861);
nor U5547 (N_5547,N_4771,N_4814);
nor U5548 (N_5548,N_4533,N_4506);
nor U5549 (N_5549,N_4124,N_4135);
xor U5550 (N_5550,N_4071,N_4429);
nand U5551 (N_5551,N_4242,N_4707);
nor U5552 (N_5552,N_4157,N_4351);
xor U5553 (N_5553,N_4618,N_4395);
xor U5554 (N_5554,N_4491,N_4550);
nand U5555 (N_5555,N_4381,N_4196);
or U5556 (N_5556,N_4601,N_4801);
nor U5557 (N_5557,N_4105,N_4742);
nor U5558 (N_5558,N_4236,N_4682);
nand U5559 (N_5559,N_4520,N_4637);
nand U5560 (N_5560,N_4732,N_4705);
nor U5561 (N_5561,N_4685,N_4080);
or U5562 (N_5562,N_4412,N_4595);
nor U5563 (N_5563,N_4861,N_4361);
nand U5564 (N_5564,N_4302,N_4718);
or U5565 (N_5565,N_4269,N_4717);
nor U5566 (N_5566,N_4749,N_4139);
nand U5567 (N_5567,N_4895,N_4020);
or U5568 (N_5568,N_4015,N_4663);
nand U5569 (N_5569,N_4158,N_4955);
nor U5570 (N_5570,N_4486,N_4506);
nor U5571 (N_5571,N_4645,N_4037);
nand U5572 (N_5572,N_4191,N_4281);
nor U5573 (N_5573,N_4161,N_4722);
nand U5574 (N_5574,N_4654,N_4518);
xnor U5575 (N_5575,N_4693,N_4610);
nor U5576 (N_5576,N_4698,N_4187);
and U5577 (N_5577,N_4215,N_4231);
and U5578 (N_5578,N_4077,N_4870);
xnor U5579 (N_5579,N_4245,N_4888);
or U5580 (N_5580,N_4689,N_4180);
or U5581 (N_5581,N_4105,N_4456);
xor U5582 (N_5582,N_4946,N_4719);
xor U5583 (N_5583,N_4125,N_4723);
and U5584 (N_5584,N_4256,N_4482);
or U5585 (N_5585,N_4003,N_4291);
and U5586 (N_5586,N_4379,N_4515);
or U5587 (N_5587,N_4313,N_4643);
xor U5588 (N_5588,N_4681,N_4567);
nand U5589 (N_5589,N_4394,N_4919);
xnor U5590 (N_5590,N_4086,N_4033);
nand U5591 (N_5591,N_4228,N_4909);
and U5592 (N_5592,N_4699,N_4493);
or U5593 (N_5593,N_4739,N_4148);
or U5594 (N_5594,N_4698,N_4545);
nor U5595 (N_5595,N_4136,N_4372);
xor U5596 (N_5596,N_4056,N_4460);
xor U5597 (N_5597,N_4880,N_4480);
or U5598 (N_5598,N_4718,N_4930);
nand U5599 (N_5599,N_4009,N_4358);
or U5600 (N_5600,N_4690,N_4132);
xor U5601 (N_5601,N_4983,N_4180);
or U5602 (N_5602,N_4766,N_4389);
or U5603 (N_5603,N_4514,N_4385);
nor U5604 (N_5604,N_4081,N_4249);
xnor U5605 (N_5605,N_4313,N_4036);
nand U5606 (N_5606,N_4382,N_4204);
and U5607 (N_5607,N_4422,N_4151);
nand U5608 (N_5608,N_4534,N_4102);
or U5609 (N_5609,N_4589,N_4038);
or U5610 (N_5610,N_4522,N_4334);
nor U5611 (N_5611,N_4064,N_4328);
and U5612 (N_5612,N_4609,N_4818);
xnor U5613 (N_5613,N_4580,N_4541);
nor U5614 (N_5614,N_4981,N_4143);
nor U5615 (N_5615,N_4133,N_4312);
nand U5616 (N_5616,N_4320,N_4740);
and U5617 (N_5617,N_4325,N_4213);
xnor U5618 (N_5618,N_4885,N_4162);
and U5619 (N_5619,N_4419,N_4982);
xnor U5620 (N_5620,N_4861,N_4084);
or U5621 (N_5621,N_4480,N_4414);
xor U5622 (N_5622,N_4315,N_4748);
or U5623 (N_5623,N_4247,N_4303);
nor U5624 (N_5624,N_4883,N_4294);
or U5625 (N_5625,N_4840,N_4276);
nand U5626 (N_5626,N_4940,N_4115);
xnor U5627 (N_5627,N_4377,N_4392);
nor U5628 (N_5628,N_4202,N_4960);
or U5629 (N_5629,N_4295,N_4457);
or U5630 (N_5630,N_4248,N_4724);
nor U5631 (N_5631,N_4613,N_4428);
xnor U5632 (N_5632,N_4517,N_4353);
or U5633 (N_5633,N_4043,N_4622);
or U5634 (N_5634,N_4414,N_4608);
and U5635 (N_5635,N_4739,N_4613);
or U5636 (N_5636,N_4511,N_4265);
nor U5637 (N_5637,N_4233,N_4460);
nand U5638 (N_5638,N_4314,N_4812);
and U5639 (N_5639,N_4430,N_4307);
or U5640 (N_5640,N_4714,N_4694);
xor U5641 (N_5641,N_4139,N_4804);
or U5642 (N_5642,N_4676,N_4443);
xnor U5643 (N_5643,N_4539,N_4247);
nand U5644 (N_5644,N_4210,N_4009);
nand U5645 (N_5645,N_4115,N_4458);
or U5646 (N_5646,N_4534,N_4510);
xor U5647 (N_5647,N_4281,N_4496);
or U5648 (N_5648,N_4025,N_4939);
nor U5649 (N_5649,N_4065,N_4764);
and U5650 (N_5650,N_4830,N_4287);
xor U5651 (N_5651,N_4928,N_4033);
or U5652 (N_5652,N_4470,N_4971);
and U5653 (N_5653,N_4546,N_4421);
or U5654 (N_5654,N_4487,N_4002);
xnor U5655 (N_5655,N_4267,N_4993);
xor U5656 (N_5656,N_4183,N_4389);
xnor U5657 (N_5657,N_4719,N_4856);
and U5658 (N_5658,N_4070,N_4107);
or U5659 (N_5659,N_4687,N_4097);
and U5660 (N_5660,N_4656,N_4550);
xnor U5661 (N_5661,N_4848,N_4046);
xor U5662 (N_5662,N_4625,N_4250);
nor U5663 (N_5663,N_4986,N_4693);
xnor U5664 (N_5664,N_4809,N_4082);
nand U5665 (N_5665,N_4388,N_4616);
or U5666 (N_5666,N_4616,N_4717);
or U5667 (N_5667,N_4270,N_4063);
nand U5668 (N_5668,N_4718,N_4527);
or U5669 (N_5669,N_4665,N_4056);
nand U5670 (N_5670,N_4620,N_4259);
or U5671 (N_5671,N_4491,N_4363);
nor U5672 (N_5672,N_4855,N_4293);
nand U5673 (N_5673,N_4144,N_4469);
nand U5674 (N_5674,N_4030,N_4492);
nor U5675 (N_5675,N_4188,N_4325);
nand U5676 (N_5676,N_4590,N_4063);
nor U5677 (N_5677,N_4902,N_4101);
xor U5678 (N_5678,N_4591,N_4906);
and U5679 (N_5679,N_4330,N_4013);
nor U5680 (N_5680,N_4840,N_4728);
xor U5681 (N_5681,N_4626,N_4991);
nand U5682 (N_5682,N_4309,N_4415);
nand U5683 (N_5683,N_4707,N_4105);
and U5684 (N_5684,N_4358,N_4804);
xnor U5685 (N_5685,N_4104,N_4684);
nor U5686 (N_5686,N_4227,N_4187);
nor U5687 (N_5687,N_4817,N_4969);
xor U5688 (N_5688,N_4424,N_4028);
or U5689 (N_5689,N_4754,N_4445);
nor U5690 (N_5690,N_4625,N_4936);
and U5691 (N_5691,N_4924,N_4136);
xor U5692 (N_5692,N_4558,N_4591);
and U5693 (N_5693,N_4499,N_4626);
nor U5694 (N_5694,N_4679,N_4226);
and U5695 (N_5695,N_4327,N_4587);
or U5696 (N_5696,N_4369,N_4540);
and U5697 (N_5697,N_4381,N_4556);
or U5698 (N_5698,N_4228,N_4039);
or U5699 (N_5699,N_4951,N_4484);
and U5700 (N_5700,N_4337,N_4529);
and U5701 (N_5701,N_4587,N_4213);
nor U5702 (N_5702,N_4854,N_4434);
xor U5703 (N_5703,N_4524,N_4334);
nor U5704 (N_5704,N_4743,N_4398);
or U5705 (N_5705,N_4222,N_4327);
xor U5706 (N_5706,N_4807,N_4953);
nand U5707 (N_5707,N_4244,N_4393);
xnor U5708 (N_5708,N_4964,N_4378);
and U5709 (N_5709,N_4956,N_4771);
or U5710 (N_5710,N_4680,N_4433);
or U5711 (N_5711,N_4602,N_4410);
or U5712 (N_5712,N_4746,N_4880);
or U5713 (N_5713,N_4217,N_4884);
xnor U5714 (N_5714,N_4703,N_4475);
or U5715 (N_5715,N_4245,N_4733);
and U5716 (N_5716,N_4464,N_4150);
nor U5717 (N_5717,N_4072,N_4677);
nor U5718 (N_5718,N_4422,N_4228);
and U5719 (N_5719,N_4961,N_4108);
nand U5720 (N_5720,N_4479,N_4691);
and U5721 (N_5721,N_4429,N_4005);
nand U5722 (N_5722,N_4940,N_4928);
and U5723 (N_5723,N_4555,N_4494);
or U5724 (N_5724,N_4903,N_4510);
nor U5725 (N_5725,N_4617,N_4645);
nand U5726 (N_5726,N_4759,N_4596);
and U5727 (N_5727,N_4707,N_4722);
and U5728 (N_5728,N_4045,N_4301);
nand U5729 (N_5729,N_4116,N_4584);
and U5730 (N_5730,N_4521,N_4524);
nand U5731 (N_5731,N_4843,N_4996);
nand U5732 (N_5732,N_4071,N_4619);
nand U5733 (N_5733,N_4287,N_4707);
nand U5734 (N_5734,N_4512,N_4018);
nand U5735 (N_5735,N_4407,N_4011);
nand U5736 (N_5736,N_4911,N_4558);
nor U5737 (N_5737,N_4398,N_4863);
or U5738 (N_5738,N_4607,N_4770);
nor U5739 (N_5739,N_4269,N_4520);
or U5740 (N_5740,N_4619,N_4562);
nand U5741 (N_5741,N_4746,N_4732);
or U5742 (N_5742,N_4590,N_4429);
nor U5743 (N_5743,N_4343,N_4095);
and U5744 (N_5744,N_4439,N_4558);
xor U5745 (N_5745,N_4582,N_4119);
nor U5746 (N_5746,N_4514,N_4961);
or U5747 (N_5747,N_4556,N_4525);
and U5748 (N_5748,N_4496,N_4859);
and U5749 (N_5749,N_4061,N_4926);
nand U5750 (N_5750,N_4053,N_4878);
nand U5751 (N_5751,N_4080,N_4415);
or U5752 (N_5752,N_4765,N_4888);
and U5753 (N_5753,N_4179,N_4905);
or U5754 (N_5754,N_4521,N_4500);
nand U5755 (N_5755,N_4293,N_4446);
or U5756 (N_5756,N_4106,N_4937);
nand U5757 (N_5757,N_4996,N_4904);
or U5758 (N_5758,N_4714,N_4262);
nor U5759 (N_5759,N_4176,N_4590);
and U5760 (N_5760,N_4162,N_4632);
or U5761 (N_5761,N_4078,N_4919);
nor U5762 (N_5762,N_4810,N_4687);
nor U5763 (N_5763,N_4723,N_4986);
or U5764 (N_5764,N_4330,N_4891);
nor U5765 (N_5765,N_4390,N_4002);
xor U5766 (N_5766,N_4097,N_4639);
and U5767 (N_5767,N_4202,N_4949);
or U5768 (N_5768,N_4451,N_4045);
or U5769 (N_5769,N_4288,N_4628);
or U5770 (N_5770,N_4971,N_4656);
nand U5771 (N_5771,N_4453,N_4119);
or U5772 (N_5772,N_4317,N_4498);
and U5773 (N_5773,N_4911,N_4840);
nor U5774 (N_5774,N_4914,N_4345);
nor U5775 (N_5775,N_4399,N_4149);
or U5776 (N_5776,N_4590,N_4420);
nor U5777 (N_5777,N_4245,N_4526);
xnor U5778 (N_5778,N_4443,N_4314);
or U5779 (N_5779,N_4971,N_4087);
or U5780 (N_5780,N_4904,N_4470);
xor U5781 (N_5781,N_4439,N_4114);
and U5782 (N_5782,N_4751,N_4244);
nand U5783 (N_5783,N_4833,N_4798);
and U5784 (N_5784,N_4881,N_4540);
and U5785 (N_5785,N_4618,N_4225);
nor U5786 (N_5786,N_4637,N_4599);
nand U5787 (N_5787,N_4818,N_4233);
nand U5788 (N_5788,N_4105,N_4177);
nor U5789 (N_5789,N_4979,N_4629);
and U5790 (N_5790,N_4546,N_4330);
nor U5791 (N_5791,N_4094,N_4465);
nand U5792 (N_5792,N_4804,N_4112);
nor U5793 (N_5793,N_4101,N_4928);
nand U5794 (N_5794,N_4506,N_4677);
nand U5795 (N_5795,N_4805,N_4349);
xor U5796 (N_5796,N_4062,N_4115);
xnor U5797 (N_5797,N_4804,N_4103);
and U5798 (N_5798,N_4466,N_4687);
xor U5799 (N_5799,N_4586,N_4117);
or U5800 (N_5800,N_4434,N_4931);
or U5801 (N_5801,N_4482,N_4167);
or U5802 (N_5802,N_4512,N_4325);
nor U5803 (N_5803,N_4982,N_4815);
xor U5804 (N_5804,N_4247,N_4664);
nand U5805 (N_5805,N_4709,N_4822);
nand U5806 (N_5806,N_4534,N_4243);
nor U5807 (N_5807,N_4207,N_4972);
nand U5808 (N_5808,N_4619,N_4278);
xor U5809 (N_5809,N_4616,N_4327);
nor U5810 (N_5810,N_4683,N_4939);
and U5811 (N_5811,N_4887,N_4612);
xnor U5812 (N_5812,N_4073,N_4159);
nor U5813 (N_5813,N_4658,N_4991);
nor U5814 (N_5814,N_4831,N_4515);
or U5815 (N_5815,N_4019,N_4818);
xnor U5816 (N_5816,N_4114,N_4787);
nor U5817 (N_5817,N_4498,N_4481);
xor U5818 (N_5818,N_4395,N_4564);
nand U5819 (N_5819,N_4537,N_4701);
nor U5820 (N_5820,N_4643,N_4303);
nand U5821 (N_5821,N_4495,N_4298);
nor U5822 (N_5822,N_4326,N_4674);
xnor U5823 (N_5823,N_4007,N_4600);
or U5824 (N_5824,N_4443,N_4623);
or U5825 (N_5825,N_4249,N_4505);
and U5826 (N_5826,N_4565,N_4481);
nand U5827 (N_5827,N_4447,N_4728);
nor U5828 (N_5828,N_4654,N_4058);
nand U5829 (N_5829,N_4417,N_4575);
and U5830 (N_5830,N_4277,N_4998);
or U5831 (N_5831,N_4143,N_4061);
and U5832 (N_5832,N_4425,N_4750);
or U5833 (N_5833,N_4915,N_4783);
and U5834 (N_5834,N_4476,N_4455);
or U5835 (N_5835,N_4461,N_4291);
and U5836 (N_5836,N_4481,N_4259);
nor U5837 (N_5837,N_4938,N_4388);
nand U5838 (N_5838,N_4827,N_4044);
and U5839 (N_5839,N_4715,N_4889);
nor U5840 (N_5840,N_4370,N_4193);
xor U5841 (N_5841,N_4255,N_4436);
nor U5842 (N_5842,N_4254,N_4178);
nand U5843 (N_5843,N_4294,N_4799);
xor U5844 (N_5844,N_4405,N_4876);
xor U5845 (N_5845,N_4464,N_4856);
nand U5846 (N_5846,N_4418,N_4942);
nor U5847 (N_5847,N_4030,N_4090);
or U5848 (N_5848,N_4972,N_4485);
and U5849 (N_5849,N_4884,N_4327);
nand U5850 (N_5850,N_4850,N_4705);
nor U5851 (N_5851,N_4595,N_4553);
xnor U5852 (N_5852,N_4771,N_4863);
or U5853 (N_5853,N_4227,N_4773);
xor U5854 (N_5854,N_4683,N_4342);
xor U5855 (N_5855,N_4085,N_4778);
xor U5856 (N_5856,N_4581,N_4633);
or U5857 (N_5857,N_4897,N_4127);
and U5858 (N_5858,N_4076,N_4930);
nand U5859 (N_5859,N_4387,N_4832);
and U5860 (N_5860,N_4478,N_4833);
xnor U5861 (N_5861,N_4459,N_4272);
xor U5862 (N_5862,N_4557,N_4988);
xor U5863 (N_5863,N_4459,N_4297);
and U5864 (N_5864,N_4473,N_4796);
and U5865 (N_5865,N_4895,N_4146);
nor U5866 (N_5866,N_4785,N_4090);
xnor U5867 (N_5867,N_4862,N_4963);
and U5868 (N_5868,N_4988,N_4598);
nand U5869 (N_5869,N_4035,N_4591);
nor U5870 (N_5870,N_4999,N_4924);
nand U5871 (N_5871,N_4640,N_4342);
nand U5872 (N_5872,N_4027,N_4524);
nor U5873 (N_5873,N_4955,N_4577);
or U5874 (N_5874,N_4762,N_4555);
nand U5875 (N_5875,N_4126,N_4761);
nand U5876 (N_5876,N_4699,N_4027);
or U5877 (N_5877,N_4490,N_4063);
nand U5878 (N_5878,N_4566,N_4151);
xnor U5879 (N_5879,N_4752,N_4934);
nand U5880 (N_5880,N_4522,N_4705);
or U5881 (N_5881,N_4292,N_4888);
nor U5882 (N_5882,N_4214,N_4843);
nand U5883 (N_5883,N_4283,N_4592);
xor U5884 (N_5884,N_4995,N_4110);
xor U5885 (N_5885,N_4724,N_4615);
nor U5886 (N_5886,N_4051,N_4406);
or U5887 (N_5887,N_4897,N_4106);
nor U5888 (N_5888,N_4208,N_4228);
nand U5889 (N_5889,N_4050,N_4955);
and U5890 (N_5890,N_4295,N_4537);
xor U5891 (N_5891,N_4822,N_4279);
and U5892 (N_5892,N_4798,N_4427);
and U5893 (N_5893,N_4079,N_4704);
nand U5894 (N_5894,N_4586,N_4305);
or U5895 (N_5895,N_4417,N_4117);
nand U5896 (N_5896,N_4587,N_4135);
nand U5897 (N_5897,N_4736,N_4431);
nand U5898 (N_5898,N_4395,N_4789);
and U5899 (N_5899,N_4603,N_4864);
nand U5900 (N_5900,N_4538,N_4411);
or U5901 (N_5901,N_4442,N_4975);
nor U5902 (N_5902,N_4007,N_4392);
nand U5903 (N_5903,N_4585,N_4308);
or U5904 (N_5904,N_4494,N_4535);
xnor U5905 (N_5905,N_4106,N_4682);
xnor U5906 (N_5906,N_4612,N_4850);
and U5907 (N_5907,N_4758,N_4696);
nand U5908 (N_5908,N_4362,N_4624);
nor U5909 (N_5909,N_4631,N_4201);
or U5910 (N_5910,N_4080,N_4526);
and U5911 (N_5911,N_4449,N_4555);
nand U5912 (N_5912,N_4204,N_4090);
nor U5913 (N_5913,N_4046,N_4796);
xor U5914 (N_5914,N_4061,N_4154);
nand U5915 (N_5915,N_4915,N_4631);
xor U5916 (N_5916,N_4242,N_4334);
nor U5917 (N_5917,N_4901,N_4425);
nor U5918 (N_5918,N_4691,N_4430);
nand U5919 (N_5919,N_4561,N_4585);
nor U5920 (N_5920,N_4623,N_4716);
and U5921 (N_5921,N_4721,N_4211);
nor U5922 (N_5922,N_4797,N_4483);
nand U5923 (N_5923,N_4609,N_4521);
nand U5924 (N_5924,N_4189,N_4054);
and U5925 (N_5925,N_4433,N_4505);
and U5926 (N_5926,N_4216,N_4562);
or U5927 (N_5927,N_4956,N_4572);
or U5928 (N_5928,N_4495,N_4920);
xor U5929 (N_5929,N_4823,N_4019);
nand U5930 (N_5930,N_4913,N_4721);
xnor U5931 (N_5931,N_4334,N_4083);
xnor U5932 (N_5932,N_4038,N_4467);
nor U5933 (N_5933,N_4488,N_4857);
nor U5934 (N_5934,N_4579,N_4226);
nor U5935 (N_5935,N_4905,N_4044);
or U5936 (N_5936,N_4068,N_4022);
xor U5937 (N_5937,N_4245,N_4563);
or U5938 (N_5938,N_4272,N_4825);
xnor U5939 (N_5939,N_4909,N_4594);
and U5940 (N_5940,N_4285,N_4841);
xor U5941 (N_5941,N_4048,N_4720);
and U5942 (N_5942,N_4684,N_4090);
xnor U5943 (N_5943,N_4582,N_4495);
xor U5944 (N_5944,N_4014,N_4184);
nor U5945 (N_5945,N_4856,N_4911);
and U5946 (N_5946,N_4385,N_4465);
nand U5947 (N_5947,N_4583,N_4536);
or U5948 (N_5948,N_4398,N_4735);
nor U5949 (N_5949,N_4008,N_4372);
and U5950 (N_5950,N_4809,N_4046);
nor U5951 (N_5951,N_4536,N_4433);
and U5952 (N_5952,N_4706,N_4041);
nand U5953 (N_5953,N_4078,N_4296);
or U5954 (N_5954,N_4190,N_4184);
nand U5955 (N_5955,N_4046,N_4235);
or U5956 (N_5956,N_4802,N_4409);
nor U5957 (N_5957,N_4593,N_4875);
and U5958 (N_5958,N_4851,N_4635);
xor U5959 (N_5959,N_4098,N_4553);
and U5960 (N_5960,N_4555,N_4736);
nor U5961 (N_5961,N_4747,N_4251);
nor U5962 (N_5962,N_4014,N_4981);
nor U5963 (N_5963,N_4370,N_4660);
and U5964 (N_5964,N_4537,N_4915);
xnor U5965 (N_5965,N_4219,N_4524);
xnor U5966 (N_5966,N_4385,N_4281);
nand U5967 (N_5967,N_4500,N_4761);
or U5968 (N_5968,N_4104,N_4956);
and U5969 (N_5969,N_4054,N_4360);
or U5970 (N_5970,N_4296,N_4627);
nor U5971 (N_5971,N_4579,N_4864);
nor U5972 (N_5972,N_4333,N_4989);
and U5973 (N_5973,N_4078,N_4409);
xnor U5974 (N_5974,N_4948,N_4190);
and U5975 (N_5975,N_4473,N_4680);
nor U5976 (N_5976,N_4999,N_4560);
nand U5977 (N_5977,N_4905,N_4489);
nor U5978 (N_5978,N_4782,N_4519);
and U5979 (N_5979,N_4477,N_4391);
or U5980 (N_5980,N_4437,N_4451);
or U5981 (N_5981,N_4579,N_4122);
nor U5982 (N_5982,N_4399,N_4465);
or U5983 (N_5983,N_4799,N_4638);
nor U5984 (N_5984,N_4969,N_4926);
nand U5985 (N_5985,N_4630,N_4373);
nor U5986 (N_5986,N_4661,N_4849);
or U5987 (N_5987,N_4650,N_4034);
or U5988 (N_5988,N_4405,N_4513);
or U5989 (N_5989,N_4600,N_4761);
nand U5990 (N_5990,N_4158,N_4405);
or U5991 (N_5991,N_4320,N_4286);
nand U5992 (N_5992,N_4454,N_4870);
nand U5993 (N_5993,N_4474,N_4683);
xor U5994 (N_5994,N_4905,N_4308);
or U5995 (N_5995,N_4198,N_4590);
or U5996 (N_5996,N_4062,N_4738);
nand U5997 (N_5997,N_4908,N_4952);
nand U5998 (N_5998,N_4436,N_4758);
or U5999 (N_5999,N_4152,N_4829);
or U6000 (N_6000,N_5363,N_5039);
nand U6001 (N_6001,N_5722,N_5399);
xnor U6002 (N_6002,N_5189,N_5266);
xor U6003 (N_6003,N_5340,N_5868);
nor U6004 (N_6004,N_5691,N_5038);
xor U6005 (N_6005,N_5646,N_5292);
xor U6006 (N_6006,N_5374,N_5098);
and U6007 (N_6007,N_5063,N_5777);
or U6008 (N_6008,N_5860,N_5336);
or U6009 (N_6009,N_5661,N_5566);
and U6010 (N_6010,N_5542,N_5889);
and U6011 (N_6011,N_5744,N_5465);
and U6012 (N_6012,N_5917,N_5931);
nand U6013 (N_6013,N_5423,N_5838);
nor U6014 (N_6014,N_5872,N_5252);
nand U6015 (N_6015,N_5182,N_5392);
or U6016 (N_6016,N_5186,N_5472);
xor U6017 (N_6017,N_5117,N_5273);
nand U6018 (N_6018,N_5065,N_5519);
and U6019 (N_6019,N_5386,N_5540);
xor U6020 (N_6020,N_5674,N_5520);
xor U6021 (N_6021,N_5298,N_5525);
xor U6022 (N_6022,N_5531,N_5832);
and U6023 (N_6023,N_5796,N_5563);
or U6024 (N_6024,N_5236,N_5496);
nor U6025 (N_6025,N_5968,N_5825);
and U6026 (N_6026,N_5573,N_5885);
xnor U6027 (N_6027,N_5651,N_5800);
or U6028 (N_6028,N_5157,N_5974);
xnor U6029 (N_6029,N_5761,N_5785);
xnor U6030 (N_6030,N_5676,N_5609);
or U6031 (N_6031,N_5263,N_5662);
and U6032 (N_6032,N_5062,N_5299);
nor U6033 (N_6033,N_5612,N_5359);
or U6034 (N_6034,N_5064,N_5242);
nand U6035 (N_6035,N_5059,N_5037);
nor U6036 (N_6036,N_5891,N_5396);
and U6037 (N_6037,N_5224,N_5258);
or U6038 (N_6038,N_5355,N_5874);
nand U6039 (N_6039,N_5094,N_5765);
nor U6040 (N_6040,N_5653,N_5394);
nor U6041 (N_6041,N_5068,N_5331);
nor U6042 (N_6042,N_5549,N_5710);
xnor U6043 (N_6043,N_5594,N_5578);
nor U6044 (N_6044,N_5920,N_5895);
nand U6045 (N_6045,N_5294,N_5639);
nor U6046 (N_6046,N_5663,N_5556);
xnor U6047 (N_6047,N_5978,N_5305);
and U6048 (N_6048,N_5339,N_5217);
and U6049 (N_6049,N_5051,N_5004);
or U6050 (N_6050,N_5324,N_5013);
and U6051 (N_6051,N_5929,N_5300);
nand U6052 (N_6052,N_5853,N_5763);
and U6053 (N_6053,N_5108,N_5364);
nand U6054 (N_6054,N_5767,N_5949);
xor U6055 (N_6055,N_5867,N_5183);
and U6056 (N_6056,N_5672,N_5600);
xnor U6057 (N_6057,N_5848,N_5577);
and U6058 (N_6058,N_5664,N_5174);
or U6059 (N_6059,N_5426,N_5124);
and U6060 (N_6060,N_5405,N_5097);
nor U6061 (N_6061,N_5367,N_5704);
nand U6062 (N_6062,N_5454,N_5192);
xnor U6063 (N_6063,N_5547,N_5541);
nor U6064 (N_6064,N_5175,N_5040);
and U6065 (N_6065,N_5981,N_5477);
xor U6066 (N_6066,N_5230,N_5781);
nor U6067 (N_6067,N_5247,N_5153);
xor U6068 (N_6068,N_5086,N_5060);
or U6069 (N_6069,N_5254,N_5003);
nand U6070 (N_6070,N_5634,N_5116);
and U6071 (N_6071,N_5738,N_5315);
nor U6072 (N_6072,N_5078,N_5162);
nand U6073 (N_6073,N_5122,N_5249);
or U6074 (N_6074,N_5746,N_5647);
nor U6075 (N_6075,N_5757,N_5128);
and U6076 (N_6076,N_5090,N_5870);
nor U6077 (N_6077,N_5479,N_5700);
nor U6078 (N_6078,N_5852,N_5089);
and U6079 (N_6079,N_5176,N_5548);
xnor U6080 (N_6080,N_5415,N_5407);
and U6081 (N_6081,N_5862,N_5512);
and U6082 (N_6082,N_5344,N_5125);
nor U6083 (N_6083,N_5989,N_5213);
nor U6084 (N_6084,N_5635,N_5136);
xnor U6085 (N_6085,N_5081,N_5311);
or U6086 (N_6086,N_5741,N_5726);
and U6087 (N_6087,N_5366,N_5864);
xnor U6088 (N_6088,N_5502,N_5421);
and U6089 (N_6089,N_5205,N_5732);
nand U6090 (N_6090,N_5554,N_5105);
xnor U6091 (N_6091,N_5383,N_5528);
and U6092 (N_6092,N_5231,N_5633);
and U6093 (N_6093,N_5952,N_5539);
or U6094 (N_6094,N_5042,N_5129);
and U6095 (N_6095,N_5202,N_5716);
or U6096 (N_6096,N_5380,N_5260);
and U6097 (N_6097,N_5018,N_5774);
xnor U6098 (N_6098,N_5666,N_5288);
nor U6099 (N_6099,N_5475,N_5518);
and U6100 (N_6100,N_5886,N_5474);
nor U6101 (N_6101,N_5375,N_5684);
xor U6102 (N_6102,N_5130,N_5131);
and U6103 (N_6103,N_5845,N_5591);
or U6104 (N_6104,N_5698,N_5026);
or U6105 (N_6105,N_5967,N_5002);
or U6106 (N_6106,N_5999,N_5717);
or U6107 (N_6107,N_5121,N_5016);
nand U6108 (N_6108,N_5986,N_5524);
nand U6109 (N_6109,N_5621,N_5842);
xnor U6110 (N_6110,N_5543,N_5028);
or U6111 (N_6111,N_5821,N_5823);
or U6112 (N_6112,N_5276,N_5836);
or U6113 (N_6113,N_5784,N_5846);
and U6114 (N_6114,N_5450,N_5576);
and U6115 (N_6115,N_5927,N_5811);
and U6116 (N_6116,N_5601,N_5087);
nand U6117 (N_6117,N_5681,N_5720);
or U6118 (N_6118,N_5526,N_5161);
xor U6119 (N_6119,N_5909,N_5899);
or U6120 (N_6120,N_5278,N_5995);
xnor U6121 (N_6121,N_5144,N_5010);
xnor U6122 (N_6122,N_5654,N_5517);
nand U6123 (N_6123,N_5951,N_5509);
and U6124 (N_6124,N_5317,N_5602);
nand U6125 (N_6125,N_5892,N_5001);
nor U6126 (N_6126,N_5873,N_5504);
nand U6127 (N_6127,N_5665,N_5679);
or U6128 (N_6128,N_5788,N_5748);
nor U6129 (N_6129,N_5753,N_5559);
nor U6130 (N_6130,N_5824,N_5023);
and U6131 (N_6131,N_5140,N_5992);
or U6132 (N_6132,N_5215,N_5962);
xor U6133 (N_6133,N_5462,N_5204);
and U6134 (N_6134,N_5341,N_5497);
or U6135 (N_6135,N_5228,N_5149);
nand U6136 (N_6136,N_5773,N_5533);
nor U6137 (N_6137,N_5277,N_5233);
or U6138 (N_6138,N_5841,N_5887);
nand U6139 (N_6139,N_5257,N_5485);
or U6140 (N_6140,N_5768,N_5812);
nand U6141 (N_6141,N_5114,N_5985);
and U6142 (N_6142,N_5072,N_5537);
nand U6143 (N_6143,N_5569,N_5043);
and U6144 (N_6144,N_5752,N_5631);
nand U6145 (N_6145,N_5077,N_5151);
and U6146 (N_6146,N_5819,N_5430);
xor U6147 (N_6147,N_5286,N_5932);
nand U6148 (N_6148,N_5431,N_5776);
and U6149 (N_6149,N_5172,N_5285);
nor U6150 (N_6150,N_5565,N_5749);
or U6151 (N_6151,N_5048,N_5201);
xnor U6152 (N_6152,N_5262,N_5088);
xnor U6153 (N_6153,N_5586,N_5483);
nand U6154 (N_6154,N_5207,N_5057);
xor U6155 (N_6155,N_5350,N_5333);
nor U6156 (N_6156,N_5314,N_5239);
nor U6157 (N_6157,N_5442,N_5027);
nand U6158 (N_6158,N_5379,N_5327);
nand U6159 (N_6159,N_5316,N_5735);
or U6160 (N_6160,N_5358,N_5181);
or U6161 (N_6161,N_5758,N_5670);
or U6162 (N_6162,N_5104,N_5325);
nand U6163 (N_6163,N_5481,N_5575);
and U6164 (N_6164,N_5850,N_5034);
nor U6165 (N_6165,N_5865,N_5851);
nand U6166 (N_6166,N_5115,N_5793);
or U6167 (N_6167,N_5582,N_5067);
and U6168 (N_6168,N_5580,N_5629);
xnor U6169 (N_6169,N_5395,N_5160);
xnor U6170 (N_6170,N_5323,N_5322);
nand U6171 (N_6171,N_5730,N_5611);
nor U6172 (N_6172,N_5342,N_5403);
xnor U6173 (N_6173,N_5268,N_5782);
nand U6174 (N_6174,N_5351,N_5253);
or U6175 (N_6175,N_5638,N_5965);
nand U6176 (N_6176,N_5771,N_5096);
or U6177 (N_6177,N_5963,N_5058);
nand U6178 (N_6178,N_5550,N_5218);
nand U6179 (N_6179,N_5925,N_5480);
or U6180 (N_6180,N_5792,N_5093);
nor U6181 (N_6181,N_5667,N_5148);
nand U6182 (N_6182,N_5269,N_5356);
xnor U6183 (N_6183,N_5282,N_5558);
nor U6184 (N_6184,N_5102,N_5076);
nand U6185 (N_6185,N_5914,N_5778);
xor U6186 (N_6186,N_5372,N_5216);
nor U6187 (N_6187,N_5424,N_5969);
and U6188 (N_6188,N_5234,N_5755);
nand U6189 (N_6189,N_5677,N_5461);
nor U6190 (N_6190,N_5113,N_5280);
nor U6191 (N_6191,N_5680,N_5604);
or U6192 (N_6192,N_5551,N_5926);
xor U6193 (N_6193,N_5420,N_5373);
and U6194 (N_6194,N_5830,N_5507);
and U6195 (N_6195,N_5417,N_5460);
xor U6196 (N_6196,N_5267,N_5107);
xnor U6197 (N_6197,N_5803,N_5588);
nand U6198 (N_6198,N_5489,N_5274);
or U6199 (N_6199,N_5406,N_5469);
and U6200 (N_6200,N_5809,N_5718);
xor U6201 (N_6201,N_5365,N_5177);
xor U6202 (N_6202,N_5046,N_5284);
xnor U6203 (N_6203,N_5139,N_5206);
xnor U6204 (N_6204,N_5400,N_5235);
xnor U6205 (N_6205,N_5522,N_5780);
or U6206 (N_6206,N_5901,N_5622);
nor U6207 (N_6207,N_5958,N_5142);
nor U6208 (N_6208,N_5956,N_5742);
nand U6209 (N_6209,N_5156,N_5100);
nand U6210 (N_6210,N_5453,N_5168);
and U6211 (N_6211,N_5011,N_5226);
nor U6212 (N_6212,N_5625,N_5238);
or U6213 (N_6213,N_5976,N_5835);
xnor U6214 (N_6214,N_5618,N_5326);
or U6215 (N_6215,N_5939,N_5593);
or U6216 (N_6216,N_5346,N_5849);
nand U6217 (N_6217,N_5291,N_5943);
nor U6218 (N_6218,N_5701,N_5227);
xor U6219 (N_6219,N_5947,N_5099);
or U6220 (N_6220,N_5402,N_5118);
or U6221 (N_6221,N_5728,N_5721);
xor U6222 (N_6222,N_5200,N_5025);
nand U6223 (N_6223,N_5246,N_5514);
and U6224 (N_6224,N_5737,N_5561);
xnor U6225 (N_6225,N_5908,N_5719);
nor U6226 (N_6226,N_5837,N_5050);
or U6227 (N_6227,N_5805,N_5476);
nor U6228 (N_6228,N_5733,N_5608);
and U6229 (N_6229,N_5219,N_5530);
nor U6230 (N_6230,N_5152,N_5434);
nand U6231 (N_6231,N_5546,N_5705);
nand U6232 (N_6232,N_5712,N_5779);
xnor U6233 (N_6233,N_5970,N_5135);
and U6234 (N_6234,N_5490,N_5723);
or U6235 (N_6235,N_5857,N_5191);
and U6236 (N_6236,N_5005,N_5378);
and U6237 (N_6237,N_5605,N_5270);
xor U6238 (N_6238,N_5132,N_5416);
or U6239 (N_6239,N_5856,N_5641);
nand U6240 (N_6240,N_5203,N_5772);
nor U6241 (N_6241,N_5673,N_5185);
nand U6242 (N_6242,N_5671,N_5134);
nand U6243 (N_6243,N_5014,N_5839);
and U6244 (N_6244,N_5789,N_5126);
and U6245 (N_6245,N_5583,N_5991);
nor U6246 (N_6246,N_5937,N_5448);
xnor U6247 (N_6247,N_5360,N_5628);
nor U6248 (N_6248,N_5880,N_5706);
nand U6249 (N_6249,N_5669,N_5008);
nand U6250 (N_6250,N_5702,N_5170);
xnor U6251 (N_6251,N_5632,N_5855);
xor U6252 (N_6252,N_5054,N_5897);
and U6253 (N_6253,N_5760,N_5387);
or U6254 (N_6254,N_5996,N_5451);
nor U6255 (N_6255,N_5523,N_5368);
nand U6256 (N_6256,N_5419,N_5119);
and U6257 (N_6257,N_5446,N_5942);
nor U6258 (N_6258,N_5210,N_5320);
nor U6259 (N_6259,N_5900,N_5345);
nand U6260 (N_6260,N_5946,N_5893);
or U6261 (N_6261,N_5815,N_5980);
nand U6262 (N_6262,N_5095,N_5281);
or U6263 (N_6263,N_5101,N_5302);
nor U6264 (N_6264,N_5377,N_5643);
nand U6265 (N_6265,N_5903,N_5869);
or U6266 (N_6266,N_5685,N_5397);
or U6267 (N_6267,N_5473,N_5188);
and U6268 (N_6268,N_5973,N_5456);
or U6269 (N_6269,N_5595,N_5686);
xor U6270 (N_6270,N_5699,N_5627);
xnor U6271 (N_6271,N_5910,N_5626);
or U6272 (N_6272,N_5499,N_5030);
nand U6273 (N_6273,N_5668,N_5173);
nor U6274 (N_6274,N_5933,N_5915);
xnor U6275 (N_6275,N_5488,N_5743);
and U6276 (N_6276,N_5391,N_5167);
or U6277 (N_6277,N_5876,N_5923);
or U6278 (N_6278,N_5944,N_5019);
xor U6279 (N_6279,N_5445,N_5179);
nor U6280 (N_6280,N_5898,N_5644);
nor U6281 (N_6281,N_5854,N_5145);
nand U6282 (N_6282,N_5906,N_5692);
xor U6283 (N_6283,N_5337,N_5560);
nand U6284 (N_6284,N_5994,N_5715);
or U6285 (N_6285,N_5388,N_5623);
and U6286 (N_6286,N_5444,N_5599);
nand U6287 (N_6287,N_5888,N_5491);
or U6288 (N_6288,N_5922,N_5052);
nor U6289 (N_6289,N_5624,N_5527);
and U6290 (N_6290,N_5979,N_5143);
nor U6291 (N_6291,N_5739,N_5301);
and U6292 (N_6292,N_5318,N_5410);
nand U6293 (N_6293,N_5637,N_5075);
xnor U6294 (N_6294,N_5930,N_5418);
nand U6295 (N_6295,N_5727,N_5801);
nor U6296 (N_6296,N_5935,N_5808);
nor U6297 (N_6297,N_5532,N_5330);
and U6298 (N_6298,N_5879,N_5658);
nand U6299 (N_6299,N_5826,N_5959);
or U6300 (N_6300,N_5357,N_5521);
nand U6301 (N_6301,N_5304,N_5552);
nand U6302 (N_6302,N_5766,N_5557);
nor U6303 (N_6303,N_5436,N_5289);
nand U6304 (N_6304,N_5581,N_5487);
and U6305 (N_6305,N_5354,N_5029);
nor U6306 (N_6306,N_5343,N_5687);
nor U6307 (N_6307,N_5615,N_5694);
and U6308 (N_6308,N_5422,N_5606);
and U6309 (N_6309,N_5572,N_5085);
and U6310 (N_6310,N_5237,N_5983);
nor U6311 (N_6311,N_5178,N_5964);
or U6312 (N_6312,N_5697,N_5412);
and U6313 (N_6313,N_5875,N_5740);
nor U6314 (N_6314,N_5443,N_5783);
nor U6315 (N_6315,N_5713,N_5287);
nor U6316 (N_6316,N_5248,N_5709);
xnor U6317 (N_6317,N_5275,N_5829);
or U6318 (N_6318,N_5180,N_5954);
nor U6319 (N_6319,N_5833,N_5494);
or U6320 (N_6320,N_5675,N_5084);
nor U6321 (N_6321,N_5660,N_5141);
and U6322 (N_6322,N_5478,N_5197);
nand U6323 (N_6323,N_5385,N_5492);
or U6324 (N_6324,N_5598,N_5938);
nand U6325 (N_6325,N_5810,N_5066);
and U6326 (N_6326,N_5907,N_5112);
nor U6327 (N_6327,N_5770,N_5847);
and U6328 (N_6328,N_5589,N_5376);
nor U6329 (N_6329,N_5321,N_5921);
and U6330 (N_6330,N_5877,N_5369);
xor U6331 (N_6331,N_5155,N_5229);
nor U6332 (N_6332,N_5871,N_5455);
or U6333 (N_6333,N_5592,N_5756);
and U6334 (N_6334,N_5017,N_5500);
nor U6335 (N_6335,N_5154,N_5120);
nand U6336 (N_6336,N_5433,N_5251);
or U6337 (N_6337,N_5564,N_5482);
xnor U6338 (N_6338,N_5225,N_5731);
or U6339 (N_6339,N_5127,N_5310);
xnor U6340 (N_6340,N_5585,N_5940);
nand U6341 (N_6341,N_5133,N_5223);
and U6342 (N_6342,N_5682,N_5069);
nand U6343 (N_6343,N_5484,N_5255);
xnor U6344 (N_6344,N_5193,N_5678);
or U6345 (N_6345,N_5147,N_5458);
or U6346 (N_6346,N_5441,N_5295);
or U6347 (N_6347,N_5306,N_5703);
xor U6348 (N_6348,N_5332,N_5381);
xor U6349 (N_6349,N_5169,N_5655);
nor U6350 (N_6350,N_5911,N_5438);
nand U6351 (N_6351,N_5813,N_5371);
nor U6352 (N_6352,N_5493,N_5389);
nor U6353 (N_6353,N_5544,N_5031);
and U6354 (N_6354,N_5505,N_5790);
xnor U6355 (N_6355,N_5998,N_5259);
xor U6356 (N_6356,N_5261,N_5409);
and U6357 (N_6357,N_5414,N_5083);
nor U6358 (N_6358,N_5022,N_5092);
nor U6359 (N_6359,N_5211,N_5972);
nor U6360 (N_6360,N_5427,N_5690);
nand U6361 (N_6361,N_5449,N_5617);
nand U6362 (N_6362,N_5882,N_5693);
and U6363 (N_6363,N_5272,N_5975);
xor U6364 (N_6364,N_5061,N_5290);
and U6365 (N_6365,N_5804,N_5109);
and U6366 (N_6366,N_5498,N_5652);
nand U6367 (N_6367,N_5074,N_5957);
and U6368 (N_6368,N_5584,N_5734);
nor U6369 (N_6369,N_5425,N_5960);
nand U6370 (N_6370,N_5787,N_5470);
and U6371 (N_6371,N_5070,N_5828);
nor U6372 (N_6372,N_5020,N_5603);
nor U6373 (N_6373,N_5948,N_5404);
nor U6374 (N_6374,N_5091,N_5645);
or U6375 (N_6375,N_5843,N_5111);
and U6376 (N_6376,N_5501,N_5918);
nor U6377 (N_6377,N_5440,N_5165);
and U6378 (N_6378,N_5199,N_5032);
or U6379 (N_6379,N_5159,N_5457);
nor U6380 (N_6380,N_5945,N_5794);
or U6381 (N_6381,N_5411,N_5607);
xnor U6382 (N_6382,N_5816,N_5319);
nand U6383 (N_6383,N_5123,N_5568);
nor U6384 (N_6384,N_5393,N_5881);
nand U6385 (N_6385,N_5764,N_5822);
or U6386 (N_6386,N_5538,N_5711);
and U6387 (N_6387,N_5007,N_5590);
xnor U6388 (N_6388,N_5171,N_5688);
nand U6389 (N_6389,N_5904,N_5799);
nor U6390 (N_6390,N_5208,N_5187);
xor U6391 (N_6391,N_5827,N_5447);
and U6392 (N_6392,N_5184,N_5035);
nor U6393 (N_6393,N_5055,N_5307);
nand U6394 (N_6394,N_5045,N_5928);
nor U6395 (N_6395,N_5265,N_5297);
or U6396 (N_6396,N_5866,N_5545);
nor U6397 (N_6397,N_5467,N_5163);
xor U6398 (N_6398,N_5630,N_5401);
nor U6399 (N_6399,N_5390,N_5640);
nor U6400 (N_6400,N_5106,N_5786);
nand U6401 (N_6401,N_5529,N_5190);
nor U6402 (N_6402,N_5913,N_5222);
nand U6403 (N_6403,N_5036,N_5814);
xor U6404 (N_6404,N_5198,N_5214);
xnor U6405 (N_6405,N_5695,N_5347);
nand U6406 (N_6406,N_5158,N_5006);
and U6407 (N_6407,N_5245,N_5831);
or U6408 (N_6408,N_5150,N_5000);
nand U6409 (N_6409,N_5110,N_5047);
or U6410 (N_6410,N_5610,N_5513);
or U6411 (N_6411,N_5049,N_5382);
and U6412 (N_6412,N_5503,N_5015);
or U6413 (N_6413,N_5240,N_5990);
xor U6414 (N_6414,N_5082,N_5437);
or U6415 (N_6415,N_5797,N_5195);
and U6416 (N_6416,N_5955,N_5890);
nor U6417 (N_6417,N_5338,N_5883);
nand U6418 (N_6418,N_5817,N_5335);
xor U6419 (N_6419,N_5614,N_5689);
and U6420 (N_6420,N_5936,N_5775);
nand U6421 (N_6421,N_5807,N_5508);
nand U6422 (N_6422,N_5353,N_5863);
or U6423 (N_6423,N_5751,N_5574);
and U6424 (N_6424,N_5009,N_5293);
nand U6425 (N_6425,N_5435,N_5243);
xor U6426 (N_6426,N_5495,N_5596);
and U6427 (N_6427,N_5619,N_5754);
nand U6428 (N_6428,N_5012,N_5279);
nor U6429 (N_6429,N_5349,N_5370);
xnor U6430 (N_6430,N_5079,N_5649);
nor U6431 (N_6431,N_5620,N_5648);
xnor U6432 (N_6432,N_5818,N_5428);
and U6433 (N_6433,N_5555,N_5264);
xor U6434 (N_6434,N_5536,N_5232);
xor U6435 (N_6435,N_5613,N_5656);
nand U6436 (N_6436,N_5724,N_5362);
or U6437 (N_6437,N_5452,N_5820);
xor U6438 (N_6438,N_5071,N_5747);
and U6439 (N_6439,N_5534,N_5736);
nand U6440 (N_6440,N_5553,N_5196);
xnor U6441 (N_6441,N_5166,N_5616);
xor U6442 (N_6442,N_5977,N_5950);
nor U6443 (N_6443,N_5636,N_5103);
and U6444 (N_6444,N_5997,N_5571);
nor U6445 (N_6445,N_5858,N_5941);
nand U6446 (N_6446,N_5516,N_5650);
and U6447 (N_6447,N_5587,N_5953);
nor U6448 (N_6448,N_5987,N_5137);
nor U6449 (N_6449,N_5221,N_5982);
and U6450 (N_6450,N_5984,N_5296);
and U6451 (N_6451,N_5313,N_5642);
xor U6452 (N_6452,N_5471,N_5510);
nand U6453 (N_6453,N_5033,N_5798);
nor U6454 (N_6454,N_5993,N_5398);
and U6455 (N_6455,N_5579,N_5861);
or U6456 (N_6456,N_5429,N_5659);
xor U6457 (N_6457,N_5146,N_5361);
xnor U6458 (N_6458,N_5802,N_5515);
or U6459 (N_6459,N_5459,N_5138);
or U6460 (N_6460,N_5657,N_5053);
xnor U6461 (N_6461,N_5073,N_5024);
nand U6462 (N_6462,N_5044,N_5329);
and U6463 (N_6463,N_5902,N_5408);
and U6464 (N_6464,N_5466,N_5309);
nor U6465 (N_6465,N_5439,N_5916);
or U6466 (N_6466,N_5283,N_5432);
and U6467 (N_6467,N_5878,N_5795);
nor U6468 (N_6468,N_5934,N_5464);
xor U6469 (N_6469,N_5971,N_5762);
nor U6470 (N_6470,N_5570,N_5256);
and U6471 (N_6471,N_5924,N_5769);
nor U6472 (N_6472,N_5334,N_5725);
or U6473 (N_6473,N_5966,N_5463);
nand U6474 (N_6474,N_5759,N_5894);
nor U6475 (N_6475,N_5750,N_5220);
nor U6476 (N_6476,N_5729,N_5988);
and U6477 (N_6477,N_5919,N_5511);
and U6478 (N_6478,N_5708,N_5250);
nand U6479 (N_6479,N_5745,N_5041);
nor U6480 (N_6480,N_5884,N_5468);
or U6481 (N_6481,N_5834,N_5021);
nand U6482 (N_6482,N_5859,N_5506);
or U6483 (N_6483,N_5844,N_5707);
and U6484 (N_6484,N_5080,N_5912);
nand U6485 (N_6485,N_5791,N_5696);
and U6486 (N_6486,N_5806,N_5896);
xor U6487 (N_6487,N_5384,N_5348);
and U6488 (N_6488,N_5328,N_5312);
or U6489 (N_6489,N_5212,N_5905);
nor U6490 (N_6490,N_5567,N_5961);
xnor U6491 (N_6491,N_5194,N_5271);
xnor U6492 (N_6492,N_5535,N_5352);
nand U6493 (N_6493,N_5244,N_5840);
nor U6494 (N_6494,N_5209,N_5413);
and U6495 (N_6495,N_5241,N_5308);
or U6496 (N_6496,N_5164,N_5683);
or U6497 (N_6497,N_5714,N_5303);
nor U6498 (N_6498,N_5486,N_5562);
and U6499 (N_6499,N_5056,N_5597);
or U6500 (N_6500,N_5234,N_5266);
or U6501 (N_6501,N_5336,N_5118);
and U6502 (N_6502,N_5283,N_5990);
nor U6503 (N_6503,N_5302,N_5040);
nor U6504 (N_6504,N_5467,N_5213);
xor U6505 (N_6505,N_5172,N_5855);
and U6506 (N_6506,N_5622,N_5733);
and U6507 (N_6507,N_5230,N_5200);
and U6508 (N_6508,N_5651,N_5431);
xnor U6509 (N_6509,N_5624,N_5732);
or U6510 (N_6510,N_5761,N_5622);
nand U6511 (N_6511,N_5856,N_5248);
xor U6512 (N_6512,N_5557,N_5301);
nand U6513 (N_6513,N_5941,N_5527);
or U6514 (N_6514,N_5953,N_5527);
or U6515 (N_6515,N_5534,N_5582);
nor U6516 (N_6516,N_5914,N_5506);
and U6517 (N_6517,N_5964,N_5790);
and U6518 (N_6518,N_5385,N_5909);
xnor U6519 (N_6519,N_5844,N_5266);
nand U6520 (N_6520,N_5275,N_5967);
and U6521 (N_6521,N_5017,N_5704);
xnor U6522 (N_6522,N_5499,N_5790);
nor U6523 (N_6523,N_5690,N_5814);
nor U6524 (N_6524,N_5379,N_5158);
or U6525 (N_6525,N_5315,N_5825);
and U6526 (N_6526,N_5214,N_5491);
and U6527 (N_6527,N_5170,N_5583);
and U6528 (N_6528,N_5084,N_5311);
or U6529 (N_6529,N_5813,N_5978);
xor U6530 (N_6530,N_5277,N_5095);
and U6531 (N_6531,N_5608,N_5360);
and U6532 (N_6532,N_5096,N_5782);
nor U6533 (N_6533,N_5745,N_5848);
or U6534 (N_6534,N_5485,N_5052);
and U6535 (N_6535,N_5711,N_5525);
and U6536 (N_6536,N_5935,N_5645);
nand U6537 (N_6537,N_5861,N_5645);
nand U6538 (N_6538,N_5826,N_5015);
and U6539 (N_6539,N_5261,N_5983);
xnor U6540 (N_6540,N_5144,N_5660);
nand U6541 (N_6541,N_5636,N_5414);
or U6542 (N_6542,N_5716,N_5397);
or U6543 (N_6543,N_5407,N_5561);
xnor U6544 (N_6544,N_5825,N_5866);
and U6545 (N_6545,N_5453,N_5565);
or U6546 (N_6546,N_5961,N_5091);
and U6547 (N_6547,N_5279,N_5989);
nand U6548 (N_6548,N_5548,N_5498);
or U6549 (N_6549,N_5745,N_5734);
and U6550 (N_6550,N_5457,N_5568);
nor U6551 (N_6551,N_5073,N_5089);
or U6552 (N_6552,N_5819,N_5970);
xor U6553 (N_6553,N_5820,N_5205);
and U6554 (N_6554,N_5056,N_5794);
xor U6555 (N_6555,N_5569,N_5657);
or U6556 (N_6556,N_5259,N_5262);
or U6557 (N_6557,N_5748,N_5767);
nor U6558 (N_6558,N_5564,N_5179);
and U6559 (N_6559,N_5845,N_5361);
nand U6560 (N_6560,N_5896,N_5136);
nor U6561 (N_6561,N_5741,N_5650);
or U6562 (N_6562,N_5327,N_5665);
or U6563 (N_6563,N_5328,N_5721);
xnor U6564 (N_6564,N_5956,N_5555);
nor U6565 (N_6565,N_5843,N_5695);
xnor U6566 (N_6566,N_5665,N_5334);
and U6567 (N_6567,N_5286,N_5962);
xnor U6568 (N_6568,N_5323,N_5168);
and U6569 (N_6569,N_5872,N_5228);
or U6570 (N_6570,N_5898,N_5449);
xor U6571 (N_6571,N_5118,N_5343);
nand U6572 (N_6572,N_5700,N_5520);
xor U6573 (N_6573,N_5603,N_5930);
and U6574 (N_6574,N_5717,N_5011);
or U6575 (N_6575,N_5032,N_5975);
xor U6576 (N_6576,N_5928,N_5681);
nor U6577 (N_6577,N_5655,N_5276);
nor U6578 (N_6578,N_5354,N_5191);
or U6579 (N_6579,N_5018,N_5444);
and U6580 (N_6580,N_5835,N_5907);
and U6581 (N_6581,N_5067,N_5331);
or U6582 (N_6582,N_5572,N_5836);
nand U6583 (N_6583,N_5597,N_5186);
nor U6584 (N_6584,N_5689,N_5009);
or U6585 (N_6585,N_5582,N_5488);
nor U6586 (N_6586,N_5957,N_5020);
and U6587 (N_6587,N_5995,N_5093);
and U6588 (N_6588,N_5979,N_5341);
nor U6589 (N_6589,N_5290,N_5162);
nor U6590 (N_6590,N_5289,N_5394);
and U6591 (N_6591,N_5864,N_5114);
and U6592 (N_6592,N_5992,N_5895);
or U6593 (N_6593,N_5387,N_5144);
or U6594 (N_6594,N_5396,N_5651);
nor U6595 (N_6595,N_5614,N_5074);
nand U6596 (N_6596,N_5389,N_5538);
and U6597 (N_6597,N_5182,N_5758);
nand U6598 (N_6598,N_5198,N_5812);
xor U6599 (N_6599,N_5929,N_5979);
or U6600 (N_6600,N_5913,N_5767);
xor U6601 (N_6601,N_5332,N_5312);
nor U6602 (N_6602,N_5093,N_5885);
or U6603 (N_6603,N_5029,N_5107);
xor U6604 (N_6604,N_5741,N_5591);
nand U6605 (N_6605,N_5792,N_5533);
and U6606 (N_6606,N_5990,N_5772);
xor U6607 (N_6607,N_5713,N_5522);
xor U6608 (N_6608,N_5417,N_5094);
nor U6609 (N_6609,N_5424,N_5965);
nor U6610 (N_6610,N_5457,N_5814);
xnor U6611 (N_6611,N_5882,N_5479);
nand U6612 (N_6612,N_5846,N_5627);
nor U6613 (N_6613,N_5886,N_5338);
xnor U6614 (N_6614,N_5157,N_5808);
nand U6615 (N_6615,N_5956,N_5539);
or U6616 (N_6616,N_5722,N_5525);
or U6617 (N_6617,N_5394,N_5157);
xnor U6618 (N_6618,N_5461,N_5934);
and U6619 (N_6619,N_5710,N_5495);
nand U6620 (N_6620,N_5609,N_5843);
xnor U6621 (N_6621,N_5120,N_5405);
and U6622 (N_6622,N_5687,N_5400);
xnor U6623 (N_6623,N_5328,N_5557);
xor U6624 (N_6624,N_5098,N_5834);
or U6625 (N_6625,N_5560,N_5786);
xor U6626 (N_6626,N_5195,N_5674);
nand U6627 (N_6627,N_5280,N_5156);
or U6628 (N_6628,N_5450,N_5873);
nand U6629 (N_6629,N_5754,N_5862);
nand U6630 (N_6630,N_5592,N_5124);
xnor U6631 (N_6631,N_5416,N_5692);
xor U6632 (N_6632,N_5144,N_5493);
xor U6633 (N_6633,N_5448,N_5172);
and U6634 (N_6634,N_5850,N_5248);
nand U6635 (N_6635,N_5957,N_5202);
xor U6636 (N_6636,N_5721,N_5841);
or U6637 (N_6637,N_5997,N_5053);
or U6638 (N_6638,N_5922,N_5021);
and U6639 (N_6639,N_5030,N_5332);
nor U6640 (N_6640,N_5508,N_5000);
nand U6641 (N_6641,N_5646,N_5152);
nor U6642 (N_6642,N_5622,N_5429);
and U6643 (N_6643,N_5069,N_5884);
or U6644 (N_6644,N_5808,N_5962);
xor U6645 (N_6645,N_5796,N_5598);
or U6646 (N_6646,N_5526,N_5383);
nor U6647 (N_6647,N_5775,N_5608);
nor U6648 (N_6648,N_5266,N_5994);
nor U6649 (N_6649,N_5072,N_5961);
nor U6650 (N_6650,N_5440,N_5128);
or U6651 (N_6651,N_5197,N_5212);
xor U6652 (N_6652,N_5885,N_5502);
and U6653 (N_6653,N_5222,N_5502);
nand U6654 (N_6654,N_5951,N_5814);
nand U6655 (N_6655,N_5702,N_5415);
and U6656 (N_6656,N_5324,N_5073);
nand U6657 (N_6657,N_5471,N_5940);
or U6658 (N_6658,N_5728,N_5154);
xor U6659 (N_6659,N_5091,N_5824);
nor U6660 (N_6660,N_5110,N_5473);
or U6661 (N_6661,N_5658,N_5983);
or U6662 (N_6662,N_5106,N_5694);
nor U6663 (N_6663,N_5264,N_5532);
nand U6664 (N_6664,N_5872,N_5145);
xnor U6665 (N_6665,N_5623,N_5378);
xor U6666 (N_6666,N_5935,N_5801);
or U6667 (N_6667,N_5091,N_5686);
nor U6668 (N_6668,N_5363,N_5397);
and U6669 (N_6669,N_5648,N_5804);
and U6670 (N_6670,N_5266,N_5301);
or U6671 (N_6671,N_5710,N_5987);
or U6672 (N_6672,N_5538,N_5180);
and U6673 (N_6673,N_5204,N_5080);
or U6674 (N_6674,N_5553,N_5195);
and U6675 (N_6675,N_5699,N_5999);
or U6676 (N_6676,N_5906,N_5294);
nor U6677 (N_6677,N_5736,N_5824);
and U6678 (N_6678,N_5018,N_5189);
and U6679 (N_6679,N_5879,N_5502);
and U6680 (N_6680,N_5123,N_5083);
xor U6681 (N_6681,N_5210,N_5032);
or U6682 (N_6682,N_5584,N_5366);
or U6683 (N_6683,N_5936,N_5581);
and U6684 (N_6684,N_5943,N_5018);
and U6685 (N_6685,N_5197,N_5237);
nor U6686 (N_6686,N_5619,N_5225);
nor U6687 (N_6687,N_5774,N_5281);
nor U6688 (N_6688,N_5443,N_5758);
nand U6689 (N_6689,N_5156,N_5411);
nor U6690 (N_6690,N_5468,N_5396);
nand U6691 (N_6691,N_5887,N_5340);
nor U6692 (N_6692,N_5433,N_5871);
nand U6693 (N_6693,N_5350,N_5592);
nand U6694 (N_6694,N_5620,N_5477);
xnor U6695 (N_6695,N_5995,N_5098);
nor U6696 (N_6696,N_5238,N_5958);
and U6697 (N_6697,N_5583,N_5337);
nand U6698 (N_6698,N_5993,N_5289);
nor U6699 (N_6699,N_5373,N_5552);
nand U6700 (N_6700,N_5594,N_5345);
nand U6701 (N_6701,N_5492,N_5444);
nand U6702 (N_6702,N_5010,N_5526);
or U6703 (N_6703,N_5498,N_5501);
nand U6704 (N_6704,N_5874,N_5398);
or U6705 (N_6705,N_5359,N_5317);
and U6706 (N_6706,N_5214,N_5679);
xnor U6707 (N_6707,N_5641,N_5570);
nor U6708 (N_6708,N_5855,N_5913);
and U6709 (N_6709,N_5018,N_5114);
and U6710 (N_6710,N_5295,N_5956);
or U6711 (N_6711,N_5499,N_5911);
nor U6712 (N_6712,N_5438,N_5272);
and U6713 (N_6713,N_5215,N_5019);
xnor U6714 (N_6714,N_5474,N_5003);
or U6715 (N_6715,N_5739,N_5753);
nand U6716 (N_6716,N_5702,N_5016);
nor U6717 (N_6717,N_5345,N_5498);
and U6718 (N_6718,N_5777,N_5286);
or U6719 (N_6719,N_5244,N_5200);
or U6720 (N_6720,N_5688,N_5954);
xor U6721 (N_6721,N_5390,N_5732);
nand U6722 (N_6722,N_5756,N_5851);
and U6723 (N_6723,N_5293,N_5470);
or U6724 (N_6724,N_5587,N_5746);
xor U6725 (N_6725,N_5007,N_5797);
and U6726 (N_6726,N_5882,N_5002);
nor U6727 (N_6727,N_5651,N_5980);
or U6728 (N_6728,N_5128,N_5648);
and U6729 (N_6729,N_5946,N_5147);
nor U6730 (N_6730,N_5262,N_5580);
nand U6731 (N_6731,N_5359,N_5115);
or U6732 (N_6732,N_5076,N_5449);
nand U6733 (N_6733,N_5029,N_5353);
or U6734 (N_6734,N_5890,N_5083);
xnor U6735 (N_6735,N_5894,N_5762);
or U6736 (N_6736,N_5355,N_5269);
nand U6737 (N_6737,N_5267,N_5136);
or U6738 (N_6738,N_5444,N_5128);
or U6739 (N_6739,N_5782,N_5984);
nand U6740 (N_6740,N_5474,N_5081);
nor U6741 (N_6741,N_5852,N_5704);
and U6742 (N_6742,N_5396,N_5265);
nand U6743 (N_6743,N_5594,N_5405);
nor U6744 (N_6744,N_5678,N_5542);
xor U6745 (N_6745,N_5131,N_5726);
and U6746 (N_6746,N_5739,N_5690);
and U6747 (N_6747,N_5904,N_5445);
or U6748 (N_6748,N_5761,N_5748);
and U6749 (N_6749,N_5901,N_5657);
or U6750 (N_6750,N_5391,N_5299);
nand U6751 (N_6751,N_5234,N_5520);
xor U6752 (N_6752,N_5297,N_5786);
xor U6753 (N_6753,N_5900,N_5207);
xor U6754 (N_6754,N_5078,N_5095);
and U6755 (N_6755,N_5700,N_5648);
xnor U6756 (N_6756,N_5734,N_5884);
nor U6757 (N_6757,N_5837,N_5414);
and U6758 (N_6758,N_5454,N_5467);
nand U6759 (N_6759,N_5502,N_5814);
nor U6760 (N_6760,N_5684,N_5056);
or U6761 (N_6761,N_5165,N_5011);
xnor U6762 (N_6762,N_5212,N_5025);
nand U6763 (N_6763,N_5140,N_5579);
nand U6764 (N_6764,N_5390,N_5092);
nor U6765 (N_6765,N_5399,N_5002);
or U6766 (N_6766,N_5511,N_5250);
or U6767 (N_6767,N_5427,N_5900);
and U6768 (N_6768,N_5446,N_5131);
or U6769 (N_6769,N_5469,N_5276);
or U6770 (N_6770,N_5053,N_5390);
xor U6771 (N_6771,N_5939,N_5514);
nor U6772 (N_6772,N_5141,N_5840);
nand U6773 (N_6773,N_5577,N_5026);
nand U6774 (N_6774,N_5674,N_5806);
or U6775 (N_6775,N_5360,N_5796);
and U6776 (N_6776,N_5555,N_5224);
xor U6777 (N_6777,N_5054,N_5711);
nor U6778 (N_6778,N_5205,N_5612);
or U6779 (N_6779,N_5696,N_5812);
nand U6780 (N_6780,N_5982,N_5003);
nand U6781 (N_6781,N_5368,N_5803);
and U6782 (N_6782,N_5308,N_5823);
nand U6783 (N_6783,N_5500,N_5936);
and U6784 (N_6784,N_5596,N_5615);
nor U6785 (N_6785,N_5077,N_5430);
nand U6786 (N_6786,N_5305,N_5499);
nand U6787 (N_6787,N_5461,N_5817);
xor U6788 (N_6788,N_5113,N_5145);
xnor U6789 (N_6789,N_5893,N_5189);
nor U6790 (N_6790,N_5436,N_5035);
and U6791 (N_6791,N_5420,N_5449);
nor U6792 (N_6792,N_5438,N_5932);
nand U6793 (N_6793,N_5951,N_5966);
and U6794 (N_6794,N_5320,N_5592);
and U6795 (N_6795,N_5245,N_5756);
nand U6796 (N_6796,N_5585,N_5621);
nor U6797 (N_6797,N_5542,N_5444);
or U6798 (N_6798,N_5961,N_5066);
xor U6799 (N_6799,N_5279,N_5369);
or U6800 (N_6800,N_5683,N_5575);
xnor U6801 (N_6801,N_5947,N_5993);
nand U6802 (N_6802,N_5195,N_5930);
nor U6803 (N_6803,N_5205,N_5015);
and U6804 (N_6804,N_5858,N_5605);
or U6805 (N_6805,N_5870,N_5552);
xor U6806 (N_6806,N_5829,N_5353);
and U6807 (N_6807,N_5609,N_5192);
or U6808 (N_6808,N_5877,N_5911);
nor U6809 (N_6809,N_5703,N_5447);
xor U6810 (N_6810,N_5367,N_5427);
nand U6811 (N_6811,N_5235,N_5840);
nand U6812 (N_6812,N_5012,N_5918);
or U6813 (N_6813,N_5263,N_5423);
nand U6814 (N_6814,N_5671,N_5347);
xor U6815 (N_6815,N_5191,N_5071);
and U6816 (N_6816,N_5614,N_5394);
and U6817 (N_6817,N_5563,N_5200);
or U6818 (N_6818,N_5772,N_5646);
nor U6819 (N_6819,N_5750,N_5559);
xor U6820 (N_6820,N_5453,N_5426);
nor U6821 (N_6821,N_5689,N_5151);
nor U6822 (N_6822,N_5494,N_5078);
nor U6823 (N_6823,N_5235,N_5790);
nand U6824 (N_6824,N_5388,N_5293);
or U6825 (N_6825,N_5249,N_5080);
nand U6826 (N_6826,N_5941,N_5616);
nand U6827 (N_6827,N_5406,N_5027);
nand U6828 (N_6828,N_5902,N_5912);
nand U6829 (N_6829,N_5116,N_5329);
nor U6830 (N_6830,N_5070,N_5122);
and U6831 (N_6831,N_5469,N_5705);
and U6832 (N_6832,N_5914,N_5532);
nor U6833 (N_6833,N_5817,N_5647);
xnor U6834 (N_6834,N_5715,N_5023);
nand U6835 (N_6835,N_5542,N_5624);
nand U6836 (N_6836,N_5495,N_5354);
nand U6837 (N_6837,N_5381,N_5784);
or U6838 (N_6838,N_5030,N_5261);
xnor U6839 (N_6839,N_5958,N_5489);
xnor U6840 (N_6840,N_5887,N_5819);
nor U6841 (N_6841,N_5676,N_5763);
or U6842 (N_6842,N_5493,N_5507);
and U6843 (N_6843,N_5643,N_5800);
and U6844 (N_6844,N_5717,N_5505);
xor U6845 (N_6845,N_5852,N_5394);
nor U6846 (N_6846,N_5156,N_5296);
nand U6847 (N_6847,N_5244,N_5786);
nor U6848 (N_6848,N_5579,N_5484);
xnor U6849 (N_6849,N_5736,N_5182);
nor U6850 (N_6850,N_5681,N_5852);
and U6851 (N_6851,N_5333,N_5710);
nand U6852 (N_6852,N_5252,N_5002);
nor U6853 (N_6853,N_5092,N_5824);
xnor U6854 (N_6854,N_5880,N_5924);
nor U6855 (N_6855,N_5927,N_5362);
nand U6856 (N_6856,N_5552,N_5828);
and U6857 (N_6857,N_5545,N_5914);
nor U6858 (N_6858,N_5116,N_5346);
or U6859 (N_6859,N_5724,N_5779);
nand U6860 (N_6860,N_5548,N_5161);
or U6861 (N_6861,N_5616,N_5860);
nand U6862 (N_6862,N_5027,N_5856);
nor U6863 (N_6863,N_5310,N_5449);
nor U6864 (N_6864,N_5855,N_5257);
nor U6865 (N_6865,N_5804,N_5104);
nor U6866 (N_6866,N_5099,N_5474);
nor U6867 (N_6867,N_5545,N_5930);
nand U6868 (N_6868,N_5063,N_5469);
or U6869 (N_6869,N_5875,N_5851);
nand U6870 (N_6870,N_5813,N_5590);
nor U6871 (N_6871,N_5553,N_5809);
nor U6872 (N_6872,N_5498,N_5947);
or U6873 (N_6873,N_5151,N_5141);
xor U6874 (N_6874,N_5471,N_5991);
and U6875 (N_6875,N_5783,N_5110);
or U6876 (N_6876,N_5551,N_5408);
or U6877 (N_6877,N_5919,N_5313);
nand U6878 (N_6878,N_5526,N_5068);
nand U6879 (N_6879,N_5068,N_5891);
nor U6880 (N_6880,N_5561,N_5796);
nand U6881 (N_6881,N_5570,N_5188);
or U6882 (N_6882,N_5965,N_5709);
xnor U6883 (N_6883,N_5407,N_5478);
xnor U6884 (N_6884,N_5412,N_5392);
and U6885 (N_6885,N_5608,N_5200);
nand U6886 (N_6886,N_5318,N_5379);
or U6887 (N_6887,N_5362,N_5538);
or U6888 (N_6888,N_5130,N_5839);
or U6889 (N_6889,N_5787,N_5142);
nor U6890 (N_6890,N_5904,N_5456);
and U6891 (N_6891,N_5036,N_5470);
nor U6892 (N_6892,N_5413,N_5682);
xor U6893 (N_6893,N_5125,N_5885);
or U6894 (N_6894,N_5849,N_5899);
or U6895 (N_6895,N_5806,N_5255);
nand U6896 (N_6896,N_5241,N_5482);
and U6897 (N_6897,N_5485,N_5085);
xor U6898 (N_6898,N_5494,N_5573);
or U6899 (N_6899,N_5622,N_5635);
and U6900 (N_6900,N_5057,N_5065);
xnor U6901 (N_6901,N_5563,N_5742);
and U6902 (N_6902,N_5328,N_5842);
nand U6903 (N_6903,N_5926,N_5916);
or U6904 (N_6904,N_5505,N_5405);
xor U6905 (N_6905,N_5521,N_5042);
xor U6906 (N_6906,N_5963,N_5442);
nor U6907 (N_6907,N_5284,N_5629);
nand U6908 (N_6908,N_5313,N_5412);
nand U6909 (N_6909,N_5159,N_5391);
xor U6910 (N_6910,N_5837,N_5132);
or U6911 (N_6911,N_5272,N_5181);
and U6912 (N_6912,N_5613,N_5128);
or U6913 (N_6913,N_5142,N_5017);
nor U6914 (N_6914,N_5556,N_5847);
or U6915 (N_6915,N_5420,N_5077);
nand U6916 (N_6916,N_5261,N_5645);
nor U6917 (N_6917,N_5576,N_5853);
nand U6918 (N_6918,N_5803,N_5666);
or U6919 (N_6919,N_5000,N_5349);
nor U6920 (N_6920,N_5295,N_5294);
or U6921 (N_6921,N_5236,N_5493);
and U6922 (N_6922,N_5797,N_5798);
and U6923 (N_6923,N_5137,N_5614);
or U6924 (N_6924,N_5716,N_5226);
xor U6925 (N_6925,N_5111,N_5689);
nor U6926 (N_6926,N_5460,N_5506);
nand U6927 (N_6927,N_5465,N_5553);
nand U6928 (N_6928,N_5874,N_5696);
nor U6929 (N_6929,N_5712,N_5468);
xnor U6930 (N_6930,N_5205,N_5547);
nor U6931 (N_6931,N_5006,N_5771);
nor U6932 (N_6932,N_5556,N_5132);
or U6933 (N_6933,N_5470,N_5099);
nor U6934 (N_6934,N_5379,N_5617);
xor U6935 (N_6935,N_5129,N_5426);
nor U6936 (N_6936,N_5939,N_5581);
nor U6937 (N_6937,N_5733,N_5934);
xor U6938 (N_6938,N_5877,N_5260);
and U6939 (N_6939,N_5550,N_5234);
and U6940 (N_6940,N_5393,N_5731);
and U6941 (N_6941,N_5869,N_5450);
nor U6942 (N_6942,N_5005,N_5322);
and U6943 (N_6943,N_5978,N_5274);
and U6944 (N_6944,N_5689,N_5910);
xor U6945 (N_6945,N_5240,N_5085);
nand U6946 (N_6946,N_5503,N_5174);
xor U6947 (N_6947,N_5843,N_5304);
and U6948 (N_6948,N_5801,N_5324);
and U6949 (N_6949,N_5120,N_5032);
nand U6950 (N_6950,N_5645,N_5490);
nand U6951 (N_6951,N_5228,N_5178);
nand U6952 (N_6952,N_5779,N_5080);
and U6953 (N_6953,N_5325,N_5727);
or U6954 (N_6954,N_5234,N_5810);
xnor U6955 (N_6955,N_5119,N_5189);
or U6956 (N_6956,N_5404,N_5453);
xor U6957 (N_6957,N_5497,N_5521);
nor U6958 (N_6958,N_5620,N_5444);
and U6959 (N_6959,N_5963,N_5980);
nor U6960 (N_6960,N_5155,N_5171);
and U6961 (N_6961,N_5652,N_5008);
and U6962 (N_6962,N_5923,N_5213);
and U6963 (N_6963,N_5967,N_5566);
xnor U6964 (N_6964,N_5512,N_5098);
nand U6965 (N_6965,N_5154,N_5622);
nor U6966 (N_6966,N_5184,N_5764);
nor U6967 (N_6967,N_5230,N_5136);
xor U6968 (N_6968,N_5578,N_5043);
or U6969 (N_6969,N_5433,N_5924);
nor U6970 (N_6970,N_5018,N_5791);
nor U6971 (N_6971,N_5723,N_5185);
nand U6972 (N_6972,N_5000,N_5430);
nand U6973 (N_6973,N_5403,N_5416);
and U6974 (N_6974,N_5449,N_5583);
nand U6975 (N_6975,N_5036,N_5483);
or U6976 (N_6976,N_5556,N_5808);
or U6977 (N_6977,N_5501,N_5185);
nor U6978 (N_6978,N_5513,N_5529);
nor U6979 (N_6979,N_5150,N_5900);
or U6980 (N_6980,N_5905,N_5616);
xor U6981 (N_6981,N_5148,N_5056);
xor U6982 (N_6982,N_5734,N_5450);
nor U6983 (N_6983,N_5940,N_5154);
nor U6984 (N_6984,N_5872,N_5858);
nor U6985 (N_6985,N_5084,N_5444);
and U6986 (N_6986,N_5010,N_5702);
and U6987 (N_6987,N_5557,N_5697);
nand U6988 (N_6988,N_5750,N_5299);
and U6989 (N_6989,N_5320,N_5817);
or U6990 (N_6990,N_5093,N_5242);
nor U6991 (N_6991,N_5464,N_5105);
or U6992 (N_6992,N_5709,N_5570);
and U6993 (N_6993,N_5490,N_5336);
nor U6994 (N_6994,N_5456,N_5868);
or U6995 (N_6995,N_5921,N_5085);
nand U6996 (N_6996,N_5172,N_5090);
and U6997 (N_6997,N_5905,N_5510);
xnor U6998 (N_6998,N_5222,N_5818);
nor U6999 (N_6999,N_5444,N_5075);
nand U7000 (N_7000,N_6456,N_6997);
or U7001 (N_7001,N_6287,N_6406);
or U7002 (N_7002,N_6946,N_6345);
and U7003 (N_7003,N_6882,N_6437);
xnor U7004 (N_7004,N_6835,N_6523);
xnor U7005 (N_7005,N_6863,N_6401);
nor U7006 (N_7006,N_6839,N_6323);
or U7007 (N_7007,N_6162,N_6051);
and U7008 (N_7008,N_6830,N_6152);
nand U7009 (N_7009,N_6365,N_6273);
or U7010 (N_7010,N_6665,N_6029);
nor U7011 (N_7011,N_6389,N_6100);
xnor U7012 (N_7012,N_6881,N_6361);
nand U7013 (N_7013,N_6897,N_6360);
and U7014 (N_7014,N_6122,N_6126);
or U7015 (N_7015,N_6074,N_6561);
and U7016 (N_7016,N_6517,N_6724);
or U7017 (N_7017,N_6104,N_6395);
nand U7018 (N_7018,N_6777,N_6818);
nor U7019 (N_7019,N_6834,N_6915);
nand U7020 (N_7020,N_6021,N_6279);
nand U7021 (N_7021,N_6901,N_6663);
nor U7022 (N_7022,N_6366,N_6786);
and U7023 (N_7023,N_6763,N_6951);
nor U7024 (N_7024,N_6566,N_6033);
xor U7025 (N_7025,N_6353,N_6433);
nand U7026 (N_7026,N_6793,N_6772);
or U7027 (N_7027,N_6283,N_6128);
xnor U7028 (N_7028,N_6813,N_6962);
nand U7029 (N_7029,N_6142,N_6933);
xor U7030 (N_7030,N_6143,N_6837);
nand U7031 (N_7031,N_6014,N_6728);
nand U7032 (N_7032,N_6003,N_6699);
or U7033 (N_7033,N_6332,N_6963);
nand U7034 (N_7034,N_6879,N_6845);
xor U7035 (N_7035,N_6269,N_6828);
or U7036 (N_7036,N_6011,N_6646);
xnor U7037 (N_7037,N_6060,N_6335);
nand U7038 (N_7038,N_6094,N_6926);
xnor U7039 (N_7039,N_6854,N_6680);
nand U7040 (N_7040,N_6722,N_6106);
xor U7041 (N_7041,N_6661,N_6423);
nor U7042 (N_7042,N_6485,N_6877);
or U7043 (N_7043,N_6864,N_6719);
or U7044 (N_7044,N_6795,N_6027);
nand U7045 (N_7045,N_6120,N_6498);
nor U7046 (N_7046,N_6270,N_6820);
nor U7047 (N_7047,N_6922,N_6377);
nand U7048 (N_7048,N_6035,N_6505);
or U7049 (N_7049,N_6072,N_6560);
xnor U7050 (N_7050,N_6618,N_6204);
nand U7051 (N_7051,N_6391,N_6535);
and U7052 (N_7052,N_6579,N_6672);
or U7053 (N_7053,N_6949,N_6427);
nand U7054 (N_7054,N_6938,N_6165);
xor U7055 (N_7055,N_6540,N_6464);
xnor U7056 (N_7056,N_6292,N_6659);
xor U7057 (N_7057,N_6337,N_6862);
and U7058 (N_7058,N_6694,N_6534);
and U7059 (N_7059,N_6848,N_6707);
and U7060 (N_7060,N_6925,N_6622);
and U7061 (N_7061,N_6931,N_6764);
or U7062 (N_7062,N_6317,N_6359);
or U7063 (N_7063,N_6978,N_6017);
xnor U7064 (N_7064,N_6826,N_6354);
nor U7065 (N_7065,N_6172,N_6343);
xor U7066 (N_7066,N_6852,N_6265);
and U7067 (N_7067,N_6836,N_6616);
or U7068 (N_7068,N_6369,N_6333);
xor U7069 (N_7069,N_6649,N_6291);
and U7070 (N_7070,N_6179,N_6264);
nor U7071 (N_7071,N_6024,N_6206);
xor U7072 (N_7072,N_6895,N_6528);
and U7073 (N_7073,N_6967,N_6001);
or U7074 (N_7074,N_6583,N_6816);
and U7075 (N_7075,N_6999,N_6198);
and U7076 (N_7076,N_6666,N_6948);
nor U7077 (N_7077,N_6441,N_6746);
xor U7078 (N_7078,N_6606,N_6544);
xnor U7079 (N_7079,N_6910,N_6714);
xor U7080 (N_7080,N_6387,N_6564);
nand U7081 (N_7081,N_6068,N_6115);
and U7082 (N_7082,N_6687,N_6689);
nand U7083 (N_7083,N_6110,N_6013);
nor U7084 (N_7084,N_6015,N_6542);
nand U7085 (N_7085,N_6934,N_6303);
or U7086 (N_7086,N_6973,N_6478);
or U7087 (N_7087,N_6809,N_6936);
and U7088 (N_7088,N_6932,N_6496);
or U7089 (N_7089,N_6415,N_6522);
nor U7090 (N_7090,N_6582,N_6298);
and U7091 (N_7091,N_6349,N_6526);
nand U7092 (N_7092,N_6116,N_6741);
and U7093 (N_7093,N_6043,N_6411);
nor U7094 (N_7094,N_6501,N_6603);
nand U7095 (N_7095,N_6161,N_6339);
xnor U7096 (N_7096,N_6675,N_6455);
nand U7097 (N_7097,N_6903,N_6892);
or U7098 (N_7098,N_6815,N_6612);
nand U7099 (N_7099,N_6420,N_6226);
nand U7100 (N_7100,N_6766,N_6945);
nand U7101 (N_7101,N_6923,N_6236);
or U7102 (N_7102,N_6151,N_6222);
nand U7103 (N_7103,N_6524,N_6040);
or U7104 (N_7104,N_6458,N_6806);
or U7105 (N_7105,N_6054,N_6907);
or U7106 (N_7106,N_6166,N_6373);
nor U7107 (N_7107,N_6443,N_6187);
or U7108 (N_7108,N_6481,N_6944);
nand U7109 (N_7109,N_6905,N_6638);
and U7110 (N_7110,N_6727,N_6444);
or U7111 (N_7111,N_6657,N_6276);
nor U7112 (N_7112,N_6911,N_6346);
nand U7113 (N_7113,N_6593,N_6733);
nor U7114 (N_7114,N_6992,N_6851);
nor U7115 (N_7115,N_6531,N_6243);
or U7116 (N_7116,N_6008,N_6121);
xor U7117 (N_7117,N_6184,N_6347);
or U7118 (N_7118,N_6701,N_6434);
nor U7119 (N_7119,N_6617,N_6843);
or U7120 (N_7120,N_6306,N_6224);
or U7121 (N_7121,N_6334,N_6867);
or U7122 (N_7122,N_6696,N_6470);
nor U7123 (N_7123,N_6518,N_6254);
and U7124 (N_7124,N_6237,N_6639);
or U7125 (N_7125,N_6284,N_6872);
nor U7126 (N_7126,N_6705,N_6408);
xnor U7127 (N_7127,N_6082,N_6249);
nand U7128 (N_7128,N_6451,N_6990);
xor U7129 (N_7129,N_6555,N_6153);
nor U7130 (N_7130,N_6201,N_6469);
or U7131 (N_7131,N_6574,N_6798);
nor U7132 (N_7132,N_6429,N_6503);
nand U7133 (N_7133,N_6147,N_6484);
xor U7134 (N_7134,N_6131,N_6796);
and U7135 (N_7135,N_6930,N_6871);
or U7136 (N_7136,N_6145,N_6846);
nand U7137 (N_7137,N_6076,N_6738);
or U7138 (N_7138,N_6969,N_6327);
or U7139 (N_7139,N_6030,N_6575);
or U7140 (N_7140,N_6278,N_6573);
nand U7141 (N_7141,N_6987,N_6554);
nor U7142 (N_7142,N_6817,N_6929);
or U7143 (N_7143,N_6866,N_6869);
and U7144 (N_7144,N_6621,N_6736);
xnor U7145 (N_7145,N_6258,N_6829);
and U7146 (N_7146,N_6776,N_6421);
nand U7147 (N_7147,N_6630,N_6611);
or U7148 (N_7148,N_6025,N_6241);
xor U7149 (N_7149,N_6239,N_6918);
or U7150 (N_7150,N_6005,N_6170);
nor U7151 (N_7151,N_6823,N_6899);
and U7152 (N_7152,N_6174,N_6957);
and U7153 (N_7153,N_6625,N_6086);
nand U7154 (N_7154,N_6487,N_6197);
nor U7155 (N_7155,N_6465,N_6779);
or U7156 (N_7156,N_6220,N_6752);
xnor U7157 (N_7157,N_6855,N_6330);
xnor U7158 (N_7158,N_6263,N_6647);
and U7159 (N_7159,N_6750,N_6304);
nand U7160 (N_7160,N_6295,N_6405);
or U7161 (N_7161,N_6381,N_6223);
nand U7162 (N_7162,N_6860,N_6362);
nor U7163 (N_7163,N_6099,N_6417);
nor U7164 (N_7164,N_6902,N_6536);
nand U7165 (N_7165,N_6340,N_6504);
xnor U7166 (N_7166,N_6130,N_6018);
or U7167 (N_7167,N_6227,N_6314);
nor U7168 (N_7168,N_6732,N_6171);
xnor U7169 (N_7169,N_6693,N_6148);
nand U7170 (N_7170,N_6608,N_6594);
xnor U7171 (N_7171,N_6403,N_6802);
and U7172 (N_7172,N_6547,N_6384);
nor U7173 (N_7173,N_6585,N_6414);
and U7174 (N_7174,N_6371,N_6486);
or U7175 (N_7175,N_6590,N_6350);
and U7176 (N_7176,N_6023,N_6471);
and U7177 (N_7177,N_6286,N_6650);
xor U7178 (N_7178,N_6702,N_6324);
nor U7179 (N_7179,N_6480,N_6970);
or U7180 (N_7180,N_6697,N_6725);
xnor U7181 (N_7181,N_6160,N_6744);
xor U7182 (N_7182,N_6510,N_6037);
xnor U7183 (N_7183,N_6662,N_6525);
xnor U7184 (N_7184,N_6438,N_6873);
nor U7185 (N_7185,N_6461,N_6424);
or U7186 (N_7186,N_6450,N_6664);
xnor U7187 (N_7187,N_6971,N_6870);
xor U7188 (N_7188,N_6896,N_6726);
xor U7189 (N_7189,N_6824,N_6259);
or U7190 (N_7190,N_6508,N_6538);
nand U7191 (N_7191,N_6352,N_6475);
nor U7192 (N_7192,N_6418,N_6208);
xnor U7193 (N_7193,N_6132,N_6158);
and U7194 (N_7194,N_6520,N_6571);
and U7195 (N_7195,N_6311,N_6740);
and U7196 (N_7196,N_6118,N_6768);
nor U7197 (N_7197,N_6898,N_6173);
nor U7198 (N_7198,N_6580,N_6095);
or U7199 (N_7199,N_6889,N_6598);
or U7200 (N_7200,N_6256,N_6681);
or U7201 (N_7201,N_6453,N_6979);
xor U7202 (N_7202,N_6202,N_6615);
xor U7203 (N_7203,N_6016,N_6445);
nor U7204 (N_7204,N_6546,N_6642);
nand U7205 (N_7205,N_6937,N_6507);
nand U7206 (N_7206,N_6770,N_6993);
and U7207 (N_7207,N_6364,N_6460);
and U7208 (N_7208,N_6838,N_6549);
and U7209 (N_7209,N_6757,N_6336);
nand U7210 (N_7210,N_6467,N_6515);
or U7211 (N_7211,N_6570,N_6038);
nand U7212 (N_7212,N_6117,N_6217);
nand U7213 (N_7213,N_6010,N_6765);
nand U7214 (N_7214,N_6888,N_6952);
nand U7215 (N_7215,N_6342,N_6568);
and U7216 (N_7216,N_6394,N_6861);
and U7217 (N_7217,N_6190,N_6294);
or U7218 (N_7218,N_6410,N_6790);
nor U7219 (N_7219,N_6998,N_6318);
xnor U7220 (N_7220,N_6183,N_6940);
nor U7221 (N_7221,N_6045,N_6755);
xnor U7222 (N_7222,N_6626,N_6974);
xor U7223 (N_7223,N_6482,N_6552);
nor U7224 (N_7224,N_6039,N_6474);
nand U7225 (N_7225,N_6532,N_6692);
and U7226 (N_7226,N_6124,N_6326);
or U7227 (N_7227,N_6009,N_6066);
or U7228 (N_7228,N_6320,N_6767);
and U7229 (N_7229,N_6632,N_6211);
nand U7230 (N_7230,N_6519,N_6609);
xnor U7231 (N_7231,N_6084,N_6840);
nor U7232 (N_7232,N_6026,N_6716);
nand U7233 (N_7233,N_6676,N_6378);
nor U7234 (N_7234,N_6799,N_6137);
nand U7235 (N_7235,N_6442,N_6466);
nand U7236 (N_7236,N_6230,N_6251);
nor U7237 (N_7237,N_6297,N_6513);
or U7238 (N_7238,N_6379,N_6723);
xnor U7239 (N_7239,N_6556,N_6706);
or U7240 (N_7240,N_6995,N_6144);
nand U7241 (N_7241,N_6966,N_6492);
and U7242 (N_7242,N_6686,N_6215);
xor U7243 (N_7243,N_6983,N_6007);
nor U7244 (N_7244,N_6180,N_6042);
and U7245 (N_7245,N_6325,N_6578);
nand U7246 (N_7246,N_6792,N_6782);
nor U7247 (N_7247,N_6409,N_6233);
nor U7248 (N_7248,N_6383,N_6261);
nand U7249 (N_7249,N_6430,N_6351);
and U7250 (N_7250,N_6956,N_6097);
xnor U7251 (N_7251,N_6964,N_6577);
or U7252 (N_7252,N_6847,N_6034);
nor U7253 (N_7253,N_6098,N_6199);
nand U7254 (N_7254,N_6169,N_6558);
or U7255 (N_7255,N_6904,N_6654);
nand U7256 (N_7256,N_6338,N_6914);
or U7257 (N_7257,N_6272,N_6288);
and U7258 (N_7258,N_6277,N_6057);
and U7259 (N_7259,N_6375,N_6473);
nand U7260 (N_7260,N_6192,N_6791);
nand U7261 (N_7261,N_6514,N_6101);
and U7262 (N_7262,N_6880,N_6900);
and U7263 (N_7263,N_6252,N_6274);
nand U7264 (N_7264,N_6168,N_6127);
or U7265 (N_7265,N_6958,N_6400);
and U7266 (N_7266,N_6628,N_6402);
or U7267 (N_7267,N_6413,N_6031);
or U7268 (N_7268,N_6022,N_6643);
xor U7269 (N_7269,N_6656,N_6396);
or U7270 (N_7270,N_6849,N_6240);
xnor U7271 (N_7271,N_6228,N_6981);
xor U7272 (N_7272,N_6113,N_6134);
or U7273 (N_7273,N_6177,N_6189);
or U7274 (N_7274,N_6246,N_6671);
and U7275 (N_7275,N_6238,N_6586);
nor U7276 (N_7276,N_6457,N_6506);
or U7277 (N_7277,N_6355,N_6404);
xor U7278 (N_7278,N_6541,N_6231);
nand U7279 (N_7279,N_6712,N_6479);
xnor U7280 (N_7280,N_6250,N_6652);
nand U7281 (N_7281,N_6368,N_6827);
xnor U7282 (N_7282,N_6089,N_6221);
nor U7283 (N_7283,N_6721,N_6613);
nand U7284 (N_7284,N_6745,N_6805);
and U7285 (N_7285,N_6913,N_6093);
or U7286 (N_7286,N_6299,N_6631);
and U7287 (N_7287,N_6698,N_6248);
xor U7288 (N_7288,N_6856,N_6602);
xor U7289 (N_7289,N_6668,N_6376);
nor U7290 (N_7290,N_6658,N_6787);
xnor U7291 (N_7291,N_6103,N_6266);
nand U7292 (N_7292,N_6502,N_6748);
nand U7293 (N_7293,N_6947,N_6703);
xor U7294 (N_7294,N_6052,N_6300);
nor U7295 (N_7295,N_6214,N_6315);
or U7296 (N_7296,N_6280,N_6077);
xor U7297 (N_7297,N_6557,N_6119);
and U7298 (N_7298,N_6439,N_6919);
nor U7299 (N_7299,N_6452,N_6186);
and U7300 (N_7300,N_6977,N_6814);
or U7301 (N_7301,N_6512,N_6419);
nor U7302 (N_7302,N_6761,N_6388);
and U7303 (N_7303,N_6012,N_6123);
and U7304 (N_7304,N_6494,N_6111);
xor U7305 (N_7305,N_6316,N_6645);
or U7306 (N_7306,N_6653,N_6185);
or U7307 (N_7307,N_6200,N_6059);
and U7308 (N_7308,N_6576,N_6071);
and U7309 (N_7309,N_6397,N_6032);
nor U7310 (N_7310,N_6150,N_6125);
nand U7311 (N_7311,N_6917,N_6623);
xnor U7312 (N_7312,N_6312,N_6812);
and U7313 (N_7313,N_6247,N_6797);
nor U7314 (N_7314,N_6521,N_6041);
or U7315 (N_7315,N_6301,N_6669);
nor U7316 (N_7316,N_6924,N_6500);
xnor U7317 (N_7317,N_6067,N_6773);
and U7318 (N_7318,N_6807,N_6942);
nor U7319 (N_7319,N_6927,N_6530);
nor U7320 (N_7320,N_6462,N_6876);
nor U7321 (N_7321,N_6019,N_6730);
nand U7322 (N_7322,N_6778,N_6313);
nand U7323 (N_7323,N_6908,N_6988);
and U7324 (N_7324,N_6894,N_6156);
nand U7325 (N_7325,N_6225,N_6372);
nand U7326 (N_7326,N_6194,N_6271);
or U7327 (N_7327,N_6390,N_6203);
and U7328 (N_7328,N_6209,N_6509);
nor U7329 (N_7329,N_6002,N_6614);
and U7330 (N_7330,N_6619,N_6293);
nor U7331 (N_7331,N_6245,N_6769);
nand U7332 (N_7332,N_6747,N_6529);
and U7333 (N_7333,N_6428,N_6363);
nor U7334 (N_7334,N_6087,N_6006);
nand U7335 (N_7335,N_6660,N_6448);
xnor U7336 (N_7336,N_6175,N_6234);
nand U7337 (N_7337,N_6685,N_6563);
and U7338 (N_7338,N_6374,N_6641);
nor U7339 (N_7339,N_6309,N_6079);
or U7340 (N_7340,N_6307,N_6348);
nand U7341 (N_7341,N_6825,N_6717);
nor U7342 (N_7342,N_6891,N_6213);
and U7343 (N_7343,N_6781,N_6961);
xor U7344 (N_7344,N_6155,N_6167);
nor U7345 (N_7345,N_6065,N_6589);
nand U7346 (N_7346,N_6785,N_6088);
nand U7347 (N_7347,N_6841,N_6588);
nor U7348 (N_7348,N_6435,N_6874);
and U7349 (N_7349,N_6921,N_6688);
nor U7350 (N_7350,N_6604,N_6794);
xor U7351 (N_7351,N_6328,N_6743);
nor U7352 (N_7352,N_6229,N_6760);
or U7353 (N_7353,N_6803,N_6296);
nand U7354 (N_7354,N_6960,N_6463);
and U7355 (N_7355,N_6302,N_6253);
and U7356 (N_7356,N_6440,N_6991);
and U7357 (N_7357,N_6488,N_6857);
xnor U7358 (N_7358,N_6610,N_6587);
nor U7359 (N_7359,N_6595,N_6046);
or U7360 (N_7360,N_6235,N_6709);
nor U7361 (N_7361,N_6633,N_6819);
xnor U7362 (N_7362,N_6984,N_6720);
nand U7363 (N_7363,N_6064,N_6446);
or U7364 (N_7364,N_6607,N_6605);
or U7365 (N_7365,N_6591,N_6928);
nand U7366 (N_7366,N_6592,N_6620);
or U7367 (N_7367,N_6020,N_6972);
or U7368 (N_7368,N_6624,N_6912);
and U7369 (N_7369,N_6762,N_6108);
nor U7370 (N_7370,N_6109,N_6141);
nand U7371 (N_7371,N_6543,N_6629);
and U7372 (N_7372,N_6050,N_6138);
nor U7373 (N_7373,N_6887,N_6062);
nand U7374 (N_7374,N_6875,N_6416);
nor U7375 (N_7375,N_6955,N_6985);
nand U7376 (N_7376,N_6426,N_6695);
nand U7377 (N_7377,N_6275,N_6735);
nand U7378 (N_7378,N_6080,N_6385);
xnor U7379 (N_7379,N_6559,N_6810);
or U7380 (N_7380,N_6893,N_6367);
and U7381 (N_7381,N_6196,N_6996);
or U7382 (N_7382,N_6562,N_6737);
nor U7383 (N_7383,N_6176,N_6454);
or U7384 (N_7384,N_6569,N_6499);
xor U7385 (N_7385,N_6449,N_6751);
or U7386 (N_7386,N_6868,N_6788);
xor U7387 (N_7387,N_6651,N_6644);
or U7388 (N_7388,N_6690,N_6154);
xor U7389 (N_7389,N_6133,N_6683);
or U7390 (N_7390,N_6447,N_6382);
xnor U7391 (N_7391,N_6193,N_6821);
and U7392 (N_7392,N_6774,N_6207);
xor U7393 (N_7393,N_6163,N_6289);
xor U7394 (N_7394,N_6597,N_6102);
or U7395 (N_7395,N_6063,N_6980);
and U7396 (N_7396,N_6159,N_6801);
nand U7397 (N_7397,N_6081,N_6178);
nand U7398 (N_7398,N_6092,N_6634);
xor U7399 (N_7399,N_6056,N_6968);
and U7400 (N_7400,N_6356,N_6731);
or U7401 (N_7401,N_6070,N_6527);
xor U7402 (N_7402,N_6670,N_6489);
or U7403 (N_7403,N_6321,N_6425);
or U7404 (N_7404,N_6036,N_6704);
xor U7405 (N_7405,N_6112,N_6358);
nor U7406 (N_7406,N_6920,N_6511);
nand U7407 (N_7407,N_6212,N_6976);
or U7408 (N_7408,N_6545,N_6885);
xnor U7409 (N_7409,N_6090,N_6939);
and U7410 (N_7410,N_6808,N_6436);
nand U7411 (N_7411,N_6599,N_6906);
and U7412 (N_7412,N_6975,N_6565);
xor U7413 (N_7413,N_6242,N_6811);
or U7414 (N_7414,N_6069,N_6865);
xor U7415 (N_7415,N_6357,N_6267);
xor U7416 (N_7416,N_6537,N_6218);
and U7417 (N_7417,N_6771,N_6677);
or U7418 (N_7418,N_6055,N_6567);
and U7419 (N_7419,N_6539,N_6477);
nand U7420 (N_7420,N_6210,N_6953);
or U7421 (N_7421,N_6048,N_6789);
and U7422 (N_7422,N_6853,N_6329);
nand U7423 (N_7423,N_6004,N_6135);
and U7424 (N_7424,N_6718,N_6000);
or U7425 (N_7425,N_6850,N_6136);
nand U7426 (N_7426,N_6553,N_6308);
or U7427 (N_7427,N_6061,N_6257);
or U7428 (N_7428,N_6640,N_6742);
or U7429 (N_7429,N_6548,N_6584);
nor U7430 (N_7430,N_6550,N_6753);
nor U7431 (N_7431,N_6916,N_6831);
xor U7432 (N_7432,N_6483,N_6713);
or U7433 (N_7433,N_6078,N_6679);
or U7434 (N_7434,N_6491,N_6468);
nor U7435 (N_7435,N_6600,N_6305);
nor U7436 (N_7436,N_6935,N_6049);
nor U7437 (N_7437,N_6216,N_6407);
nand U7438 (N_7438,N_6859,N_6710);
nor U7439 (N_7439,N_6729,N_6804);
and U7440 (N_7440,N_6581,N_6832);
nor U7441 (N_7441,N_6341,N_6516);
nor U7442 (N_7442,N_6954,N_6627);
nand U7443 (N_7443,N_6244,N_6322);
nor U7444 (N_7444,N_6290,N_6886);
and U7445 (N_7445,N_6982,N_6191);
nor U7446 (N_7446,N_6884,N_6493);
nor U7447 (N_7447,N_6959,N_6422);
nand U7448 (N_7448,N_6380,N_6386);
nor U7449 (N_7449,N_6459,N_6533);
xnor U7450 (N_7450,N_6637,N_6994);
nor U7451 (N_7451,N_6195,N_6684);
nor U7452 (N_7452,N_6047,N_6682);
and U7453 (N_7453,N_6572,N_6319);
nor U7454 (N_7454,N_6673,N_6083);
or U7455 (N_7455,N_6219,N_6310);
and U7456 (N_7456,N_6085,N_6596);
or U7457 (N_7457,N_6648,N_6398);
nor U7458 (N_7458,N_6495,N_6800);
nor U7459 (N_7459,N_6399,N_6096);
and U7460 (N_7460,N_6708,N_6476);
and U7461 (N_7461,N_6497,N_6105);
nor U7462 (N_7462,N_6943,N_6667);
and U7463 (N_7463,N_6344,N_6181);
and U7464 (N_7464,N_6188,N_6490);
nand U7465 (N_7465,N_6053,N_6883);
and U7466 (N_7466,N_6833,N_6551);
nand U7467 (N_7467,N_6678,N_6044);
nand U7468 (N_7468,N_6775,N_6139);
xnor U7469 (N_7469,N_6655,N_6232);
or U7470 (N_7470,N_6331,N_6989);
nor U7471 (N_7471,N_6734,N_6950);
xor U7472 (N_7472,N_6073,N_6756);
nand U7473 (N_7473,N_6146,N_6844);
nand U7474 (N_7474,N_6075,N_6635);
and U7475 (N_7475,N_6370,N_6715);
nor U7476 (N_7476,N_6754,N_6674);
and U7477 (N_7477,N_6107,N_6091);
and U7478 (N_7478,N_6129,N_6986);
xnor U7479 (N_7479,N_6636,N_6431);
and U7480 (N_7480,N_6941,N_6739);
nand U7481 (N_7481,N_6157,N_6691);
and U7482 (N_7482,N_6255,N_6182);
nand U7483 (N_7483,N_6262,N_6393);
xnor U7484 (N_7484,N_6601,N_6392);
or U7485 (N_7485,N_6758,N_6784);
nor U7486 (N_7486,N_6890,N_6822);
and U7487 (N_7487,N_6260,N_6780);
xnor U7488 (N_7488,N_6281,N_6909);
and U7489 (N_7489,N_6759,N_6783);
xnor U7490 (N_7490,N_6749,N_6432);
and U7491 (N_7491,N_6965,N_6412);
xnor U7492 (N_7492,N_6285,N_6028);
or U7493 (N_7493,N_6282,N_6114);
xor U7494 (N_7494,N_6711,N_6858);
xnor U7495 (N_7495,N_6058,N_6164);
xnor U7496 (N_7496,N_6878,N_6842);
nor U7497 (N_7497,N_6268,N_6700);
xnor U7498 (N_7498,N_6149,N_6140);
nor U7499 (N_7499,N_6205,N_6472);
nor U7500 (N_7500,N_6281,N_6201);
xnor U7501 (N_7501,N_6533,N_6190);
nor U7502 (N_7502,N_6326,N_6147);
xnor U7503 (N_7503,N_6681,N_6342);
nand U7504 (N_7504,N_6600,N_6479);
nand U7505 (N_7505,N_6983,N_6611);
or U7506 (N_7506,N_6596,N_6485);
xor U7507 (N_7507,N_6678,N_6880);
nor U7508 (N_7508,N_6958,N_6427);
nor U7509 (N_7509,N_6662,N_6852);
nand U7510 (N_7510,N_6897,N_6099);
nand U7511 (N_7511,N_6036,N_6978);
nand U7512 (N_7512,N_6150,N_6464);
nor U7513 (N_7513,N_6135,N_6640);
or U7514 (N_7514,N_6141,N_6103);
nor U7515 (N_7515,N_6266,N_6268);
and U7516 (N_7516,N_6235,N_6784);
nand U7517 (N_7517,N_6516,N_6152);
or U7518 (N_7518,N_6152,N_6587);
and U7519 (N_7519,N_6000,N_6279);
and U7520 (N_7520,N_6853,N_6006);
xnor U7521 (N_7521,N_6912,N_6926);
and U7522 (N_7522,N_6755,N_6228);
xor U7523 (N_7523,N_6289,N_6930);
nor U7524 (N_7524,N_6851,N_6548);
nor U7525 (N_7525,N_6034,N_6079);
and U7526 (N_7526,N_6055,N_6894);
nand U7527 (N_7527,N_6420,N_6288);
nand U7528 (N_7528,N_6117,N_6473);
nor U7529 (N_7529,N_6860,N_6444);
or U7530 (N_7530,N_6451,N_6789);
nor U7531 (N_7531,N_6766,N_6671);
or U7532 (N_7532,N_6186,N_6818);
xor U7533 (N_7533,N_6871,N_6163);
xnor U7534 (N_7534,N_6513,N_6021);
nand U7535 (N_7535,N_6277,N_6687);
nand U7536 (N_7536,N_6696,N_6350);
or U7537 (N_7537,N_6439,N_6146);
xor U7538 (N_7538,N_6922,N_6071);
nor U7539 (N_7539,N_6197,N_6686);
nand U7540 (N_7540,N_6338,N_6641);
nor U7541 (N_7541,N_6504,N_6278);
and U7542 (N_7542,N_6565,N_6215);
xor U7543 (N_7543,N_6171,N_6301);
xnor U7544 (N_7544,N_6734,N_6210);
and U7545 (N_7545,N_6542,N_6574);
nand U7546 (N_7546,N_6327,N_6515);
and U7547 (N_7547,N_6621,N_6912);
nand U7548 (N_7548,N_6894,N_6425);
or U7549 (N_7549,N_6865,N_6371);
nor U7550 (N_7550,N_6919,N_6928);
and U7551 (N_7551,N_6056,N_6750);
nor U7552 (N_7552,N_6644,N_6117);
nor U7553 (N_7553,N_6029,N_6394);
xor U7554 (N_7554,N_6560,N_6887);
or U7555 (N_7555,N_6203,N_6815);
xor U7556 (N_7556,N_6442,N_6876);
nand U7557 (N_7557,N_6640,N_6188);
nor U7558 (N_7558,N_6785,N_6843);
xnor U7559 (N_7559,N_6830,N_6274);
or U7560 (N_7560,N_6354,N_6218);
nand U7561 (N_7561,N_6862,N_6695);
xor U7562 (N_7562,N_6579,N_6387);
xor U7563 (N_7563,N_6472,N_6365);
or U7564 (N_7564,N_6043,N_6739);
and U7565 (N_7565,N_6164,N_6657);
xnor U7566 (N_7566,N_6143,N_6024);
xnor U7567 (N_7567,N_6169,N_6048);
or U7568 (N_7568,N_6683,N_6945);
nor U7569 (N_7569,N_6470,N_6698);
or U7570 (N_7570,N_6316,N_6860);
nand U7571 (N_7571,N_6427,N_6807);
nand U7572 (N_7572,N_6382,N_6861);
or U7573 (N_7573,N_6772,N_6463);
or U7574 (N_7574,N_6667,N_6467);
xnor U7575 (N_7575,N_6687,N_6264);
and U7576 (N_7576,N_6406,N_6985);
nor U7577 (N_7577,N_6628,N_6239);
or U7578 (N_7578,N_6381,N_6847);
xnor U7579 (N_7579,N_6857,N_6947);
nand U7580 (N_7580,N_6691,N_6847);
xnor U7581 (N_7581,N_6320,N_6269);
and U7582 (N_7582,N_6224,N_6243);
and U7583 (N_7583,N_6560,N_6898);
nor U7584 (N_7584,N_6334,N_6411);
or U7585 (N_7585,N_6832,N_6398);
nor U7586 (N_7586,N_6813,N_6354);
or U7587 (N_7587,N_6055,N_6492);
nor U7588 (N_7588,N_6496,N_6691);
nor U7589 (N_7589,N_6952,N_6361);
and U7590 (N_7590,N_6046,N_6037);
xnor U7591 (N_7591,N_6855,N_6361);
and U7592 (N_7592,N_6098,N_6593);
and U7593 (N_7593,N_6379,N_6633);
xnor U7594 (N_7594,N_6296,N_6239);
nand U7595 (N_7595,N_6941,N_6388);
and U7596 (N_7596,N_6148,N_6676);
xor U7597 (N_7597,N_6903,N_6914);
xor U7598 (N_7598,N_6171,N_6960);
or U7599 (N_7599,N_6504,N_6324);
nor U7600 (N_7600,N_6057,N_6447);
and U7601 (N_7601,N_6661,N_6893);
xnor U7602 (N_7602,N_6789,N_6919);
or U7603 (N_7603,N_6075,N_6713);
or U7604 (N_7604,N_6823,N_6488);
or U7605 (N_7605,N_6733,N_6204);
and U7606 (N_7606,N_6788,N_6882);
xor U7607 (N_7607,N_6104,N_6948);
and U7608 (N_7608,N_6715,N_6893);
xnor U7609 (N_7609,N_6352,N_6795);
xor U7610 (N_7610,N_6714,N_6099);
or U7611 (N_7611,N_6426,N_6814);
and U7612 (N_7612,N_6312,N_6785);
and U7613 (N_7613,N_6478,N_6281);
nor U7614 (N_7614,N_6647,N_6870);
xor U7615 (N_7615,N_6816,N_6266);
xnor U7616 (N_7616,N_6761,N_6504);
xnor U7617 (N_7617,N_6763,N_6208);
and U7618 (N_7618,N_6484,N_6423);
nand U7619 (N_7619,N_6152,N_6726);
or U7620 (N_7620,N_6539,N_6239);
xor U7621 (N_7621,N_6650,N_6639);
nand U7622 (N_7622,N_6318,N_6603);
or U7623 (N_7623,N_6561,N_6940);
xnor U7624 (N_7624,N_6858,N_6074);
xor U7625 (N_7625,N_6359,N_6274);
nor U7626 (N_7626,N_6043,N_6655);
nor U7627 (N_7627,N_6088,N_6709);
and U7628 (N_7628,N_6336,N_6278);
xnor U7629 (N_7629,N_6737,N_6006);
nor U7630 (N_7630,N_6769,N_6279);
and U7631 (N_7631,N_6276,N_6427);
nor U7632 (N_7632,N_6502,N_6417);
nor U7633 (N_7633,N_6141,N_6427);
and U7634 (N_7634,N_6056,N_6321);
xor U7635 (N_7635,N_6300,N_6318);
nor U7636 (N_7636,N_6391,N_6350);
nor U7637 (N_7637,N_6294,N_6947);
nor U7638 (N_7638,N_6185,N_6935);
xnor U7639 (N_7639,N_6937,N_6552);
or U7640 (N_7640,N_6226,N_6224);
or U7641 (N_7641,N_6989,N_6484);
nor U7642 (N_7642,N_6665,N_6737);
or U7643 (N_7643,N_6954,N_6919);
xnor U7644 (N_7644,N_6453,N_6715);
nand U7645 (N_7645,N_6738,N_6388);
or U7646 (N_7646,N_6349,N_6148);
xor U7647 (N_7647,N_6427,N_6266);
or U7648 (N_7648,N_6304,N_6474);
nand U7649 (N_7649,N_6162,N_6811);
nand U7650 (N_7650,N_6625,N_6642);
nand U7651 (N_7651,N_6458,N_6733);
nand U7652 (N_7652,N_6392,N_6305);
xnor U7653 (N_7653,N_6336,N_6308);
nand U7654 (N_7654,N_6332,N_6784);
and U7655 (N_7655,N_6563,N_6406);
and U7656 (N_7656,N_6485,N_6326);
or U7657 (N_7657,N_6531,N_6379);
nor U7658 (N_7658,N_6936,N_6637);
nor U7659 (N_7659,N_6655,N_6031);
nand U7660 (N_7660,N_6506,N_6602);
nand U7661 (N_7661,N_6162,N_6341);
nand U7662 (N_7662,N_6362,N_6514);
xnor U7663 (N_7663,N_6210,N_6051);
nor U7664 (N_7664,N_6138,N_6736);
nor U7665 (N_7665,N_6341,N_6063);
xnor U7666 (N_7666,N_6044,N_6607);
nand U7667 (N_7667,N_6478,N_6762);
nor U7668 (N_7668,N_6993,N_6896);
xor U7669 (N_7669,N_6833,N_6999);
nor U7670 (N_7670,N_6312,N_6825);
nor U7671 (N_7671,N_6488,N_6250);
or U7672 (N_7672,N_6529,N_6559);
or U7673 (N_7673,N_6050,N_6110);
nor U7674 (N_7674,N_6116,N_6827);
nand U7675 (N_7675,N_6878,N_6308);
nor U7676 (N_7676,N_6790,N_6491);
and U7677 (N_7677,N_6260,N_6176);
xnor U7678 (N_7678,N_6637,N_6342);
nor U7679 (N_7679,N_6894,N_6366);
nor U7680 (N_7680,N_6772,N_6981);
and U7681 (N_7681,N_6291,N_6389);
and U7682 (N_7682,N_6221,N_6113);
or U7683 (N_7683,N_6015,N_6318);
or U7684 (N_7684,N_6604,N_6515);
nor U7685 (N_7685,N_6453,N_6487);
xor U7686 (N_7686,N_6287,N_6766);
and U7687 (N_7687,N_6243,N_6542);
or U7688 (N_7688,N_6367,N_6016);
nand U7689 (N_7689,N_6664,N_6283);
and U7690 (N_7690,N_6445,N_6321);
or U7691 (N_7691,N_6584,N_6445);
nor U7692 (N_7692,N_6468,N_6815);
and U7693 (N_7693,N_6078,N_6769);
nor U7694 (N_7694,N_6058,N_6342);
nand U7695 (N_7695,N_6604,N_6862);
and U7696 (N_7696,N_6540,N_6057);
and U7697 (N_7697,N_6668,N_6752);
nor U7698 (N_7698,N_6670,N_6756);
nor U7699 (N_7699,N_6112,N_6810);
or U7700 (N_7700,N_6358,N_6920);
xor U7701 (N_7701,N_6629,N_6053);
nand U7702 (N_7702,N_6098,N_6657);
xor U7703 (N_7703,N_6375,N_6738);
nand U7704 (N_7704,N_6242,N_6500);
nor U7705 (N_7705,N_6173,N_6138);
nor U7706 (N_7706,N_6257,N_6681);
or U7707 (N_7707,N_6413,N_6476);
and U7708 (N_7708,N_6983,N_6343);
xor U7709 (N_7709,N_6535,N_6438);
nor U7710 (N_7710,N_6854,N_6412);
or U7711 (N_7711,N_6321,N_6962);
xnor U7712 (N_7712,N_6181,N_6718);
xnor U7713 (N_7713,N_6457,N_6841);
nor U7714 (N_7714,N_6403,N_6963);
xor U7715 (N_7715,N_6469,N_6623);
and U7716 (N_7716,N_6438,N_6466);
nand U7717 (N_7717,N_6418,N_6190);
or U7718 (N_7718,N_6149,N_6536);
and U7719 (N_7719,N_6015,N_6605);
and U7720 (N_7720,N_6831,N_6372);
xnor U7721 (N_7721,N_6667,N_6958);
xnor U7722 (N_7722,N_6325,N_6977);
nand U7723 (N_7723,N_6596,N_6566);
nor U7724 (N_7724,N_6767,N_6181);
xor U7725 (N_7725,N_6574,N_6230);
nor U7726 (N_7726,N_6241,N_6583);
or U7727 (N_7727,N_6127,N_6991);
or U7728 (N_7728,N_6373,N_6914);
xor U7729 (N_7729,N_6846,N_6606);
nand U7730 (N_7730,N_6559,N_6077);
or U7731 (N_7731,N_6209,N_6223);
nand U7732 (N_7732,N_6394,N_6568);
nand U7733 (N_7733,N_6761,N_6427);
and U7734 (N_7734,N_6051,N_6045);
xor U7735 (N_7735,N_6678,N_6893);
xnor U7736 (N_7736,N_6882,N_6583);
and U7737 (N_7737,N_6403,N_6734);
xnor U7738 (N_7738,N_6691,N_6784);
and U7739 (N_7739,N_6558,N_6216);
and U7740 (N_7740,N_6844,N_6907);
xnor U7741 (N_7741,N_6390,N_6609);
and U7742 (N_7742,N_6068,N_6197);
nor U7743 (N_7743,N_6650,N_6217);
or U7744 (N_7744,N_6920,N_6997);
nor U7745 (N_7745,N_6673,N_6858);
or U7746 (N_7746,N_6601,N_6503);
or U7747 (N_7747,N_6807,N_6509);
and U7748 (N_7748,N_6107,N_6213);
nand U7749 (N_7749,N_6684,N_6770);
and U7750 (N_7750,N_6745,N_6341);
or U7751 (N_7751,N_6452,N_6362);
nand U7752 (N_7752,N_6754,N_6244);
and U7753 (N_7753,N_6006,N_6413);
or U7754 (N_7754,N_6366,N_6185);
and U7755 (N_7755,N_6221,N_6432);
nand U7756 (N_7756,N_6191,N_6522);
or U7757 (N_7757,N_6712,N_6142);
nand U7758 (N_7758,N_6626,N_6273);
nand U7759 (N_7759,N_6871,N_6964);
and U7760 (N_7760,N_6031,N_6201);
xor U7761 (N_7761,N_6542,N_6252);
xor U7762 (N_7762,N_6431,N_6166);
nor U7763 (N_7763,N_6920,N_6682);
xor U7764 (N_7764,N_6964,N_6488);
and U7765 (N_7765,N_6186,N_6400);
or U7766 (N_7766,N_6572,N_6531);
nor U7767 (N_7767,N_6207,N_6785);
and U7768 (N_7768,N_6784,N_6258);
nor U7769 (N_7769,N_6820,N_6926);
or U7770 (N_7770,N_6972,N_6255);
or U7771 (N_7771,N_6877,N_6848);
and U7772 (N_7772,N_6041,N_6373);
xor U7773 (N_7773,N_6501,N_6951);
nand U7774 (N_7774,N_6856,N_6962);
or U7775 (N_7775,N_6375,N_6040);
or U7776 (N_7776,N_6137,N_6513);
xnor U7777 (N_7777,N_6478,N_6684);
or U7778 (N_7778,N_6272,N_6954);
nor U7779 (N_7779,N_6187,N_6704);
nand U7780 (N_7780,N_6725,N_6009);
nand U7781 (N_7781,N_6466,N_6717);
nor U7782 (N_7782,N_6536,N_6876);
and U7783 (N_7783,N_6376,N_6771);
and U7784 (N_7784,N_6224,N_6963);
xnor U7785 (N_7785,N_6147,N_6313);
nor U7786 (N_7786,N_6007,N_6589);
xor U7787 (N_7787,N_6760,N_6510);
nand U7788 (N_7788,N_6624,N_6878);
or U7789 (N_7789,N_6241,N_6058);
and U7790 (N_7790,N_6345,N_6925);
and U7791 (N_7791,N_6876,N_6547);
xor U7792 (N_7792,N_6953,N_6340);
and U7793 (N_7793,N_6990,N_6782);
or U7794 (N_7794,N_6582,N_6448);
or U7795 (N_7795,N_6837,N_6866);
or U7796 (N_7796,N_6511,N_6313);
nand U7797 (N_7797,N_6026,N_6494);
nand U7798 (N_7798,N_6419,N_6129);
xnor U7799 (N_7799,N_6581,N_6420);
xor U7800 (N_7800,N_6259,N_6850);
and U7801 (N_7801,N_6198,N_6372);
and U7802 (N_7802,N_6744,N_6179);
nor U7803 (N_7803,N_6640,N_6143);
xor U7804 (N_7804,N_6946,N_6890);
and U7805 (N_7805,N_6880,N_6600);
or U7806 (N_7806,N_6965,N_6977);
xor U7807 (N_7807,N_6424,N_6514);
or U7808 (N_7808,N_6661,N_6220);
nand U7809 (N_7809,N_6868,N_6640);
nor U7810 (N_7810,N_6451,N_6820);
or U7811 (N_7811,N_6556,N_6318);
xor U7812 (N_7812,N_6000,N_6201);
nand U7813 (N_7813,N_6199,N_6186);
nor U7814 (N_7814,N_6262,N_6464);
nand U7815 (N_7815,N_6189,N_6825);
and U7816 (N_7816,N_6562,N_6471);
and U7817 (N_7817,N_6846,N_6455);
xor U7818 (N_7818,N_6135,N_6508);
and U7819 (N_7819,N_6307,N_6161);
or U7820 (N_7820,N_6593,N_6949);
nand U7821 (N_7821,N_6967,N_6582);
and U7822 (N_7822,N_6410,N_6542);
xnor U7823 (N_7823,N_6885,N_6192);
nand U7824 (N_7824,N_6566,N_6153);
and U7825 (N_7825,N_6383,N_6698);
xor U7826 (N_7826,N_6064,N_6352);
or U7827 (N_7827,N_6941,N_6814);
nand U7828 (N_7828,N_6548,N_6748);
nor U7829 (N_7829,N_6266,N_6952);
and U7830 (N_7830,N_6132,N_6114);
nor U7831 (N_7831,N_6291,N_6503);
or U7832 (N_7832,N_6132,N_6511);
or U7833 (N_7833,N_6169,N_6796);
xor U7834 (N_7834,N_6408,N_6634);
or U7835 (N_7835,N_6057,N_6258);
or U7836 (N_7836,N_6672,N_6890);
and U7837 (N_7837,N_6927,N_6622);
xnor U7838 (N_7838,N_6098,N_6900);
xnor U7839 (N_7839,N_6316,N_6386);
and U7840 (N_7840,N_6534,N_6296);
and U7841 (N_7841,N_6655,N_6644);
or U7842 (N_7842,N_6962,N_6542);
nand U7843 (N_7843,N_6724,N_6936);
xor U7844 (N_7844,N_6447,N_6797);
and U7845 (N_7845,N_6896,N_6784);
and U7846 (N_7846,N_6510,N_6285);
or U7847 (N_7847,N_6146,N_6563);
or U7848 (N_7848,N_6359,N_6707);
or U7849 (N_7849,N_6341,N_6017);
nand U7850 (N_7850,N_6175,N_6108);
nand U7851 (N_7851,N_6956,N_6828);
or U7852 (N_7852,N_6210,N_6238);
nand U7853 (N_7853,N_6146,N_6575);
nand U7854 (N_7854,N_6213,N_6218);
xnor U7855 (N_7855,N_6879,N_6491);
nand U7856 (N_7856,N_6599,N_6262);
nor U7857 (N_7857,N_6153,N_6621);
nor U7858 (N_7858,N_6024,N_6438);
or U7859 (N_7859,N_6978,N_6630);
and U7860 (N_7860,N_6331,N_6475);
xnor U7861 (N_7861,N_6941,N_6514);
nor U7862 (N_7862,N_6256,N_6641);
xor U7863 (N_7863,N_6211,N_6653);
or U7864 (N_7864,N_6270,N_6052);
xnor U7865 (N_7865,N_6250,N_6785);
nand U7866 (N_7866,N_6482,N_6798);
nor U7867 (N_7867,N_6529,N_6744);
nand U7868 (N_7868,N_6901,N_6967);
or U7869 (N_7869,N_6110,N_6099);
and U7870 (N_7870,N_6562,N_6752);
nor U7871 (N_7871,N_6440,N_6926);
nand U7872 (N_7872,N_6566,N_6137);
xor U7873 (N_7873,N_6547,N_6497);
nand U7874 (N_7874,N_6561,N_6535);
nor U7875 (N_7875,N_6561,N_6637);
nand U7876 (N_7876,N_6563,N_6565);
or U7877 (N_7877,N_6893,N_6834);
or U7878 (N_7878,N_6517,N_6678);
nand U7879 (N_7879,N_6559,N_6187);
and U7880 (N_7880,N_6788,N_6500);
nand U7881 (N_7881,N_6059,N_6725);
xor U7882 (N_7882,N_6767,N_6058);
nor U7883 (N_7883,N_6363,N_6832);
nand U7884 (N_7884,N_6967,N_6665);
nand U7885 (N_7885,N_6815,N_6854);
or U7886 (N_7886,N_6758,N_6142);
or U7887 (N_7887,N_6680,N_6147);
and U7888 (N_7888,N_6999,N_6837);
xor U7889 (N_7889,N_6974,N_6656);
nand U7890 (N_7890,N_6505,N_6644);
nor U7891 (N_7891,N_6854,N_6991);
nand U7892 (N_7892,N_6803,N_6256);
nand U7893 (N_7893,N_6783,N_6917);
xnor U7894 (N_7894,N_6957,N_6748);
and U7895 (N_7895,N_6389,N_6023);
xor U7896 (N_7896,N_6863,N_6188);
and U7897 (N_7897,N_6335,N_6257);
nand U7898 (N_7898,N_6733,N_6214);
nand U7899 (N_7899,N_6121,N_6513);
nor U7900 (N_7900,N_6715,N_6457);
and U7901 (N_7901,N_6554,N_6042);
nand U7902 (N_7902,N_6047,N_6333);
xor U7903 (N_7903,N_6011,N_6908);
nand U7904 (N_7904,N_6633,N_6386);
or U7905 (N_7905,N_6517,N_6948);
nand U7906 (N_7906,N_6425,N_6437);
nand U7907 (N_7907,N_6567,N_6237);
nand U7908 (N_7908,N_6965,N_6752);
xnor U7909 (N_7909,N_6281,N_6421);
nand U7910 (N_7910,N_6510,N_6630);
and U7911 (N_7911,N_6236,N_6650);
nand U7912 (N_7912,N_6381,N_6368);
or U7913 (N_7913,N_6351,N_6492);
and U7914 (N_7914,N_6928,N_6745);
xnor U7915 (N_7915,N_6957,N_6250);
nand U7916 (N_7916,N_6262,N_6041);
xor U7917 (N_7917,N_6957,N_6381);
or U7918 (N_7918,N_6648,N_6325);
or U7919 (N_7919,N_6783,N_6344);
nand U7920 (N_7920,N_6042,N_6864);
nor U7921 (N_7921,N_6322,N_6590);
nor U7922 (N_7922,N_6484,N_6798);
nand U7923 (N_7923,N_6683,N_6480);
or U7924 (N_7924,N_6161,N_6640);
nor U7925 (N_7925,N_6621,N_6008);
xor U7926 (N_7926,N_6286,N_6507);
nor U7927 (N_7927,N_6001,N_6640);
and U7928 (N_7928,N_6721,N_6028);
and U7929 (N_7929,N_6998,N_6489);
nand U7930 (N_7930,N_6319,N_6670);
or U7931 (N_7931,N_6506,N_6174);
or U7932 (N_7932,N_6609,N_6629);
or U7933 (N_7933,N_6849,N_6455);
xnor U7934 (N_7934,N_6276,N_6571);
nand U7935 (N_7935,N_6781,N_6194);
or U7936 (N_7936,N_6152,N_6448);
nor U7937 (N_7937,N_6298,N_6763);
and U7938 (N_7938,N_6124,N_6948);
nand U7939 (N_7939,N_6840,N_6818);
and U7940 (N_7940,N_6180,N_6031);
and U7941 (N_7941,N_6876,N_6793);
nand U7942 (N_7942,N_6750,N_6333);
xor U7943 (N_7943,N_6657,N_6775);
nor U7944 (N_7944,N_6371,N_6731);
and U7945 (N_7945,N_6361,N_6188);
nor U7946 (N_7946,N_6551,N_6514);
or U7947 (N_7947,N_6781,N_6727);
nor U7948 (N_7948,N_6889,N_6347);
nor U7949 (N_7949,N_6078,N_6252);
or U7950 (N_7950,N_6316,N_6590);
or U7951 (N_7951,N_6482,N_6530);
nor U7952 (N_7952,N_6157,N_6706);
xor U7953 (N_7953,N_6781,N_6841);
nand U7954 (N_7954,N_6644,N_6319);
xor U7955 (N_7955,N_6599,N_6820);
nand U7956 (N_7956,N_6575,N_6579);
or U7957 (N_7957,N_6889,N_6661);
xnor U7958 (N_7958,N_6666,N_6780);
nand U7959 (N_7959,N_6804,N_6789);
and U7960 (N_7960,N_6244,N_6933);
nand U7961 (N_7961,N_6622,N_6740);
nand U7962 (N_7962,N_6598,N_6581);
nor U7963 (N_7963,N_6276,N_6138);
and U7964 (N_7964,N_6390,N_6557);
nor U7965 (N_7965,N_6190,N_6068);
nand U7966 (N_7966,N_6494,N_6330);
nor U7967 (N_7967,N_6612,N_6942);
or U7968 (N_7968,N_6929,N_6864);
xor U7969 (N_7969,N_6007,N_6260);
or U7970 (N_7970,N_6605,N_6271);
xor U7971 (N_7971,N_6839,N_6737);
or U7972 (N_7972,N_6611,N_6014);
nor U7973 (N_7973,N_6115,N_6497);
nand U7974 (N_7974,N_6684,N_6312);
xor U7975 (N_7975,N_6649,N_6677);
xnor U7976 (N_7976,N_6189,N_6673);
or U7977 (N_7977,N_6514,N_6129);
or U7978 (N_7978,N_6595,N_6497);
and U7979 (N_7979,N_6477,N_6478);
nand U7980 (N_7980,N_6428,N_6462);
or U7981 (N_7981,N_6167,N_6924);
nand U7982 (N_7982,N_6196,N_6081);
xnor U7983 (N_7983,N_6812,N_6250);
xnor U7984 (N_7984,N_6332,N_6402);
and U7985 (N_7985,N_6165,N_6362);
nand U7986 (N_7986,N_6099,N_6039);
xnor U7987 (N_7987,N_6285,N_6865);
and U7988 (N_7988,N_6224,N_6086);
nor U7989 (N_7989,N_6686,N_6534);
nor U7990 (N_7990,N_6355,N_6726);
and U7991 (N_7991,N_6730,N_6660);
nor U7992 (N_7992,N_6045,N_6952);
xnor U7993 (N_7993,N_6620,N_6327);
nor U7994 (N_7994,N_6855,N_6455);
and U7995 (N_7995,N_6456,N_6236);
xor U7996 (N_7996,N_6120,N_6207);
nand U7997 (N_7997,N_6781,N_6906);
xor U7998 (N_7998,N_6708,N_6734);
nand U7999 (N_7999,N_6390,N_6487);
nand U8000 (N_8000,N_7147,N_7861);
xnor U8001 (N_8001,N_7282,N_7600);
or U8002 (N_8002,N_7107,N_7416);
and U8003 (N_8003,N_7124,N_7409);
nand U8004 (N_8004,N_7126,N_7224);
or U8005 (N_8005,N_7621,N_7995);
or U8006 (N_8006,N_7618,N_7752);
nand U8007 (N_8007,N_7673,N_7211);
and U8008 (N_8008,N_7572,N_7963);
xor U8009 (N_8009,N_7472,N_7777);
xor U8010 (N_8010,N_7164,N_7766);
nand U8011 (N_8011,N_7907,N_7510);
and U8012 (N_8012,N_7095,N_7424);
nand U8013 (N_8013,N_7445,N_7437);
or U8014 (N_8014,N_7238,N_7976);
nand U8015 (N_8015,N_7143,N_7878);
and U8016 (N_8016,N_7674,N_7578);
and U8017 (N_8017,N_7084,N_7082);
and U8018 (N_8018,N_7473,N_7832);
xor U8019 (N_8019,N_7079,N_7257);
nand U8020 (N_8020,N_7531,N_7936);
or U8021 (N_8021,N_7867,N_7940);
nor U8022 (N_8022,N_7225,N_7688);
and U8023 (N_8023,N_7060,N_7313);
xor U8024 (N_8024,N_7213,N_7251);
and U8025 (N_8025,N_7876,N_7717);
nand U8026 (N_8026,N_7817,N_7194);
xor U8027 (N_8027,N_7722,N_7958);
nor U8028 (N_8028,N_7807,N_7274);
nand U8029 (N_8029,N_7675,N_7949);
nand U8030 (N_8030,N_7197,N_7347);
and U8031 (N_8031,N_7353,N_7410);
or U8032 (N_8032,N_7507,N_7430);
nor U8033 (N_8033,N_7522,N_7452);
xnor U8034 (N_8034,N_7054,N_7074);
xor U8035 (N_8035,N_7707,N_7318);
and U8036 (N_8036,N_7287,N_7567);
xnor U8037 (N_8037,N_7484,N_7778);
xnor U8038 (N_8038,N_7253,N_7063);
xnor U8039 (N_8039,N_7177,N_7924);
xnor U8040 (N_8040,N_7261,N_7072);
or U8041 (N_8041,N_7064,N_7818);
nor U8042 (N_8042,N_7889,N_7863);
xnor U8043 (N_8043,N_7358,N_7683);
nor U8044 (N_8044,N_7000,N_7456);
nor U8045 (N_8045,N_7679,N_7432);
or U8046 (N_8046,N_7880,N_7462);
and U8047 (N_8047,N_7773,N_7231);
nand U8048 (N_8048,N_7067,N_7560);
nand U8049 (N_8049,N_7024,N_7512);
nor U8050 (N_8050,N_7299,N_7178);
or U8051 (N_8051,N_7721,N_7202);
or U8052 (N_8052,N_7938,N_7041);
and U8053 (N_8053,N_7615,N_7801);
nor U8054 (N_8054,N_7302,N_7397);
nor U8055 (N_8055,N_7638,N_7737);
or U8056 (N_8056,N_7981,N_7919);
nand U8057 (N_8057,N_7341,N_7290);
and U8058 (N_8058,N_7874,N_7731);
or U8059 (N_8059,N_7839,N_7639);
nor U8060 (N_8060,N_7712,N_7451);
and U8061 (N_8061,N_7168,N_7622);
and U8062 (N_8062,N_7400,N_7393);
and U8063 (N_8063,N_7923,N_7463);
xnor U8064 (N_8064,N_7101,N_7086);
xnor U8065 (N_8065,N_7258,N_7118);
and U8066 (N_8066,N_7846,N_7561);
or U8067 (N_8067,N_7191,N_7285);
nand U8068 (N_8068,N_7853,N_7009);
and U8069 (N_8069,N_7031,N_7659);
or U8070 (N_8070,N_7726,N_7188);
nor U8071 (N_8071,N_7797,N_7189);
and U8072 (N_8072,N_7661,N_7080);
nand U8073 (N_8073,N_7687,N_7383);
or U8074 (N_8074,N_7127,N_7154);
nor U8075 (N_8075,N_7992,N_7155);
and U8076 (N_8076,N_7539,N_7325);
nand U8077 (N_8077,N_7911,N_7681);
nand U8078 (N_8078,N_7392,N_7888);
and U8079 (N_8079,N_7740,N_7957);
and U8080 (N_8080,N_7742,N_7983);
nand U8081 (N_8081,N_7803,N_7042);
nor U8082 (N_8082,N_7134,N_7511);
xnor U8083 (N_8083,N_7950,N_7401);
nand U8084 (N_8084,N_7623,N_7743);
xnor U8085 (N_8085,N_7331,N_7736);
nor U8086 (N_8086,N_7948,N_7152);
nor U8087 (N_8087,N_7144,N_7214);
xor U8088 (N_8088,N_7344,N_7799);
nand U8089 (N_8089,N_7279,N_7204);
and U8090 (N_8090,N_7866,N_7577);
xor U8091 (N_8091,N_7943,N_7075);
nand U8092 (N_8092,N_7402,N_7771);
xnor U8093 (N_8093,N_7720,N_7209);
and U8094 (N_8094,N_7944,N_7809);
nor U8095 (N_8095,N_7912,N_7482);
or U8096 (N_8096,N_7808,N_7614);
xor U8097 (N_8097,N_7269,N_7027);
nor U8098 (N_8098,N_7723,N_7488);
or U8099 (N_8099,N_7449,N_7881);
and U8100 (N_8100,N_7730,N_7763);
and U8101 (N_8101,N_7732,N_7230);
nand U8102 (N_8102,N_7148,N_7120);
xnor U8103 (N_8103,N_7094,N_7062);
or U8104 (N_8104,N_7423,N_7457);
nand U8105 (N_8105,N_7394,N_7046);
or U8106 (N_8106,N_7844,N_7099);
xnor U8107 (N_8107,N_7671,N_7527);
or U8108 (N_8108,N_7796,N_7317);
and U8109 (N_8109,N_7926,N_7904);
xor U8110 (N_8110,N_7403,N_7974);
nand U8111 (N_8111,N_7216,N_7085);
and U8112 (N_8112,N_7929,N_7444);
or U8113 (N_8113,N_7010,N_7529);
xor U8114 (N_8114,N_7083,N_7309);
or U8115 (N_8115,N_7635,N_7658);
and U8116 (N_8116,N_7055,N_7613);
and U8117 (N_8117,N_7634,N_7350);
nand U8118 (N_8118,N_7518,N_7192);
nor U8119 (N_8119,N_7422,N_7713);
and U8120 (N_8120,N_7965,N_7089);
and U8121 (N_8121,N_7336,N_7377);
nand U8122 (N_8122,N_7654,N_7665);
nand U8123 (N_8123,N_7185,N_7495);
nor U8124 (N_8124,N_7002,N_7479);
nor U8125 (N_8125,N_7369,N_7859);
or U8126 (N_8126,N_7921,N_7235);
and U8127 (N_8127,N_7241,N_7543);
and U8128 (N_8128,N_7714,N_7092);
or U8129 (N_8129,N_7110,N_7985);
or U8130 (N_8130,N_7745,N_7286);
and U8131 (N_8131,N_7343,N_7190);
xor U8132 (N_8132,N_7744,N_7619);
and U8133 (N_8133,N_7651,N_7153);
or U8134 (N_8134,N_7032,N_7415);
nor U8135 (N_8135,N_7770,N_7852);
and U8136 (N_8136,N_7215,N_7691);
xor U8137 (N_8137,N_7012,N_7052);
nand U8138 (N_8138,N_7509,N_7291);
or U8139 (N_8139,N_7583,N_7239);
xnor U8140 (N_8140,N_7454,N_7245);
nor U8141 (N_8141,N_7829,N_7709);
and U8142 (N_8142,N_7129,N_7895);
and U8143 (N_8143,N_7698,N_7990);
nor U8144 (N_8144,N_7066,N_7374);
xor U8145 (N_8145,N_7738,N_7301);
nand U8146 (N_8146,N_7334,N_7916);
nand U8147 (N_8147,N_7977,N_7340);
and U8148 (N_8148,N_7946,N_7151);
or U8149 (N_8149,N_7428,N_7708);
nor U8150 (N_8150,N_7648,N_7812);
and U8151 (N_8151,N_7856,N_7486);
nand U8152 (N_8152,N_7303,N_7324);
and U8153 (N_8153,N_7642,N_7956);
nand U8154 (N_8154,N_7953,N_7868);
nand U8155 (N_8155,N_7321,N_7264);
xor U8156 (N_8156,N_7232,N_7598);
or U8157 (N_8157,N_7588,N_7920);
or U8158 (N_8158,N_7203,N_7775);
and U8159 (N_8159,N_7696,N_7398);
nor U8160 (N_8160,N_7467,N_7487);
or U8161 (N_8161,N_7800,N_7972);
or U8162 (N_8162,N_7987,N_7597);
xor U8163 (N_8163,N_7112,N_7632);
and U8164 (N_8164,N_7033,N_7308);
nand U8165 (N_8165,N_7333,N_7991);
nor U8166 (N_8166,N_7186,N_7751);
or U8167 (N_8167,N_7364,N_7833);
nor U8168 (N_8168,N_7959,N_7806);
or U8169 (N_8169,N_7821,N_7975);
and U8170 (N_8170,N_7447,N_7813);
nand U8171 (N_8171,N_7898,N_7494);
nor U8172 (N_8172,N_7768,N_7469);
and U8173 (N_8173,N_7246,N_7076);
or U8174 (N_8174,N_7237,N_7128);
or U8175 (N_8175,N_7779,N_7755);
nand U8176 (N_8176,N_7969,N_7049);
and U8177 (N_8177,N_7592,N_7030);
nand U8178 (N_8178,N_7694,N_7565);
and U8179 (N_8179,N_7116,N_7657);
nand U8180 (N_8180,N_7701,N_7998);
nand U8181 (N_8181,N_7762,N_7882);
or U8182 (N_8182,N_7625,N_7090);
and U8183 (N_8183,N_7633,N_7865);
xnor U8184 (N_8184,N_7540,N_7058);
nor U8185 (N_8185,N_7794,N_7326);
nand U8186 (N_8186,N_7200,N_7157);
and U8187 (N_8187,N_7716,N_7073);
or U8188 (N_8188,N_7142,N_7133);
and U8189 (N_8189,N_7193,N_7875);
xor U8190 (N_8190,N_7906,N_7433);
nand U8191 (N_8191,N_7620,N_7414);
nor U8192 (N_8192,N_7014,N_7320);
xor U8193 (N_8193,N_7373,N_7908);
and U8194 (N_8194,N_7071,N_7163);
nand U8195 (N_8195,N_7585,N_7700);
or U8196 (N_8196,N_7589,N_7001);
xor U8197 (N_8197,N_7259,N_7551);
xnor U8198 (N_8198,N_7695,N_7478);
nand U8199 (N_8199,N_7396,N_7418);
xor U8200 (N_8200,N_7439,N_7604);
and U8201 (N_8201,N_7984,N_7108);
nor U8202 (N_8202,N_7043,N_7175);
xor U8203 (N_8203,N_7660,N_7069);
nand U8204 (N_8204,N_7728,N_7004);
xor U8205 (N_8205,N_7506,N_7897);
or U8206 (N_8206,N_7363,N_7294);
nand U8207 (N_8207,N_7616,N_7431);
and U8208 (N_8208,N_7901,N_7823);
or U8209 (N_8209,N_7917,N_7986);
and U8210 (N_8210,N_7774,N_7146);
or U8211 (N_8211,N_7173,N_7420);
or U8212 (N_8212,N_7162,N_7425);
nor U8213 (N_8213,N_7220,N_7886);
and U8214 (N_8214,N_7212,N_7640);
and U8215 (N_8215,N_7117,N_7464);
or U8216 (N_8216,N_7339,N_7316);
nand U8217 (N_8217,N_7769,N_7370);
or U8218 (N_8218,N_7195,N_7485);
or U8219 (N_8219,N_7971,N_7169);
nor U8220 (N_8220,N_7574,N_7161);
or U8221 (N_8221,N_7524,N_7367);
nor U8222 (N_8222,N_7968,N_7349);
nand U8223 (N_8223,N_7421,N_7593);
nor U8224 (N_8224,N_7413,N_7692);
nor U8225 (N_8225,N_7606,N_7646);
and U8226 (N_8226,N_7820,N_7980);
and U8227 (N_8227,N_7300,N_7653);
or U8228 (N_8228,N_7182,N_7450);
and U8229 (N_8229,N_7902,N_7571);
xnor U8230 (N_8230,N_7749,N_7180);
nand U8231 (N_8231,N_7525,N_7405);
and U8232 (N_8232,N_7670,N_7504);
nand U8233 (N_8233,N_7103,N_7379);
nand U8234 (N_8234,N_7429,N_7480);
or U8235 (N_8235,N_7375,N_7997);
nor U8236 (N_8236,N_7492,N_7140);
or U8237 (N_8237,N_7244,N_7711);
and U8238 (N_8238,N_7952,N_7523);
xnor U8239 (N_8239,N_7727,N_7669);
xnor U8240 (N_8240,N_7008,N_7758);
nor U8241 (N_8241,N_7909,N_7475);
nand U8242 (N_8242,N_7955,N_7227);
nand U8243 (N_8243,N_7121,N_7057);
nand U8244 (N_8244,N_7263,N_7434);
nand U8245 (N_8245,N_7158,N_7939);
xnor U8246 (N_8246,N_7704,N_7159);
nor U8247 (N_8247,N_7252,N_7647);
nand U8248 (N_8248,N_7575,N_7276);
nand U8249 (N_8249,N_7855,N_7724);
or U8250 (N_8250,N_7372,N_7217);
and U8251 (N_8251,N_7044,N_7526);
nor U8252 (N_8252,N_7787,N_7490);
or U8253 (N_8253,N_7021,N_7885);
nand U8254 (N_8254,N_7590,N_7077);
or U8255 (N_8255,N_7022,N_7115);
xnor U8256 (N_8256,N_7003,N_7656);
or U8257 (N_8257,N_7840,N_7254);
xor U8258 (N_8258,N_7275,N_7061);
and U8259 (N_8259,N_7236,N_7877);
and U8260 (N_8260,N_7627,N_7649);
or U8261 (N_8261,N_7547,N_7130);
nand U8262 (N_8262,N_7139,N_7699);
nor U8263 (N_8263,N_7160,N_7546);
nor U8264 (N_8264,N_7862,N_7378);
xor U8265 (N_8265,N_7453,N_7757);
xor U8266 (N_8266,N_7608,N_7441);
xor U8267 (N_8267,N_7739,N_7240);
or U8268 (N_8268,N_7825,N_7248);
nand U8269 (N_8269,N_7038,N_7382);
or U8270 (N_8270,N_7172,N_7229);
nand U8271 (N_8271,N_7491,N_7366);
nor U8272 (N_8272,N_7964,N_7930);
or U8273 (N_8273,N_7489,N_7978);
nand U8274 (N_8274,N_7636,N_7208);
and U8275 (N_8275,N_7284,N_7360);
or U8276 (N_8276,N_7942,N_7555);
nand U8277 (N_8277,N_7776,N_7903);
nand U8278 (N_8278,N_7481,N_7804);
or U8279 (N_8279,N_7689,N_7498);
nand U8280 (N_8280,N_7493,N_7270);
nor U8281 (N_8281,N_7497,N_7470);
or U8282 (N_8282,N_7748,N_7884);
nor U8283 (N_8283,N_7747,N_7932);
xor U8284 (N_8284,N_7690,N_7267);
and U8285 (N_8285,N_7156,N_7788);
nor U8286 (N_8286,N_7871,N_7772);
or U8287 (N_8287,N_7918,N_7179);
and U8288 (N_8288,N_7205,N_7780);
nand U8289 (N_8289,N_7365,N_7947);
nand U8290 (N_8290,N_7563,N_7548);
xnor U8291 (N_8291,N_7684,N_7584);
or U8292 (N_8292,N_7686,N_7097);
nand U8293 (N_8293,N_7537,N_7719);
and U8294 (N_8294,N_7322,N_7315);
nor U8295 (N_8295,N_7328,N_7521);
or U8296 (N_8296,N_7337,N_7011);
xnor U8297 (N_8297,N_7219,N_7676);
nand U8298 (N_8298,N_7234,N_7273);
xnor U8299 (N_8299,N_7078,N_7292);
and U8300 (N_8300,N_7680,N_7811);
xor U8301 (N_8301,N_7532,N_7138);
and U8302 (N_8302,N_7296,N_7581);
and U8303 (N_8303,N_7982,N_7357);
xor U8304 (N_8304,N_7017,N_7123);
and U8305 (N_8305,N_7937,N_7994);
xor U8306 (N_8306,N_7715,N_7725);
nand U8307 (N_8307,N_7544,N_7386);
xor U8308 (N_8308,N_7280,N_7734);
or U8309 (N_8309,N_7650,N_7081);
nand U8310 (N_8310,N_7858,N_7198);
and U8311 (N_8311,N_7132,N_7048);
or U8312 (N_8312,N_7517,N_7376);
nor U8313 (N_8313,N_7233,N_7816);
and U8314 (N_8314,N_7915,N_7999);
or U8315 (N_8315,N_7104,N_7387);
and U8316 (N_8316,N_7102,N_7354);
nand U8317 (N_8317,N_7570,N_7388);
nand U8318 (N_8318,N_7568,N_7542);
or U8319 (N_8319,N_7093,N_7760);
or U8320 (N_8320,N_7471,N_7528);
nand U8321 (N_8321,N_7834,N_7652);
nand U8322 (N_8322,N_7533,N_7283);
xor U8323 (N_8323,N_7256,N_7289);
or U8324 (N_8324,N_7566,N_7474);
or U8325 (N_8325,N_7925,N_7399);
or U8326 (N_8326,N_7789,N_7281);
or U8327 (N_8327,N_7136,N_7891);
or U8328 (N_8328,N_7013,N_7458);
nor U8329 (N_8329,N_7247,N_7890);
nand U8330 (N_8330,N_7557,N_7672);
and U8331 (N_8331,N_7838,N_7556);
or U8332 (N_8332,N_7666,N_7814);
nand U8333 (N_8333,N_7206,N_7065);
nor U8334 (N_8334,N_7174,N_7166);
nor U8335 (N_8335,N_7607,N_7352);
nand U8336 (N_8336,N_7602,N_7667);
nor U8337 (N_8337,N_7199,N_7795);
nand U8338 (N_8338,N_7595,N_7201);
nor U8339 (N_8339,N_7662,N_7643);
xnor U8340 (N_8340,N_7710,N_7966);
xnor U8341 (N_8341,N_7020,N_7831);
nor U8342 (N_8342,N_7345,N_7056);
and U8343 (N_8343,N_7266,N_7631);
nor U8344 (N_8344,N_7466,N_7609);
nand U8345 (N_8345,N_7872,N_7626);
or U8346 (N_8346,N_7242,N_7305);
nor U8347 (N_8347,N_7016,N_7552);
and U8348 (N_8348,N_7187,N_7860);
nand U8349 (N_8349,N_7426,N_7149);
nor U8350 (N_8350,N_7945,N_7873);
or U8351 (N_8351,N_7312,N_7226);
or U8352 (N_8352,N_7176,N_7693);
and U8353 (N_8353,N_7845,N_7167);
or U8354 (N_8354,N_7591,N_7135);
xnor U8355 (N_8355,N_7798,N_7573);
xor U8356 (N_8356,N_7419,N_7905);
nand U8357 (N_8357,N_7356,N_7603);
or U8358 (N_8358,N_7535,N_7288);
nand U8359 (N_8359,N_7465,N_7790);
nand U8360 (N_8360,N_7023,N_7554);
and U8361 (N_8361,N_7477,N_7348);
xnor U8362 (N_8362,N_7131,N_7541);
or U8363 (N_8363,N_7951,N_7849);
nand U8364 (N_8364,N_7989,N_7307);
or U8365 (N_8365,N_7436,N_7756);
nor U8366 (N_8366,N_7781,N_7822);
nand U8367 (N_8367,N_7265,N_7828);
xnor U8368 (N_8368,N_7207,N_7501);
or U8369 (N_8369,N_7842,N_7059);
nand U8370 (N_8370,N_7096,N_7141);
or U8371 (N_8371,N_7594,N_7767);
and U8372 (N_8372,N_7703,N_7848);
nand U8373 (N_8373,N_7854,N_7610);
nand U8374 (N_8374,N_7782,N_7934);
nor U8375 (N_8375,N_7784,N_7268);
or U8376 (N_8376,N_7505,N_7677);
nor U8377 (N_8377,N_7922,N_7534);
xnor U8378 (N_8378,N_7754,N_7508);
xnor U8379 (N_8379,N_7304,N_7819);
xor U8380 (N_8380,N_7050,N_7408);
nand U8381 (N_8381,N_7165,N_7028);
nor U8382 (N_8382,N_7815,N_7841);
or U8383 (N_8383,N_7183,N_7034);
xor U8384 (N_8384,N_7483,N_7323);
and U8385 (N_8385,N_7617,N_7630);
nand U8386 (N_8386,N_7655,N_7900);
xor U8387 (N_8387,N_7440,N_7025);
xnor U8388 (N_8388,N_7850,N_7894);
and U8389 (N_8389,N_7298,N_7390);
and U8390 (N_8390,N_7810,N_7601);
and U8391 (N_8391,N_7996,N_7791);
xnor U8392 (N_8392,N_7786,N_7122);
nand U8393 (N_8393,N_7765,N_7870);
or U8394 (N_8394,N_7805,N_7330);
xnor U8395 (N_8395,N_7438,N_7582);
xor U8396 (N_8396,N_7836,N_7411);
or U8397 (N_8397,N_7362,N_7035);
nand U8398 (N_8398,N_7664,N_7928);
and U8399 (N_8399,N_7380,N_7218);
or U8400 (N_8400,N_7500,N_7586);
xor U8401 (N_8401,N_7476,N_7255);
nor U8402 (N_8402,N_7053,N_7015);
or U8403 (N_8403,N_7029,N_7697);
xor U8404 (N_8404,N_7558,N_7857);
nand U8405 (N_8405,N_7896,N_7040);
or U8406 (N_8406,N_7037,N_7329);
and U8407 (N_8407,N_7406,N_7047);
and U8408 (N_8408,N_7931,N_7459);
nor U8409 (N_8409,N_7297,N_7802);
and U8410 (N_8410,N_7611,N_7468);
nand U8411 (N_8411,N_7222,N_7106);
nor U8412 (N_8412,N_7088,N_7549);
xnor U8413 (N_8413,N_7612,N_7105);
and U8414 (N_8414,N_7914,N_7579);
or U8415 (N_8415,N_7068,N_7513);
xor U8416 (N_8416,N_7087,N_7039);
nand U8417 (N_8417,N_7249,N_7962);
nor U8418 (N_8418,N_7407,N_7051);
nor U8419 (N_8419,N_7170,N_7368);
nor U8420 (N_8420,N_7927,N_7272);
or U8421 (N_8421,N_7070,N_7442);
xnor U8422 (N_8422,N_7883,N_7536);
nor U8423 (N_8423,N_7278,N_7530);
nand U8424 (N_8424,N_7435,N_7006);
or U8425 (N_8425,N_7210,N_7830);
xnor U8426 (N_8426,N_7792,N_7913);
nor U8427 (N_8427,N_7783,N_7113);
xnor U8428 (N_8428,N_7385,N_7843);
or U8429 (N_8429,N_7718,N_7091);
nor U8430 (N_8430,N_7935,N_7007);
nor U8431 (N_8431,N_7005,N_7538);
nand U8432 (N_8432,N_7851,N_7705);
xor U8433 (N_8433,N_7346,N_7682);
nand U8434 (N_8434,N_7970,N_7384);
xor U8435 (N_8435,N_7306,N_7759);
nand U8436 (N_8436,N_7559,N_7520);
nand U8437 (N_8437,N_7446,N_7260);
or U8438 (N_8438,N_7553,N_7184);
xnor U8439 (N_8439,N_7824,N_7026);
xor U8440 (N_8440,N_7395,N_7599);
xnor U8441 (N_8441,N_7564,N_7150);
nand U8442 (N_8442,N_7271,N_7644);
nor U8443 (N_8443,N_7496,N_7761);
nand U8444 (N_8444,N_7637,N_7746);
nor U8445 (N_8445,N_7645,N_7685);
nor U8446 (N_8446,N_7355,N_7277);
nor U8447 (N_8447,N_7837,N_7018);
or U8448 (N_8448,N_7111,N_7295);
nor U8449 (N_8449,N_7893,N_7733);
nor U8450 (N_8450,N_7351,N_7335);
nand U8451 (N_8451,N_7338,N_7181);
xor U8452 (N_8452,N_7221,N_7741);
nand U8453 (N_8453,N_7826,N_7847);
xor U8454 (N_8454,N_7404,N_7391);
or U8455 (N_8455,N_7448,N_7332);
xor U8456 (N_8456,N_7735,N_7311);
xnor U8457 (N_8457,N_7036,N_7993);
nand U8458 (N_8458,N_7359,N_7514);
or U8459 (N_8459,N_7460,N_7461);
and U8460 (N_8460,N_7519,N_7381);
or U8461 (N_8461,N_7145,N_7764);
nor U8462 (N_8462,N_7933,N_7979);
xor U8463 (N_8463,N_7417,N_7785);
and U8464 (N_8464,N_7098,N_7550);
and U8465 (N_8465,N_7628,N_7753);
nor U8466 (N_8466,N_7596,N_7605);
xnor U8467 (N_8467,N_7125,N_7389);
or U8468 (N_8468,N_7171,N_7100);
or U8469 (N_8469,N_7910,N_7887);
and U8470 (N_8470,N_7954,N_7502);
or U8471 (N_8471,N_7293,N_7706);
and U8472 (N_8472,N_7702,N_7892);
nor U8473 (N_8473,N_7443,N_7668);
nor U8474 (N_8474,N_7678,N_7427);
or U8475 (N_8475,N_7864,N_7342);
xor U8476 (N_8476,N_7624,N_7988);
nor U8477 (N_8477,N_7663,N_7114);
or U8478 (N_8478,N_7045,N_7973);
and U8479 (N_8479,N_7729,N_7899);
or U8480 (N_8480,N_7371,N_7119);
xnor U8481 (N_8481,N_7243,N_7869);
nor U8482 (N_8482,N_7827,N_7109);
nand U8483 (N_8483,N_7562,N_7516);
or U8484 (N_8484,N_7941,N_7750);
nand U8485 (N_8485,N_7793,N_7545);
nand U8486 (N_8486,N_7961,N_7580);
and U8487 (N_8487,N_7262,N_7569);
xor U8488 (N_8488,N_7960,N_7499);
or U8489 (N_8489,N_7327,N_7310);
or U8490 (N_8490,N_7319,N_7629);
nand U8491 (N_8491,N_7879,N_7967);
or U8492 (N_8492,N_7361,N_7019);
or U8493 (N_8493,N_7137,N_7412);
and U8494 (N_8494,N_7250,N_7196);
nand U8495 (N_8495,N_7223,N_7228);
nand U8496 (N_8496,N_7641,N_7835);
nor U8497 (N_8497,N_7587,N_7455);
and U8498 (N_8498,N_7314,N_7576);
and U8499 (N_8499,N_7503,N_7515);
nand U8500 (N_8500,N_7223,N_7311);
and U8501 (N_8501,N_7701,N_7103);
xnor U8502 (N_8502,N_7865,N_7657);
nor U8503 (N_8503,N_7673,N_7953);
or U8504 (N_8504,N_7157,N_7645);
and U8505 (N_8505,N_7983,N_7147);
and U8506 (N_8506,N_7156,N_7543);
xor U8507 (N_8507,N_7075,N_7335);
and U8508 (N_8508,N_7152,N_7905);
xnor U8509 (N_8509,N_7228,N_7426);
and U8510 (N_8510,N_7431,N_7177);
or U8511 (N_8511,N_7410,N_7136);
or U8512 (N_8512,N_7903,N_7328);
nand U8513 (N_8513,N_7195,N_7514);
nor U8514 (N_8514,N_7640,N_7606);
or U8515 (N_8515,N_7127,N_7247);
xor U8516 (N_8516,N_7905,N_7039);
or U8517 (N_8517,N_7640,N_7129);
nor U8518 (N_8518,N_7057,N_7315);
nor U8519 (N_8519,N_7647,N_7445);
nor U8520 (N_8520,N_7284,N_7338);
xor U8521 (N_8521,N_7350,N_7198);
nor U8522 (N_8522,N_7569,N_7895);
nor U8523 (N_8523,N_7945,N_7329);
or U8524 (N_8524,N_7669,N_7400);
nor U8525 (N_8525,N_7384,N_7958);
nand U8526 (N_8526,N_7382,N_7001);
or U8527 (N_8527,N_7628,N_7691);
nand U8528 (N_8528,N_7302,N_7587);
nand U8529 (N_8529,N_7815,N_7311);
nor U8530 (N_8530,N_7842,N_7180);
or U8531 (N_8531,N_7234,N_7867);
nor U8532 (N_8532,N_7032,N_7927);
nor U8533 (N_8533,N_7458,N_7910);
and U8534 (N_8534,N_7922,N_7011);
or U8535 (N_8535,N_7999,N_7950);
nand U8536 (N_8536,N_7749,N_7966);
or U8537 (N_8537,N_7054,N_7130);
nand U8538 (N_8538,N_7438,N_7703);
or U8539 (N_8539,N_7981,N_7929);
or U8540 (N_8540,N_7584,N_7901);
and U8541 (N_8541,N_7832,N_7468);
xor U8542 (N_8542,N_7314,N_7251);
or U8543 (N_8543,N_7744,N_7476);
nor U8544 (N_8544,N_7118,N_7767);
and U8545 (N_8545,N_7714,N_7268);
and U8546 (N_8546,N_7531,N_7872);
and U8547 (N_8547,N_7892,N_7303);
nor U8548 (N_8548,N_7689,N_7735);
nand U8549 (N_8549,N_7576,N_7646);
nand U8550 (N_8550,N_7434,N_7843);
or U8551 (N_8551,N_7012,N_7533);
or U8552 (N_8552,N_7349,N_7974);
and U8553 (N_8553,N_7153,N_7414);
nand U8554 (N_8554,N_7659,N_7384);
xor U8555 (N_8555,N_7161,N_7424);
or U8556 (N_8556,N_7842,N_7110);
xor U8557 (N_8557,N_7108,N_7324);
nand U8558 (N_8558,N_7527,N_7930);
and U8559 (N_8559,N_7943,N_7700);
xor U8560 (N_8560,N_7747,N_7715);
nand U8561 (N_8561,N_7602,N_7651);
or U8562 (N_8562,N_7442,N_7183);
nor U8563 (N_8563,N_7219,N_7063);
nor U8564 (N_8564,N_7557,N_7937);
xnor U8565 (N_8565,N_7469,N_7460);
nor U8566 (N_8566,N_7476,N_7241);
xor U8567 (N_8567,N_7943,N_7616);
or U8568 (N_8568,N_7422,N_7706);
nand U8569 (N_8569,N_7018,N_7740);
or U8570 (N_8570,N_7657,N_7578);
nand U8571 (N_8571,N_7908,N_7759);
xnor U8572 (N_8572,N_7895,N_7726);
xor U8573 (N_8573,N_7285,N_7624);
xnor U8574 (N_8574,N_7137,N_7804);
or U8575 (N_8575,N_7637,N_7337);
or U8576 (N_8576,N_7962,N_7905);
and U8577 (N_8577,N_7548,N_7658);
or U8578 (N_8578,N_7405,N_7692);
nor U8579 (N_8579,N_7842,N_7078);
nand U8580 (N_8580,N_7754,N_7465);
or U8581 (N_8581,N_7871,N_7771);
xnor U8582 (N_8582,N_7784,N_7092);
nand U8583 (N_8583,N_7949,N_7792);
nand U8584 (N_8584,N_7778,N_7220);
and U8585 (N_8585,N_7387,N_7436);
xnor U8586 (N_8586,N_7154,N_7909);
and U8587 (N_8587,N_7253,N_7537);
nor U8588 (N_8588,N_7744,N_7445);
nand U8589 (N_8589,N_7862,N_7443);
and U8590 (N_8590,N_7731,N_7930);
xor U8591 (N_8591,N_7885,N_7572);
or U8592 (N_8592,N_7075,N_7565);
nand U8593 (N_8593,N_7147,N_7411);
and U8594 (N_8594,N_7557,N_7709);
nor U8595 (N_8595,N_7465,N_7771);
xnor U8596 (N_8596,N_7205,N_7528);
xor U8597 (N_8597,N_7221,N_7688);
xor U8598 (N_8598,N_7106,N_7954);
and U8599 (N_8599,N_7196,N_7784);
xor U8600 (N_8600,N_7011,N_7620);
xor U8601 (N_8601,N_7981,N_7850);
and U8602 (N_8602,N_7711,N_7275);
or U8603 (N_8603,N_7738,N_7586);
and U8604 (N_8604,N_7041,N_7716);
nor U8605 (N_8605,N_7453,N_7139);
and U8606 (N_8606,N_7693,N_7961);
and U8607 (N_8607,N_7277,N_7866);
and U8608 (N_8608,N_7211,N_7048);
nor U8609 (N_8609,N_7936,N_7370);
and U8610 (N_8610,N_7993,N_7922);
or U8611 (N_8611,N_7717,N_7671);
xnor U8612 (N_8612,N_7565,N_7166);
xor U8613 (N_8613,N_7480,N_7833);
xnor U8614 (N_8614,N_7833,N_7535);
or U8615 (N_8615,N_7267,N_7947);
xnor U8616 (N_8616,N_7487,N_7728);
xor U8617 (N_8617,N_7055,N_7323);
nor U8618 (N_8618,N_7904,N_7751);
xnor U8619 (N_8619,N_7370,N_7330);
or U8620 (N_8620,N_7599,N_7941);
and U8621 (N_8621,N_7001,N_7614);
xnor U8622 (N_8622,N_7858,N_7261);
or U8623 (N_8623,N_7169,N_7473);
or U8624 (N_8624,N_7217,N_7232);
xor U8625 (N_8625,N_7049,N_7099);
nand U8626 (N_8626,N_7862,N_7136);
xnor U8627 (N_8627,N_7479,N_7347);
or U8628 (N_8628,N_7175,N_7111);
nand U8629 (N_8629,N_7158,N_7314);
and U8630 (N_8630,N_7548,N_7315);
nor U8631 (N_8631,N_7095,N_7438);
nand U8632 (N_8632,N_7646,N_7666);
nor U8633 (N_8633,N_7982,N_7442);
nand U8634 (N_8634,N_7273,N_7473);
nor U8635 (N_8635,N_7287,N_7945);
nand U8636 (N_8636,N_7844,N_7500);
or U8637 (N_8637,N_7834,N_7699);
nor U8638 (N_8638,N_7387,N_7566);
xor U8639 (N_8639,N_7220,N_7550);
nor U8640 (N_8640,N_7451,N_7508);
xor U8641 (N_8641,N_7578,N_7666);
nand U8642 (N_8642,N_7949,N_7547);
or U8643 (N_8643,N_7826,N_7422);
nor U8644 (N_8644,N_7509,N_7749);
and U8645 (N_8645,N_7250,N_7816);
nand U8646 (N_8646,N_7823,N_7440);
or U8647 (N_8647,N_7764,N_7565);
xnor U8648 (N_8648,N_7820,N_7365);
nand U8649 (N_8649,N_7084,N_7658);
nand U8650 (N_8650,N_7823,N_7610);
nand U8651 (N_8651,N_7605,N_7135);
xnor U8652 (N_8652,N_7994,N_7047);
nor U8653 (N_8653,N_7698,N_7991);
nor U8654 (N_8654,N_7998,N_7069);
or U8655 (N_8655,N_7618,N_7443);
and U8656 (N_8656,N_7250,N_7476);
nor U8657 (N_8657,N_7485,N_7204);
or U8658 (N_8658,N_7348,N_7196);
and U8659 (N_8659,N_7496,N_7611);
or U8660 (N_8660,N_7363,N_7743);
nand U8661 (N_8661,N_7718,N_7685);
and U8662 (N_8662,N_7875,N_7367);
nor U8663 (N_8663,N_7773,N_7149);
xor U8664 (N_8664,N_7263,N_7800);
and U8665 (N_8665,N_7016,N_7098);
or U8666 (N_8666,N_7029,N_7231);
or U8667 (N_8667,N_7064,N_7221);
and U8668 (N_8668,N_7041,N_7873);
nand U8669 (N_8669,N_7920,N_7638);
nor U8670 (N_8670,N_7966,N_7612);
xnor U8671 (N_8671,N_7655,N_7184);
nor U8672 (N_8672,N_7484,N_7603);
xor U8673 (N_8673,N_7253,N_7698);
nand U8674 (N_8674,N_7947,N_7721);
and U8675 (N_8675,N_7205,N_7689);
and U8676 (N_8676,N_7741,N_7797);
xor U8677 (N_8677,N_7059,N_7677);
xor U8678 (N_8678,N_7745,N_7518);
nor U8679 (N_8679,N_7821,N_7593);
xor U8680 (N_8680,N_7276,N_7567);
and U8681 (N_8681,N_7042,N_7253);
or U8682 (N_8682,N_7842,N_7255);
nand U8683 (N_8683,N_7018,N_7797);
or U8684 (N_8684,N_7763,N_7614);
or U8685 (N_8685,N_7674,N_7671);
and U8686 (N_8686,N_7589,N_7407);
nand U8687 (N_8687,N_7258,N_7911);
or U8688 (N_8688,N_7545,N_7933);
xnor U8689 (N_8689,N_7004,N_7587);
nor U8690 (N_8690,N_7985,N_7658);
nor U8691 (N_8691,N_7675,N_7138);
or U8692 (N_8692,N_7935,N_7723);
or U8693 (N_8693,N_7558,N_7646);
and U8694 (N_8694,N_7440,N_7405);
nand U8695 (N_8695,N_7269,N_7002);
and U8696 (N_8696,N_7031,N_7205);
and U8697 (N_8697,N_7878,N_7047);
nor U8698 (N_8698,N_7497,N_7029);
nor U8699 (N_8699,N_7580,N_7898);
xor U8700 (N_8700,N_7243,N_7943);
xor U8701 (N_8701,N_7864,N_7558);
or U8702 (N_8702,N_7297,N_7288);
or U8703 (N_8703,N_7208,N_7722);
xor U8704 (N_8704,N_7766,N_7439);
or U8705 (N_8705,N_7944,N_7920);
or U8706 (N_8706,N_7243,N_7667);
xor U8707 (N_8707,N_7991,N_7347);
xnor U8708 (N_8708,N_7511,N_7391);
nor U8709 (N_8709,N_7529,N_7867);
or U8710 (N_8710,N_7522,N_7787);
or U8711 (N_8711,N_7313,N_7301);
or U8712 (N_8712,N_7802,N_7847);
xnor U8713 (N_8713,N_7870,N_7052);
and U8714 (N_8714,N_7056,N_7779);
and U8715 (N_8715,N_7705,N_7378);
or U8716 (N_8716,N_7609,N_7248);
and U8717 (N_8717,N_7993,N_7341);
or U8718 (N_8718,N_7000,N_7046);
nor U8719 (N_8719,N_7359,N_7509);
and U8720 (N_8720,N_7980,N_7572);
nand U8721 (N_8721,N_7686,N_7328);
xnor U8722 (N_8722,N_7796,N_7472);
or U8723 (N_8723,N_7609,N_7699);
and U8724 (N_8724,N_7458,N_7489);
xor U8725 (N_8725,N_7711,N_7170);
nor U8726 (N_8726,N_7779,N_7115);
xnor U8727 (N_8727,N_7851,N_7876);
or U8728 (N_8728,N_7491,N_7768);
and U8729 (N_8729,N_7879,N_7788);
nand U8730 (N_8730,N_7904,N_7026);
xor U8731 (N_8731,N_7035,N_7280);
and U8732 (N_8732,N_7004,N_7749);
or U8733 (N_8733,N_7702,N_7744);
nand U8734 (N_8734,N_7054,N_7224);
nand U8735 (N_8735,N_7250,N_7644);
nand U8736 (N_8736,N_7827,N_7337);
xnor U8737 (N_8737,N_7521,N_7028);
xor U8738 (N_8738,N_7137,N_7288);
xor U8739 (N_8739,N_7063,N_7166);
or U8740 (N_8740,N_7594,N_7096);
and U8741 (N_8741,N_7750,N_7543);
nand U8742 (N_8742,N_7859,N_7622);
and U8743 (N_8743,N_7805,N_7212);
nor U8744 (N_8744,N_7427,N_7384);
xor U8745 (N_8745,N_7747,N_7858);
nand U8746 (N_8746,N_7628,N_7424);
and U8747 (N_8747,N_7506,N_7284);
and U8748 (N_8748,N_7111,N_7272);
nor U8749 (N_8749,N_7093,N_7015);
nor U8750 (N_8750,N_7524,N_7646);
nor U8751 (N_8751,N_7176,N_7547);
and U8752 (N_8752,N_7741,N_7342);
xor U8753 (N_8753,N_7749,N_7859);
xor U8754 (N_8754,N_7936,N_7283);
nor U8755 (N_8755,N_7025,N_7554);
and U8756 (N_8756,N_7581,N_7914);
and U8757 (N_8757,N_7374,N_7307);
and U8758 (N_8758,N_7333,N_7565);
or U8759 (N_8759,N_7815,N_7073);
and U8760 (N_8760,N_7807,N_7270);
or U8761 (N_8761,N_7659,N_7468);
or U8762 (N_8762,N_7517,N_7388);
xnor U8763 (N_8763,N_7046,N_7461);
and U8764 (N_8764,N_7364,N_7018);
or U8765 (N_8765,N_7075,N_7454);
nor U8766 (N_8766,N_7936,N_7960);
or U8767 (N_8767,N_7431,N_7887);
nand U8768 (N_8768,N_7417,N_7423);
xor U8769 (N_8769,N_7811,N_7304);
or U8770 (N_8770,N_7984,N_7829);
nand U8771 (N_8771,N_7290,N_7242);
nor U8772 (N_8772,N_7510,N_7188);
nor U8773 (N_8773,N_7406,N_7396);
or U8774 (N_8774,N_7783,N_7256);
or U8775 (N_8775,N_7652,N_7585);
or U8776 (N_8776,N_7451,N_7749);
nand U8777 (N_8777,N_7978,N_7677);
xor U8778 (N_8778,N_7686,N_7651);
nor U8779 (N_8779,N_7997,N_7393);
or U8780 (N_8780,N_7184,N_7303);
nand U8781 (N_8781,N_7492,N_7293);
nand U8782 (N_8782,N_7615,N_7673);
and U8783 (N_8783,N_7069,N_7945);
and U8784 (N_8784,N_7689,N_7244);
and U8785 (N_8785,N_7061,N_7449);
xnor U8786 (N_8786,N_7303,N_7215);
xor U8787 (N_8787,N_7077,N_7857);
xor U8788 (N_8788,N_7143,N_7184);
nand U8789 (N_8789,N_7281,N_7204);
nand U8790 (N_8790,N_7788,N_7824);
nand U8791 (N_8791,N_7126,N_7112);
or U8792 (N_8792,N_7686,N_7756);
xor U8793 (N_8793,N_7367,N_7622);
nand U8794 (N_8794,N_7232,N_7810);
and U8795 (N_8795,N_7168,N_7687);
nand U8796 (N_8796,N_7918,N_7801);
nand U8797 (N_8797,N_7414,N_7614);
nor U8798 (N_8798,N_7589,N_7440);
or U8799 (N_8799,N_7853,N_7386);
xnor U8800 (N_8800,N_7365,N_7199);
or U8801 (N_8801,N_7268,N_7351);
nor U8802 (N_8802,N_7818,N_7065);
nand U8803 (N_8803,N_7871,N_7004);
nor U8804 (N_8804,N_7119,N_7256);
or U8805 (N_8805,N_7490,N_7100);
nor U8806 (N_8806,N_7360,N_7268);
and U8807 (N_8807,N_7653,N_7723);
xor U8808 (N_8808,N_7908,N_7971);
or U8809 (N_8809,N_7370,N_7139);
nor U8810 (N_8810,N_7487,N_7717);
xor U8811 (N_8811,N_7987,N_7587);
xor U8812 (N_8812,N_7836,N_7370);
or U8813 (N_8813,N_7591,N_7780);
nor U8814 (N_8814,N_7337,N_7709);
or U8815 (N_8815,N_7159,N_7777);
nor U8816 (N_8816,N_7341,N_7530);
nand U8817 (N_8817,N_7398,N_7695);
or U8818 (N_8818,N_7303,N_7204);
nor U8819 (N_8819,N_7747,N_7036);
xnor U8820 (N_8820,N_7848,N_7801);
nand U8821 (N_8821,N_7419,N_7012);
or U8822 (N_8822,N_7735,N_7752);
nand U8823 (N_8823,N_7378,N_7695);
and U8824 (N_8824,N_7353,N_7634);
nor U8825 (N_8825,N_7534,N_7784);
xnor U8826 (N_8826,N_7176,N_7147);
and U8827 (N_8827,N_7664,N_7481);
or U8828 (N_8828,N_7275,N_7570);
xnor U8829 (N_8829,N_7921,N_7587);
and U8830 (N_8830,N_7243,N_7828);
and U8831 (N_8831,N_7395,N_7690);
and U8832 (N_8832,N_7231,N_7704);
xor U8833 (N_8833,N_7301,N_7308);
nor U8834 (N_8834,N_7325,N_7994);
xnor U8835 (N_8835,N_7743,N_7315);
xor U8836 (N_8836,N_7480,N_7234);
or U8837 (N_8837,N_7554,N_7688);
nand U8838 (N_8838,N_7259,N_7310);
nor U8839 (N_8839,N_7772,N_7462);
or U8840 (N_8840,N_7126,N_7767);
and U8841 (N_8841,N_7890,N_7117);
or U8842 (N_8842,N_7289,N_7890);
nor U8843 (N_8843,N_7111,N_7240);
xnor U8844 (N_8844,N_7964,N_7182);
or U8845 (N_8845,N_7836,N_7932);
nand U8846 (N_8846,N_7516,N_7376);
nand U8847 (N_8847,N_7275,N_7749);
xnor U8848 (N_8848,N_7688,N_7186);
and U8849 (N_8849,N_7659,N_7788);
or U8850 (N_8850,N_7302,N_7740);
and U8851 (N_8851,N_7254,N_7994);
xnor U8852 (N_8852,N_7826,N_7153);
or U8853 (N_8853,N_7744,N_7434);
nand U8854 (N_8854,N_7094,N_7911);
nand U8855 (N_8855,N_7905,N_7828);
and U8856 (N_8856,N_7482,N_7352);
and U8857 (N_8857,N_7720,N_7881);
and U8858 (N_8858,N_7052,N_7409);
nand U8859 (N_8859,N_7482,N_7309);
nor U8860 (N_8860,N_7887,N_7423);
and U8861 (N_8861,N_7481,N_7494);
and U8862 (N_8862,N_7712,N_7384);
nor U8863 (N_8863,N_7387,N_7352);
nand U8864 (N_8864,N_7391,N_7463);
or U8865 (N_8865,N_7375,N_7214);
or U8866 (N_8866,N_7889,N_7348);
or U8867 (N_8867,N_7142,N_7496);
nor U8868 (N_8868,N_7158,N_7192);
and U8869 (N_8869,N_7426,N_7445);
nand U8870 (N_8870,N_7223,N_7352);
xnor U8871 (N_8871,N_7236,N_7441);
nand U8872 (N_8872,N_7526,N_7936);
nor U8873 (N_8873,N_7606,N_7913);
or U8874 (N_8874,N_7086,N_7850);
and U8875 (N_8875,N_7921,N_7771);
xor U8876 (N_8876,N_7518,N_7760);
or U8877 (N_8877,N_7756,N_7940);
nor U8878 (N_8878,N_7714,N_7466);
and U8879 (N_8879,N_7477,N_7110);
xor U8880 (N_8880,N_7726,N_7100);
or U8881 (N_8881,N_7070,N_7887);
or U8882 (N_8882,N_7840,N_7606);
nor U8883 (N_8883,N_7682,N_7545);
nor U8884 (N_8884,N_7680,N_7877);
and U8885 (N_8885,N_7077,N_7700);
or U8886 (N_8886,N_7010,N_7955);
and U8887 (N_8887,N_7763,N_7278);
and U8888 (N_8888,N_7756,N_7810);
or U8889 (N_8889,N_7340,N_7696);
and U8890 (N_8890,N_7786,N_7788);
or U8891 (N_8891,N_7164,N_7738);
nand U8892 (N_8892,N_7967,N_7265);
and U8893 (N_8893,N_7127,N_7584);
and U8894 (N_8894,N_7094,N_7416);
xor U8895 (N_8895,N_7981,N_7000);
nor U8896 (N_8896,N_7019,N_7453);
nand U8897 (N_8897,N_7714,N_7957);
and U8898 (N_8898,N_7724,N_7683);
nor U8899 (N_8899,N_7435,N_7468);
nand U8900 (N_8900,N_7085,N_7938);
xnor U8901 (N_8901,N_7293,N_7423);
or U8902 (N_8902,N_7000,N_7558);
xnor U8903 (N_8903,N_7753,N_7991);
nor U8904 (N_8904,N_7198,N_7749);
or U8905 (N_8905,N_7226,N_7801);
and U8906 (N_8906,N_7865,N_7905);
and U8907 (N_8907,N_7631,N_7965);
or U8908 (N_8908,N_7625,N_7608);
and U8909 (N_8909,N_7638,N_7425);
nand U8910 (N_8910,N_7937,N_7137);
or U8911 (N_8911,N_7519,N_7253);
nand U8912 (N_8912,N_7105,N_7521);
nor U8913 (N_8913,N_7935,N_7271);
and U8914 (N_8914,N_7498,N_7684);
and U8915 (N_8915,N_7040,N_7193);
xnor U8916 (N_8916,N_7359,N_7504);
nand U8917 (N_8917,N_7353,N_7627);
nand U8918 (N_8918,N_7692,N_7962);
and U8919 (N_8919,N_7416,N_7682);
nand U8920 (N_8920,N_7674,N_7004);
nor U8921 (N_8921,N_7997,N_7276);
nor U8922 (N_8922,N_7387,N_7155);
nand U8923 (N_8923,N_7237,N_7401);
and U8924 (N_8924,N_7540,N_7451);
and U8925 (N_8925,N_7751,N_7660);
nand U8926 (N_8926,N_7937,N_7095);
nand U8927 (N_8927,N_7984,N_7767);
and U8928 (N_8928,N_7371,N_7285);
nand U8929 (N_8929,N_7293,N_7700);
nand U8930 (N_8930,N_7053,N_7960);
nand U8931 (N_8931,N_7704,N_7776);
nand U8932 (N_8932,N_7149,N_7479);
or U8933 (N_8933,N_7404,N_7121);
and U8934 (N_8934,N_7270,N_7059);
xnor U8935 (N_8935,N_7879,N_7842);
or U8936 (N_8936,N_7181,N_7581);
nand U8937 (N_8937,N_7081,N_7354);
xnor U8938 (N_8938,N_7389,N_7474);
or U8939 (N_8939,N_7652,N_7818);
or U8940 (N_8940,N_7621,N_7548);
or U8941 (N_8941,N_7751,N_7464);
or U8942 (N_8942,N_7451,N_7603);
xor U8943 (N_8943,N_7914,N_7014);
and U8944 (N_8944,N_7171,N_7555);
nand U8945 (N_8945,N_7025,N_7683);
nor U8946 (N_8946,N_7174,N_7968);
nor U8947 (N_8947,N_7613,N_7822);
xor U8948 (N_8948,N_7763,N_7802);
and U8949 (N_8949,N_7245,N_7446);
nand U8950 (N_8950,N_7827,N_7603);
nor U8951 (N_8951,N_7879,N_7618);
or U8952 (N_8952,N_7990,N_7113);
and U8953 (N_8953,N_7486,N_7513);
or U8954 (N_8954,N_7710,N_7467);
and U8955 (N_8955,N_7109,N_7759);
or U8956 (N_8956,N_7298,N_7860);
or U8957 (N_8957,N_7801,N_7412);
xnor U8958 (N_8958,N_7192,N_7358);
xnor U8959 (N_8959,N_7171,N_7778);
nand U8960 (N_8960,N_7332,N_7784);
xnor U8961 (N_8961,N_7407,N_7550);
nor U8962 (N_8962,N_7692,N_7724);
and U8963 (N_8963,N_7433,N_7006);
nor U8964 (N_8964,N_7042,N_7801);
nand U8965 (N_8965,N_7926,N_7976);
nor U8966 (N_8966,N_7408,N_7359);
and U8967 (N_8967,N_7029,N_7841);
nor U8968 (N_8968,N_7259,N_7866);
or U8969 (N_8969,N_7235,N_7837);
nor U8970 (N_8970,N_7654,N_7461);
or U8971 (N_8971,N_7894,N_7710);
xor U8972 (N_8972,N_7563,N_7928);
xor U8973 (N_8973,N_7178,N_7556);
nand U8974 (N_8974,N_7286,N_7709);
or U8975 (N_8975,N_7323,N_7388);
or U8976 (N_8976,N_7985,N_7143);
xor U8977 (N_8977,N_7861,N_7298);
or U8978 (N_8978,N_7148,N_7916);
nand U8979 (N_8979,N_7667,N_7457);
and U8980 (N_8980,N_7674,N_7842);
xnor U8981 (N_8981,N_7597,N_7832);
nand U8982 (N_8982,N_7286,N_7122);
or U8983 (N_8983,N_7615,N_7359);
xor U8984 (N_8984,N_7397,N_7541);
nor U8985 (N_8985,N_7610,N_7388);
and U8986 (N_8986,N_7237,N_7011);
nor U8987 (N_8987,N_7359,N_7649);
nand U8988 (N_8988,N_7384,N_7515);
nand U8989 (N_8989,N_7793,N_7646);
xnor U8990 (N_8990,N_7577,N_7845);
and U8991 (N_8991,N_7247,N_7352);
nor U8992 (N_8992,N_7145,N_7668);
xor U8993 (N_8993,N_7729,N_7478);
xnor U8994 (N_8994,N_7896,N_7239);
xnor U8995 (N_8995,N_7587,N_7020);
xnor U8996 (N_8996,N_7420,N_7179);
nand U8997 (N_8997,N_7243,N_7256);
nor U8998 (N_8998,N_7525,N_7632);
nand U8999 (N_8999,N_7138,N_7988);
or U9000 (N_9000,N_8718,N_8901);
nand U9001 (N_9001,N_8754,N_8424);
nand U9002 (N_9002,N_8951,N_8411);
or U9003 (N_9003,N_8750,N_8657);
nand U9004 (N_9004,N_8073,N_8071);
and U9005 (N_9005,N_8059,N_8868);
nand U9006 (N_9006,N_8114,N_8092);
xor U9007 (N_9007,N_8282,N_8061);
xnor U9008 (N_9008,N_8892,N_8500);
or U9009 (N_9009,N_8139,N_8262);
nand U9010 (N_9010,N_8453,N_8415);
nor U9011 (N_9011,N_8172,N_8514);
and U9012 (N_9012,N_8375,N_8221);
nand U9013 (N_9013,N_8460,N_8769);
nand U9014 (N_9014,N_8461,N_8349);
nand U9015 (N_9015,N_8843,N_8604);
and U9016 (N_9016,N_8010,N_8060);
or U9017 (N_9017,N_8708,N_8354);
and U9018 (N_9018,N_8988,N_8076);
nand U9019 (N_9019,N_8249,N_8021);
and U9020 (N_9020,N_8519,N_8985);
or U9021 (N_9021,N_8789,N_8326);
xor U9022 (N_9022,N_8701,N_8904);
or U9023 (N_9023,N_8751,N_8456);
xor U9024 (N_9024,N_8558,N_8940);
or U9025 (N_9025,N_8556,N_8016);
nor U9026 (N_9026,N_8767,N_8089);
or U9027 (N_9027,N_8648,N_8723);
xor U9028 (N_9028,N_8703,N_8573);
xor U9029 (N_9029,N_8385,N_8119);
xor U9030 (N_9030,N_8711,N_8809);
nand U9031 (N_9031,N_8852,N_8917);
nor U9032 (N_9032,N_8002,N_8559);
nand U9033 (N_9033,N_8834,N_8271);
nor U9034 (N_9034,N_8108,N_8664);
nand U9035 (N_9035,N_8142,N_8782);
and U9036 (N_9036,N_8839,N_8749);
nand U9037 (N_9037,N_8737,N_8196);
or U9038 (N_9038,N_8726,N_8134);
nand U9039 (N_9039,N_8105,N_8106);
and U9040 (N_9040,N_8536,N_8584);
xor U9041 (N_9041,N_8979,N_8020);
nand U9042 (N_9042,N_8548,N_8619);
xnor U9043 (N_9043,N_8111,N_8659);
nand U9044 (N_9044,N_8379,N_8990);
nand U9045 (N_9045,N_8964,N_8296);
and U9046 (N_9046,N_8308,N_8642);
xnor U9047 (N_9047,N_8116,N_8425);
or U9048 (N_9048,N_8420,N_8608);
or U9049 (N_9049,N_8913,N_8862);
and U9050 (N_9050,N_8314,N_8126);
xnor U9051 (N_9051,N_8128,N_8431);
or U9052 (N_9052,N_8035,N_8094);
or U9053 (N_9053,N_8077,N_8840);
nor U9054 (N_9054,N_8051,N_8045);
nor U9055 (N_9055,N_8147,N_8978);
or U9056 (N_9056,N_8710,N_8476);
xor U9057 (N_9057,N_8881,N_8747);
or U9058 (N_9058,N_8992,N_8507);
and U9059 (N_9059,N_8575,N_8733);
nor U9060 (N_9060,N_8003,N_8110);
xor U9061 (N_9061,N_8074,N_8104);
nand U9062 (N_9062,N_8755,N_8890);
nor U9063 (N_9063,N_8325,N_8005);
nand U9064 (N_9064,N_8407,N_8595);
nand U9065 (N_9065,N_8129,N_8593);
xnor U9066 (N_9066,N_8182,N_8403);
or U9067 (N_9067,N_8240,N_8958);
nand U9068 (N_9068,N_8390,N_8309);
nor U9069 (N_9069,N_8540,N_8874);
and U9070 (N_9070,N_8631,N_8138);
and U9071 (N_9071,N_8564,N_8870);
nand U9072 (N_9072,N_8223,N_8253);
xor U9073 (N_9073,N_8009,N_8788);
xor U9074 (N_9074,N_8357,N_8144);
xor U9075 (N_9075,N_8423,N_8658);
and U9076 (N_9076,N_8472,N_8479);
nor U9077 (N_9077,N_8374,N_8683);
xnor U9078 (N_9078,N_8096,N_8184);
nor U9079 (N_9079,N_8932,N_8724);
and U9080 (N_9080,N_8239,N_8083);
or U9081 (N_9081,N_8865,N_8275);
xnor U9082 (N_9082,N_8444,N_8669);
and U9083 (N_9083,N_8891,N_8458);
nor U9084 (N_9084,N_8638,N_8900);
nand U9085 (N_9085,N_8580,N_8705);
xnor U9086 (N_9086,N_8244,N_8033);
nor U9087 (N_9087,N_8712,N_8494);
xor U9088 (N_9088,N_8023,N_8534);
xor U9089 (N_9089,N_8607,N_8136);
and U9090 (N_9090,N_8827,N_8081);
nor U9091 (N_9091,N_8360,N_8482);
nand U9092 (N_9092,N_8412,N_8930);
xor U9093 (N_9093,N_8250,N_8406);
and U9094 (N_9094,N_8836,N_8471);
xnor U9095 (N_9095,N_8384,N_8149);
nor U9096 (N_9096,N_8270,N_8690);
and U9097 (N_9097,N_8831,N_8915);
xor U9098 (N_9098,N_8161,N_8084);
nand U9099 (N_9099,N_8307,N_8195);
xor U9100 (N_9100,N_8920,N_8222);
and U9101 (N_9101,N_8004,N_8748);
and U9102 (N_9102,N_8306,N_8049);
nor U9103 (N_9103,N_8273,N_8905);
and U9104 (N_9104,N_8447,N_8246);
nand U9105 (N_9105,N_8473,N_8700);
nor U9106 (N_9106,N_8510,N_8995);
xnor U9107 (N_9107,N_8800,N_8893);
or U9108 (N_9108,N_8395,N_8762);
xnor U9109 (N_9109,N_8457,N_8070);
and U9110 (N_9110,N_8392,N_8511);
nor U9111 (N_9111,N_8770,N_8961);
and U9112 (N_9112,N_8833,N_8280);
and U9113 (N_9113,N_8744,N_8466);
nand U9114 (N_9114,N_8435,N_8135);
nor U9115 (N_9115,N_8886,N_8611);
xor U9116 (N_9116,N_8630,N_8159);
nand U9117 (N_9117,N_8842,N_8605);
nand U9118 (N_9118,N_8968,N_8826);
nor U9119 (N_9119,N_8670,N_8557);
nand U9120 (N_9120,N_8037,N_8947);
and U9121 (N_9121,N_8328,N_8140);
xor U9122 (N_9122,N_8288,N_8481);
and U9123 (N_9123,N_8409,N_8168);
nor U9124 (N_9124,N_8332,N_8602);
nand U9125 (N_9125,N_8313,N_8696);
or U9126 (N_9126,N_8102,N_8957);
nand U9127 (N_9127,N_8706,N_8192);
or U9128 (N_9128,N_8676,N_8151);
nand U9129 (N_9129,N_8279,N_8614);
or U9130 (N_9130,N_8987,N_8794);
and U9131 (N_9131,N_8449,N_8115);
nand U9132 (N_9132,N_8480,N_8633);
xnor U9133 (N_9133,N_8428,N_8819);
nor U9134 (N_9134,N_8418,N_8721);
xnor U9135 (N_9135,N_8908,N_8329);
or U9136 (N_9136,N_8936,N_8967);
nand U9137 (N_9137,N_8627,N_8372);
nand U9138 (N_9138,N_8066,N_8505);
xnor U9139 (N_9139,N_8207,N_8430);
or U9140 (N_9140,N_8509,N_8512);
or U9141 (N_9141,N_8739,N_8764);
nor U9142 (N_9142,N_8345,N_8014);
nand U9143 (N_9143,N_8441,N_8224);
or U9144 (N_9144,N_8731,N_8955);
nor U9145 (N_9145,N_8613,N_8561);
xnor U9146 (N_9146,N_8274,N_8822);
and U9147 (N_9147,N_8860,N_8760);
and U9148 (N_9148,N_8846,N_8465);
and U9149 (N_9149,N_8956,N_8260);
xnor U9150 (N_9150,N_8953,N_8067);
xor U9151 (N_9151,N_8885,N_8871);
nor U9152 (N_9152,N_8553,N_8966);
or U9153 (N_9153,N_8130,N_8784);
nand U9154 (N_9154,N_8335,N_8585);
nor U9155 (N_9155,N_8637,N_8365);
nor U9156 (N_9156,N_8729,N_8927);
and U9157 (N_9157,N_8436,N_8590);
or U9158 (N_9158,N_8327,N_8685);
nand U9159 (N_9159,N_8208,N_8623);
nor U9160 (N_9160,N_8888,N_8996);
xor U9161 (N_9161,N_8263,N_8790);
xor U9162 (N_9162,N_8983,N_8422);
and U9163 (N_9163,N_8232,N_8463);
nor U9164 (N_9164,N_8591,N_8233);
nor U9165 (N_9165,N_8245,N_8228);
xor U9166 (N_9166,N_8455,N_8334);
xnor U9167 (N_9167,N_8668,N_8048);
and U9168 (N_9168,N_8267,N_8587);
nor U9169 (N_9169,N_8153,N_8662);
nand U9170 (N_9170,N_8171,N_8187);
or U9171 (N_9171,N_8941,N_8351);
and U9172 (N_9172,N_8167,N_8880);
or U9173 (N_9173,N_8516,N_8903);
nand U9174 (N_9174,N_8715,N_8554);
and U9175 (N_9175,N_8298,N_8364);
or U9176 (N_9176,N_8856,N_8916);
xor U9177 (N_9177,N_8524,N_8474);
nand U9178 (N_9178,N_8699,N_8205);
nand U9179 (N_9179,N_8198,N_8889);
and U9180 (N_9180,N_8419,N_8186);
and U9181 (N_9181,N_8937,N_8997);
and U9182 (N_9182,N_8707,N_8709);
and U9183 (N_9183,N_8717,N_8165);
nand U9184 (N_9184,N_8738,N_8193);
xor U9185 (N_9185,N_8062,N_8017);
or U9186 (N_9186,N_8853,N_8811);
nor U9187 (N_9187,N_8746,N_8399);
nand U9188 (N_9188,N_8867,N_8068);
nand U9189 (N_9189,N_8291,N_8719);
xor U9190 (N_9190,N_8363,N_8179);
xnor U9191 (N_9191,N_8100,N_8620);
and U9192 (N_9192,N_8347,N_8145);
xor U9193 (N_9193,N_8396,N_8157);
and U9194 (N_9194,N_8798,N_8121);
nor U9195 (N_9195,N_8649,N_8072);
nand U9196 (N_9196,N_8495,N_8948);
or U9197 (N_9197,N_8772,N_8213);
or U9198 (N_9198,N_8214,N_8301);
or U9199 (N_9199,N_8634,N_8022);
nor U9200 (N_9200,N_8497,N_8655);
nand U9201 (N_9201,N_8535,N_8356);
nand U9202 (N_9202,N_8973,N_8621);
or U9203 (N_9203,N_8131,N_8727);
nand U9204 (N_9204,N_8231,N_8303);
nor U9205 (N_9205,N_8615,N_8169);
and U9206 (N_9206,N_8692,N_8487);
or U9207 (N_9207,N_8448,N_8506);
or U9208 (N_9208,N_8366,N_8938);
xor U9209 (N_9209,N_8043,N_8148);
and U9210 (N_9210,N_8854,N_8687);
nor U9211 (N_9211,N_8146,N_8065);
xor U9212 (N_9212,N_8923,N_8226);
nor U9213 (N_9213,N_8380,N_8109);
and U9214 (N_9214,N_8910,N_8626);
nor U9215 (N_9215,N_8432,N_8610);
xor U9216 (N_9216,N_8799,N_8663);
or U9217 (N_9217,N_8498,N_8993);
nand U9218 (N_9218,N_8359,N_8440);
and U9219 (N_9219,N_8319,N_8736);
and U9220 (N_9220,N_8013,N_8786);
or U9221 (N_9221,N_8277,N_8918);
nand U9222 (N_9222,N_8484,N_8323);
or U9223 (N_9223,N_8123,N_8776);
xor U9224 (N_9224,N_8625,N_8581);
and U9225 (N_9225,N_8814,N_8999);
or U9226 (N_9226,N_8684,N_8376);
and U9227 (N_9227,N_8241,N_8030);
or U9228 (N_9228,N_8079,N_8039);
or U9229 (N_9229,N_8644,N_8050);
xor U9230 (N_9230,N_8493,N_8370);
and U9231 (N_9231,N_8686,N_8041);
xnor U9232 (N_9232,N_8008,N_8928);
xnor U9233 (N_9233,N_8518,N_8882);
and U9234 (N_9234,N_8302,N_8829);
nor U9235 (N_9235,N_8001,N_8256);
xor U9236 (N_9236,N_8740,N_8266);
nand U9237 (N_9237,N_8522,N_8765);
nor U9238 (N_9238,N_8531,N_8855);
and U9239 (N_9239,N_8550,N_8693);
nand U9240 (N_9240,N_8785,N_8792);
and U9241 (N_9241,N_8780,N_8287);
or U9242 (N_9242,N_8551,N_8489);
and U9243 (N_9243,N_8097,N_8906);
xnor U9244 (N_9244,N_8572,N_8952);
nor U9245 (N_9245,N_8775,N_8201);
and U9246 (N_9246,N_8181,N_8416);
nor U9247 (N_9247,N_8215,N_8219);
and U9248 (N_9248,N_8160,N_8872);
xor U9249 (N_9249,N_8803,N_8289);
and U9250 (N_9250,N_8849,N_8503);
and U9251 (N_9251,N_8791,N_8174);
and U9252 (N_9252,N_8237,N_8098);
nand U9253 (N_9253,N_8210,N_8646);
nand U9254 (N_9254,N_8211,N_8156);
and U9255 (N_9255,N_8725,N_8338);
or U9256 (N_9256,N_8353,N_8133);
or U9257 (N_9257,N_8317,N_8688);
or U9258 (N_9258,N_8469,N_8342);
nand U9259 (N_9259,N_8645,N_8450);
nor U9260 (N_9260,N_8774,N_8445);
xor U9261 (N_9261,N_8653,N_8166);
xnor U9262 (N_9262,N_8824,N_8568);
or U9263 (N_9263,N_8838,N_8925);
xnor U9264 (N_9264,N_8386,N_8589);
and U9265 (N_9265,N_8802,N_8694);
and U9266 (N_9266,N_8029,N_8227);
or U9267 (N_9267,N_8962,N_8355);
or U9268 (N_9268,N_8285,N_8485);
xor U9269 (N_9269,N_8348,N_8099);
and U9270 (N_9270,N_8875,N_8333);
and U9271 (N_9271,N_8031,N_8869);
nor U9272 (N_9272,N_8741,N_8204);
nor U9273 (N_9273,N_8124,N_8527);
nand U9274 (N_9274,N_8127,N_8235);
xnor U9275 (N_9275,N_8592,N_8082);
xor U9276 (N_9276,N_8722,N_8197);
nand U9277 (N_9277,N_8055,N_8596);
nand U9278 (N_9278,N_8815,N_8178);
and U9279 (N_9279,N_8520,N_8426);
nor U9280 (N_9280,N_8768,N_8290);
or U9281 (N_9281,N_8758,N_8264);
xnor U9282 (N_9282,N_8299,N_8341);
nor U9283 (N_9283,N_8152,N_8742);
xnor U9284 (N_9284,N_8477,N_8054);
nand U9285 (N_9285,N_8000,N_8896);
xor U9286 (N_9286,N_8622,N_8177);
nor U9287 (N_9287,N_8191,N_8678);
and U9288 (N_9288,N_8808,N_8340);
and U9289 (N_9289,N_8796,N_8414);
xnor U9290 (N_9290,N_8281,N_8753);
nor U9291 (N_9291,N_8851,N_8806);
or U9292 (N_9292,N_8636,N_8137);
or U9293 (N_9293,N_8141,N_8562);
nand U9294 (N_9294,N_8857,N_8297);
or U9295 (N_9295,N_8574,N_8080);
xor U9296 (N_9296,N_8528,N_8743);
and U9297 (N_9297,N_8994,N_8929);
nand U9298 (N_9298,N_8063,N_8011);
nand U9299 (N_9299,N_8960,N_8845);
and U9300 (N_9300,N_8609,N_8583);
xor U9301 (N_9301,N_8661,N_8783);
or U9302 (N_9302,N_8442,N_8702);
or U9303 (N_9303,N_8118,N_8502);
nor U9304 (N_9304,N_8597,N_8006);
xnor U9305 (N_9305,N_8897,N_8909);
or U9306 (N_9306,N_8276,N_8984);
xor U9307 (N_9307,N_8439,N_8294);
nor U9308 (N_9308,N_8599,N_8866);
nand U9309 (N_9309,N_8499,N_8337);
nor U9310 (N_9310,N_8057,N_8781);
and U9311 (N_9311,N_8976,N_8251);
and U9312 (N_9312,N_8367,N_8513);
or U9313 (N_9313,N_8268,N_8624);
xor U9314 (N_9314,N_8847,N_8939);
and U9315 (N_9315,N_8443,N_8405);
xor U9316 (N_9316,N_8926,N_8336);
xor U9317 (N_9317,N_8606,N_8427);
nor U9318 (N_9318,N_8209,N_8086);
xnor U9319 (N_9319,N_8292,N_8488);
xnor U9320 (N_9320,N_8848,N_8389);
xnor U9321 (N_9321,N_8601,N_8438);
and U9322 (N_9322,N_8734,N_8508);
nor U9323 (N_9323,N_8258,N_8413);
nand U9324 (N_9324,N_8566,N_8504);
nand U9325 (N_9325,N_8943,N_8640);
xnor U9326 (N_9326,N_8408,N_8394);
xor U9327 (N_9327,N_8828,N_8162);
nor U9328 (N_9328,N_8628,N_8681);
xnor U9329 (N_9329,N_8199,N_8286);
nor U9330 (N_9330,N_8745,N_8931);
nand U9331 (N_9331,N_8539,N_8761);
nor U9332 (N_9332,N_8899,N_8989);
xnor U9333 (N_9333,N_8026,N_8907);
xor U9334 (N_9334,N_8042,N_8818);
nand U9335 (N_9335,N_8969,N_8612);
nand U9336 (N_9336,N_8038,N_8019);
and U9337 (N_9337,N_8069,N_8346);
and U9338 (N_9338,N_8887,N_8052);
xnor U9339 (N_9339,N_8567,N_8651);
nand U9340 (N_9340,N_8844,N_8183);
nand U9341 (N_9341,N_8015,N_8486);
nor U9342 (N_9342,N_8521,N_8234);
xnor U9343 (N_9343,N_8577,N_8689);
nand U9344 (N_9344,N_8821,N_8933);
xor U9345 (N_9345,N_8085,N_8437);
or U9346 (N_9346,N_8823,N_8185);
or U9347 (N_9347,N_8565,N_8537);
and U9348 (N_9348,N_8344,N_8491);
and U9349 (N_9349,N_8180,N_8830);
xnor U9350 (N_9350,N_8470,N_8578);
and U9351 (N_9351,N_8720,N_8666);
nand U9352 (N_9352,N_8944,N_8189);
and U9353 (N_9353,N_8804,N_8991);
or U9354 (N_9354,N_8934,N_8058);
nor U9355 (N_9355,N_8036,N_8714);
nand U9356 (N_9356,N_8837,N_8813);
and U9357 (N_9357,N_8877,N_8401);
or U9358 (N_9358,N_8752,N_8588);
nand U9359 (N_9359,N_8257,N_8667);
and U9360 (N_9360,N_8778,N_8218);
xor U9361 (N_9361,N_8242,N_8093);
xor U9362 (N_9362,N_8552,N_8368);
nor U9363 (N_9363,N_8586,N_8305);
nor U9364 (N_9364,N_8555,N_8523);
nand U9365 (N_9365,N_8143,N_8674);
and U9366 (N_9366,N_8315,N_8028);
or U9367 (N_9367,N_8654,N_8970);
nor U9368 (N_9368,N_8324,N_8265);
and U9369 (N_9369,N_8377,N_8120);
xnor U9370 (N_9370,N_8680,N_8350);
xnor U9371 (N_9371,N_8388,N_8571);
and U9372 (N_9372,N_8295,N_8475);
or U9373 (N_9373,N_8248,N_8200);
xor U9374 (N_9374,N_8810,N_8569);
nand U9375 (N_9375,N_8950,N_8873);
xnor U9376 (N_9376,N_8155,N_8795);
xnor U9377 (N_9377,N_8361,N_8787);
nor U9378 (N_9378,N_8330,N_8697);
nand U9379 (N_9379,N_8091,N_8496);
nor U9380 (N_9380,N_8695,N_8618);
and U9381 (N_9381,N_8236,N_8598);
nor U9382 (N_9382,N_8641,N_8032);
nor U9383 (N_9383,N_8616,N_8454);
nand U9384 (N_9384,N_8793,N_8492);
nand U9385 (N_9385,N_8304,N_8047);
or U9386 (N_9386,N_8912,N_8490);
or U9387 (N_9387,N_8850,N_8600);
xor U9388 (N_9388,N_8170,N_8816);
or U9389 (N_9389,N_8378,N_8369);
or U9390 (N_9390,N_8190,N_8164);
and U9391 (N_9391,N_8398,N_8858);
nor U9392 (N_9392,N_8320,N_8173);
and U9393 (N_9393,N_8980,N_8300);
nand U9394 (N_9394,N_8293,N_8805);
xnor U9395 (N_9395,N_8704,N_8763);
nor U9396 (N_9396,N_8464,N_8371);
or U9397 (N_9397,N_8515,N_8922);
and U9398 (N_9398,N_8238,N_8773);
nand U9399 (N_9399,N_8194,N_8635);
and U9400 (N_9400,N_8639,N_8252);
and U9401 (N_9401,N_8312,N_8797);
and U9402 (N_9402,N_8397,N_8971);
xnor U9403 (N_9403,N_8671,N_8945);
and U9404 (N_9404,N_8629,N_8501);
or U9405 (N_9405,N_8576,N_8981);
nor U9406 (N_9406,N_8665,N_8087);
xnor U9407 (N_9407,N_8462,N_8217);
and U9408 (N_9408,N_8986,N_8541);
and U9409 (N_9409,N_8381,N_8698);
nor U9410 (N_9410,N_8358,N_8088);
nand U9411 (N_9411,N_8544,N_8113);
and U9412 (N_9412,N_8362,N_8545);
nor U9413 (N_9413,N_8339,N_8677);
or U9414 (N_9414,N_8283,N_8863);
xnor U9415 (N_9415,N_8911,N_8716);
and U9416 (N_9416,N_8570,N_8163);
and U9417 (N_9417,N_8459,N_8650);
and U9418 (N_9418,N_8977,N_8660);
and U9419 (N_9419,N_8533,N_8269);
or U9420 (N_9420,N_8421,N_8876);
or U9421 (N_9421,N_8040,N_8756);
and U9422 (N_9422,N_8975,N_8034);
or U9423 (N_9423,N_8543,N_8779);
xnor U9424 (N_9424,N_8206,N_8322);
nor U9425 (N_9425,N_8582,N_8216);
nor U9426 (N_9426,N_8202,N_8526);
and U9427 (N_9427,N_8924,N_8825);
nor U9428 (N_9428,N_8046,N_8451);
xor U9429 (N_9429,N_8402,N_8383);
nor U9430 (N_9430,N_8603,N_8898);
nor U9431 (N_9431,N_8064,N_8652);
and U9432 (N_9432,N_8272,N_8643);
nor U9433 (N_9433,N_8965,N_8012);
xor U9434 (N_9434,N_8027,N_8579);
xnor U9435 (N_9435,N_8018,N_8914);
and U9436 (N_9436,N_8467,N_8730);
or U9437 (N_9437,N_8117,N_8954);
xor U9438 (N_9438,N_8254,N_8343);
xnor U9439 (N_9439,N_8759,N_8154);
nand U9440 (N_9440,N_8679,N_8150);
nor U9441 (N_9441,N_8230,N_8563);
xor U9442 (N_9442,N_8942,N_8517);
or U9443 (N_9443,N_8807,N_8247);
and U9444 (N_9444,N_8766,N_8452);
and U9445 (N_9445,N_8125,N_8243);
xor U9446 (N_9446,N_8546,N_8777);
nand U9447 (N_9447,N_8434,N_8542);
and U9448 (N_9448,N_8538,N_8732);
nor U9449 (N_9449,N_8919,N_8728);
nand U9450 (N_9450,N_8894,N_8675);
xor U9451 (N_9451,N_8529,N_8560);
or U9452 (N_9452,N_8175,N_8547);
nand U9453 (N_9453,N_8203,N_8921);
nor U9454 (N_9454,N_8656,N_8284);
nand U9455 (N_9455,N_8053,N_8255);
xnor U9456 (N_9456,N_8158,N_8417);
nand U9457 (N_9457,N_8404,N_8832);
nor U9458 (N_9458,N_8884,N_8982);
xnor U9459 (N_9459,N_8122,N_8095);
or U9460 (N_9460,N_8902,N_8817);
nor U9461 (N_9461,N_8393,N_8673);
nor U9462 (N_9462,N_8532,N_8935);
nor U9463 (N_9463,N_8278,N_8107);
and U9464 (N_9464,N_8321,N_8410);
xor U9465 (N_9465,N_8101,N_8525);
nand U9466 (N_9466,N_8078,N_8632);
xnor U9467 (N_9467,N_8895,N_8103);
xnor U9468 (N_9468,N_8672,N_8044);
nor U9469 (N_9469,N_8025,N_8949);
or U9470 (N_9470,N_8311,N_8878);
nor U9471 (N_9471,N_8735,N_8859);
and U9472 (N_9472,N_8841,N_8429);
nor U9473 (N_9473,N_8220,N_8812);
xnor U9474 (N_9474,N_8757,N_8530);
and U9475 (N_9475,N_8382,N_8261);
xnor U9476 (N_9476,N_8446,N_8820);
and U9477 (N_9477,N_8549,N_8188);
nand U9478 (N_9478,N_8112,N_8974);
and U9479 (N_9479,N_8963,N_8387);
or U9480 (N_9480,N_8132,N_8691);
or U9481 (N_9481,N_8259,N_8713);
xor U9482 (N_9482,N_8331,N_8959);
nand U9483 (N_9483,N_8946,N_8176);
and U9484 (N_9484,N_8483,N_8310);
nor U9485 (N_9485,N_8225,N_8771);
or U9486 (N_9486,N_8433,N_8647);
nand U9487 (N_9487,N_8864,N_8373);
or U9488 (N_9488,N_8400,N_8316);
nand U9489 (N_9489,N_8090,N_8801);
nand U9490 (N_9490,N_8007,N_8391);
nand U9491 (N_9491,N_8879,N_8352);
nor U9492 (N_9492,N_8212,N_8318);
and U9493 (N_9493,N_8861,N_8056);
nand U9494 (N_9494,N_8024,N_8478);
xnor U9495 (N_9495,N_8883,N_8468);
xnor U9496 (N_9496,N_8617,N_8682);
nand U9497 (N_9497,N_8972,N_8229);
and U9498 (N_9498,N_8594,N_8835);
nor U9499 (N_9499,N_8075,N_8998);
xor U9500 (N_9500,N_8206,N_8819);
xor U9501 (N_9501,N_8031,N_8231);
nand U9502 (N_9502,N_8849,N_8087);
nor U9503 (N_9503,N_8027,N_8515);
nand U9504 (N_9504,N_8161,N_8983);
nand U9505 (N_9505,N_8129,N_8347);
nand U9506 (N_9506,N_8146,N_8980);
or U9507 (N_9507,N_8151,N_8917);
or U9508 (N_9508,N_8008,N_8355);
or U9509 (N_9509,N_8203,N_8224);
and U9510 (N_9510,N_8070,N_8325);
and U9511 (N_9511,N_8390,N_8742);
and U9512 (N_9512,N_8310,N_8683);
or U9513 (N_9513,N_8681,N_8617);
and U9514 (N_9514,N_8591,N_8070);
or U9515 (N_9515,N_8872,N_8112);
xnor U9516 (N_9516,N_8960,N_8461);
nand U9517 (N_9517,N_8989,N_8102);
nand U9518 (N_9518,N_8392,N_8565);
or U9519 (N_9519,N_8851,N_8519);
and U9520 (N_9520,N_8050,N_8605);
and U9521 (N_9521,N_8843,N_8971);
nand U9522 (N_9522,N_8774,N_8309);
nor U9523 (N_9523,N_8956,N_8503);
and U9524 (N_9524,N_8747,N_8726);
xor U9525 (N_9525,N_8239,N_8817);
nand U9526 (N_9526,N_8138,N_8355);
nor U9527 (N_9527,N_8838,N_8217);
nand U9528 (N_9528,N_8658,N_8362);
xor U9529 (N_9529,N_8009,N_8134);
and U9530 (N_9530,N_8765,N_8866);
xor U9531 (N_9531,N_8841,N_8122);
nor U9532 (N_9532,N_8879,N_8309);
or U9533 (N_9533,N_8809,N_8129);
nand U9534 (N_9534,N_8718,N_8917);
nand U9535 (N_9535,N_8066,N_8780);
nand U9536 (N_9536,N_8582,N_8529);
or U9537 (N_9537,N_8528,N_8097);
nand U9538 (N_9538,N_8479,N_8892);
nand U9539 (N_9539,N_8408,N_8771);
or U9540 (N_9540,N_8309,N_8620);
and U9541 (N_9541,N_8318,N_8382);
and U9542 (N_9542,N_8087,N_8813);
xnor U9543 (N_9543,N_8900,N_8849);
or U9544 (N_9544,N_8106,N_8415);
xor U9545 (N_9545,N_8761,N_8496);
xor U9546 (N_9546,N_8383,N_8468);
or U9547 (N_9547,N_8154,N_8460);
nand U9548 (N_9548,N_8455,N_8997);
xnor U9549 (N_9549,N_8404,N_8219);
xnor U9550 (N_9550,N_8063,N_8463);
or U9551 (N_9551,N_8985,N_8540);
nor U9552 (N_9552,N_8225,N_8571);
and U9553 (N_9553,N_8469,N_8782);
or U9554 (N_9554,N_8863,N_8520);
and U9555 (N_9555,N_8312,N_8093);
nor U9556 (N_9556,N_8863,N_8116);
and U9557 (N_9557,N_8868,N_8135);
nor U9558 (N_9558,N_8245,N_8607);
nor U9559 (N_9559,N_8032,N_8310);
xnor U9560 (N_9560,N_8578,N_8122);
xor U9561 (N_9561,N_8479,N_8017);
or U9562 (N_9562,N_8603,N_8472);
nand U9563 (N_9563,N_8517,N_8984);
and U9564 (N_9564,N_8032,N_8692);
xor U9565 (N_9565,N_8243,N_8169);
or U9566 (N_9566,N_8176,N_8056);
nand U9567 (N_9567,N_8247,N_8026);
and U9568 (N_9568,N_8921,N_8687);
nor U9569 (N_9569,N_8290,N_8055);
xor U9570 (N_9570,N_8016,N_8007);
or U9571 (N_9571,N_8434,N_8747);
xor U9572 (N_9572,N_8097,N_8687);
and U9573 (N_9573,N_8562,N_8556);
xor U9574 (N_9574,N_8360,N_8946);
nand U9575 (N_9575,N_8714,N_8892);
nand U9576 (N_9576,N_8835,N_8118);
and U9577 (N_9577,N_8081,N_8189);
nand U9578 (N_9578,N_8988,N_8587);
xor U9579 (N_9579,N_8331,N_8192);
nand U9580 (N_9580,N_8049,N_8168);
nor U9581 (N_9581,N_8230,N_8950);
xor U9582 (N_9582,N_8927,N_8910);
nor U9583 (N_9583,N_8316,N_8514);
or U9584 (N_9584,N_8714,N_8904);
xnor U9585 (N_9585,N_8664,N_8902);
and U9586 (N_9586,N_8344,N_8454);
xnor U9587 (N_9587,N_8017,N_8746);
and U9588 (N_9588,N_8516,N_8031);
nor U9589 (N_9589,N_8582,N_8631);
xnor U9590 (N_9590,N_8470,N_8633);
xor U9591 (N_9591,N_8277,N_8187);
xor U9592 (N_9592,N_8061,N_8546);
or U9593 (N_9593,N_8839,N_8634);
xnor U9594 (N_9594,N_8791,N_8844);
nand U9595 (N_9595,N_8604,N_8141);
xnor U9596 (N_9596,N_8357,N_8662);
and U9597 (N_9597,N_8384,N_8989);
xor U9598 (N_9598,N_8182,N_8793);
or U9599 (N_9599,N_8125,N_8704);
nand U9600 (N_9600,N_8313,N_8422);
nor U9601 (N_9601,N_8268,N_8677);
nand U9602 (N_9602,N_8713,N_8383);
or U9603 (N_9603,N_8295,N_8690);
and U9604 (N_9604,N_8107,N_8003);
nor U9605 (N_9605,N_8291,N_8555);
nand U9606 (N_9606,N_8681,N_8858);
or U9607 (N_9607,N_8851,N_8101);
nor U9608 (N_9608,N_8919,N_8873);
nand U9609 (N_9609,N_8658,N_8540);
nor U9610 (N_9610,N_8920,N_8990);
or U9611 (N_9611,N_8567,N_8467);
or U9612 (N_9612,N_8836,N_8006);
or U9613 (N_9613,N_8792,N_8528);
nand U9614 (N_9614,N_8960,N_8936);
or U9615 (N_9615,N_8917,N_8219);
nor U9616 (N_9616,N_8373,N_8288);
nand U9617 (N_9617,N_8269,N_8145);
or U9618 (N_9618,N_8893,N_8674);
xnor U9619 (N_9619,N_8732,N_8593);
nor U9620 (N_9620,N_8913,N_8004);
and U9621 (N_9621,N_8467,N_8081);
xnor U9622 (N_9622,N_8252,N_8985);
and U9623 (N_9623,N_8272,N_8766);
and U9624 (N_9624,N_8945,N_8643);
nand U9625 (N_9625,N_8750,N_8171);
and U9626 (N_9626,N_8158,N_8924);
xnor U9627 (N_9627,N_8964,N_8895);
xnor U9628 (N_9628,N_8594,N_8325);
and U9629 (N_9629,N_8946,N_8620);
nand U9630 (N_9630,N_8390,N_8950);
nor U9631 (N_9631,N_8092,N_8474);
nor U9632 (N_9632,N_8587,N_8703);
nor U9633 (N_9633,N_8316,N_8757);
xor U9634 (N_9634,N_8604,N_8508);
xor U9635 (N_9635,N_8604,N_8036);
xnor U9636 (N_9636,N_8392,N_8275);
nor U9637 (N_9637,N_8575,N_8507);
and U9638 (N_9638,N_8116,N_8626);
or U9639 (N_9639,N_8421,N_8680);
and U9640 (N_9640,N_8660,N_8727);
nand U9641 (N_9641,N_8626,N_8134);
nor U9642 (N_9642,N_8103,N_8688);
xnor U9643 (N_9643,N_8054,N_8006);
xor U9644 (N_9644,N_8561,N_8904);
xor U9645 (N_9645,N_8307,N_8470);
and U9646 (N_9646,N_8198,N_8679);
or U9647 (N_9647,N_8912,N_8733);
or U9648 (N_9648,N_8652,N_8115);
and U9649 (N_9649,N_8191,N_8450);
and U9650 (N_9650,N_8130,N_8069);
and U9651 (N_9651,N_8141,N_8250);
xor U9652 (N_9652,N_8977,N_8106);
and U9653 (N_9653,N_8297,N_8410);
xor U9654 (N_9654,N_8692,N_8745);
or U9655 (N_9655,N_8862,N_8127);
nand U9656 (N_9656,N_8845,N_8594);
xor U9657 (N_9657,N_8779,N_8453);
nand U9658 (N_9658,N_8965,N_8031);
xor U9659 (N_9659,N_8925,N_8262);
nand U9660 (N_9660,N_8176,N_8514);
or U9661 (N_9661,N_8454,N_8545);
nand U9662 (N_9662,N_8902,N_8291);
nor U9663 (N_9663,N_8579,N_8555);
nor U9664 (N_9664,N_8191,N_8451);
nor U9665 (N_9665,N_8992,N_8989);
or U9666 (N_9666,N_8175,N_8332);
or U9667 (N_9667,N_8560,N_8734);
or U9668 (N_9668,N_8371,N_8783);
or U9669 (N_9669,N_8937,N_8840);
xor U9670 (N_9670,N_8723,N_8526);
nor U9671 (N_9671,N_8747,N_8401);
nor U9672 (N_9672,N_8877,N_8975);
xor U9673 (N_9673,N_8761,N_8555);
and U9674 (N_9674,N_8467,N_8517);
xor U9675 (N_9675,N_8420,N_8488);
and U9676 (N_9676,N_8855,N_8587);
xnor U9677 (N_9677,N_8211,N_8376);
or U9678 (N_9678,N_8942,N_8139);
or U9679 (N_9679,N_8171,N_8641);
xor U9680 (N_9680,N_8983,N_8601);
and U9681 (N_9681,N_8405,N_8455);
xor U9682 (N_9682,N_8994,N_8168);
or U9683 (N_9683,N_8795,N_8741);
and U9684 (N_9684,N_8454,N_8988);
xnor U9685 (N_9685,N_8354,N_8126);
or U9686 (N_9686,N_8855,N_8581);
or U9687 (N_9687,N_8208,N_8369);
nand U9688 (N_9688,N_8010,N_8712);
and U9689 (N_9689,N_8197,N_8110);
xnor U9690 (N_9690,N_8615,N_8085);
or U9691 (N_9691,N_8074,N_8448);
and U9692 (N_9692,N_8488,N_8294);
xor U9693 (N_9693,N_8458,N_8367);
and U9694 (N_9694,N_8026,N_8718);
nor U9695 (N_9695,N_8741,N_8301);
or U9696 (N_9696,N_8565,N_8883);
nand U9697 (N_9697,N_8172,N_8870);
and U9698 (N_9698,N_8172,N_8553);
nand U9699 (N_9699,N_8031,N_8763);
or U9700 (N_9700,N_8409,N_8361);
nor U9701 (N_9701,N_8282,N_8142);
nand U9702 (N_9702,N_8593,N_8669);
xor U9703 (N_9703,N_8027,N_8449);
nand U9704 (N_9704,N_8032,N_8223);
nor U9705 (N_9705,N_8878,N_8673);
xnor U9706 (N_9706,N_8324,N_8013);
nor U9707 (N_9707,N_8451,N_8709);
nand U9708 (N_9708,N_8304,N_8619);
nand U9709 (N_9709,N_8930,N_8971);
nor U9710 (N_9710,N_8513,N_8574);
nor U9711 (N_9711,N_8794,N_8554);
xor U9712 (N_9712,N_8006,N_8322);
nand U9713 (N_9713,N_8367,N_8818);
xnor U9714 (N_9714,N_8998,N_8203);
nor U9715 (N_9715,N_8032,N_8293);
nor U9716 (N_9716,N_8055,N_8171);
and U9717 (N_9717,N_8014,N_8924);
and U9718 (N_9718,N_8374,N_8822);
nand U9719 (N_9719,N_8900,N_8367);
nand U9720 (N_9720,N_8793,N_8923);
nand U9721 (N_9721,N_8641,N_8418);
xor U9722 (N_9722,N_8736,N_8246);
nor U9723 (N_9723,N_8595,N_8312);
and U9724 (N_9724,N_8942,N_8809);
xor U9725 (N_9725,N_8954,N_8585);
and U9726 (N_9726,N_8986,N_8667);
or U9727 (N_9727,N_8374,N_8910);
or U9728 (N_9728,N_8564,N_8296);
or U9729 (N_9729,N_8766,N_8343);
and U9730 (N_9730,N_8629,N_8971);
or U9731 (N_9731,N_8369,N_8975);
nand U9732 (N_9732,N_8575,N_8046);
nand U9733 (N_9733,N_8780,N_8840);
nor U9734 (N_9734,N_8042,N_8790);
or U9735 (N_9735,N_8244,N_8787);
xor U9736 (N_9736,N_8113,N_8911);
nor U9737 (N_9737,N_8439,N_8343);
or U9738 (N_9738,N_8662,N_8328);
and U9739 (N_9739,N_8264,N_8639);
and U9740 (N_9740,N_8956,N_8723);
and U9741 (N_9741,N_8499,N_8614);
nand U9742 (N_9742,N_8473,N_8479);
nand U9743 (N_9743,N_8889,N_8536);
and U9744 (N_9744,N_8473,N_8173);
or U9745 (N_9745,N_8587,N_8382);
nor U9746 (N_9746,N_8558,N_8397);
xnor U9747 (N_9747,N_8915,N_8857);
or U9748 (N_9748,N_8638,N_8023);
or U9749 (N_9749,N_8701,N_8512);
nor U9750 (N_9750,N_8482,N_8225);
nor U9751 (N_9751,N_8924,N_8148);
or U9752 (N_9752,N_8658,N_8450);
nand U9753 (N_9753,N_8124,N_8779);
and U9754 (N_9754,N_8854,N_8233);
nor U9755 (N_9755,N_8587,N_8440);
xnor U9756 (N_9756,N_8130,N_8404);
xor U9757 (N_9757,N_8145,N_8148);
and U9758 (N_9758,N_8766,N_8865);
xor U9759 (N_9759,N_8607,N_8384);
nor U9760 (N_9760,N_8718,N_8823);
nor U9761 (N_9761,N_8149,N_8336);
nand U9762 (N_9762,N_8371,N_8288);
nand U9763 (N_9763,N_8549,N_8993);
xor U9764 (N_9764,N_8199,N_8083);
xor U9765 (N_9765,N_8742,N_8133);
or U9766 (N_9766,N_8847,N_8707);
xor U9767 (N_9767,N_8979,N_8948);
nor U9768 (N_9768,N_8877,N_8283);
xor U9769 (N_9769,N_8674,N_8996);
xnor U9770 (N_9770,N_8144,N_8998);
xnor U9771 (N_9771,N_8943,N_8710);
or U9772 (N_9772,N_8745,N_8281);
nand U9773 (N_9773,N_8083,N_8968);
nand U9774 (N_9774,N_8748,N_8597);
xnor U9775 (N_9775,N_8373,N_8334);
xnor U9776 (N_9776,N_8524,N_8614);
and U9777 (N_9777,N_8235,N_8939);
nand U9778 (N_9778,N_8687,N_8816);
and U9779 (N_9779,N_8264,N_8714);
or U9780 (N_9780,N_8239,N_8444);
nand U9781 (N_9781,N_8937,N_8501);
nor U9782 (N_9782,N_8513,N_8264);
xnor U9783 (N_9783,N_8081,N_8571);
nor U9784 (N_9784,N_8590,N_8639);
and U9785 (N_9785,N_8042,N_8431);
nand U9786 (N_9786,N_8198,N_8170);
or U9787 (N_9787,N_8768,N_8085);
and U9788 (N_9788,N_8963,N_8172);
and U9789 (N_9789,N_8636,N_8176);
xnor U9790 (N_9790,N_8079,N_8577);
xor U9791 (N_9791,N_8442,N_8206);
nand U9792 (N_9792,N_8822,N_8263);
nand U9793 (N_9793,N_8835,N_8613);
nor U9794 (N_9794,N_8597,N_8536);
xnor U9795 (N_9795,N_8137,N_8713);
and U9796 (N_9796,N_8251,N_8526);
and U9797 (N_9797,N_8635,N_8028);
xor U9798 (N_9798,N_8418,N_8681);
nand U9799 (N_9799,N_8146,N_8653);
and U9800 (N_9800,N_8994,N_8802);
or U9801 (N_9801,N_8568,N_8139);
nor U9802 (N_9802,N_8663,N_8367);
and U9803 (N_9803,N_8600,N_8736);
nor U9804 (N_9804,N_8025,N_8989);
xnor U9805 (N_9805,N_8933,N_8960);
and U9806 (N_9806,N_8913,N_8931);
nand U9807 (N_9807,N_8979,N_8010);
xor U9808 (N_9808,N_8675,N_8712);
or U9809 (N_9809,N_8962,N_8976);
nand U9810 (N_9810,N_8181,N_8132);
nand U9811 (N_9811,N_8506,N_8415);
and U9812 (N_9812,N_8652,N_8775);
nor U9813 (N_9813,N_8365,N_8654);
xnor U9814 (N_9814,N_8924,N_8999);
nor U9815 (N_9815,N_8813,N_8886);
nand U9816 (N_9816,N_8515,N_8846);
xnor U9817 (N_9817,N_8727,N_8526);
and U9818 (N_9818,N_8453,N_8820);
nor U9819 (N_9819,N_8985,N_8942);
or U9820 (N_9820,N_8166,N_8007);
nor U9821 (N_9821,N_8536,N_8622);
and U9822 (N_9822,N_8441,N_8988);
xor U9823 (N_9823,N_8958,N_8564);
nor U9824 (N_9824,N_8733,N_8466);
and U9825 (N_9825,N_8665,N_8555);
and U9826 (N_9826,N_8926,N_8934);
nand U9827 (N_9827,N_8568,N_8438);
or U9828 (N_9828,N_8173,N_8151);
nand U9829 (N_9829,N_8251,N_8130);
or U9830 (N_9830,N_8643,N_8086);
or U9831 (N_9831,N_8696,N_8024);
or U9832 (N_9832,N_8095,N_8802);
xor U9833 (N_9833,N_8166,N_8370);
nor U9834 (N_9834,N_8955,N_8460);
nand U9835 (N_9835,N_8878,N_8100);
nor U9836 (N_9836,N_8790,N_8152);
or U9837 (N_9837,N_8203,N_8622);
xor U9838 (N_9838,N_8608,N_8097);
or U9839 (N_9839,N_8686,N_8742);
or U9840 (N_9840,N_8132,N_8169);
and U9841 (N_9841,N_8519,N_8448);
and U9842 (N_9842,N_8973,N_8051);
and U9843 (N_9843,N_8790,N_8524);
nor U9844 (N_9844,N_8543,N_8987);
and U9845 (N_9845,N_8538,N_8849);
and U9846 (N_9846,N_8520,N_8072);
or U9847 (N_9847,N_8658,N_8129);
or U9848 (N_9848,N_8011,N_8732);
and U9849 (N_9849,N_8850,N_8604);
nand U9850 (N_9850,N_8507,N_8314);
xnor U9851 (N_9851,N_8682,N_8627);
nor U9852 (N_9852,N_8217,N_8495);
nor U9853 (N_9853,N_8725,N_8431);
nand U9854 (N_9854,N_8555,N_8675);
nand U9855 (N_9855,N_8746,N_8888);
nor U9856 (N_9856,N_8753,N_8619);
or U9857 (N_9857,N_8167,N_8757);
nand U9858 (N_9858,N_8968,N_8508);
or U9859 (N_9859,N_8436,N_8840);
xnor U9860 (N_9860,N_8508,N_8100);
nor U9861 (N_9861,N_8127,N_8352);
and U9862 (N_9862,N_8061,N_8675);
xnor U9863 (N_9863,N_8569,N_8115);
and U9864 (N_9864,N_8440,N_8397);
nand U9865 (N_9865,N_8426,N_8462);
nand U9866 (N_9866,N_8950,N_8595);
and U9867 (N_9867,N_8264,N_8578);
and U9868 (N_9868,N_8611,N_8916);
nor U9869 (N_9869,N_8101,N_8464);
and U9870 (N_9870,N_8938,N_8600);
nand U9871 (N_9871,N_8496,N_8692);
or U9872 (N_9872,N_8870,N_8511);
xor U9873 (N_9873,N_8570,N_8629);
and U9874 (N_9874,N_8386,N_8802);
nand U9875 (N_9875,N_8866,N_8428);
nand U9876 (N_9876,N_8264,N_8056);
xor U9877 (N_9877,N_8613,N_8382);
nand U9878 (N_9878,N_8529,N_8164);
nor U9879 (N_9879,N_8192,N_8650);
nor U9880 (N_9880,N_8953,N_8360);
xor U9881 (N_9881,N_8095,N_8375);
nor U9882 (N_9882,N_8826,N_8105);
nor U9883 (N_9883,N_8174,N_8679);
nor U9884 (N_9884,N_8766,N_8375);
xor U9885 (N_9885,N_8811,N_8114);
xor U9886 (N_9886,N_8374,N_8606);
and U9887 (N_9887,N_8336,N_8477);
xor U9888 (N_9888,N_8810,N_8220);
or U9889 (N_9889,N_8175,N_8823);
nor U9890 (N_9890,N_8045,N_8068);
nand U9891 (N_9891,N_8915,N_8024);
xor U9892 (N_9892,N_8905,N_8806);
nand U9893 (N_9893,N_8537,N_8992);
xor U9894 (N_9894,N_8908,N_8759);
nor U9895 (N_9895,N_8767,N_8376);
xor U9896 (N_9896,N_8938,N_8678);
and U9897 (N_9897,N_8550,N_8269);
nor U9898 (N_9898,N_8142,N_8838);
nor U9899 (N_9899,N_8263,N_8922);
and U9900 (N_9900,N_8927,N_8057);
or U9901 (N_9901,N_8753,N_8445);
nand U9902 (N_9902,N_8043,N_8445);
nand U9903 (N_9903,N_8297,N_8097);
xor U9904 (N_9904,N_8589,N_8899);
or U9905 (N_9905,N_8293,N_8627);
and U9906 (N_9906,N_8454,N_8214);
or U9907 (N_9907,N_8551,N_8900);
and U9908 (N_9908,N_8972,N_8015);
nand U9909 (N_9909,N_8197,N_8432);
nor U9910 (N_9910,N_8932,N_8895);
or U9911 (N_9911,N_8548,N_8831);
and U9912 (N_9912,N_8491,N_8914);
or U9913 (N_9913,N_8594,N_8319);
nand U9914 (N_9914,N_8575,N_8942);
nand U9915 (N_9915,N_8329,N_8781);
xnor U9916 (N_9916,N_8784,N_8395);
nand U9917 (N_9917,N_8940,N_8254);
xnor U9918 (N_9918,N_8194,N_8467);
and U9919 (N_9919,N_8424,N_8173);
and U9920 (N_9920,N_8502,N_8399);
xor U9921 (N_9921,N_8144,N_8731);
xnor U9922 (N_9922,N_8974,N_8014);
and U9923 (N_9923,N_8056,N_8569);
and U9924 (N_9924,N_8750,N_8488);
nand U9925 (N_9925,N_8055,N_8917);
nand U9926 (N_9926,N_8183,N_8749);
and U9927 (N_9927,N_8580,N_8129);
xnor U9928 (N_9928,N_8559,N_8720);
nor U9929 (N_9929,N_8012,N_8593);
and U9930 (N_9930,N_8232,N_8727);
nand U9931 (N_9931,N_8029,N_8362);
or U9932 (N_9932,N_8017,N_8142);
or U9933 (N_9933,N_8604,N_8842);
nor U9934 (N_9934,N_8279,N_8232);
nand U9935 (N_9935,N_8636,N_8067);
nand U9936 (N_9936,N_8115,N_8921);
or U9937 (N_9937,N_8341,N_8993);
nor U9938 (N_9938,N_8424,N_8772);
xor U9939 (N_9939,N_8256,N_8665);
or U9940 (N_9940,N_8436,N_8641);
nor U9941 (N_9941,N_8078,N_8847);
nand U9942 (N_9942,N_8050,N_8196);
nor U9943 (N_9943,N_8301,N_8105);
and U9944 (N_9944,N_8894,N_8660);
and U9945 (N_9945,N_8101,N_8823);
nor U9946 (N_9946,N_8661,N_8362);
nand U9947 (N_9947,N_8145,N_8425);
and U9948 (N_9948,N_8596,N_8266);
or U9949 (N_9949,N_8368,N_8765);
nor U9950 (N_9950,N_8231,N_8162);
xnor U9951 (N_9951,N_8469,N_8273);
nand U9952 (N_9952,N_8633,N_8015);
nand U9953 (N_9953,N_8876,N_8417);
nand U9954 (N_9954,N_8585,N_8866);
or U9955 (N_9955,N_8684,N_8694);
nand U9956 (N_9956,N_8245,N_8082);
and U9957 (N_9957,N_8531,N_8195);
nand U9958 (N_9958,N_8108,N_8377);
or U9959 (N_9959,N_8875,N_8580);
xor U9960 (N_9960,N_8754,N_8438);
and U9961 (N_9961,N_8964,N_8625);
nand U9962 (N_9962,N_8305,N_8408);
or U9963 (N_9963,N_8860,N_8230);
nand U9964 (N_9964,N_8878,N_8123);
nand U9965 (N_9965,N_8655,N_8672);
or U9966 (N_9966,N_8624,N_8854);
nand U9967 (N_9967,N_8113,N_8697);
nor U9968 (N_9968,N_8817,N_8440);
nor U9969 (N_9969,N_8800,N_8194);
xnor U9970 (N_9970,N_8254,N_8630);
nor U9971 (N_9971,N_8945,N_8814);
and U9972 (N_9972,N_8385,N_8288);
or U9973 (N_9973,N_8918,N_8534);
xnor U9974 (N_9974,N_8925,N_8186);
xor U9975 (N_9975,N_8231,N_8826);
nand U9976 (N_9976,N_8024,N_8022);
nor U9977 (N_9977,N_8168,N_8666);
xor U9978 (N_9978,N_8675,N_8691);
and U9979 (N_9979,N_8902,N_8064);
xnor U9980 (N_9980,N_8429,N_8439);
nand U9981 (N_9981,N_8965,N_8151);
nand U9982 (N_9982,N_8475,N_8421);
and U9983 (N_9983,N_8140,N_8432);
nand U9984 (N_9984,N_8196,N_8603);
and U9985 (N_9985,N_8156,N_8524);
and U9986 (N_9986,N_8428,N_8522);
nand U9987 (N_9987,N_8647,N_8334);
or U9988 (N_9988,N_8568,N_8876);
xor U9989 (N_9989,N_8414,N_8160);
nor U9990 (N_9990,N_8626,N_8522);
and U9991 (N_9991,N_8558,N_8394);
or U9992 (N_9992,N_8234,N_8111);
nand U9993 (N_9993,N_8973,N_8022);
nand U9994 (N_9994,N_8048,N_8727);
xnor U9995 (N_9995,N_8889,N_8745);
nor U9996 (N_9996,N_8279,N_8989);
xor U9997 (N_9997,N_8150,N_8479);
nand U9998 (N_9998,N_8653,N_8168);
xnor U9999 (N_9999,N_8976,N_8942);
nor U10000 (N_10000,N_9102,N_9639);
and U10001 (N_10001,N_9426,N_9301);
nor U10002 (N_10002,N_9405,N_9083);
or U10003 (N_10003,N_9131,N_9836);
xnor U10004 (N_10004,N_9975,N_9423);
nor U10005 (N_10005,N_9759,N_9197);
or U10006 (N_10006,N_9464,N_9659);
xnor U10007 (N_10007,N_9498,N_9284);
and U10008 (N_10008,N_9551,N_9000);
and U10009 (N_10009,N_9973,N_9809);
and U10010 (N_10010,N_9762,N_9242);
and U10011 (N_10011,N_9654,N_9957);
nor U10012 (N_10012,N_9215,N_9448);
or U10013 (N_10013,N_9271,N_9731);
and U10014 (N_10014,N_9704,N_9564);
or U10015 (N_10015,N_9141,N_9336);
nand U10016 (N_10016,N_9670,N_9646);
or U10017 (N_10017,N_9502,N_9875);
or U10018 (N_10018,N_9992,N_9458);
xnor U10019 (N_10019,N_9989,N_9770);
xnor U10020 (N_10020,N_9800,N_9283);
and U10021 (N_10021,N_9309,N_9560);
or U10022 (N_10022,N_9016,N_9643);
xnor U10023 (N_10023,N_9999,N_9298);
xnor U10024 (N_10024,N_9287,N_9549);
xnor U10025 (N_10025,N_9321,N_9281);
and U10026 (N_10026,N_9700,N_9982);
nand U10027 (N_10027,N_9915,N_9447);
nand U10028 (N_10028,N_9419,N_9618);
and U10029 (N_10029,N_9246,N_9668);
and U10030 (N_10030,N_9760,N_9345);
nand U10031 (N_10031,N_9615,N_9944);
nor U10032 (N_10032,N_9289,N_9100);
and U10033 (N_10033,N_9075,N_9721);
or U10034 (N_10034,N_9471,N_9767);
xor U10035 (N_10035,N_9182,N_9825);
nand U10036 (N_10036,N_9511,N_9185);
xor U10037 (N_10037,N_9755,N_9389);
xnor U10038 (N_10038,N_9358,N_9941);
nand U10039 (N_10039,N_9793,N_9814);
nand U10040 (N_10040,N_9877,N_9276);
nor U10041 (N_10041,N_9572,N_9997);
xor U10042 (N_10042,N_9217,N_9592);
and U10043 (N_10043,N_9586,N_9637);
nand U10044 (N_10044,N_9921,N_9372);
xnor U10045 (N_10045,N_9487,N_9407);
nor U10046 (N_10046,N_9557,N_9077);
nand U10047 (N_10047,N_9518,N_9398);
and U10048 (N_10048,N_9765,N_9106);
or U10049 (N_10049,N_9418,N_9459);
or U10050 (N_10050,N_9203,N_9369);
or U10051 (N_10051,N_9515,N_9051);
or U10052 (N_10052,N_9621,N_9208);
nand U10053 (N_10053,N_9319,N_9130);
and U10054 (N_10054,N_9853,N_9881);
nor U10055 (N_10055,N_9323,N_9155);
xor U10056 (N_10056,N_9935,N_9544);
nor U10057 (N_10057,N_9777,N_9865);
and U10058 (N_10058,N_9540,N_9421);
and U10059 (N_10059,N_9678,N_9286);
xnor U10060 (N_10060,N_9085,N_9552);
nor U10061 (N_10061,N_9681,N_9205);
and U10062 (N_10062,N_9055,N_9375);
xnor U10063 (N_10063,N_9893,N_9521);
nor U10064 (N_10064,N_9835,N_9121);
nor U10065 (N_10065,N_9053,N_9742);
or U10066 (N_10066,N_9177,N_9348);
nand U10067 (N_10067,N_9711,N_9612);
and U10068 (N_10068,N_9910,N_9249);
nand U10069 (N_10069,N_9524,N_9829);
or U10070 (N_10070,N_9265,N_9847);
nand U10071 (N_10071,N_9917,N_9716);
nor U10072 (N_10072,N_9206,N_9529);
nand U10073 (N_10073,N_9134,N_9780);
nor U10074 (N_10074,N_9489,N_9707);
nand U10075 (N_10075,N_9382,N_9616);
nor U10076 (N_10076,N_9142,N_9124);
nor U10077 (N_10077,N_9528,N_9980);
nand U10078 (N_10078,N_9011,N_9555);
xor U10079 (N_10079,N_9280,N_9132);
or U10080 (N_10080,N_9031,N_9933);
nand U10081 (N_10081,N_9326,N_9725);
and U10082 (N_10082,N_9679,N_9923);
nand U10083 (N_10083,N_9516,N_9320);
nand U10084 (N_10084,N_9046,N_9505);
nand U10085 (N_10085,N_9173,N_9337);
and U10086 (N_10086,N_9507,N_9672);
or U10087 (N_10087,N_9532,N_9222);
and U10088 (N_10088,N_9066,N_9054);
nor U10089 (N_10089,N_9439,N_9690);
xnor U10090 (N_10090,N_9950,N_9786);
nand U10091 (N_10091,N_9109,N_9408);
nand U10092 (N_10092,N_9306,N_9894);
nand U10093 (N_10093,N_9671,N_9437);
xnor U10094 (N_10094,N_9480,N_9118);
or U10095 (N_10095,N_9037,N_9525);
or U10096 (N_10096,N_9484,N_9191);
or U10097 (N_10097,N_9390,N_9161);
xnor U10098 (N_10098,N_9949,N_9015);
nor U10099 (N_10099,N_9868,N_9261);
and U10100 (N_10100,N_9606,N_9899);
nor U10101 (N_10101,N_9019,N_9022);
or U10102 (N_10102,N_9535,N_9071);
xnor U10103 (N_10103,N_9684,N_9856);
nand U10104 (N_10104,N_9905,N_9870);
nor U10105 (N_10105,N_9597,N_9994);
nor U10106 (N_10106,N_9201,N_9329);
xnor U10107 (N_10107,N_9436,N_9682);
nand U10108 (N_10108,N_9635,N_9351);
or U10109 (N_10109,N_9137,N_9067);
nand U10110 (N_10110,N_9686,N_9673);
nand U10111 (N_10111,N_9582,N_9244);
or U10112 (N_10112,N_9932,N_9315);
nand U10113 (N_10113,N_9730,N_9526);
and U10114 (N_10114,N_9154,N_9479);
or U10115 (N_10115,N_9900,N_9955);
nand U10116 (N_10116,N_9231,N_9113);
nor U10117 (N_10117,N_9744,N_9602);
or U10118 (N_10118,N_9661,N_9338);
nor U10119 (N_10119,N_9769,N_9070);
nor U10120 (N_10120,N_9831,N_9514);
nor U10121 (N_10121,N_9429,N_9775);
nand U10122 (N_10122,N_9928,N_9198);
nand U10123 (N_10123,N_9709,N_9761);
nor U10124 (N_10124,N_9939,N_9539);
and U10125 (N_10125,N_9773,N_9492);
and U10126 (N_10126,N_9237,N_9962);
nor U10127 (N_10127,N_9171,N_9813);
or U10128 (N_10128,N_9743,N_9675);
nand U10129 (N_10129,N_9463,N_9342);
xnor U10130 (N_10130,N_9963,N_9209);
nor U10131 (N_10131,N_9260,N_9702);
nand U10132 (N_10132,N_9974,N_9397);
and U10133 (N_10133,N_9501,N_9895);
nand U10134 (N_10134,N_9359,N_9763);
and U10135 (N_10135,N_9826,N_9241);
xor U10136 (N_10136,N_9849,N_9293);
and U10137 (N_10137,N_9512,N_9680);
or U10138 (N_10138,N_9566,N_9772);
and U10139 (N_10139,N_9435,N_9629);
nor U10140 (N_10140,N_9691,N_9737);
xor U10141 (N_10141,N_9259,N_9354);
and U10142 (N_10142,N_9032,N_9490);
or U10143 (N_10143,N_9753,N_9158);
or U10144 (N_10144,N_9757,N_9713);
or U10145 (N_10145,N_9240,N_9416);
or U10146 (N_10146,N_9993,N_9936);
or U10147 (N_10147,N_9349,N_9653);
and U10148 (N_10148,N_9537,N_9225);
nand U10149 (N_10149,N_9114,N_9656);
xor U10150 (N_10150,N_9530,N_9050);
and U10151 (N_10151,N_9004,N_9147);
nor U10152 (N_10152,N_9491,N_9331);
or U10153 (N_10153,N_9367,N_9876);
xor U10154 (N_10154,N_9655,N_9802);
nor U10155 (N_10155,N_9285,N_9837);
nor U10156 (N_10156,N_9226,N_9676);
or U10157 (N_10157,N_9563,N_9127);
nor U10158 (N_10158,N_9495,N_9277);
nand U10159 (N_10159,N_9882,N_9396);
xnor U10160 (N_10160,N_9091,N_9860);
and U10161 (N_10161,N_9116,N_9694);
nand U10162 (N_10162,N_9040,N_9228);
nor U10163 (N_10163,N_9609,N_9219);
nand U10164 (N_10164,N_9985,N_9726);
or U10165 (N_10165,N_9090,N_9188);
nand U10166 (N_10166,N_9181,N_9698);
xnor U10167 (N_10167,N_9977,N_9754);
xnor U10168 (N_10168,N_9043,N_9454);
xnor U10169 (N_10169,N_9446,N_9749);
nor U10170 (N_10170,N_9376,N_9233);
or U10171 (N_10171,N_9048,N_9556);
or U10172 (N_10172,N_9189,N_9162);
or U10173 (N_10173,N_9916,N_9787);
and U10174 (N_10174,N_9522,N_9169);
or U10175 (N_10175,N_9801,N_9630);
nor U10176 (N_10176,N_9662,N_9224);
xnor U10177 (N_10177,N_9442,N_9045);
nand U10178 (N_10178,N_9862,N_9341);
nor U10179 (N_10179,N_9821,N_9604);
nand U10180 (N_10180,N_9568,N_9449);
xor U10181 (N_10181,N_9776,N_9445);
nand U10182 (N_10182,N_9105,N_9346);
or U10183 (N_10183,N_9677,N_9569);
and U10184 (N_10184,N_9632,N_9296);
nor U10185 (N_10185,N_9290,N_9715);
or U10186 (N_10186,N_9558,N_9039);
and U10187 (N_10187,N_9506,N_9892);
or U10188 (N_10188,N_9305,N_9194);
or U10189 (N_10189,N_9256,N_9424);
xnor U10190 (N_10190,N_9819,N_9510);
or U10191 (N_10191,N_9650,N_9006);
nand U10192 (N_10192,N_9692,N_9781);
nand U10193 (N_10193,N_9697,N_9545);
nor U10194 (N_10194,N_9712,N_9808);
and U10195 (N_10195,N_9991,N_9804);
or U10196 (N_10196,N_9144,N_9394);
nor U10197 (N_10197,N_9660,N_9574);
nor U10198 (N_10198,N_9546,N_9473);
nor U10199 (N_10199,N_9764,N_9842);
xor U10200 (N_10200,N_9029,N_9168);
nor U10201 (N_10201,N_9232,N_9968);
nor U10202 (N_10202,N_9014,N_9462);
or U10203 (N_10203,N_9561,N_9990);
or U10204 (N_10204,N_9806,N_9403);
nor U10205 (N_10205,N_9184,N_9344);
nor U10206 (N_10206,N_9562,N_9373);
or U10207 (N_10207,N_9214,N_9410);
nand U10208 (N_10208,N_9095,N_9746);
or U10209 (N_10209,N_9890,N_9844);
xnor U10210 (N_10210,N_9828,N_9385);
nand U10211 (N_10211,N_9701,N_9363);
or U10212 (N_10212,N_9607,N_9553);
nor U10213 (N_10213,N_9135,N_9380);
nor U10214 (N_10214,N_9140,N_9571);
nand U10215 (N_10215,N_9911,N_9057);
and U10216 (N_10216,N_9620,N_9047);
nor U10217 (N_10217,N_9628,N_9428);
or U10218 (N_10218,N_9115,N_9976);
and U10219 (N_10219,N_9878,N_9583);
and U10220 (N_10220,N_9024,N_9758);
or U10221 (N_10221,N_9797,N_9611);
xor U10222 (N_10222,N_9920,N_9509);
nand U10223 (N_10223,N_9248,N_9598);
xnor U10224 (N_10224,N_9013,N_9883);
or U10225 (N_10225,N_9745,N_9710);
and U10226 (N_10226,N_9961,N_9603);
and U10227 (N_10227,N_9782,N_9577);
or U10228 (N_10228,N_9379,N_9295);
nor U10229 (N_10229,N_9404,N_9978);
nor U10230 (N_10230,N_9665,N_9347);
and U10231 (N_10231,N_9596,N_9508);
xor U10232 (N_10232,N_9452,N_9120);
or U10233 (N_10233,N_9239,N_9266);
xnor U10234 (N_10234,N_9401,N_9695);
nand U10235 (N_10235,N_9001,N_9311);
xor U10236 (N_10236,N_9064,N_9584);
and U10237 (N_10237,N_9438,N_9310);
or U10238 (N_10238,N_9388,N_9093);
nand U10239 (N_10239,N_9965,N_9898);
or U10240 (N_10240,N_9523,N_9970);
xor U10241 (N_10241,N_9366,N_9693);
xor U10242 (N_10242,N_9417,N_9030);
or U10243 (N_10243,N_9934,N_9183);
or U10244 (N_10244,N_9420,N_9292);
and U10245 (N_10245,N_9250,N_9617);
or U10246 (N_10246,N_9807,N_9193);
nor U10247 (N_10247,N_9778,N_9061);
xor U10248 (N_10248,N_9475,N_9128);
and U10249 (N_10249,N_9003,N_9470);
nand U10250 (N_10250,N_9841,N_9930);
nand U10251 (N_10251,N_9430,N_9392);
and U10252 (N_10252,N_9187,N_9444);
or U10253 (N_10253,N_9575,N_9111);
xor U10254 (N_10254,N_9062,N_9307);
nand U10255 (N_10255,N_9594,N_9328);
and U10256 (N_10256,N_9204,N_9322);
nor U10257 (N_10257,N_9925,N_9335);
and U10258 (N_10258,N_9815,N_9790);
and U10259 (N_10259,N_9708,N_9145);
nor U10260 (N_10260,N_9059,N_9488);
or U10261 (N_10261,N_9149,N_9952);
nand U10262 (N_10262,N_9631,N_9822);
nand U10263 (N_10263,N_9267,N_9441);
nor U10264 (N_10264,N_9610,N_9263);
nor U10265 (N_10265,N_9252,N_9588);
nor U10266 (N_10266,N_9496,N_9967);
nor U10267 (N_10267,N_9199,N_9723);
and U10268 (N_10268,N_9550,N_9919);
or U10269 (N_10269,N_9450,N_9159);
xor U10270 (N_10270,N_9986,N_9590);
xor U10271 (N_10271,N_9247,N_9794);
nor U10272 (N_10272,N_9235,N_9689);
or U10273 (N_10273,N_9422,N_9908);
xor U10274 (N_10274,N_9025,N_9133);
or U10275 (N_10275,N_9089,N_9626);
xor U10276 (N_10276,N_9481,N_9129);
xor U10277 (N_10277,N_9954,N_9174);
and U10278 (N_10278,N_9034,N_9350);
and U10279 (N_10279,N_9839,N_9356);
xor U10280 (N_10280,N_9288,N_9150);
nand U10281 (N_10281,N_9669,N_9112);
or U10282 (N_10282,N_9705,N_9042);
or U10283 (N_10283,N_9666,N_9579);
nor U10284 (N_10284,N_9190,N_9352);
and U10285 (N_10285,N_9735,N_9451);
and U10286 (N_10286,N_9472,N_9827);
nand U10287 (N_10287,N_9431,N_9327);
or U10288 (N_10288,N_9078,N_9859);
nor U10289 (N_10289,N_9253,N_9624);
nand U10290 (N_10290,N_9212,N_9258);
and U10291 (N_10291,N_9278,N_9068);
nand U10292 (N_10292,N_9645,N_9817);
nand U10293 (N_10293,N_9768,N_9370);
nand U10294 (N_10294,N_9541,N_9476);
nor U10295 (N_10295,N_9573,N_9732);
nor U10296 (N_10296,N_9805,N_9803);
or U10297 (N_10297,N_9152,N_9866);
nor U10298 (N_10298,N_9427,N_9474);
nor U10299 (N_10299,N_9838,N_9160);
xnor U10300 (N_10300,N_9519,N_9361);
or U10301 (N_10301,N_9718,N_9937);
xnor U10302 (N_10302,N_9383,N_9414);
or U10303 (N_10303,N_9196,N_9663);
nor U10304 (N_10304,N_9657,N_9387);
xor U10305 (N_10305,N_9739,N_9503);
and U10306 (N_10306,N_9736,N_9172);
or U10307 (N_10307,N_9056,N_9374);
nor U10308 (N_10308,N_9642,N_9227);
or U10309 (N_10309,N_9845,N_9833);
and U10310 (N_10310,N_9084,N_9906);
or U10311 (N_10311,N_9931,N_9125);
or U10312 (N_10312,N_9180,N_9334);
nor U10313 (N_10313,N_9998,N_9789);
xnor U10314 (N_10314,N_9685,N_9909);
nand U10315 (N_10315,N_9904,N_9981);
xor U10316 (N_10316,N_9148,N_9362);
nor U10317 (N_10317,N_9186,N_9852);
nand U10318 (N_10318,N_9343,N_9581);
xor U10319 (N_10319,N_9493,N_9094);
nand U10320 (N_10320,N_9696,N_9411);
nand U10321 (N_10321,N_9948,N_9634);
and U10322 (N_10322,N_9674,N_9072);
or U10323 (N_10323,N_9297,N_9733);
nand U10324 (N_10324,N_9080,N_9706);
or U10325 (N_10325,N_9220,N_9213);
nand U10326 (N_10326,N_9126,N_9221);
nor U10327 (N_10327,N_9440,N_9167);
and U10328 (N_10328,N_9254,N_9086);
nor U10329 (N_10329,N_9783,N_9457);
and U10330 (N_10330,N_9924,N_9536);
xor U10331 (N_10331,N_9947,N_9069);
nor U10332 (N_10332,N_9399,N_9863);
nor U10333 (N_10333,N_9216,N_9966);
nand U10334 (N_10334,N_9302,N_9339);
nand U10335 (N_10335,N_9156,N_9432);
xor U10336 (N_10336,N_9104,N_9547);
xnor U10337 (N_10337,N_9779,N_9896);
and U10338 (N_10338,N_9262,N_9243);
and U10339 (N_10339,N_9751,N_9058);
or U10340 (N_10340,N_9230,N_9840);
or U10341 (N_10341,N_9788,N_9103);
nor U10342 (N_10342,N_9887,N_9644);
or U10343 (N_10343,N_9945,N_9633);
nand U10344 (N_10344,N_9638,N_9035);
xnor U10345 (N_10345,N_9591,N_9163);
and U10346 (N_10346,N_9625,N_9282);
xnor U10347 (N_10347,N_9494,N_9752);
nor U10348 (N_10348,N_9667,N_9333);
and U10349 (N_10349,N_9500,N_9409);
nor U10350 (N_10350,N_9640,N_9088);
nor U10351 (N_10351,N_9018,N_9810);
and U10352 (N_10352,N_9234,N_9874);
or U10353 (N_10353,N_9303,N_9818);
xor U10354 (N_10354,N_9122,N_9565);
and U10355 (N_10355,N_9504,N_9720);
nor U10356 (N_10356,N_9060,N_9143);
nand U10357 (N_10357,N_9812,N_9867);
or U10358 (N_10358,N_9178,N_9330);
xnor U10359 (N_10359,N_9273,N_9959);
and U10360 (N_10360,N_9792,N_9434);
and U10361 (N_10361,N_9317,N_9264);
and U10362 (N_10362,N_9005,N_9593);
or U10363 (N_10363,N_9741,N_9082);
nand U10364 (N_10364,N_9117,N_9938);
xnor U10365 (N_10365,N_9728,N_9613);
nand U10366 (N_10366,N_9360,N_9649);
xnor U10367 (N_10367,N_9605,N_9533);
nand U10368 (N_10368,N_9497,N_9846);
nor U10369 (N_10369,N_9798,N_9049);
nor U10370 (N_10370,N_9785,N_9983);
nor U10371 (N_10371,N_9008,N_9795);
nand U10372 (N_10372,N_9816,N_9651);
and U10373 (N_10373,N_9926,N_9869);
or U10374 (N_10374,N_9984,N_9520);
or U10375 (N_10375,N_9554,N_9052);
and U10376 (N_10376,N_9110,N_9195);
xnor U10377 (N_10377,N_9517,N_9873);
or U10378 (N_10378,N_9238,N_9272);
and U10379 (N_10379,N_9340,N_9157);
nor U10380 (N_10380,N_9477,N_9153);
and U10381 (N_10381,N_9857,N_9542);
xnor U10382 (N_10382,N_9799,N_9165);
xnor U10383 (N_10383,N_9766,N_9922);
nor U10384 (N_10384,N_9063,N_9461);
nand U10385 (N_10385,N_9811,N_9318);
nand U10386 (N_10386,N_9466,N_9848);
xnor U10387 (N_10387,N_9903,N_9325);
and U10388 (N_10388,N_9996,N_9960);
or U10389 (N_10389,N_9146,N_9969);
nor U10390 (N_10390,N_9824,N_9176);
and U10391 (N_10391,N_9026,N_9384);
or U10392 (N_10392,N_9096,N_9245);
or U10393 (N_10393,N_9854,N_9534);
and U10394 (N_10394,N_9098,N_9527);
nor U10395 (N_10395,N_9608,N_9717);
xor U10396 (N_10396,N_9170,N_9038);
nand U10397 (N_10397,N_9433,N_9559);
or U10398 (N_10398,N_9740,N_9469);
or U10399 (N_10399,N_9299,N_9028);
and U10400 (N_10400,N_9951,N_9714);
or U10401 (N_10401,N_9478,N_9304);
and U10402 (N_10402,N_9294,N_9099);
or U10403 (N_10403,N_9291,N_9179);
xor U10404 (N_10404,N_9065,N_9907);
nand U10405 (N_10405,N_9738,N_9465);
nand U10406 (N_10406,N_9269,N_9901);
xor U10407 (N_10407,N_9499,N_9332);
and U10408 (N_10408,N_9929,N_9614);
nand U10409 (N_10409,N_9316,N_9368);
xnor U10410 (N_10410,N_9017,N_9097);
nor U10411 (N_10411,N_9223,N_9324);
or U10412 (N_10412,N_9425,N_9402);
or U10413 (N_10413,N_9871,N_9943);
or U10414 (N_10414,N_9381,N_9756);
and U10415 (N_10415,N_9688,N_9400);
and U10416 (N_10416,N_9884,N_9192);
xor U10417 (N_10417,N_9988,N_9007);
or U10418 (N_10418,N_9886,N_9257);
nor U10419 (N_10419,N_9880,N_9636);
and U10420 (N_10420,N_9371,N_9207);
xor U10421 (N_10421,N_9995,N_9843);
xor U10422 (N_10422,N_9851,N_9251);
or U10423 (N_10423,N_9164,N_9543);
xnor U10424 (N_10424,N_9531,N_9119);
and U10425 (N_10425,N_9589,N_9443);
nand U10426 (N_10426,N_9601,N_9580);
or U10427 (N_10427,N_9623,N_9699);
nand U10428 (N_10428,N_9958,N_9734);
nor U10429 (N_10429,N_9724,N_9964);
nand U10430 (N_10430,N_9002,N_9748);
nand U10431 (N_10431,N_9079,N_9455);
xnor U10432 (N_10432,N_9619,N_9622);
nor U10433 (N_10433,N_9912,N_9771);
nor U10434 (N_10434,N_9585,N_9703);
nor U10435 (N_10435,N_9483,N_9010);
xor U10436 (N_10436,N_9942,N_9467);
nor U10437 (N_10437,N_9415,N_9312);
or U10438 (N_10438,N_9485,N_9855);
xor U10439 (N_10439,N_9888,N_9365);
or U10440 (N_10440,N_9940,N_9587);
or U10441 (N_10441,N_9274,N_9138);
and U10442 (N_10442,N_9123,N_9393);
nor U10443 (N_10443,N_9953,N_9395);
or U10444 (N_10444,N_9687,N_9987);
nand U10445 (N_10445,N_9576,N_9861);
and U10446 (N_10446,N_9313,N_9073);
and U10447 (N_10447,N_9600,N_9979);
or U10448 (N_10448,N_9377,N_9453);
xor U10449 (N_10449,N_9486,N_9664);
and U10450 (N_10450,N_9791,N_9218);
or U10451 (N_10451,N_9850,N_9567);
xor U10452 (N_10452,N_9044,N_9750);
nand U10453 (N_10453,N_9236,N_9784);
xnor U10454 (N_10454,N_9482,N_9308);
and U10455 (N_10455,N_9413,N_9041);
and U10456 (N_10456,N_9087,N_9971);
and U10457 (N_10457,N_9175,N_9074);
and U10458 (N_10458,N_9027,N_9627);
or U10459 (N_10459,N_9012,N_9658);
nand U10460 (N_10460,N_9946,N_9020);
xnor U10461 (N_10461,N_9747,N_9683);
nor U10462 (N_10462,N_9139,N_9364);
xnor U10463 (N_10463,N_9823,N_9548);
nor U10464 (N_10464,N_9538,N_9355);
and U10465 (N_10465,N_9647,N_9386);
nand U10466 (N_10466,N_9889,N_9009);
nor U10467 (N_10467,N_9151,N_9595);
xnor U10468 (N_10468,N_9719,N_9406);
and U10469 (N_10469,N_9314,N_9864);
or U10470 (N_10470,N_9202,N_9200);
or U10471 (N_10471,N_9378,N_9972);
nand U10472 (N_10472,N_9460,N_9641);
nor U10473 (N_10473,N_9570,N_9108);
and U10474 (N_10474,N_9210,N_9820);
xor U10475 (N_10475,N_9101,N_9391);
nand U10476 (N_10476,N_9902,N_9353);
nand U10477 (N_10477,N_9913,N_9255);
or U10478 (N_10478,N_9578,N_9107);
nand U10479 (N_10479,N_9357,N_9796);
nand U10480 (N_10480,N_9279,N_9858);
nor U10481 (N_10481,N_9023,N_9136);
nand U10482 (N_10482,N_9648,N_9918);
and U10483 (N_10483,N_9456,N_9897);
nand U10484 (N_10484,N_9081,N_9832);
nand U10485 (N_10485,N_9727,N_9033);
or U10486 (N_10486,N_9872,N_9891);
nor U10487 (N_10487,N_9275,N_9599);
or U10488 (N_10488,N_9300,N_9722);
or U10489 (N_10489,N_9036,N_9076);
xnor U10490 (N_10490,N_9412,N_9834);
nor U10491 (N_10491,N_9885,N_9774);
or U10492 (N_10492,N_9211,N_9268);
nand U10493 (N_10493,N_9956,N_9166);
and U10494 (N_10494,N_9513,N_9229);
nor U10495 (N_10495,N_9092,N_9468);
and U10496 (N_10496,N_9021,N_9830);
and U10497 (N_10497,N_9652,N_9270);
and U10498 (N_10498,N_9879,N_9729);
or U10499 (N_10499,N_9914,N_9927);
and U10500 (N_10500,N_9574,N_9882);
nand U10501 (N_10501,N_9915,N_9686);
nand U10502 (N_10502,N_9324,N_9381);
nor U10503 (N_10503,N_9491,N_9425);
nor U10504 (N_10504,N_9834,N_9340);
nand U10505 (N_10505,N_9412,N_9352);
and U10506 (N_10506,N_9121,N_9621);
nor U10507 (N_10507,N_9191,N_9902);
or U10508 (N_10508,N_9435,N_9863);
and U10509 (N_10509,N_9737,N_9254);
xor U10510 (N_10510,N_9370,N_9944);
nand U10511 (N_10511,N_9044,N_9770);
nand U10512 (N_10512,N_9549,N_9114);
nand U10513 (N_10513,N_9127,N_9182);
or U10514 (N_10514,N_9797,N_9253);
or U10515 (N_10515,N_9916,N_9289);
and U10516 (N_10516,N_9090,N_9314);
nand U10517 (N_10517,N_9059,N_9327);
nor U10518 (N_10518,N_9810,N_9833);
nand U10519 (N_10519,N_9098,N_9597);
and U10520 (N_10520,N_9709,N_9233);
or U10521 (N_10521,N_9954,N_9372);
and U10522 (N_10522,N_9641,N_9611);
or U10523 (N_10523,N_9779,N_9970);
nand U10524 (N_10524,N_9229,N_9577);
and U10525 (N_10525,N_9623,N_9875);
nor U10526 (N_10526,N_9934,N_9331);
nand U10527 (N_10527,N_9008,N_9625);
nor U10528 (N_10528,N_9217,N_9469);
xnor U10529 (N_10529,N_9883,N_9288);
nand U10530 (N_10530,N_9793,N_9243);
nand U10531 (N_10531,N_9050,N_9645);
nand U10532 (N_10532,N_9189,N_9891);
and U10533 (N_10533,N_9821,N_9497);
or U10534 (N_10534,N_9556,N_9540);
or U10535 (N_10535,N_9340,N_9694);
nor U10536 (N_10536,N_9979,N_9174);
xor U10537 (N_10537,N_9456,N_9885);
and U10538 (N_10538,N_9073,N_9701);
nand U10539 (N_10539,N_9346,N_9762);
nand U10540 (N_10540,N_9885,N_9924);
xor U10541 (N_10541,N_9141,N_9879);
or U10542 (N_10542,N_9233,N_9673);
nand U10543 (N_10543,N_9922,N_9737);
or U10544 (N_10544,N_9681,N_9528);
and U10545 (N_10545,N_9615,N_9398);
or U10546 (N_10546,N_9330,N_9087);
nor U10547 (N_10547,N_9981,N_9736);
and U10548 (N_10548,N_9184,N_9476);
and U10549 (N_10549,N_9878,N_9988);
or U10550 (N_10550,N_9591,N_9791);
and U10551 (N_10551,N_9967,N_9415);
and U10552 (N_10552,N_9350,N_9259);
xnor U10553 (N_10553,N_9375,N_9639);
or U10554 (N_10554,N_9620,N_9533);
and U10555 (N_10555,N_9526,N_9356);
nor U10556 (N_10556,N_9890,N_9901);
nand U10557 (N_10557,N_9292,N_9129);
or U10558 (N_10558,N_9217,N_9507);
nand U10559 (N_10559,N_9797,N_9351);
xor U10560 (N_10560,N_9381,N_9904);
xor U10561 (N_10561,N_9332,N_9149);
xor U10562 (N_10562,N_9750,N_9781);
nand U10563 (N_10563,N_9820,N_9520);
xnor U10564 (N_10564,N_9042,N_9288);
nand U10565 (N_10565,N_9344,N_9895);
nor U10566 (N_10566,N_9814,N_9739);
or U10567 (N_10567,N_9611,N_9031);
and U10568 (N_10568,N_9272,N_9153);
xor U10569 (N_10569,N_9349,N_9607);
nand U10570 (N_10570,N_9781,N_9992);
or U10571 (N_10571,N_9027,N_9024);
nor U10572 (N_10572,N_9313,N_9143);
nand U10573 (N_10573,N_9791,N_9906);
or U10574 (N_10574,N_9484,N_9701);
xor U10575 (N_10575,N_9790,N_9488);
nand U10576 (N_10576,N_9682,N_9080);
nand U10577 (N_10577,N_9046,N_9655);
xnor U10578 (N_10578,N_9498,N_9254);
or U10579 (N_10579,N_9083,N_9912);
nor U10580 (N_10580,N_9235,N_9007);
nand U10581 (N_10581,N_9750,N_9141);
xnor U10582 (N_10582,N_9916,N_9548);
and U10583 (N_10583,N_9671,N_9473);
or U10584 (N_10584,N_9418,N_9474);
nand U10585 (N_10585,N_9924,N_9753);
nor U10586 (N_10586,N_9557,N_9368);
nand U10587 (N_10587,N_9226,N_9126);
xnor U10588 (N_10588,N_9365,N_9501);
nand U10589 (N_10589,N_9136,N_9761);
and U10590 (N_10590,N_9491,N_9930);
xnor U10591 (N_10591,N_9024,N_9230);
nor U10592 (N_10592,N_9158,N_9917);
xor U10593 (N_10593,N_9020,N_9386);
or U10594 (N_10594,N_9576,N_9768);
and U10595 (N_10595,N_9589,N_9008);
or U10596 (N_10596,N_9252,N_9225);
and U10597 (N_10597,N_9465,N_9194);
nand U10598 (N_10598,N_9416,N_9336);
nand U10599 (N_10599,N_9915,N_9375);
nor U10600 (N_10600,N_9427,N_9328);
xnor U10601 (N_10601,N_9430,N_9611);
nand U10602 (N_10602,N_9622,N_9728);
and U10603 (N_10603,N_9881,N_9907);
nor U10604 (N_10604,N_9558,N_9780);
xor U10605 (N_10605,N_9156,N_9700);
xor U10606 (N_10606,N_9092,N_9810);
xnor U10607 (N_10607,N_9088,N_9631);
xor U10608 (N_10608,N_9576,N_9429);
nand U10609 (N_10609,N_9947,N_9513);
or U10610 (N_10610,N_9015,N_9034);
nor U10611 (N_10611,N_9141,N_9499);
nor U10612 (N_10612,N_9439,N_9676);
xor U10613 (N_10613,N_9661,N_9258);
nor U10614 (N_10614,N_9187,N_9189);
xor U10615 (N_10615,N_9400,N_9412);
and U10616 (N_10616,N_9275,N_9824);
and U10617 (N_10617,N_9867,N_9393);
nand U10618 (N_10618,N_9348,N_9411);
xnor U10619 (N_10619,N_9255,N_9367);
nor U10620 (N_10620,N_9235,N_9194);
nand U10621 (N_10621,N_9140,N_9685);
nand U10622 (N_10622,N_9197,N_9672);
nor U10623 (N_10623,N_9983,N_9561);
or U10624 (N_10624,N_9933,N_9495);
xnor U10625 (N_10625,N_9801,N_9269);
nand U10626 (N_10626,N_9601,N_9756);
and U10627 (N_10627,N_9376,N_9958);
and U10628 (N_10628,N_9960,N_9078);
xor U10629 (N_10629,N_9187,N_9143);
nor U10630 (N_10630,N_9124,N_9696);
and U10631 (N_10631,N_9981,N_9646);
and U10632 (N_10632,N_9492,N_9103);
and U10633 (N_10633,N_9263,N_9822);
and U10634 (N_10634,N_9357,N_9714);
nor U10635 (N_10635,N_9148,N_9587);
or U10636 (N_10636,N_9182,N_9826);
nor U10637 (N_10637,N_9670,N_9349);
nand U10638 (N_10638,N_9539,N_9973);
nor U10639 (N_10639,N_9720,N_9472);
or U10640 (N_10640,N_9397,N_9979);
and U10641 (N_10641,N_9633,N_9932);
and U10642 (N_10642,N_9751,N_9664);
nor U10643 (N_10643,N_9182,N_9121);
and U10644 (N_10644,N_9568,N_9308);
nor U10645 (N_10645,N_9484,N_9536);
or U10646 (N_10646,N_9829,N_9154);
and U10647 (N_10647,N_9552,N_9087);
and U10648 (N_10648,N_9187,N_9845);
xor U10649 (N_10649,N_9039,N_9902);
nand U10650 (N_10650,N_9332,N_9925);
nand U10651 (N_10651,N_9854,N_9051);
or U10652 (N_10652,N_9276,N_9014);
nand U10653 (N_10653,N_9476,N_9934);
and U10654 (N_10654,N_9497,N_9831);
xor U10655 (N_10655,N_9340,N_9382);
nor U10656 (N_10656,N_9298,N_9958);
and U10657 (N_10657,N_9200,N_9303);
or U10658 (N_10658,N_9046,N_9992);
and U10659 (N_10659,N_9963,N_9250);
nand U10660 (N_10660,N_9621,N_9700);
nand U10661 (N_10661,N_9885,N_9843);
or U10662 (N_10662,N_9332,N_9673);
xnor U10663 (N_10663,N_9776,N_9418);
xor U10664 (N_10664,N_9345,N_9662);
nor U10665 (N_10665,N_9781,N_9137);
nor U10666 (N_10666,N_9385,N_9763);
nor U10667 (N_10667,N_9773,N_9572);
or U10668 (N_10668,N_9502,N_9062);
and U10669 (N_10669,N_9933,N_9261);
and U10670 (N_10670,N_9138,N_9130);
and U10671 (N_10671,N_9554,N_9364);
and U10672 (N_10672,N_9202,N_9486);
or U10673 (N_10673,N_9514,N_9499);
and U10674 (N_10674,N_9273,N_9005);
xnor U10675 (N_10675,N_9293,N_9007);
and U10676 (N_10676,N_9240,N_9875);
nand U10677 (N_10677,N_9788,N_9113);
nor U10678 (N_10678,N_9087,N_9423);
nor U10679 (N_10679,N_9317,N_9078);
nor U10680 (N_10680,N_9124,N_9567);
and U10681 (N_10681,N_9949,N_9650);
nand U10682 (N_10682,N_9714,N_9943);
xor U10683 (N_10683,N_9026,N_9227);
or U10684 (N_10684,N_9816,N_9287);
or U10685 (N_10685,N_9867,N_9794);
nand U10686 (N_10686,N_9218,N_9201);
nand U10687 (N_10687,N_9699,N_9598);
nor U10688 (N_10688,N_9269,N_9468);
and U10689 (N_10689,N_9694,N_9578);
and U10690 (N_10690,N_9539,N_9330);
and U10691 (N_10691,N_9838,N_9733);
or U10692 (N_10692,N_9313,N_9695);
nor U10693 (N_10693,N_9318,N_9178);
or U10694 (N_10694,N_9527,N_9589);
nor U10695 (N_10695,N_9369,N_9946);
xnor U10696 (N_10696,N_9425,N_9462);
or U10697 (N_10697,N_9941,N_9873);
xor U10698 (N_10698,N_9095,N_9119);
xnor U10699 (N_10699,N_9648,N_9035);
or U10700 (N_10700,N_9791,N_9787);
xnor U10701 (N_10701,N_9669,N_9270);
nor U10702 (N_10702,N_9762,N_9855);
and U10703 (N_10703,N_9862,N_9066);
or U10704 (N_10704,N_9935,N_9554);
xnor U10705 (N_10705,N_9445,N_9766);
nor U10706 (N_10706,N_9266,N_9878);
xnor U10707 (N_10707,N_9812,N_9130);
nor U10708 (N_10708,N_9420,N_9429);
nor U10709 (N_10709,N_9130,N_9956);
or U10710 (N_10710,N_9911,N_9791);
nand U10711 (N_10711,N_9310,N_9072);
nor U10712 (N_10712,N_9212,N_9668);
and U10713 (N_10713,N_9280,N_9633);
nor U10714 (N_10714,N_9458,N_9302);
and U10715 (N_10715,N_9668,N_9793);
or U10716 (N_10716,N_9957,N_9045);
or U10717 (N_10717,N_9961,N_9277);
nand U10718 (N_10718,N_9018,N_9601);
or U10719 (N_10719,N_9644,N_9775);
nor U10720 (N_10720,N_9328,N_9688);
and U10721 (N_10721,N_9143,N_9800);
and U10722 (N_10722,N_9259,N_9677);
or U10723 (N_10723,N_9303,N_9645);
xor U10724 (N_10724,N_9875,N_9282);
nor U10725 (N_10725,N_9032,N_9438);
nor U10726 (N_10726,N_9238,N_9172);
nor U10727 (N_10727,N_9162,N_9944);
or U10728 (N_10728,N_9868,N_9998);
or U10729 (N_10729,N_9983,N_9901);
nand U10730 (N_10730,N_9725,N_9066);
xor U10731 (N_10731,N_9521,N_9225);
and U10732 (N_10732,N_9815,N_9980);
nand U10733 (N_10733,N_9277,N_9320);
and U10734 (N_10734,N_9512,N_9758);
xor U10735 (N_10735,N_9454,N_9400);
nand U10736 (N_10736,N_9534,N_9364);
xnor U10737 (N_10737,N_9229,N_9137);
and U10738 (N_10738,N_9055,N_9607);
xor U10739 (N_10739,N_9213,N_9938);
xnor U10740 (N_10740,N_9825,N_9850);
xor U10741 (N_10741,N_9191,N_9827);
nor U10742 (N_10742,N_9191,N_9772);
nor U10743 (N_10743,N_9351,N_9235);
xnor U10744 (N_10744,N_9025,N_9874);
nor U10745 (N_10745,N_9592,N_9678);
and U10746 (N_10746,N_9545,N_9286);
and U10747 (N_10747,N_9142,N_9545);
nand U10748 (N_10748,N_9204,N_9782);
or U10749 (N_10749,N_9667,N_9960);
nand U10750 (N_10750,N_9289,N_9468);
nand U10751 (N_10751,N_9251,N_9218);
or U10752 (N_10752,N_9915,N_9948);
or U10753 (N_10753,N_9558,N_9463);
nand U10754 (N_10754,N_9575,N_9396);
and U10755 (N_10755,N_9391,N_9907);
xnor U10756 (N_10756,N_9509,N_9739);
and U10757 (N_10757,N_9653,N_9469);
and U10758 (N_10758,N_9572,N_9919);
nand U10759 (N_10759,N_9436,N_9153);
xnor U10760 (N_10760,N_9270,N_9269);
nor U10761 (N_10761,N_9368,N_9107);
xnor U10762 (N_10762,N_9322,N_9845);
nand U10763 (N_10763,N_9942,N_9851);
or U10764 (N_10764,N_9788,N_9844);
xnor U10765 (N_10765,N_9329,N_9370);
xnor U10766 (N_10766,N_9035,N_9533);
or U10767 (N_10767,N_9467,N_9868);
or U10768 (N_10768,N_9607,N_9911);
nor U10769 (N_10769,N_9969,N_9858);
or U10770 (N_10770,N_9373,N_9314);
xnor U10771 (N_10771,N_9135,N_9021);
or U10772 (N_10772,N_9713,N_9703);
nor U10773 (N_10773,N_9897,N_9375);
and U10774 (N_10774,N_9966,N_9421);
nor U10775 (N_10775,N_9378,N_9887);
nand U10776 (N_10776,N_9920,N_9646);
nor U10777 (N_10777,N_9255,N_9172);
nand U10778 (N_10778,N_9952,N_9686);
xor U10779 (N_10779,N_9961,N_9242);
nand U10780 (N_10780,N_9706,N_9319);
or U10781 (N_10781,N_9479,N_9494);
xnor U10782 (N_10782,N_9379,N_9772);
nand U10783 (N_10783,N_9793,N_9688);
and U10784 (N_10784,N_9036,N_9582);
or U10785 (N_10785,N_9177,N_9722);
nor U10786 (N_10786,N_9497,N_9724);
and U10787 (N_10787,N_9028,N_9841);
xor U10788 (N_10788,N_9781,N_9134);
xor U10789 (N_10789,N_9605,N_9590);
or U10790 (N_10790,N_9526,N_9049);
and U10791 (N_10791,N_9896,N_9163);
and U10792 (N_10792,N_9983,N_9593);
and U10793 (N_10793,N_9882,N_9414);
nor U10794 (N_10794,N_9105,N_9348);
nand U10795 (N_10795,N_9082,N_9952);
nor U10796 (N_10796,N_9686,N_9089);
nor U10797 (N_10797,N_9652,N_9650);
xnor U10798 (N_10798,N_9061,N_9303);
or U10799 (N_10799,N_9792,N_9001);
xnor U10800 (N_10800,N_9805,N_9836);
and U10801 (N_10801,N_9937,N_9626);
nand U10802 (N_10802,N_9765,N_9312);
nand U10803 (N_10803,N_9610,N_9494);
or U10804 (N_10804,N_9805,N_9957);
xor U10805 (N_10805,N_9906,N_9846);
or U10806 (N_10806,N_9104,N_9818);
nand U10807 (N_10807,N_9237,N_9828);
xnor U10808 (N_10808,N_9347,N_9509);
nand U10809 (N_10809,N_9418,N_9264);
and U10810 (N_10810,N_9868,N_9498);
nand U10811 (N_10811,N_9422,N_9381);
nand U10812 (N_10812,N_9491,N_9956);
nor U10813 (N_10813,N_9090,N_9250);
and U10814 (N_10814,N_9427,N_9833);
xnor U10815 (N_10815,N_9480,N_9856);
or U10816 (N_10816,N_9230,N_9996);
nor U10817 (N_10817,N_9441,N_9009);
and U10818 (N_10818,N_9748,N_9667);
or U10819 (N_10819,N_9453,N_9704);
and U10820 (N_10820,N_9078,N_9041);
nand U10821 (N_10821,N_9016,N_9490);
xor U10822 (N_10822,N_9922,N_9779);
and U10823 (N_10823,N_9423,N_9306);
and U10824 (N_10824,N_9598,N_9720);
or U10825 (N_10825,N_9764,N_9850);
nand U10826 (N_10826,N_9501,N_9872);
or U10827 (N_10827,N_9792,N_9549);
nand U10828 (N_10828,N_9532,N_9745);
or U10829 (N_10829,N_9072,N_9800);
nor U10830 (N_10830,N_9119,N_9480);
nand U10831 (N_10831,N_9668,N_9339);
xor U10832 (N_10832,N_9973,N_9091);
nand U10833 (N_10833,N_9446,N_9625);
or U10834 (N_10834,N_9371,N_9087);
or U10835 (N_10835,N_9387,N_9806);
nor U10836 (N_10836,N_9333,N_9172);
nor U10837 (N_10837,N_9516,N_9641);
and U10838 (N_10838,N_9493,N_9386);
or U10839 (N_10839,N_9863,N_9917);
nor U10840 (N_10840,N_9462,N_9983);
xor U10841 (N_10841,N_9027,N_9125);
nand U10842 (N_10842,N_9280,N_9344);
xor U10843 (N_10843,N_9522,N_9937);
and U10844 (N_10844,N_9881,N_9809);
and U10845 (N_10845,N_9871,N_9361);
nor U10846 (N_10846,N_9675,N_9731);
nor U10847 (N_10847,N_9818,N_9508);
and U10848 (N_10848,N_9924,N_9509);
and U10849 (N_10849,N_9137,N_9876);
or U10850 (N_10850,N_9574,N_9444);
or U10851 (N_10851,N_9141,N_9894);
and U10852 (N_10852,N_9122,N_9855);
and U10853 (N_10853,N_9944,N_9599);
nor U10854 (N_10854,N_9249,N_9340);
and U10855 (N_10855,N_9662,N_9737);
and U10856 (N_10856,N_9031,N_9555);
and U10857 (N_10857,N_9841,N_9837);
or U10858 (N_10858,N_9246,N_9225);
or U10859 (N_10859,N_9193,N_9247);
and U10860 (N_10860,N_9347,N_9274);
or U10861 (N_10861,N_9728,N_9616);
nand U10862 (N_10862,N_9989,N_9175);
xnor U10863 (N_10863,N_9558,N_9636);
xor U10864 (N_10864,N_9651,N_9993);
or U10865 (N_10865,N_9370,N_9265);
and U10866 (N_10866,N_9877,N_9378);
nor U10867 (N_10867,N_9356,N_9495);
and U10868 (N_10868,N_9585,N_9467);
nand U10869 (N_10869,N_9711,N_9577);
xnor U10870 (N_10870,N_9710,N_9327);
and U10871 (N_10871,N_9571,N_9520);
or U10872 (N_10872,N_9459,N_9558);
nand U10873 (N_10873,N_9249,N_9958);
or U10874 (N_10874,N_9786,N_9082);
xor U10875 (N_10875,N_9545,N_9588);
xnor U10876 (N_10876,N_9359,N_9535);
nand U10877 (N_10877,N_9636,N_9186);
xnor U10878 (N_10878,N_9093,N_9133);
xor U10879 (N_10879,N_9129,N_9511);
or U10880 (N_10880,N_9593,N_9764);
or U10881 (N_10881,N_9056,N_9021);
and U10882 (N_10882,N_9209,N_9165);
and U10883 (N_10883,N_9710,N_9134);
xor U10884 (N_10884,N_9033,N_9276);
xnor U10885 (N_10885,N_9160,N_9024);
or U10886 (N_10886,N_9705,N_9224);
or U10887 (N_10887,N_9114,N_9563);
nor U10888 (N_10888,N_9716,N_9281);
nor U10889 (N_10889,N_9775,N_9417);
and U10890 (N_10890,N_9617,N_9134);
nor U10891 (N_10891,N_9432,N_9922);
and U10892 (N_10892,N_9237,N_9988);
nand U10893 (N_10893,N_9956,N_9348);
or U10894 (N_10894,N_9897,N_9363);
or U10895 (N_10895,N_9230,N_9813);
and U10896 (N_10896,N_9210,N_9601);
and U10897 (N_10897,N_9578,N_9217);
or U10898 (N_10898,N_9291,N_9795);
nor U10899 (N_10899,N_9970,N_9337);
nor U10900 (N_10900,N_9514,N_9507);
and U10901 (N_10901,N_9425,N_9235);
nand U10902 (N_10902,N_9763,N_9029);
xor U10903 (N_10903,N_9916,N_9602);
or U10904 (N_10904,N_9650,N_9065);
nor U10905 (N_10905,N_9651,N_9160);
nor U10906 (N_10906,N_9045,N_9320);
nand U10907 (N_10907,N_9678,N_9450);
and U10908 (N_10908,N_9718,N_9379);
or U10909 (N_10909,N_9119,N_9464);
nand U10910 (N_10910,N_9416,N_9449);
and U10911 (N_10911,N_9095,N_9575);
xnor U10912 (N_10912,N_9161,N_9521);
or U10913 (N_10913,N_9055,N_9869);
nand U10914 (N_10914,N_9919,N_9263);
xnor U10915 (N_10915,N_9229,N_9481);
or U10916 (N_10916,N_9045,N_9803);
and U10917 (N_10917,N_9530,N_9167);
xor U10918 (N_10918,N_9638,N_9577);
or U10919 (N_10919,N_9530,N_9991);
xor U10920 (N_10920,N_9521,N_9434);
nand U10921 (N_10921,N_9712,N_9604);
xor U10922 (N_10922,N_9805,N_9115);
or U10923 (N_10923,N_9197,N_9881);
nor U10924 (N_10924,N_9869,N_9073);
nand U10925 (N_10925,N_9201,N_9117);
nor U10926 (N_10926,N_9521,N_9314);
or U10927 (N_10927,N_9966,N_9905);
and U10928 (N_10928,N_9158,N_9596);
xor U10929 (N_10929,N_9111,N_9703);
or U10930 (N_10930,N_9055,N_9045);
and U10931 (N_10931,N_9505,N_9342);
nor U10932 (N_10932,N_9905,N_9951);
xnor U10933 (N_10933,N_9885,N_9452);
xnor U10934 (N_10934,N_9991,N_9889);
nand U10935 (N_10935,N_9869,N_9552);
or U10936 (N_10936,N_9510,N_9173);
and U10937 (N_10937,N_9332,N_9238);
nand U10938 (N_10938,N_9168,N_9282);
nor U10939 (N_10939,N_9376,N_9531);
xnor U10940 (N_10940,N_9064,N_9507);
xor U10941 (N_10941,N_9864,N_9131);
or U10942 (N_10942,N_9804,N_9439);
and U10943 (N_10943,N_9659,N_9475);
or U10944 (N_10944,N_9908,N_9032);
xor U10945 (N_10945,N_9303,N_9594);
and U10946 (N_10946,N_9170,N_9779);
nor U10947 (N_10947,N_9581,N_9018);
xor U10948 (N_10948,N_9339,N_9653);
xnor U10949 (N_10949,N_9568,N_9401);
or U10950 (N_10950,N_9719,N_9859);
nor U10951 (N_10951,N_9834,N_9804);
or U10952 (N_10952,N_9637,N_9935);
nor U10953 (N_10953,N_9371,N_9092);
xnor U10954 (N_10954,N_9085,N_9159);
nor U10955 (N_10955,N_9331,N_9199);
nand U10956 (N_10956,N_9762,N_9757);
nand U10957 (N_10957,N_9412,N_9828);
nand U10958 (N_10958,N_9738,N_9283);
xor U10959 (N_10959,N_9423,N_9980);
xor U10960 (N_10960,N_9562,N_9403);
nand U10961 (N_10961,N_9717,N_9236);
or U10962 (N_10962,N_9937,N_9609);
or U10963 (N_10963,N_9524,N_9986);
or U10964 (N_10964,N_9180,N_9788);
nor U10965 (N_10965,N_9908,N_9652);
or U10966 (N_10966,N_9455,N_9628);
and U10967 (N_10967,N_9601,N_9503);
or U10968 (N_10968,N_9706,N_9952);
or U10969 (N_10969,N_9474,N_9083);
and U10970 (N_10970,N_9917,N_9721);
and U10971 (N_10971,N_9387,N_9220);
nand U10972 (N_10972,N_9889,N_9791);
or U10973 (N_10973,N_9420,N_9568);
or U10974 (N_10974,N_9901,N_9951);
and U10975 (N_10975,N_9554,N_9016);
nand U10976 (N_10976,N_9888,N_9077);
and U10977 (N_10977,N_9489,N_9717);
and U10978 (N_10978,N_9019,N_9461);
or U10979 (N_10979,N_9154,N_9365);
nor U10980 (N_10980,N_9097,N_9637);
xor U10981 (N_10981,N_9339,N_9281);
nor U10982 (N_10982,N_9963,N_9578);
nand U10983 (N_10983,N_9726,N_9773);
nor U10984 (N_10984,N_9625,N_9271);
nor U10985 (N_10985,N_9397,N_9869);
xnor U10986 (N_10986,N_9586,N_9334);
or U10987 (N_10987,N_9584,N_9047);
xor U10988 (N_10988,N_9705,N_9995);
or U10989 (N_10989,N_9430,N_9562);
nand U10990 (N_10990,N_9154,N_9878);
nor U10991 (N_10991,N_9905,N_9994);
nand U10992 (N_10992,N_9773,N_9528);
or U10993 (N_10993,N_9050,N_9356);
nor U10994 (N_10994,N_9742,N_9913);
xnor U10995 (N_10995,N_9584,N_9284);
xor U10996 (N_10996,N_9014,N_9152);
and U10997 (N_10997,N_9221,N_9080);
and U10998 (N_10998,N_9431,N_9866);
nand U10999 (N_10999,N_9761,N_9110);
nand U11000 (N_11000,N_10544,N_10454);
xor U11001 (N_11001,N_10655,N_10829);
and U11002 (N_11002,N_10137,N_10850);
nand U11003 (N_11003,N_10141,N_10372);
nand U11004 (N_11004,N_10112,N_10576);
nand U11005 (N_11005,N_10092,N_10469);
and U11006 (N_11006,N_10941,N_10170);
xnor U11007 (N_11007,N_10106,N_10684);
and U11008 (N_11008,N_10316,N_10640);
nor U11009 (N_11009,N_10858,N_10784);
nor U11010 (N_11010,N_10256,N_10658);
xor U11011 (N_11011,N_10215,N_10455);
xnor U11012 (N_11012,N_10002,N_10633);
nand U11013 (N_11013,N_10262,N_10935);
nand U11014 (N_11014,N_10641,N_10887);
or U11015 (N_11015,N_10798,N_10390);
nand U11016 (N_11016,N_10615,N_10078);
nand U11017 (N_11017,N_10878,N_10360);
xnor U11018 (N_11018,N_10160,N_10443);
or U11019 (N_11019,N_10029,N_10644);
and U11020 (N_11020,N_10118,N_10163);
nor U11021 (N_11021,N_10569,N_10770);
or U11022 (N_11022,N_10343,N_10621);
nand U11023 (N_11023,N_10032,N_10169);
nand U11024 (N_11024,N_10760,N_10425);
nand U11025 (N_11025,N_10147,N_10749);
nand U11026 (N_11026,N_10442,N_10797);
xor U11027 (N_11027,N_10845,N_10364);
nand U11028 (N_11028,N_10752,N_10435);
nand U11029 (N_11029,N_10335,N_10586);
nor U11030 (N_11030,N_10448,N_10235);
and U11031 (N_11031,N_10445,N_10605);
nor U11032 (N_11032,N_10253,N_10421);
xor U11033 (N_11033,N_10715,N_10489);
nand U11034 (N_11034,N_10942,N_10254);
or U11035 (N_11035,N_10243,N_10102);
nand U11036 (N_11036,N_10242,N_10209);
or U11037 (N_11037,N_10963,N_10165);
xnor U11038 (N_11038,N_10894,N_10440);
nor U11039 (N_11039,N_10525,N_10076);
nand U11040 (N_11040,N_10562,N_10266);
and U11041 (N_11041,N_10532,N_10350);
nand U11042 (N_11042,N_10050,N_10116);
nor U11043 (N_11043,N_10258,N_10999);
nand U11044 (N_11044,N_10089,N_10152);
or U11045 (N_11045,N_10195,N_10593);
nand U11046 (N_11046,N_10328,N_10914);
xor U11047 (N_11047,N_10302,N_10902);
or U11048 (N_11048,N_10986,N_10074);
and U11049 (N_11049,N_10475,N_10545);
and U11050 (N_11050,N_10984,N_10844);
nor U11051 (N_11051,N_10547,N_10300);
or U11052 (N_11052,N_10663,N_10675);
nor U11053 (N_11053,N_10368,N_10166);
nor U11054 (N_11054,N_10721,N_10402);
or U11055 (N_11055,N_10765,N_10769);
or U11056 (N_11056,N_10654,N_10090);
xnor U11057 (N_11057,N_10107,N_10714);
nand U11058 (N_11058,N_10276,N_10538);
xor U11059 (N_11059,N_10839,N_10954);
xnor U11060 (N_11060,N_10724,N_10874);
nand U11061 (N_11061,N_10702,N_10818);
xnor U11062 (N_11062,N_10397,N_10950);
xnor U11063 (N_11063,N_10557,N_10125);
nor U11064 (N_11064,N_10059,N_10778);
or U11065 (N_11065,N_10503,N_10225);
nor U11066 (N_11066,N_10711,N_10167);
nand U11067 (N_11067,N_10139,N_10071);
or U11068 (N_11068,N_10953,N_10685);
and U11069 (N_11069,N_10244,N_10960);
nand U11070 (N_11070,N_10229,N_10404);
and U11071 (N_11071,N_10301,N_10245);
nand U11072 (N_11072,N_10776,N_10862);
and U11073 (N_11073,N_10136,N_10661);
nand U11074 (N_11074,N_10896,N_10533);
nand U11075 (N_11075,N_10738,N_10851);
or U11076 (N_11076,N_10321,N_10819);
or U11077 (N_11077,N_10487,N_10021);
nor U11078 (N_11078,N_10358,N_10337);
and U11079 (N_11079,N_10155,N_10647);
and U11080 (N_11080,N_10635,N_10808);
nand U11081 (N_11081,N_10252,N_10510);
nand U11082 (N_11082,N_10117,N_10591);
or U11083 (N_11083,N_10413,N_10634);
and U11084 (N_11084,N_10520,N_10824);
nand U11085 (N_11085,N_10671,N_10476);
or U11086 (N_11086,N_10471,N_10860);
or U11087 (N_11087,N_10188,N_10474);
or U11088 (N_11088,N_10062,N_10294);
nand U11089 (N_11089,N_10524,N_10535);
nand U11090 (N_11090,N_10648,N_10053);
xor U11091 (N_11091,N_10465,N_10676);
or U11092 (N_11092,N_10590,N_10747);
nor U11093 (N_11093,N_10745,N_10701);
nor U11094 (N_11094,N_10279,N_10666);
xnor U11095 (N_11095,N_10436,N_10405);
nand U11096 (N_11096,N_10363,N_10961);
nand U11097 (N_11097,N_10791,N_10908);
nor U11098 (N_11098,N_10728,N_10036);
or U11099 (N_11099,N_10846,N_10101);
and U11100 (N_11100,N_10563,N_10929);
or U11101 (N_11101,N_10656,N_10354);
nor U11102 (N_11102,N_10437,N_10610);
xnor U11103 (N_11103,N_10452,N_10055);
nand U11104 (N_11104,N_10431,N_10997);
and U11105 (N_11105,N_10611,N_10542);
nor U11106 (N_11106,N_10028,N_10864);
and U11107 (N_11107,N_10859,N_10956);
xnor U11108 (N_11108,N_10239,N_10907);
nand U11109 (N_11109,N_10973,N_10286);
or U11110 (N_11110,N_10378,N_10073);
nor U11111 (N_11111,N_10131,N_10067);
or U11112 (N_11112,N_10297,N_10216);
and U11113 (N_11113,N_10324,N_10810);
nor U11114 (N_11114,N_10081,N_10504);
xnor U11115 (N_11115,N_10758,N_10947);
xnor U11116 (N_11116,N_10650,N_10678);
nor U11117 (N_11117,N_10462,N_10522);
nor U11118 (N_11118,N_10628,N_10889);
and U11119 (N_11119,N_10150,N_10599);
xor U11120 (N_11120,N_10096,N_10821);
nor U11121 (N_11121,N_10505,N_10339);
xnor U11122 (N_11122,N_10237,N_10497);
nand U11123 (N_11123,N_10660,N_10260);
and U11124 (N_11124,N_10008,N_10744);
xnor U11125 (N_11125,N_10553,N_10554);
and U11126 (N_11126,N_10441,N_10406);
nand U11127 (N_11127,N_10417,N_10004);
xor U11128 (N_11128,N_10317,N_10273);
and U11129 (N_11129,N_10700,N_10298);
or U11130 (N_11130,N_10494,N_10045);
nor U11131 (N_11131,N_10897,N_10222);
xnor U11132 (N_11132,N_10458,N_10380);
nor U11133 (N_11133,N_10828,N_10456);
xnor U11134 (N_11134,N_10699,N_10022);
or U11135 (N_11135,N_10149,N_10221);
and U11136 (N_11136,N_10540,N_10341);
and U11137 (N_11137,N_10578,N_10756);
or U11138 (N_11138,N_10636,N_10624);
nor U11139 (N_11139,N_10501,N_10584);
xor U11140 (N_11140,N_10781,N_10970);
nand U11141 (N_11141,N_10867,N_10126);
xnor U11142 (N_11142,N_10793,N_10541);
xor U11143 (N_11143,N_10282,N_10065);
xnor U11144 (N_11144,N_10697,N_10401);
nor U11145 (N_11145,N_10592,N_10679);
xor U11146 (N_11146,N_10991,N_10607);
nor U11147 (N_11147,N_10575,N_10792);
or U11148 (N_11148,N_10861,N_10043);
nor U11149 (N_11149,N_10733,N_10771);
nor U11150 (N_11150,N_10519,N_10052);
nor U11151 (N_11151,N_10355,N_10919);
and U11152 (N_11152,N_10395,N_10882);
or U11153 (N_11153,N_10945,N_10038);
or U11154 (N_11154,N_10827,N_10723);
or U11155 (N_11155,N_10737,N_10367);
xor U11156 (N_11156,N_10375,N_10098);
xnor U11157 (N_11157,N_10289,N_10162);
nor U11158 (N_11158,N_10938,N_10691);
or U11159 (N_11159,N_10911,N_10472);
or U11160 (N_11160,N_10681,N_10764);
and U11161 (N_11161,N_10531,N_10854);
nor U11162 (N_11162,N_10171,N_10534);
nand U11163 (N_11163,N_10842,N_10080);
or U11164 (N_11164,N_10075,N_10825);
nand U11165 (N_11165,N_10849,N_10414);
nor U11166 (N_11166,N_10602,N_10114);
nor U11167 (N_11167,N_10247,N_10426);
nand U11168 (N_11168,N_10461,N_10852);
xnor U11169 (N_11169,N_10399,N_10928);
nor U11170 (N_11170,N_10492,N_10670);
and U11171 (N_11171,N_10937,N_10526);
nor U11172 (N_11172,N_10976,N_10969);
xor U11173 (N_11173,N_10523,N_10453);
xor U11174 (N_11174,N_10909,N_10037);
nor U11175 (N_11175,N_10359,N_10352);
nor U11176 (N_11176,N_10483,N_10416);
nand U11177 (N_11177,N_10275,N_10201);
or U11178 (N_11178,N_10285,N_10659);
xor U11179 (N_11179,N_10690,N_10233);
and U11180 (N_11180,N_10370,N_10313);
nand U11181 (N_11181,N_10795,N_10948);
or U11182 (N_11182,N_10608,N_10891);
xor U11183 (N_11183,N_10391,N_10934);
nor U11184 (N_11184,N_10609,N_10966);
nor U11185 (N_11185,N_10603,N_10299);
nand U11186 (N_11186,N_10159,N_10259);
xnor U11187 (N_11187,N_10091,N_10044);
nand U11188 (N_11188,N_10134,N_10692);
or U11189 (N_11189,N_10151,N_10987);
xor U11190 (N_11190,N_10645,N_10383);
or U11191 (N_11191,N_10552,N_10047);
xor U11192 (N_11192,N_10652,N_10020);
xnor U11193 (N_11193,N_10268,N_10411);
nand U11194 (N_11194,N_10172,N_10119);
or U11195 (N_11195,N_10823,N_10992);
or U11196 (N_11196,N_10001,N_10853);
nand U11197 (N_11197,N_10287,N_10408);
or U11198 (N_11198,N_10351,N_10122);
and U11199 (N_11199,N_10600,N_10802);
nor U11200 (N_11200,N_10093,N_10910);
xnor U11201 (N_11201,N_10365,N_10288);
nand U11202 (N_11202,N_10312,N_10251);
nand U11203 (N_11203,N_10333,N_10572);
xor U11204 (N_11204,N_10872,N_10639);
xor U11205 (N_11205,N_10972,N_10479);
and U11206 (N_11206,N_10869,N_10855);
or U11207 (N_11207,N_10186,N_10110);
and U11208 (N_11208,N_10493,N_10508);
and U11209 (N_11209,N_10975,N_10280);
xor U11210 (N_11210,N_10498,N_10241);
and U11211 (N_11211,N_10174,N_10310);
xor U11212 (N_11212,N_10318,N_10530);
or U11213 (N_11213,N_10587,N_10816);
xor U11214 (N_11214,N_10528,N_10631);
or U11215 (N_11215,N_10228,N_10274);
nor U11216 (N_11216,N_10079,N_10786);
and U11217 (N_11217,N_10627,N_10782);
nor U11218 (N_11218,N_10742,N_10396);
or U11219 (N_11219,N_10295,N_10665);
nand U11220 (N_11220,N_10511,N_10129);
nor U11221 (N_11221,N_10521,N_10703);
nand U11222 (N_11222,N_10732,N_10250);
nor U11223 (N_11223,N_10293,N_10133);
xor U11224 (N_11224,N_10653,N_10207);
xnor U11225 (N_11225,N_10181,N_10261);
and U11226 (N_11226,N_10084,N_10218);
and U11227 (N_11227,N_10704,N_10277);
nand U11228 (N_11228,N_10672,N_10673);
nor U11229 (N_11229,N_10594,N_10955);
or U11230 (N_11230,N_10546,N_10807);
or U11231 (N_11231,N_10019,N_10979);
nor U11232 (N_11232,N_10817,N_10693);
or U11233 (N_11233,N_10922,N_10667);
and U11234 (N_11234,N_10625,N_10898);
or U11235 (N_11235,N_10481,N_10024);
nand U11236 (N_11236,N_10198,N_10227);
nand U11237 (N_11237,N_10757,N_10529);
and U11238 (N_11238,N_10264,N_10006);
nor U11239 (N_11239,N_10993,N_10649);
or U11240 (N_11240,N_10464,N_10143);
nor U11241 (N_11241,N_10236,N_10622);
xor U11242 (N_11242,N_10377,N_10951);
and U11243 (N_11243,N_10637,N_10041);
xor U11244 (N_11244,N_10034,N_10495);
or U11245 (N_11245,N_10613,N_10446);
nor U11246 (N_11246,N_10774,N_10589);
or U11247 (N_11247,N_10000,N_10196);
and U11248 (N_11248,N_10304,N_10559);
and U11249 (N_11249,N_10780,N_10226);
xnor U11250 (N_11250,N_10866,N_10932);
xnor U11251 (N_11251,N_10574,N_10877);
or U11252 (N_11252,N_10556,N_10187);
or U11253 (N_11253,N_10459,N_10601);
or U11254 (N_11254,N_10176,N_10499);
nand U11255 (N_11255,N_10183,N_10596);
nand U11256 (N_11256,N_10430,N_10104);
xnor U11257 (N_11257,N_10729,N_10582);
nor U11258 (N_11258,N_10224,N_10381);
nor U11259 (N_11259,N_10686,N_10392);
nor U11260 (N_11260,N_10863,N_10959);
xnor U11261 (N_11261,N_10912,N_10856);
nand U11262 (N_11262,N_10980,N_10799);
or U11263 (N_11263,N_10148,N_10031);
or U11264 (N_11264,N_10389,N_10952);
xor U11265 (N_11265,N_10219,N_10070);
xor U11266 (N_11266,N_10832,N_10964);
and U11267 (N_11267,N_10130,N_10192);
nand U11268 (N_11268,N_10933,N_10892);
xor U11269 (N_11269,N_10315,N_10361);
xor U11270 (N_11270,N_10467,N_10876);
xnor U11271 (N_11271,N_10265,N_10347);
and U11272 (N_11272,N_10680,N_10357);
xor U11273 (N_11273,N_10323,N_10706);
xnor U11274 (N_11274,N_10039,N_10595);
xnor U11275 (N_11275,N_10881,N_10451);
nand U11276 (N_11276,N_10974,N_10349);
xnor U11277 (N_11277,N_10127,N_10717);
nand U11278 (N_11278,N_10433,N_10329);
nand U11279 (N_11279,N_10549,N_10583);
xor U11280 (N_11280,N_10895,N_10138);
and U11281 (N_11281,N_10722,N_10868);
nand U11282 (N_11282,N_10924,N_10826);
and U11283 (N_11283,N_10906,N_10146);
or U11284 (N_11284,N_10135,N_10629);
nand U11285 (N_11285,N_10257,N_10580);
xnor U11286 (N_11286,N_10886,N_10468);
xor U11287 (N_11287,N_10620,N_10082);
nor U11288 (N_11288,N_10536,N_10168);
or U11289 (N_11289,N_10812,N_10835);
nor U11290 (N_11290,N_10353,N_10449);
xnor U11291 (N_11291,N_10834,N_10838);
nor U11292 (N_11292,N_10916,N_10736);
xnor U11293 (N_11293,N_10657,N_10386);
nand U11294 (N_11294,N_10178,N_10988);
and U11295 (N_11295,N_10409,N_10766);
or U11296 (N_11296,N_10971,N_10438);
nand U11297 (N_11297,N_10925,N_10154);
xnor U11298 (N_11298,N_10346,N_10398);
xnor U11299 (N_11299,N_10290,N_10427);
or U11300 (N_11300,N_10128,N_10439);
and U11301 (N_11301,N_10083,N_10164);
or U11302 (N_11302,N_10687,N_10783);
xor U11303 (N_11303,N_10840,N_10263);
xor U11304 (N_11304,N_10689,N_10651);
nor U11305 (N_11305,N_10026,N_10412);
xor U11306 (N_11306,N_10103,N_10695);
and U11307 (N_11307,N_10210,N_10767);
xor U11308 (N_11308,N_10674,N_10040);
nand U11309 (N_11309,N_10132,N_10308);
or U11310 (N_11310,N_10843,N_10801);
and U11311 (N_11311,N_10551,N_10223);
xnor U11312 (N_11312,N_10967,N_10848);
nor U11313 (N_11313,N_10617,N_10108);
and U11314 (N_11314,N_10056,N_10057);
nor U11315 (N_11315,N_10027,N_10836);
nand U11316 (N_11316,N_10214,N_10113);
xnor U11317 (N_11317,N_10063,N_10800);
xnor U11318 (N_11318,N_10213,N_10725);
or U11319 (N_11319,N_10669,N_10326);
or U11320 (N_11320,N_10158,N_10199);
nor U11321 (N_11321,N_10124,N_10913);
nand U11322 (N_11322,N_10485,N_10957);
nor U11323 (N_11323,N_10457,N_10698);
nand U11324 (N_11324,N_10720,N_10012);
xnor U11325 (N_11325,N_10502,N_10005);
or U11326 (N_11326,N_10741,N_10332);
nor U11327 (N_11327,N_10014,N_10272);
xnor U11328 (N_11328,N_10708,N_10173);
xor U11329 (N_11329,N_10470,N_10958);
or U11330 (N_11330,N_10623,N_10517);
or U11331 (N_11331,N_10156,N_10918);
and U11332 (N_11332,N_10643,N_10018);
or U11333 (N_11333,N_10734,N_10208);
or U11334 (N_11334,N_10748,N_10344);
xor U11335 (N_11335,N_10565,N_10115);
nor U11336 (N_11336,N_10182,N_10820);
or U11337 (N_11337,N_10120,N_10204);
and U11338 (N_11338,N_10618,N_10884);
nand U11339 (N_11339,N_10804,N_10585);
or U11340 (N_11340,N_10785,N_10726);
or U11341 (N_11341,N_10775,N_10255);
xor U11342 (N_11342,N_10930,N_10978);
nand U11343 (N_11343,N_10473,N_10345);
nand U11344 (N_11344,N_10616,N_10746);
and U11345 (N_11345,N_10177,N_10400);
nand U11346 (N_11346,N_10190,N_10619);
nand U11347 (N_11347,N_10140,N_10509);
xor U11348 (N_11348,N_10477,N_10191);
or U11349 (N_11349,N_10570,N_10809);
xor U11350 (N_11350,N_10870,N_10314);
xnor U11351 (N_11351,N_10338,N_10931);
or U11352 (N_11352,N_10292,N_10915);
nand U11353 (N_11353,N_10217,N_10566);
nor U11354 (N_11354,N_10482,N_10995);
and U11355 (N_11355,N_10768,N_10269);
or U11356 (N_11356,N_10831,N_10777);
nor U11357 (N_11357,N_10990,N_10923);
nor U11358 (N_11358,N_10200,N_10612);
and U11359 (N_11359,N_10754,N_10322);
or U11360 (N_11360,N_10206,N_10598);
nand U11361 (N_11361,N_10144,N_10841);
nand U11362 (N_11362,N_10944,N_10054);
xor U11363 (N_11363,N_10926,N_10284);
and U11364 (N_11364,N_10983,N_10588);
and U11365 (N_11365,N_10805,N_10900);
nor U11366 (N_11366,N_10813,N_10384);
or U11367 (N_11367,N_10905,N_10240);
or U11368 (N_11368,N_10560,N_10705);
nor U11369 (N_11369,N_10539,N_10016);
xor U11370 (N_11370,N_10638,N_10248);
and U11371 (N_11371,N_10989,N_10373);
or U11372 (N_11372,N_10371,N_10205);
nor U11373 (N_11373,N_10042,N_10283);
and U11374 (N_11374,N_10901,N_10920);
nand U11375 (N_11375,N_10366,N_10007);
nor U11376 (N_11376,N_10822,N_10307);
and U11377 (N_11377,N_10561,N_10048);
nand U11378 (N_11378,N_10606,N_10415);
xnor U11379 (N_11379,N_10010,N_10403);
nand U11380 (N_11380,N_10664,N_10085);
xnor U11381 (N_11381,N_10419,N_10490);
or U11382 (N_11382,N_10463,N_10046);
nor U11383 (N_11383,N_10753,N_10334);
or U11384 (N_11384,N_10998,N_10727);
and U11385 (N_11385,N_10815,N_10374);
or U11386 (N_11386,N_10121,N_10880);
or U11387 (N_11387,N_10903,N_10712);
or U11388 (N_11388,N_10197,N_10420);
and U11389 (N_11389,N_10193,N_10696);
nand U11390 (N_11390,N_10740,N_10837);
nand U11391 (N_11391,N_10994,N_10030);
nor U11392 (N_11392,N_10220,N_10231);
nor U11393 (N_11393,N_10939,N_10743);
nand U11394 (N_11394,N_10362,N_10632);
nor U11395 (N_11395,N_10682,N_10794);
and U11396 (N_11396,N_10890,N_10100);
nand U11397 (N_11397,N_10230,N_10506);
nand U11398 (N_11398,N_10460,N_10105);
nor U11399 (N_11399,N_10211,N_10094);
nand U11400 (N_11400,N_10677,N_10086);
nor U11401 (N_11401,N_10614,N_10604);
nor U11402 (N_11402,N_10888,N_10893);
nand U11403 (N_11403,N_10796,N_10803);
xnor U11404 (N_11404,N_10066,N_10394);
xnor U11405 (N_11405,N_10646,N_10996);
and U11406 (N_11406,N_10331,N_10773);
xor U11407 (N_11407,N_10875,N_10418);
or U11408 (N_11408,N_10157,N_10883);
xor U11409 (N_11409,N_10202,N_10683);
or U11410 (N_11410,N_10145,N_10719);
nor U11411 (N_11411,N_10049,N_10977);
nand U11412 (N_11412,N_10713,N_10123);
or U11413 (N_11413,N_10833,N_10422);
nand U11414 (N_11414,N_10514,N_10051);
or U11415 (N_11415,N_10885,N_10234);
xor U11416 (N_11416,N_10630,N_10095);
xnor U11417 (N_11417,N_10484,N_10194);
nor U11418 (N_11418,N_10111,N_10087);
and U11419 (N_11419,N_10303,N_10466);
xor U11420 (N_11420,N_10291,N_10904);
nor U11421 (N_11421,N_10577,N_10642);
nand U11422 (N_11422,N_10755,N_10385);
nand U11423 (N_11423,N_10873,N_10434);
nand U11424 (N_11424,N_10278,N_10790);
nor U11425 (N_11425,N_10662,N_10548);
or U11426 (N_11426,N_10025,N_10537);
nand U11427 (N_11427,N_10342,N_10330);
and U11428 (N_11428,N_10035,N_10189);
and U11429 (N_11429,N_10626,N_10946);
and U11430 (N_11430,N_10212,N_10480);
nor U11431 (N_11431,N_10962,N_10949);
nand U11432 (N_11432,N_10555,N_10788);
nand U11433 (N_11433,N_10573,N_10762);
nor U11434 (N_11434,N_10142,N_10444);
nand U11435 (N_11435,N_10428,N_10936);
and U11436 (N_11436,N_10017,N_10387);
and U11437 (N_11437,N_10527,N_10011);
or U11438 (N_11438,N_10061,N_10311);
nand U11439 (N_11439,N_10735,N_10789);
and U11440 (N_11440,N_10718,N_10968);
or U11441 (N_11441,N_10232,N_10376);
and U11442 (N_11442,N_10806,N_10985);
or U11443 (N_11443,N_10750,N_10981);
nor U11444 (N_11444,N_10558,N_10568);
or U11445 (N_11445,N_10423,N_10410);
nand U11446 (N_11446,N_10319,N_10306);
and U11447 (N_11447,N_10109,N_10579);
nand U11448 (N_11448,N_10927,N_10309);
xnor U11449 (N_11449,N_10759,N_10153);
and U11450 (N_11450,N_10486,N_10271);
nand U11451 (N_11451,N_10488,N_10382);
nand U11452 (N_11452,N_10921,N_10899);
or U11453 (N_11453,N_10814,N_10175);
xnor U11454 (N_11454,N_10099,N_10281);
nand U11455 (N_11455,N_10917,N_10238);
nand U11456 (N_11456,N_10710,N_10068);
nor U11457 (N_11457,N_10507,N_10320);
nor U11458 (N_11458,N_10491,N_10772);
nand U11459 (N_11459,N_10943,N_10336);
or U11460 (N_11460,N_10379,N_10077);
nand U11461 (N_11461,N_10327,N_10388);
nor U11462 (N_11462,N_10550,N_10180);
nand U11463 (N_11463,N_10246,N_10581);
nor U11464 (N_11464,N_10830,N_10203);
and U11465 (N_11465,N_10249,N_10694);
xor U11466 (N_11466,N_10688,N_10088);
or U11467 (N_11467,N_10450,N_10348);
and U11468 (N_11468,N_10567,N_10072);
or U11469 (N_11469,N_10707,N_10407);
nand U11470 (N_11470,N_10060,N_10023);
and U11471 (N_11471,N_10296,N_10013);
or U11472 (N_11472,N_10811,N_10564);
nor U11473 (N_11473,N_10015,N_10518);
xor U11474 (N_11474,N_10515,N_10879);
or U11475 (N_11475,N_10730,N_10393);
nor U11476 (N_11476,N_10871,N_10857);
or U11477 (N_11477,N_10500,N_10543);
xnor U11478 (N_11478,N_10940,N_10496);
nand U11479 (N_11479,N_10432,N_10513);
nor U11480 (N_11480,N_10270,N_10716);
nand U11481 (N_11481,N_10761,N_10429);
or U11482 (N_11482,N_10739,N_10763);
and U11483 (N_11483,N_10058,N_10069);
xor U11484 (N_11484,N_10356,N_10571);
nand U11485 (N_11485,N_10179,N_10516);
nor U11486 (N_11486,N_10424,N_10447);
nor U11487 (N_11487,N_10668,N_10340);
nand U11488 (N_11488,N_10305,N_10325);
xor U11489 (N_11489,N_10865,N_10478);
xor U11490 (N_11490,N_10512,N_10731);
or U11491 (N_11491,N_10161,N_10597);
xnor U11492 (N_11492,N_10982,N_10267);
or U11493 (N_11493,N_10185,N_10097);
and U11494 (N_11494,N_10787,N_10064);
nor U11495 (N_11495,N_10709,N_10184);
and U11496 (N_11496,N_10847,N_10369);
or U11497 (N_11497,N_10779,N_10751);
nor U11498 (N_11498,N_10009,N_10033);
or U11499 (N_11499,N_10003,N_10965);
or U11500 (N_11500,N_10013,N_10433);
nand U11501 (N_11501,N_10831,N_10933);
xor U11502 (N_11502,N_10542,N_10815);
nor U11503 (N_11503,N_10909,N_10956);
nor U11504 (N_11504,N_10077,N_10816);
nand U11505 (N_11505,N_10503,N_10571);
xnor U11506 (N_11506,N_10316,N_10018);
nand U11507 (N_11507,N_10891,N_10988);
and U11508 (N_11508,N_10318,N_10029);
xor U11509 (N_11509,N_10416,N_10562);
and U11510 (N_11510,N_10049,N_10721);
or U11511 (N_11511,N_10844,N_10905);
xor U11512 (N_11512,N_10474,N_10149);
nor U11513 (N_11513,N_10526,N_10508);
and U11514 (N_11514,N_10130,N_10607);
nand U11515 (N_11515,N_10083,N_10032);
nand U11516 (N_11516,N_10895,N_10064);
nor U11517 (N_11517,N_10427,N_10041);
nor U11518 (N_11518,N_10264,N_10765);
or U11519 (N_11519,N_10826,N_10890);
nand U11520 (N_11520,N_10553,N_10833);
nor U11521 (N_11521,N_10228,N_10837);
or U11522 (N_11522,N_10488,N_10621);
nand U11523 (N_11523,N_10686,N_10585);
xnor U11524 (N_11524,N_10297,N_10496);
nor U11525 (N_11525,N_10531,N_10627);
xor U11526 (N_11526,N_10487,N_10366);
nor U11527 (N_11527,N_10000,N_10325);
and U11528 (N_11528,N_10250,N_10036);
and U11529 (N_11529,N_10901,N_10597);
or U11530 (N_11530,N_10637,N_10877);
nor U11531 (N_11531,N_10627,N_10217);
nand U11532 (N_11532,N_10784,N_10886);
or U11533 (N_11533,N_10856,N_10783);
nor U11534 (N_11534,N_10662,N_10260);
nand U11535 (N_11535,N_10701,N_10030);
nand U11536 (N_11536,N_10417,N_10846);
and U11537 (N_11537,N_10545,N_10331);
nand U11538 (N_11538,N_10981,N_10143);
or U11539 (N_11539,N_10339,N_10220);
nand U11540 (N_11540,N_10807,N_10216);
nand U11541 (N_11541,N_10707,N_10253);
or U11542 (N_11542,N_10585,N_10773);
xor U11543 (N_11543,N_10969,N_10766);
nor U11544 (N_11544,N_10928,N_10841);
nand U11545 (N_11545,N_10466,N_10243);
nor U11546 (N_11546,N_10636,N_10615);
or U11547 (N_11547,N_10268,N_10970);
or U11548 (N_11548,N_10215,N_10722);
and U11549 (N_11549,N_10013,N_10805);
nand U11550 (N_11550,N_10495,N_10491);
nand U11551 (N_11551,N_10113,N_10883);
xnor U11552 (N_11552,N_10792,N_10839);
or U11553 (N_11553,N_10681,N_10588);
nand U11554 (N_11554,N_10660,N_10719);
or U11555 (N_11555,N_10571,N_10318);
nor U11556 (N_11556,N_10636,N_10988);
xnor U11557 (N_11557,N_10748,N_10696);
nor U11558 (N_11558,N_10418,N_10541);
xnor U11559 (N_11559,N_10151,N_10109);
or U11560 (N_11560,N_10003,N_10112);
nand U11561 (N_11561,N_10717,N_10909);
xnor U11562 (N_11562,N_10687,N_10023);
nor U11563 (N_11563,N_10156,N_10247);
xnor U11564 (N_11564,N_10490,N_10516);
xnor U11565 (N_11565,N_10004,N_10577);
nand U11566 (N_11566,N_10072,N_10071);
xnor U11567 (N_11567,N_10583,N_10164);
nor U11568 (N_11568,N_10913,N_10297);
and U11569 (N_11569,N_10457,N_10745);
xnor U11570 (N_11570,N_10435,N_10047);
nand U11571 (N_11571,N_10569,N_10256);
and U11572 (N_11572,N_10300,N_10279);
or U11573 (N_11573,N_10556,N_10129);
nand U11574 (N_11574,N_10642,N_10491);
and U11575 (N_11575,N_10736,N_10552);
and U11576 (N_11576,N_10576,N_10325);
nand U11577 (N_11577,N_10886,N_10423);
nor U11578 (N_11578,N_10770,N_10255);
xor U11579 (N_11579,N_10082,N_10086);
nand U11580 (N_11580,N_10040,N_10845);
xor U11581 (N_11581,N_10961,N_10793);
xnor U11582 (N_11582,N_10894,N_10908);
nor U11583 (N_11583,N_10869,N_10722);
nand U11584 (N_11584,N_10840,N_10907);
nor U11585 (N_11585,N_10607,N_10878);
xor U11586 (N_11586,N_10744,N_10404);
nor U11587 (N_11587,N_10034,N_10991);
nor U11588 (N_11588,N_10245,N_10264);
or U11589 (N_11589,N_10343,N_10354);
xor U11590 (N_11590,N_10805,N_10971);
nor U11591 (N_11591,N_10582,N_10678);
and U11592 (N_11592,N_10221,N_10165);
xor U11593 (N_11593,N_10905,N_10890);
or U11594 (N_11594,N_10886,N_10679);
or U11595 (N_11595,N_10910,N_10568);
or U11596 (N_11596,N_10782,N_10346);
xor U11597 (N_11597,N_10352,N_10526);
xnor U11598 (N_11598,N_10866,N_10144);
and U11599 (N_11599,N_10174,N_10147);
nor U11600 (N_11600,N_10494,N_10570);
nand U11601 (N_11601,N_10340,N_10102);
xor U11602 (N_11602,N_10906,N_10426);
or U11603 (N_11603,N_10771,N_10498);
or U11604 (N_11604,N_10992,N_10998);
nand U11605 (N_11605,N_10862,N_10253);
or U11606 (N_11606,N_10309,N_10166);
nor U11607 (N_11607,N_10226,N_10938);
and U11608 (N_11608,N_10096,N_10483);
or U11609 (N_11609,N_10697,N_10002);
nor U11610 (N_11610,N_10711,N_10501);
nor U11611 (N_11611,N_10116,N_10157);
nor U11612 (N_11612,N_10413,N_10442);
or U11613 (N_11613,N_10616,N_10909);
or U11614 (N_11614,N_10810,N_10247);
nor U11615 (N_11615,N_10368,N_10209);
or U11616 (N_11616,N_10612,N_10998);
xnor U11617 (N_11617,N_10553,N_10633);
nor U11618 (N_11618,N_10759,N_10687);
xor U11619 (N_11619,N_10647,N_10852);
xor U11620 (N_11620,N_10593,N_10305);
and U11621 (N_11621,N_10845,N_10381);
xnor U11622 (N_11622,N_10765,N_10587);
and U11623 (N_11623,N_10462,N_10586);
nor U11624 (N_11624,N_10756,N_10728);
or U11625 (N_11625,N_10860,N_10208);
nand U11626 (N_11626,N_10722,N_10083);
or U11627 (N_11627,N_10554,N_10760);
xnor U11628 (N_11628,N_10205,N_10604);
nor U11629 (N_11629,N_10977,N_10363);
nand U11630 (N_11630,N_10853,N_10481);
or U11631 (N_11631,N_10021,N_10519);
and U11632 (N_11632,N_10932,N_10908);
nor U11633 (N_11633,N_10947,N_10902);
nand U11634 (N_11634,N_10566,N_10451);
xnor U11635 (N_11635,N_10087,N_10544);
xor U11636 (N_11636,N_10533,N_10589);
xnor U11637 (N_11637,N_10218,N_10200);
nor U11638 (N_11638,N_10241,N_10249);
or U11639 (N_11639,N_10022,N_10662);
xor U11640 (N_11640,N_10869,N_10427);
nand U11641 (N_11641,N_10980,N_10374);
xnor U11642 (N_11642,N_10419,N_10717);
or U11643 (N_11643,N_10711,N_10461);
or U11644 (N_11644,N_10681,N_10034);
nand U11645 (N_11645,N_10563,N_10399);
nor U11646 (N_11646,N_10752,N_10604);
nor U11647 (N_11647,N_10800,N_10964);
and U11648 (N_11648,N_10930,N_10392);
and U11649 (N_11649,N_10802,N_10726);
nand U11650 (N_11650,N_10882,N_10087);
xnor U11651 (N_11651,N_10687,N_10952);
nand U11652 (N_11652,N_10252,N_10468);
xnor U11653 (N_11653,N_10968,N_10134);
or U11654 (N_11654,N_10459,N_10850);
nand U11655 (N_11655,N_10905,N_10271);
nand U11656 (N_11656,N_10225,N_10591);
nand U11657 (N_11657,N_10992,N_10516);
or U11658 (N_11658,N_10965,N_10604);
or U11659 (N_11659,N_10327,N_10037);
and U11660 (N_11660,N_10269,N_10195);
or U11661 (N_11661,N_10937,N_10501);
or U11662 (N_11662,N_10284,N_10303);
and U11663 (N_11663,N_10212,N_10052);
nand U11664 (N_11664,N_10548,N_10430);
xnor U11665 (N_11665,N_10139,N_10803);
nand U11666 (N_11666,N_10092,N_10384);
xor U11667 (N_11667,N_10102,N_10899);
or U11668 (N_11668,N_10559,N_10566);
or U11669 (N_11669,N_10358,N_10354);
or U11670 (N_11670,N_10491,N_10221);
or U11671 (N_11671,N_10463,N_10762);
xnor U11672 (N_11672,N_10282,N_10043);
or U11673 (N_11673,N_10168,N_10006);
nand U11674 (N_11674,N_10214,N_10325);
and U11675 (N_11675,N_10492,N_10266);
nand U11676 (N_11676,N_10578,N_10291);
xnor U11677 (N_11677,N_10634,N_10757);
or U11678 (N_11678,N_10290,N_10218);
nand U11679 (N_11679,N_10463,N_10516);
nand U11680 (N_11680,N_10868,N_10765);
nand U11681 (N_11681,N_10083,N_10541);
nand U11682 (N_11682,N_10372,N_10045);
and U11683 (N_11683,N_10681,N_10054);
nand U11684 (N_11684,N_10531,N_10155);
nand U11685 (N_11685,N_10377,N_10582);
nor U11686 (N_11686,N_10712,N_10427);
and U11687 (N_11687,N_10389,N_10614);
and U11688 (N_11688,N_10882,N_10372);
nor U11689 (N_11689,N_10348,N_10746);
or U11690 (N_11690,N_10166,N_10377);
nor U11691 (N_11691,N_10187,N_10685);
or U11692 (N_11692,N_10287,N_10231);
and U11693 (N_11693,N_10504,N_10547);
nor U11694 (N_11694,N_10724,N_10853);
xnor U11695 (N_11695,N_10845,N_10758);
nand U11696 (N_11696,N_10884,N_10452);
nand U11697 (N_11697,N_10665,N_10877);
or U11698 (N_11698,N_10904,N_10528);
nand U11699 (N_11699,N_10536,N_10952);
nand U11700 (N_11700,N_10142,N_10196);
and U11701 (N_11701,N_10253,N_10876);
and U11702 (N_11702,N_10441,N_10594);
and U11703 (N_11703,N_10061,N_10214);
and U11704 (N_11704,N_10555,N_10178);
nand U11705 (N_11705,N_10748,N_10479);
nor U11706 (N_11706,N_10086,N_10358);
nor U11707 (N_11707,N_10469,N_10218);
or U11708 (N_11708,N_10998,N_10207);
nor U11709 (N_11709,N_10337,N_10945);
nor U11710 (N_11710,N_10618,N_10412);
nor U11711 (N_11711,N_10927,N_10882);
nor U11712 (N_11712,N_10738,N_10360);
xor U11713 (N_11713,N_10887,N_10483);
and U11714 (N_11714,N_10687,N_10174);
or U11715 (N_11715,N_10513,N_10507);
nand U11716 (N_11716,N_10179,N_10470);
nor U11717 (N_11717,N_10690,N_10820);
and U11718 (N_11718,N_10044,N_10668);
nor U11719 (N_11719,N_10790,N_10872);
xor U11720 (N_11720,N_10641,N_10623);
nand U11721 (N_11721,N_10326,N_10363);
nor U11722 (N_11722,N_10156,N_10093);
nor U11723 (N_11723,N_10259,N_10282);
nor U11724 (N_11724,N_10424,N_10647);
nand U11725 (N_11725,N_10005,N_10066);
xnor U11726 (N_11726,N_10880,N_10304);
nand U11727 (N_11727,N_10290,N_10307);
and U11728 (N_11728,N_10939,N_10009);
xnor U11729 (N_11729,N_10165,N_10167);
nor U11730 (N_11730,N_10376,N_10890);
xor U11731 (N_11731,N_10654,N_10548);
nor U11732 (N_11732,N_10747,N_10937);
xor U11733 (N_11733,N_10449,N_10671);
xor U11734 (N_11734,N_10327,N_10203);
or U11735 (N_11735,N_10562,N_10274);
nor U11736 (N_11736,N_10347,N_10844);
nor U11737 (N_11737,N_10829,N_10720);
or U11738 (N_11738,N_10321,N_10244);
or U11739 (N_11739,N_10622,N_10632);
nand U11740 (N_11740,N_10523,N_10414);
nor U11741 (N_11741,N_10391,N_10040);
xnor U11742 (N_11742,N_10379,N_10715);
or U11743 (N_11743,N_10402,N_10622);
and U11744 (N_11744,N_10443,N_10977);
xor U11745 (N_11745,N_10140,N_10531);
or U11746 (N_11746,N_10754,N_10533);
nor U11747 (N_11747,N_10550,N_10596);
and U11748 (N_11748,N_10961,N_10608);
nand U11749 (N_11749,N_10329,N_10937);
xor U11750 (N_11750,N_10226,N_10703);
nand U11751 (N_11751,N_10078,N_10706);
and U11752 (N_11752,N_10668,N_10993);
nor U11753 (N_11753,N_10846,N_10666);
nor U11754 (N_11754,N_10926,N_10763);
or U11755 (N_11755,N_10617,N_10442);
xnor U11756 (N_11756,N_10166,N_10033);
or U11757 (N_11757,N_10659,N_10753);
or U11758 (N_11758,N_10632,N_10553);
or U11759 (N_11759,N_10346,N_10883);
xor U11760 (N_11760,N_10640,N_10880);
nor U11761 (N_11761,N_10661,N_10207);
and U11762 (N_11762,N_10266,N_10270);
or U11763 (N_11763,N_10730,N_10503);
and U11764 (N_11764,N_10328,N_10097);
xnor U11765 (N_11765,N_10435,N_10512);
xor U11766 (N_11766,N_10385,N_10186);
or U11767 (N_11767,N_10802,N_10456);
nor U11768 (N_11768,N_10763,N_10513);
or U11769 (N_11769,N_10215,N_10622);
xnor U11770 (N_11770,N_10699,N_10320);
xor U11771 (N_11771,N_10440,N_10203);
or U11772 (N_11772,N_10411,N_10357);
nor U11773 (N_11773,N_10464,N_10914);
nor U11774 (N_11774,N_10593,N_10569);
nand U11775 (N_11775,N_10290,N_10027);
nor U11776 (N_11776,N_10662,N_10116);
xnor U11777 (N_11777,N_10241,N_10422);
or U11778 (N_11778,N_10193,N_10639);
xnor U11779 (N_11779,N_10886,N_10116);
or U11780 (N_11780,N_10258,N_10539);
or U11781 (N_11781,N_10111,N_10983);
or U11782 (N_11782,N_10586,N_10777);
and U11783 (N_11783,N_10001,N_10905);
nor U11784 (N_11784,N_10714,N_10218);
or U11785 (N_11785,N_10353,N_10472);
nor U11786 (N_11786,N_10447,N_10102);
and U11787 (N_11787,N_10826,N_10789);
and U11788 (N_11788,N_10848,N_10025);
and U11789 (N_11789,N_10488,N_10261);
and U11790 (N_11790,N_10671,N_10089);
and U11791 (N_11791,N_10039,N_10757);
or U11792 (N_11792,N_10323,N_10348);
or U11793 (N_11793,N_10785,N_10194);
xnor U11794 (N_11794,N_10781,N_10767);
nand U11795 (N_11795,N_10034,N_10547);
nand U11796 (N_11796,N_10004,N_10126);
xor U11797 (N_11797,N_10656,N_10457);
or U11798 (N_11798,N_10225,N_10061);
xnor U11799 (N_11799,N_10771,N_10070);
nand U11800 (N_11800,N_10403,N_10603);
or U11801 (N_11801,N_10878,N_10232);
xor U11802 (N_11802,N_10196,N_10170);
and U11803 (N_11803,N_10967,N_10477);
and U11804 (N_11804,N_10588,N_10836);
xor U11805 (N_11805,N_10666,N_10627);
nand U11806 (N_11806,N_10276,N_10433);
nand U11807 (N_11807,N_10008,N_10687);
nor U11808 (N_11808,N_10152,N_10559);
or U11809 (N_11809,N_10848,N_10095);
nor U11810 (N_11810,N_10214,N_10223);
nand U11811 (N_11811,N_10274,N_10671);
and U11812 (N_11812,N_10345,N_10279);
or U11813 (N_11813,N_10742,N_10669);
and U11814 (N_11814,N_10599,N_10534);
nor U11815 (N_11815,N_10304,N_10248);
nand U11816 (N_11816,N_10742,N_10273);
nand U11817 (N_11817,N_10643,N_10378);
nand U11818 (N_11818,N_10196,N_10023);
xor U11819 (N_11819,N_10003,N_10773);
or U11820 (N_11820,N_10766,N_10299);
nand U11821 (N_11821,N_10364,N_10283);
nor U11822 (N_11822,N_10469,N_10171);
or U11823 (N_11823,N_10586,N_10245);
and U11824 (N_11824,N_10617,N_10068);
or U11825 (N_11825,N_10561,N_10739);
and U11826 (N_11826,N_10790,N_10742);
and U11827 (N_11827,N_10352,N_10402);
nand U11828 (N_11828,N_10165,N_10538);
nand U11829 (N_11829,N_10353,N_10743);
nor U11830 (N_11830,N_10473,N_10676);
and U11831 (N_11831,N_10463,N_10208);
and U11832 (N_11832,N_10220,N_10395);
xor U11833 (N_11833,N_10596,N_10730);
and U11834 (N_11834,N_10878,N_10695);
and U11835 (N_11835,N_10392,N_10282);
and U11836 (N_11836,N_10920,N_10733);
xor U11837 (N_11837,N_10328,N_10061);
xor U11838 (N_11838,N_10598,N_10624);
or U11839 (N_11839,N_10498,N_10233);
and U11840 (N_11840,N_10097,N_10354);
xor U11841 (N_11841,N_10225,N_10357);
xnor U11842 (N_11842,N_10813,N_10141);
and U11843 (N_11843,N_10675,N_10331);
and U11844 (N_11844,N_10400,N_10913);
or U11845 (N_11845,N_10259,N_10463);
xnor U11846 (N_11846,N_10510,N_10747);
nor U11847 (N_11847,N_10724,N_10272);
nand U11848 (N_11848,N_10170,N_10875);
nand U11849 (N_11849,N_10617,N_10594);
xor U11850 (N_11850,N_10831,N_10634);
and U11851 (N_11851,N_10136,N_10005);
xnor U11852 (N_11852,N_10178,N_10312);
and U11853 (N_11853,N_10103,N_10990);
or U11854 (N_11854,N_10848,N_10468);
nand U11855 (N_11855,N_10248,N_10251);
nand U11856 (N_11856,N_10084,N_10176);
or U11857 (N_11857,N_10506,N_10338);
or U11858 (N_11858,N_10649,N_10512);
and U11859 (N_11859,N_10753,N_10711);
nand U11860 (N_11860,N_10759,N_10206);
nand U11861 (N_11861,N_10236,N_10154);
nor U11862 (N_11862,N_10175,N_10414);
and U11863 (N_11863,N_10123,N_10188);
nand U11864 (N_11864,N_10863,N_10138);
nor U11865 (N_11865,N_10276,N_10997);
nor U11866 (N_11866,N_10924,N_10692);
and U11867 (N_11867,N_10779,N_10289);
and U11868 (N_11868,N_10577,N_10088);
or U11869 (N_11869,N_10917,N_10807);
nand U11870 (N_11870,N_10889,N_10044);
nor U11871 (N_11871,N_10253,N_10798);
nor U11872 (N_11872,N_10042,N_10023);
xor U11873 (N_11873,N_10514,N_10664);
and U11874 (N_11874,N_10627,N_10386);
nor U11875 (N_11875,N_10233,N_10142);
nand U11876 (N_11876,N_10158,N_10127);
and U11877 (N_11877,N_10305,N_10811);
nor U11878 (N_11878,N_10713,N_10673);
nor U11879 (N_11879,N_10597,N_10908);
and U11880 (N_11880,N_10707,N_10505);
or U11881 (N_11881,N_10756,N_10325);
nor U11882 (N_11882,N_10220,N_10775);
and U11883 (N_11883,N_10837,N_10010);
and U11884 (N_11884,N_10664,N_10755);
nand U11885 (N_11885,N_10808,N_10430);
xnor U11886 (N_11886,N_10474,N_10796);
xor U11887 (N_11887,N_10333,N_10141);
or U11888 (N_11888,N_10897,N_10178);
and U11889 (N_11889,N_10426,N_10935);
and U11890 (N_11890,N_10181,N_10487);
nor U11891 (N_11891,N_10528,N_10935);
or U11892 (N_11892,N_10460,N_10063);
and U11893 (N_11893,N_10665,N_10459);
nor U11894 (N_11894,N_10337,N_10009);
nor U11895 (N_11895,N_10363,N_10888);
and U11896 (N_11896,N_10166,N_10536);
or U11897 (N_11897,N_10448,N_10008);
xor U11898 (N_11898,N_10661,N_10949);
nor U11899 (N_11899,N_10626,N_10104);
xnor U11900 (N_11900,N_10294,N_10790);
xnor U11901 (N_11901,N_10895,N_10544);
and U11902 (N_11902,N_10917,N_10307);
xor U11903 (N_11903,N_10221,N_10950);
xnor U11904 (N_11904,N_10742,N_10082);
nand U11905 (N_11905,N_10211,N_10703);
nand U11906 (N_11906,N_10192,N_10744);
nand U11907 (N_11907,N_10005,N_10299);
and U11908 (N_11908,N_10045,N_10677);
xor U11909 (N_11909,N_10695,N_10443);
and U11910 (N_11910,N_10379,N_10864);
xnor U11911 (N_11911,N_10308,N_10402);
xnor U11912 (N_11912,N_10080,N_10107);
or U11913 (N_11913,N_10700,N_10650);
or U11914 (N_11914,N_10033,N_10241);
nor U11915 (N_11915,N_10905,N_10886);
nor U11916 (N_11916,N_10509,N_10529);
nand U11917 (N_11917,N_10780,N_10985);
xnor U11918 (N_11918,N_10607,N_10086);
nand U11919 (N_11919,N_10404,N_10587);
nor U11920 (N_11920,N_10623,N_10918);
xnor U11921 (N_11921,N_10501,N_10639);
nor U11922 (N_11922,N_10777,N_10404);
nor U11923 (N_11923,N_10585,N_10359);
and U11924 (N_11924,N_10700,N_10588);
and U11925 (N_11925,N_10718,N_10169);
nor U11926 (N_11926,N_10283,N_10774);
nor U11927 (N_11927,N_10460,N_10682);
xor U11928 (N_11928,N_10981,N_10542);
xnor U11929 (N_11929,N_10574,N_10084);
nor U11930 (N_11930,N_10511,N_10582);
or U11931 (N_11931,N_10027,N_10044);
or U11932 (N_11932,N_10524,N_10997);
nor U11933 (N_11933,N_10351,N_10591);
or U11934 (N_11934,N_10321,N_10833);
xnor U11935 (N_11935,N_10922,N_10836);
nand U11936 (N_11936,N_10321,N_10344);
nand U11937 (N_11937,N_10018,N_10071);
or U11938 (N_11938,N_10986,N_10244);
and U11939 (N_11939,N_10362,N_10986);
and U11940 (N_11940,N_10313,N_10303);
xor U11941 (N_11941,N_10730,N_10281);
nor U11942 (N_11942,N_10420,N_10474);
and U11943 (N_11943,N_10286,N_10152);
xor U11944 (N_11944,N_10888,N_10225);
and U11945 (N_11945,N_10291,N_10058);
or U11946 (N_11946,N_10914,N_10445);
nand U11947 (N_11947,N_10302,N_10862);
nand U11948 (N_11948,N_10224,N_10792);
nor U11949 (N_11949,N_10582,N_10013);
or U11950 (N_11950,N_10467,N_10638);
and U11951 (N_11951,N_10484,N_10300);
xnor U11952 (N_11952,N_10346,N_10982);
xor U11953 (N_11953,N_10429,N_10040);
nor U11954 (N_11954,N_10845,N_10478);
nor U11955 (N_11955,N_10640,N_10220);
xnor U11956 (N_11956,N_10305,N_10051);
or U11957 (N_11957,N_10585,N_10324);
and U11958 (N_11958,N_10493,N_10856);
xor U11959 (N_11959,N_10455,N_10616);
nand U11960 (N_11960,N_10304,N_10694);
or U11961 (N_11961,N_10145,N_10473);
or U11962 (N_11962,N_10019,N_10558);
nor U11963 (N_11963,N_10251,N_10351);
nand U11964 (N_11964,N_10111,N_10985);
nor U11965 (N_11965,N_10212,N_10669);
or U11966 (N_11966,N_10640,N_10489);
xnor U11967 (N_11967,N_10352,N_10838);
nand U11968 (N_11968,N_10467,N_10523);
nor U11969 (N_11969,N_10575,N_10431);
nand U11970 (N_11970,N_10340,N_10687);
nor U11971 (N_11971,N_10123,N_10883);
nor U11972 (N_11972,N_10507,N_10318);
nor U11973 (N_11973,N_10205,N_10541);
nand U11974 (N_11974,N_10510,N_10794);
nor U11975 (N_11975,N_10803,N_10761);
nand U11976 (N_11976,N_10463,N_10973);
nor U11977 (N_11977,N_10637,N_10967);
nand U11978 (N_11978,N_10813,N_10569);
or U11979 (N_11979,N_10979,N_10541);
or U11980 (N_11980,N_10329,N_10548);
or U11981 (N_11981,N_10969,N_10900);
or U11982 (N_11982,N_10107,N_10167);
nor U11983 (N_11983,N_10181,N_10056);
or U11984 (N_11984,N_10714,N_10017);
nor U11985 (N_11985,N_10114,N_10810);
xor U11986 (N_11986,N_10283,N_10147);
xnor U11987 (N_11987,N_10183,N_10281);
xnor U11988 (N_11988,N_10947,N_10991);
or U11989 (N_11989,N_10867,N_10020);
nor U11990 (N_11990,N_10054,N_10541);
nor U11991 (N_11991,N_10027,N_10764);
nand U11992 (N_11992,N_10836,N_10740);
and U11993 (N_11993,N_10015,N_10288);
xnor U11994 (N_11994,N_10169,N_10137);
and U11995 (N_11995,N_10291,N_10388);
or U11996 (N_11996,N_10705,N_10118);
and U11997 (N_11997,N_10997,N_10319);
or U11998 (N_11998,N_10733,N_10996);
and U11999 (N_11999,N_10037,N_10968);
and U12000 (N_12000,N_11201,N_11507);
nor U12001 (N_12001,N_11819,N_11967);
nand U12002 (N_12002,N_11028,N_11412);
or U12003 (N_12003,N_11980,N_11692);
or U12004 (N_12004,N_11287,N_11673);
nor U12005 (N_12005,N_11568,N_11422);
and U12006 (N_12006,N_11892,N_11738);
nor U12007 (N_12007,N_11853,N_11563);
and U12008 (N_12008,N_11255,N_11119);
nand U12009 (N_12009,N_11319,N_11887);
or U12010 (N_12010,N_11624,N_11452);
nand U12011 (N_12011,N_11803,N_11053);
or U12012 (N_12012,N_11664,N_11289);
nand U12013 (N_12013,N_11597,N_11162);
nand U12014 (N_12014,N_11812,N_11654);
nor U12015 (N_12015,N_11868,N_11690);
nor U12016 (N_12016,N_11665,N_11639);
nand U12017 (N_12017,N_11847,N_11099);
or U12018 (N_12018,N_11310,N_11503);
nor U12019 (N_12019,N_11703,N_11098);
xnor U12020 (N_12020,N_11934,N_11519);
xor U12021 (N_12021,N_11882,N_11033);
nand U12022 (N_12022,N_11547,N_11916);
or U12023 (N_12023,N_11393,N_11727);
and U12024 (N_12024,N_11689,N_11527);
and U12025 (N_12025,N_11754,N_11094);
xnor U12026 (N_12026,N_11675,N_11408);
and U12027 (N_12027,N_11591,N_11721);
nand U12028 (N_12028,N_11757,N_11249);
nand U12029 (N_12029,N_11062,N_11686);
xor U12030 (N_12030,N_11663,N_11891);
xnor U12031 (N_12031,N_11797,N_11630);
or U12032 (N_12032,N_11950,N_11961);
and U12033 (N_12033,N_11962,N_11268);
nor U12034 (N_12034,N_11646,N_11065);
and U12035 (N_12035,N_11500,N_11359);
nor U12036 (N_12036,N_11341,N_11533);
xnor U12037 (N_12037,N_11383,N_11059);
or U12038 (N_12038,N_11538,N_11279);
nor U12039 (N_12039,N_11171,N_11710);
or U12040 (N_12040,N_11859,N_11518);
and U12041 (N_12041,N_11904,N_11340);
nor U12042 (N_12042,N_11571,N_11264);
nor U12043 (N_12043,N_11579,N_11331);
nor U12044 (N_12044,N_11946,N_11873);
nor U12045 (N_12045,N_11282,N_11932);
and U12046 (N_12046,N_11574,N_11076);
or U12047 (N_12047,N_11577,N_11292);
nor U12048 (N_12048,N_11371,N_11169);
nor U12049 (N_12049,N_11894,N_11149);
nand U12050 (N_12050,N_11970,N_11711);
or U12051 (N_12051,N_11130,N_11650);
and U12052 (N_12052,N_11242,N_11016);
nor U12053 (N_12053,N_11203,N_11875);
xnor U12054 (N_12054,N_11040,N_11036);
nor U12055 (N_12055,N_11862,N_11318);
and U12056 (N_12056,N_11281,N_11800);
or U12057 (N_12057,N_11725,N_11479);
or U12058 (N_12058,N_11958,N_11813);
nor U12059 (N_12059,N_11621,N_11253);
nand U12060 (N_12060,N_11517,N_11442);
and U12061 (N_12061,N_11489,N_11768);
xor U12062 (N_12062,N_11009,N_11481);
nor U12063 (N_12063,N_11222,N_11997);
nand U12064 (N_12064,N_11746,N_11155);
or U12065 (N_12065,N_11845,N_11039);
xor U12066 (N_12066,N_11349,N_11783);
xor U12067 (N_12067,N_11638,N_11485);
or U12068 (N_12068,N_11974,N_11909);
nand U12069 (N_12069,N_11532,N_11267);
nor U12070 (N_12070,N_11195,N_11251);
nand U12071 (N_12071,N_11214,N_11930);
xnor U12072 (N_12072,N_11590,N_11271);
and U12073 (N_12073,N_11756,N_11976);
xor U12074 (N_12074,N_11414,N_11122);
and U12075 (N_12075,N_11830,N_11573);
xnor U12076 (N_12076,N_11776,N_11954);
or U12077 (N_12077,N_11594,N_11304);
or U12078 (N_12078,N_11717,N_11982);
and U12079 (N_12079,N_11323,N_11258);
xor U12080 (N_12080,N_11123,N_11805);
nor U12081 (N_12081,N_11933,N_11101);
and U12082 (N_12082,N_11668,N_11430);
and U12083 (N_12083,N_11494,N_11669);
and U12084 (N_12084,N_11620,N_11990);
nand U12085 (N_12085,N_11237,N_11838);
nand U12086 (N_12086,N_11354,N_11188);
and U12087 (N_12087,N_11248,N_11491);
nor U12088 (N_12088,N_11213,N_11423);
nand U12089 (N_12089,N_11993,N_11132);
nand U12090 (N_12090,N_11178,N_11615);
nor U12091 (N_12091,N_11666,N_11938);
nor U12092 (N_12092,N_11870,N_11957);
nor U12093 (N_12093,N_11534,N_11295);
and U12094 (N_12094,N_11326,N_11339);
or U12095 (N_12095,N_11513,N_11739);
nand U12096 (N_12096,N_11150,N_11045);
or U12097 (N_12097,N_11157,N_11451);
or U12098 (N_12098,N_11308,N_11979);
nor U12099 (N_12099,N_11667,N_11566);
and U12100 (N_12100,N_11476,N_11345);
and U12101 (N_12101,N_11823,N_11029);
nand U12102 (N_12102,N_11587,N_11885);
nor U12103 (N_12103,N_11828,N_11385);
and U12104 (N_12104,N_11198,N_11161);
and U12105 (N_12105,N_11632,N_11735);
xor U12106 (N_12106,N_11469,N_11225);
xor U12107 (N_12107,N_11116,N_11083);
and U12108 (N_12108,N_11761,N_11606);
and U12109 (N_12109,N_11484,N_11762);
or U12110 (N_12110,N_11593,N_11411);
and U12111 (N_12111,N_11835,N_11963);
and U12112 (N_12112,N_11454,N_11866);
nor U12113 (N_12113,N_11680,N_11113);
nand U12114 (N_12114,N_11899,N_11446);
nand U12115 (N_12115,N_11081,N_11205);
or U12116 (N_12116,N_11917,N_11370);
and U12117 (N_12117,N_11473,N_11106);
xor U12118 (N_12118,N_11181,N_11030);
nor U12119 (N_12119,N_11978,N_11464);
xor U12120 (N_12120,N_11733,N_11086);
and U12121 (N_12121,N_11965,N_11775);
nor U12122 (N_12122,N_11625,N_11269);
nor U12123 (N_12123,N_11512,N_11701);
and U12124 (N_12124,N_11350,N_11804);
xnor U12125 (N_12125,N_11325,N_11855);
and U12126 (N_12126,N_11937,N_11832);
nand U12127 (N_12127,N_11501,N_11005);
xor U12128 (N_12128,N_11023,N_11296);
nand U12129 (N_12129,N_11444,N_11784);
or U12130 (N_12130,N_11802,N_11709);
nor U12131 (N_12131,N_11228,N_11170);
or U12132 (N_12132,N_11063,N_11025);
xor U12133 (N_12133,N_11031,N_11392);
nand U12134 (N_12134,N_11960,N_11004);
or U12135 (N_12135,N_11037,N_11440);
or U12136 (N_12136,N_11107,N_11486);
nand U12137 (N_12137,N_11343,N_11187);
xnor U12138 (N_12138,N_11857,N_11194);
or U12139 (N_12139,N_11315,N_11402);
nand U12140 (N_12140,N_11604,N_11919);
nor U12141 (N_12141,N_11043,N_11889);
or U12142 (N_12142,N_11372,N_11927);
nand U12143 (N_12143,N_11439,N_11944);
nand U12144 (N_12144,N_11276,N_11151);
xor U12145 (N_12145,N_11089,N_11854);
nand U12146 (N_12146,N_11897,N_11660);
and U12147 (N_12147,N_11105,N_11619);
and U12148 (N_12148,N_11360,N_11312);
nor U12149 (N_12149,N_11229,N_11344);
xnor U12150 (N_12150,N_11219,N_11465);
xor U12151 (N_12151,N_11626,N_11734);
nor U12152 (N_12152,N_11273,N_11376);
nor U12153 (N_12153,N_11696,N_11796);
nor U12154 (N_12154,N_11285,N_11262);
nand U12155 (N_12155,N_11226,N_11000);
xor U12156 (N_12156,N_11693,N_11139);
xnor U12157 (N_12157,N_11061,N_11699);
xor U12158 (N_12158,N_11453,N_11792);
and U12159 (N_12159,N_11850,N_11495);
nor U12160 (N_12160,N_11069,N_11910);
nor U12161 (N_12161,N_11760,N_11233);
and U12162 (N_12162,N_11147,N_11881);
nand U12163 (N_12163,N_11208,N_11247);
nand U12164 (N_12164,N_11833,N_11179);
or U12165 (N_12165,N_11541,N_11622);
nand U12166 (N_12166,N_11490,N_11871);
and U12167 (N_12167,N_11841,N_11070);
nor U12168 (N_12168,N_11723,N_11457);
nand U12169 (N_12169,N_11763,N_11002);
and U12170 (N_12170,N_11988,N_11297);
nand U12171 (N_12171,N_11911,N_11348);
or U12172 (N_12172,N_11715,N_11356);
xor U12173 (N_12173,N_11460,N_11050);
xnor U12174 (N_12174,N_11006,N_11462);
nand U12175 (N_12175,N_11896,N_11102);
and U12176 (N_12176,N_11562,N_11731);
nand U12177 (N_12177,N_11096,N_11567);
nor U12178 (N_12178,N_11018,N_11218);
and U12179 (N_12179,N_11280,N_11821);
or U12180 (N_12180,N_11900,N_11172);
or U12181 (N_12181,N_11288,N_11653);
nand U12182 (N_12182,N_11959,N_11134);
and U12183 (N_12183,N_11051,N_11516);
nand U12184 (N_12184,N_11397,N_11243);
nand U12185 (N_12185,N_11546,N_11109);
nor U12186 (N_12186,N_11623,N_11712);
nor U12187 (N_12187,N_11921,N_11261);
and U12188 (N_12188,N_11421,N_11694);
nand U12189 (N_12189,N_11374,N_11953);
nand U12190 (N_12190,N_11092,N_11608);
xnor U12191 (N_12191,N_11918,N_11191);
or U12192 (N_12192,N_11683,N_11972);
and U12193 (N_12193,N_11366,N_11022);
and U12194 (N_12194,N_11656,N_11770);
or U12195 (N_12195,N_11060,N_11324);
xor U12196 (N_12196,N_11379,N_11508);
xor U12197 (N_12197,N_11204,N_11111);
or U12198 (N_12198,N_11174,N_11284);
nand U12199 (N_12199,N_11613,N_11415);
xnor U12200 (N_12200,N_11886,N_11940);
nor U12201 (N_12201,N_11521,N_11795);
xor U12202 (N_12202,N_11555,N_11975);
xnor U12203 (N_12203,N_11466,N_11215);
nand U12204 (N_12204,N_11766,N_11554);
and U12205 (N_12205,N_11759,N_11011);
nand U12206 (N_12206,N_11601,N_11017);
or U12207 (N_12207,N_11245,N_11814);
xor U12208 (N_12208,N_11498,N_11322);
and U12209 (N_12209,N_11265,N_11286);
and U12210 (N_12210,N_11544,N_11396);
and U12211 (N_12211,N_11952,N_11382);
nand U12212 (N_12212,N_11945,N_11335);
nor U12213 (N_12213,N_11742,N_11448);
nand U12214 (N_12214,N_11391,N_11274);
and U12215 (N_12215,N_11337,N_11266);
xor U12216 (N_12216,N_11614,N_11584);
and U12217 (N_12217,N_11145,N_11216);
and U12218 (N_12218,N_11649,N_11071);
nor U12219 (N_12219,N_11394,N_11112);
nor U12220 (N_12220,N_11144,N_11263);
or U12221 (N_12221,N_11244,N_11200);
nor U12222 (N_12222,N_11920,N_11605);
nor U12223 (N_12223,N_11082,N_11472);
nand U12224 (N_12224,N_11865,N_11941);
nor U12225 (N_12225,N_11458,N_11015);
nor U12226 (N_12226,N_11407,N_11642);
xor U12227 (N_12227,N_11602,N_11674);
nand U12228 (N_12228,N_11774,N_11552);
nor U12229 (N_12229,N_11992,N_11038);
and U12230 (N_12230,N_11809,N_11557);
and U12231 (N_12231,N_11852,N_11403);
xnor U12232 (N_12232,N_11152,N_11585);
nor U12233 (N_12233,N_11588,N_11332);
nand U12234 (N_12234,N_11596,N_11115);
and U12235 (N_12235,N_11902,N_11177);
or U12236 (N_12236,N_11915,N_11592);
xnor U12237 (N_12237,N_11589,N_11197);
or U12238 (N_12238,N_11781,N_11504);
and U12239 (N_12239,N_11133,N_11603);
and U12240 (N_12240,N_11355,N_11879);
nand U12241 (N_12241,N_11166,N_11232);
xnor U12242 (N_12242,N_11073,N_11328);
nand U12243 (N_12243,N_11939,N_11629);
or U12244 (N_12244,N_11316,N_11861);
xor U12245 (N_12245,N_11126,N_11008);
and U12246 (N_12246,N_11450,N_11931);
nor U12247 (N_12247,N_11925,N_11492);
and U12248 (N_12248,N_11075,N_11447);
xnor U12249 (N_12249,N_11836,N_11146);
nor U12250 (N_12250,N_11272,N_11235);
nor U12251 (N_12251,N_11578,N_11309);
and U12252 (N_12252,N_11353,N_11346);
nor U12253 (N_12253,N_11523,N_11640);
nor U12254 (N_12254,N_11505,N_11388);
xor U12255 (N_12255,N_11260,N_11080);
or U12256 (N_12256,N_11032,N_11072);
or U12257 (N_12257,N_11026,N_11951);
or U12258 (N_12258,N_11670,N_11685);
nor U12259 (N_12259,N_11704,N_11947);
xnor U12260 (N_12260,N_11118,N_11807);
nand U12261 (N_12261,N_11750,N_11810);
and U12262 (N_12262,N_11645,N_11510);
nand U12263 (N_12263,N_11236,N_11455);
nand U12264 (N_12264,N_11129,N_11981);
and U12265 (N_12265,N_11483,N_11676);
or U12266 (N_12266,N_11827,N_11820);
xnor U12267 (N_12267,N_11404,N_11419);
nand U12268 (N_12268,N_11661,N_11067);
and U12269 (N_12269,N_11747,N_11793);
nor U12270 (N_12270,N_11336,N_11048);
or U12271 (N_12271,N_11124,N_11636);
xor U12272 (N_12272,N_11773,N_11365);
nand U12273 (N_12273,N_11684,N_11426);
xnor U12274 (N_12274,N_11716,N_11375);
and U12275 (N_12275,N_11856,N_11443);
or U12276 (N_12276,N_11876,N_11586);
and U12277 (N_12277,N_11330,N_11878);
nand U12278 (N_12278,N_11390,N_11502);
or U12279 (N_12279,N_11429,N_11358);
xor U12280 (N_12280,N_11138,N_11548);
nand U12281 (N_12281,N_11436,N_11190);
nand U12282 (N_12282,N_11474,N_11764);
nor U12283 (N_12283,N_11782,N_11074);
xor U12284 (N_12284,N_11068,N_11829);
xor U12285 (N_12285,N_11173,N_11539);
and U12286 (N_12286,N_11482,N_11989);
or U12287 (N_12287,N_11987,N_11041);
or U12288 (N_12288,N_11186,N_11908);
nand U12289 (N_12289,N_11700,N_11837);
xnor U12290 (N_12290,N_11751,N_11313);
or U12291 (N_12291,N_11769,N_11561);
or U12292 (N_12292,N_11898,N_11884);
nor U12293 (N_12293,N_11305,N_11826);
xor U12294 (N_12294,N_11445,N_11798);
xor U12295 (N_12295,N_11140,N_11831);
nand U12296 (N_12296,N_11034,N_11655);
xor U12297 (N_12297,N_11314,N_11175);
and U12298 (N_12298,N_11231,N_11565);
or U12299 (N_12299,N_11078,N_11535);
nand U12300 (N_12300,N_11991,N_11609);
and U12301 (N_12301,N_11895,N_11583);
nand U12302 (N_12302,N_11478,N_11634);
nor U12303 (N_12303,N_11434,N_11558);
xor U12304 (N_12304,N_11526,N_11441);
xor U12305 (N_12305,N_11432,N_11955);
xor U12306 (N_12306,N_11531,N_11816);
nor U12307 (N_12307,N_11706,N_11400);
nand U12308 (N_12308,N_11525,N_11199);
and U12309 (N_12309,N_11867,N_11298);
and U12310 (N_12310,N_11128,N_11291);
or U12311 (N_12311,N_11327,N_11643);
nand U12312 (N_12312,N_11611,N_11748);
nor U12313 (N_12313,N_11582,N_11801);
and U12314 (N_12314,N_11506,N_11347);
nand U12315 (N_12315,N_11741,N_11737);
xnor U12316 (N_12316,N_11057,N_11097);
xnor U12317 (N_12317,N_11671,N_11020);
nand U12318 (N_12318,N_11651,N_11914);
nor U12319 (N_12319,N_11822,N_11467);
xor U12320 (N_12320,N_11368,N_11277);
xor U12321 (N_12321,N_11872,N_11743);
and U12322 (N_12322,N_11406,N_11311);
nand U12323 (N_12323,N_11695,N_11007);
nand U12324 (N_12324,N_11220,N_11688);
nor U12325 (N_12325,N_11417,N_11569);
xnor U12326 (N_12326,N_11389,N_11117);
and U12327 (N_12327,N_11787,N_11752);
nor U12328 (N_12328,N_11035,N_11163);
nand U12329 (N_12329,N_11252,N_11104);
xor U12330 (N_12330,N_11398,N_11806);
or U12331 (N_12331,N_11905,N_11536);
nand U12332 (N_12332,N_11079,N_11405);
nor U12333 (N_12333,N_11681,N_11647);
xor U12334 (N_12334,N_11087,N_11021);
xnor U12335 (N_12335,N_11321,N_11811);
xor U12336 (N_12336,N_11736,N_11256);
and U12337 (N_12337,N_11424,N_11046);
and U12338 (N_12338,N_11241,N_11913);
xor U12339 (N_12339,N_11682,N_11209);
xor U12340 (N_12340,N_11928,N_11010);
or U12341 (N_12341,N_11851,N_11246);
or U12342 (N_12342,N_11493,N_11628);
xor U12343 (N_12343,N_11788,N_11912);
nand U12344 (N_12344,N_11869,N_11984);
and U12345 (N_12345,N_11511,N_11942);
nor U12346 (N_12346,N_11014,N_11637);
nand U12347 (N_12347,N_11713,N_11409);
or U12348 (N_12348,N_11641,N_11719);
xor U12349 (N_12349,N_11238,N_11250);
xor U12350 (N_12350,N_11848,N_11860);
and U12351 (N_12351,N_11054,N_11971);
and U12352 (N_12352,N_11528,N_11672);
and U12353 (N_12353,N_11790,N_11537);
nor U12354 (N_12354,N_11027,N_11202);
nor U12355 (N_12355,N_11658,N_11329);
nand U12356 (N_12356,N_11758,N_11165);
nand U12357 (N_12357,N_11189,N_11791);
nor U12358 (N_12358,N_11223,N_11679);
nor U12359 (N_12359,N_11459,N_11019);
xnor U12360 (N_12360,N_11088,N_11293);
nor U12361 (N_12361,N_11294,N_11678);
nand U12362 (N_12362,N_11572,N_11652);
nand U12363 (N_12363,N_11948,N_11283);
nand U12364 (N_12364,N_11732,N_11996);
nand U12365 (N_12365,N_11581,N_11120);
or U12366 (N_12366,N_11718,N_11413);
nand U12367 (N_12367,N_11141,N_11143);
and U12368 (N_12368,N_11530,N_11363);
xor U12369 (N_12369,N_11488,N_11299);
nand U12370 (N_12370,N_11817,N_11730);
and U12371 (N_12371,N_11771,N_11167);
nand U12372 (N_12372,N_11224,N_11985);
xnor U12373 (N_12373,N_11131,N_11598);
and U12374 (N_12374,N_11239,N_11780);
or U12375 (N_12375,N_11342,N_11212);
nand U12376 (N_12376,N_11786,N_11923);
xor U12377 (N_12377,N_11983,N_11744);
or U12378 (N_12378,N_11003,N_11777);
and U12379 (N_12379,N_11617,N_11001);
nand U12380 (N_12380,N_11657,N_11595);
or U12381 (N_12381,N_11399,N_11425);
and U12382 (N_12382,N_11509,N_11883);
xnor U12383 (N_12383,N_11922,N_11153);
and U12384 (N_12384,N_11351,N_11352);
and U12385 (N_12385,N_11367,N_11556);
nor U12386 (N_12386,N_11480,N_11522);
xor U12387 (N_12387,N_11290,N_11275);
nand U12388 (N_12388,N_11749,N_11825);
or U12389 (N_12389,N_11612,N_11077);
and U12390 (N_12390,N_11728,N_11843);
or U12391 (N_12391,N_11049,N_11977);
and U12392 (N_12392,N_11994,N_11986);
nand U12393 (N_12393,N_11168,N_11785);
nor U12394 (N_12394,N_11844,N_11789);
and U12395 (N_12395,N_11999,N_11100);
nor U12396 (N_12396,N_11906,N_11697);
nand U12397 (N_12397,N_11520,N_11599);
nand U12398 (N_12398,N_11013,N_11230);
or U12399 (N_12399,N_11470,N_11137);
or U12400 (N_12400,N_11936,N_11576);
or U12401 (N_12401,N_11193,N_11560);
or U12402 (N_12402,N_11012,N_11477);
xnor U12403 (N_12403,N_11499,N_11745);
nor U12404 (N_12404,N_11184,N_11303);
nor U12405 (N_12405,N_11160,N_11420);
or U12406 (N_12406,N_11361,N_11461);
nor U12407 (N_12407,N_11257,N_11708);
and U12408 (N_12408,N_11127,N_11090);
or U12409 (N_12409,N_11755,N_11540);
and U12410 (N_12410,N_11427,N_11818);
xor U12411 (N_12411,N_11618,N_11926);
and U12412 (N_12412,N_11549,N_11369);
xor U12413 (N_12413,N_11362,N_11156);
nand U12414 (N_12414,N_11206,N_11475);
and U12415 (N_12415,N_11108,N_11428);
nand U12416 (N_12416,N_11091,N_11136);
xnor U12417 (N_12417,N_11395,N_11471);
nor U12418 (N_12418,N_11627,N_11438);
nor U12419 (N_12419,N_11767,N_11164);
nand U12420 (N_12420,N_11468,N_11373);
and U12421 (N_12421,N_11888,N_11211);
or U12422 (N_12422,N_11662,N_11949);
xor U12423 (N_12423,N_11648,N_11705);
nor U12424 (N_12424,N_11024,N_11416);
xnor U12425 (N_12425,N_11564,N_11207);
or U12426 (N_12426,N_11724,N_11142);
nor U12427 (N_12427,N_11877,N_11056);
nor U12428 (N_12428,N_11559,N_11765);
nand U12429 (N_12429,N_11995,N_11874);
xnor U12430 (N_12430,N_11497,N_11553);
xnor U12431 (N_12431,N_11514,N_11772);
nor U12432 (N_12432,N_11616,N_11924);
xnor U12433 (N_12433,N_11047,N_11095);
and U12434 (N_12434,N_11846,N_11306);
nand U12435 (N_12435,N_11066,N_11148);
or U12436 (N_12436,N_11550,N_11720);
and U12437 (N_12437,N_11815,N_11487);
or U12438 (N_12438,N_11698,N_11435);
and U12439 (N_12439,N_11176,N_11042);
nand U12440 (N_12440,N_11158,N_11849);
nand U12441 (N_12441,N_11259,N_11159);
nand U12442 (N_12442,N_11307,N_11890);
and U12443 (N_12443,N_11357,N_11956);
nor U12444 (N_12444,N_11935,N_11384);
or U12445 (N_12445,N_11180,N_11210);
or U12446 (N_12446,N_11515,N_11707);
and U12447 (N_12447,N_11110,N_11794);
and U12448 (N_12448,N_11114,N_11691);
or U12449 (N_12449,N_11799,N_11320);
xor U12450 (N_12450,N_11125,N_11687);
nand U12451 (N_12451,N_11901,N_11880);
and U12452 (N_12452,N_11183,N_11401);
or U12453 (N_12453,N_11824,N_11570);
nor U12454 (N_12454,N_11387,N_11726);
and U12455 (N_12455,N_11302,N_11052);
xor U12456 (N_12456,N_11386,N_11633);
nor U12457 (N_12457,N_11103,N_11381);
nand U12458 (N_12458,N_11964,N_11364);
nor U12459 (N_12459,N_11496,N_11410);
or U12460 (N_12460,N_11575,N_11433);
nand U12461 (N_12461,N_11437,N_11064);
and U12462 (N_12462,N_11702,N_11234);
nor U12463 (N_12463,N_11893,N_11449);
nor U12464 (N_12464,N_11093,N_11929);
xnor U12465 (N_12465,N_11580,N_11610);
nor U12466 (N_12466,N_11842,N_11185);
and U12467 (N_12467,N_11300,N_11966);
xor U12468 (N_12468,N_11431,N_11968);
or U12469 (N_12469,N_11753,N_11524);
nor U12470 (N_12470,N_11192,N_11377);
or U12471 (N_12471,N_11722,N_11121);
nand U12472 (N_12472,N_11154,N_11529);
or U12473 (N_12473,N_11644,N_11864);
nand U12474 (N_12474,N_11714,N_11631);
or U12475 (N_12475,N_11545,N_11227);
xor U12476 (N_12476,N_11317,N_11196);
and U12477 (N_12477,N_11903,N_11542);
nand U12478 (N_12478,N_11182,N_11378);
and U12479 (N_12479,N_11270,N_11085);
nand U12480 (N_12480,N_11334,N_11221);
nor U12481 (N_12481,N_11973,N_11418);
nand U12482 (N_12482,N_11858,N_11778);
and U12483 (N_12483,N_11779,N_11740);
nand U12484 (N_12484,N_11333,N_11463);
or U12485 (N_12485,N_11044,N_11808);
or U12486 (N_12486,N_11863,N_11635);
and U12487 (N_12487,N_11380,N_11839);
xnor U12488 (N_12488,N_11301,N_11729);
xnor U12489 (N_12489,N_11217,N_11677);
nand U12490 (N_12490,N_11278,N_11456);
and U12491 (N_12491,N_11055,N_11338);
nor U12492 (N_12492,N_11907,N_11551);
nand U12493 (N_12493,N_11998,N_11840);
and U12494 (N_12494,N_11058,N_11135);
nor U12495 (N_12495,N_11943,N_11254);
xnor U12496 (N_12496,N_11607,N_11834);
and U12497 (N_12497,N_11240,N_11543);
xor U12498 (N_12498,N_11969,N_11659);
and U12499 (N_12499,N_11600,N_11084);
and U12500 (N_12500,N_11974,N_11246);
nand U12501 (N_12501,N_11421,N_11900);
and U12502 (N_12502,N_11521,N_11745);
nor U12503 (N_12503,N_11639,N_11917);
nand U12504 (N_12504,N_11191,N_11033);
nor U12505 (N_12505,N_11955,N_11011);
xor U12506 (N_12506,N_11129,N_11670);
nand U12507 (N_12507,N_11595,N_11497);
nand U12508 (N_12508,N_11296,N_11730);
nor U12509 (N_12509,N_11458,N_11238);
or U12510 (N_12510,N_11741,N_11723);
nand U12511 (N_12511,N_11854,N_11407);
nand U12512 (N_12512,N_11534,N_11872);
nand U12513 (N_12513,N_11605,N_11116);
nand U12514 (N_12514,N_11922,N_11441);
and U12515 (N_12515,N_11071,N_11918);
nor U12516 (N_12516,N_11183,N_11625);
nor U12517 (N_12517,N_11733,N_11878);
nand U12518 (N_12518,N_11068,N_11535);
nor U12519 (N_12519,N_11722,N_11713);
xnor U12520 (N_12520,N_11524,N_11590);
xnor U12521 (N_12521,N_11950,N_11885);
nand U12522 (N_12522,N_11047,N_11309);
or U12523 (N_12523,N_11712,N_11372);
and U12524 (N_12524,N_11716,N_11541);
nand U12525 (N_12525,N_11688,N_11402);
and U12526 (N_12526,N_11626,N_11453);
nor U12527 (N_12527,N_11731,N_11564);
nand U12528 (N_12528,N_11022,N_11559);
and U12529 (N_12529,N_11706,N_11666);
nand U12530 (N_12530,N_11195,N_11003);
and U12531 (N_12531,N_11845,N_11290);
or U12532 (N_12532,N_11515,N_11815);
or U12533 (N_12533,N_11428,N_11343);
nor U12534 (N_12534,N_11194,N_11756);
or U12535 (N_12535,N_11060,N_11737);
nand U12536 (N_12536,N_11038,N_11462);
nand U12537 (N_12537,N_11045,N_11183);
xor U12538 (N_12538,N_11500,N_11953);
nor U12539 (N_12539,N_11479,N_11372);
nand U12540 (N_12540,N_11322,N_11456);
nor U12541 (N_12541,N_11760,N_11898);
and U12542 (N_12542,N_11906,N_11304);
or U12543 (N_12543,N_11963,N_11276);
nor U12544 (N_12544,N_11260,N_11504);
nor U12545 (N_12545,N_11126,N_11717);
xor U12546 (N_12546,N_11275,N_11565);
nor U12547 (N_12547,N_11012,N_11752);
xnor U12548 (N_12548,N_11705,N_11931);
or U12549 (N_12549,N_11020,N_11994);
nor U12550 (N_12550,N_11228,N_11715);
xor U12551 (N_12551,N_11614,N_11458);
nor U12552 (N_12552,N_11179,N_11876);
and U12553 (N_12553,N_11729,N_11118);
and U12554 (N_12554,N_11827,N_11291);
xnor U12555 (N_12555,N_11553,N_11915);
xor U12556 (N_12556,N_11678,N_11806);
or U12557 (N_12557,N_11252,N_11722);
nor U12558 (N_12558,N_11997,N_11104);
nand U12559 (N_12559,N_11258,N_11014);
or U12560 (N_12560,N_11365,N_11636);
or U12561 (N_12561,N_11630,N_11221);
xnor U12562 (N_12562,N_11754,N_11202);
nor U12563 (N_12563,N_11373,N_11386);
and U12564 (N_12564,N_11034,N_11406);
nor U12565 (N_12565,N_11701,N_11656);
and U12566 (N_12566,N_11689,N_11143);
nand U12567 (N_12567,N_11507,N_11720);
nor U12568 (N_12568,N_11706,N_11538);
xor U12569 (N_12569,N_11485,N_11795);
nor U12570 (N_12570,N_11117,N_11875);
or U12571 (N_12571,N_11419,N_11909);
nand U12572 (N_12572,N_11307,N_11951);
nor U12573 (N_12573,N_11901,N_11222);
or U12574 (N_12574,N_11797,N_11528);
nand U12575 (N_12575,N_11794,N_11239);
or U12576 (N_12576,N_11091,N_11237);
and U12577 (N_12577,N_11120,N_11718);
nor U12578 (N_12578,N_11237,N_11573);
nand U12579 (N_12579,N_11482,N_11496);
nand U12580 (N_12580,N_11858,N_11189);
and U12581 (N_12581,N_11760,N_11169);
nor U12582 (N_12582,N_11943,N_11172);
nor U12583 (N_12583,N_11835,N_11186);
xnor U12584 (N_12584,N_11842,N_11367);
xor U12585 (N_12585,N_11508,N_11622);
xor U12586 (N_12586,N_11781,N_11334);
and U12587 (N_12587,N_11121,N_11097);
nor U12588 (N_12588,N_11922,N_11981);
nand U12589 (N_12589,N_11052,N_11162);
and U12590 (N_12590,N_11048,N_11914);
nor U12591 (N_12591,N_11636,N_11662);
nor U12592 (N_12592,N_11262,N_11125);
nor U12593 (N_12593,N_11653,N_11953);
xnor U12594 (N_12594,N_11590,N_11934);
nand U12595 (N_12595,N_11786,N_11825);
and U12596 (N_12596,N_11414,N_11107);
nand U12597 (N_12597,N_11804,N_11437);
or U12598 (N_12598,N_11571,N_11188);
nand U12599 (N_12599,N_11569,N_11045);
nor U12600 (N_12600,N_11950,N_11095);
nor U12601 (N_12601,N_11383,N_11262);
nor U12602 (N_12602,N_11726,N_11887);
and U12603 (N_12603,N_11951,N_11753);
or U12604 (N_12604,N_11932,N_11217);
or U12605 (N_12605,N_11858,N_11170);
nand U12606 (N_12606,N_11481,N_11288);
or U12607 (N_12607,N_11223,N_11886);
nand U12608 (N_12608,N_11572,N_11642);
nand U12609 (N_12609,N_11486,N_11037);
xnor U12610 (N_12610,N_11810,N_11183);
and U12611 (N_12611,N_11886,N_11305);
or U12612 (N_12612,N_11964,N_11644);
nor U12613 (N_12613,N_11166,N_11894);
and U12614 (N_12614,N_11453,N_11900);
nand U12615 (N_12615,N_11152,N_11967);
xnor U12616 (N_12616,N_11695,N_11544);
or U12617 (N_12617,N_11768,N_11698);
or U12618 (N_12618,N_11741,N_11027);
nor U12619 (N_12619,N_11577,N_11174);
xor U12620 (N_12620,N_11101,N_11469);
nand U12621 (N_12621,N_11872,N_11875);
or U12622 (N_12622,N_11169,N_11515);
and U12623 (N_12623,N_11950,N_11531);
nor U12624 (N_12624,N_11159,N_11742);
and U12625 (N_12625,N_11066,N_11811);
nand U12626 (N_12626,N_11932,N_11068);
and U12627 (N_12627,N_11641,N_11373);
xor U12628 (N_12628,N_11678,N_11709);
nor U12629 (N_12629,N_11031,N_11747);
nor U12630 (N_12630,N_11126,N_11079);
nand U12631 (N_12631,N_11012,N_11871);
and U12632 (N_12632,N_11631,N_11691);
or U12633 (N_12633,N_11204,N_11957);
nor U12634 (N_12634,N_11638,N_11034);
and U12635 (N_12635,N_11867,N_11159);
or U12636 (N_12636,N_11540,N_11000);
or U12637 (N_12637,N_11419,N_11725);
nand U12638 (N_12638,N_11179,N_11880);
xor U12639 (N_12639,N_11968,N_11561);
nor U12640 (N_12640,N_11599,N_11284);
nand U12641 (N_12641,N_11757,N_11292);
xnor U12642 (N_12642,N_11386,N_11218);
or U12643 (N_12643,N_11024,N_11696);
nor U12644 (N_12644,N_11304,N_11104);
and U12645 (N_12645,N_11469,N_11489);
nor U12646 (N_12646,N_11347,N_11964);
and U12647 (N_12647,N_11923,N_11974);
or U12648 (N_12648,N_11590,N_11814);
nor U12649 (N_12649,N_11396,N_11783);
or U12650 (N_12650,N_11471,N_11033);
nor U12651 (N_12651,N_11446,N_11555);
xnor U12652 (N_12652,N_11963,N_11188);
xor U12653 (N_12653,N_11695,N_11624);
and U12654 (N_12654,N_11655,N_11853);
or U12655 (N_12655,N_11007,N_11979);
xnor U12656 (N_12656,N_11016,N_11920);
and U12657 (N_12657,N_11154,N_11143);
and U12658 (N_12658,N_11247,N_11626);
nand U12659 (N_12659,N_11201,N_11062);
nor U12660 (N_12660,N_11146,N_11181);
or U12661 (N_12661,N_11892,N_11633);
and U12662 (N_12662,N_11950,N_11233);
or U12663 (N_12663,N_11544,N_11318);
xnor U12664 (N_12664,N_11909,N_11377);
nor U12665 (N_12665,N_11177,N_11509);
or U12666 (N_12666,N_11985,N_11396);
nor U12667 (N_12667,N_11370,N_11102);
or U12668 (N_12668,N_11333,N_11746);
nand U12669 (N_12669,N_11500,N_11050);
and U12670 (N_12670,N_11104,N_11664);
nor U12671 (N_12671,N_11136,N_11169);
nand U12672 (N_12672,N_11052,N_11299);
nor U12673 (N_12673,N_11293,N_11176);
or U12674 (N_12674,N_11731,N_11876);
xnor U12675 (N_12675,N_11640,N_11971);
nand U12676 (N_12676,N_11022,N_11786);
nand U12677 (N_12677,N_11690,N_11835);
nand U12678 (N_12678,N_11084,N_11461);
nor U12679 (N_12679,N_11618,N_11507);
and U12680 (N_12680,N_11416,N_11032);
or U12681 (N_12681,N_11905,N_11077);
nand U12682 (N_12682,N_11799,N_11067);
nor U12683 (N_12683,N_11935,N_11612);
xor U12684 (N_12684,N_11367,N_11900);
or U12685 (N_12685,N_11783,N_11717);
or U12686 (N_12686,N_11863,N_11868);
nor U12687 (N_12687,N_11676,N_11509);
nand U12688 (N_12688,N_11137,N_11467);
nand U12689 (N_12689,N_11729,N_11924);
or U12690 (N_12690,N_11870,N_11123);
nand U12691 (N_12691,N_11029,N_11568);
and U12692 (N_12692,N_11940,N_11151);
nor U12693 (N_12693,N_11115,N_11256);
nand U12694 (N_12694,N_11217,N_11644);
or U12695 (N_12695,N_11542,N_11812);
and U12696 (N_12696,N_11134,N_11214);
xor U12697 (N_12697,N_11664,N_11861);
nand U12698 (N_12698,N_11207,N_11641);
or U12699 (N_12699,N_11166,N_11072);
nand U12700 (N_12700,N_11306,N_11677);
nand U12701 (N_12701,N_11618,N_11351);
nor U12702 (N_12702,N_11720,N_11420);
nor U12703 (N_12703,N_11230,N_11141);
and U12704 (N_12704,N_11329,N_11410);
and U12705 (N_12705,N_11572,N_11503);
or U12706 (N_12706,N_11594,N_11666);
nand U12707 (N_12707,N_11968,N_11925);
and U12708 (N_12708,N_11884,N_11062);
and U12709 (N_12709,N_11458,N_11794);
xnor U12710 (N_12710,N_11986,N_11904);
xor U12711 (N_12711,N_11927,N_11475);
xor U12712 (N_12712,N_11720,N_11643);
nand U12713 (N_12713,N_11082,N_11593);
nand U12714 (N_12714,N_11414,N_11084);
nor U12715 (N_12715,N_11158,N_11798);
and U12716 (N_12716,N_11339,N_11480);
xnor U12717 (N_12717,N_11652,N_11545);
nor U12718 (N_12718,N_11238,N_11959);
nor U12719 (N_12719,N_11419,N_11749);
and U12720 (N_12720,N_11850,N_11310);
or U12721 (N_12721,N_11964,N_11796);
nand U12722 (N_12722,N_11357,N_11312);
or U12723 (N_12723,N_11297,N_11899);
nor U12724 (N_12724,N_11847,N_11532);
or U12725 (N_12725,N_11665,N_11058);
xnor U12726 (N_12726,N_11553,N_11522);
or U12727 (N_12727,N_11743,N_11561);
nor U12728 (N_12728,N_11546,N_11427);
nor U12729 (N_12729,N_11689,N_11660);
xor U12730 (N_12730,N_11689,N_11459);
or U12731 (N_12731,N_11724,N_11884);
xor U12732 (N_12732,N_11039,N_11596);
nand U12733 (N_12733,N_11557,N_11856);
nand U12734 (N_12734,N_11480,N_11776);
nor U12735 (N_12735,N_11006,N_11280);
and U12736 (N_12736,N_11531,N_11560);
and U12737 (N_12737,N_11008,N_11916);
nor U12738 (N_12738,N_11498,N_11995);
and U12739 (N_12739,N_11557,N_11124);
nand U12740 (N_12740,N_11893,N_11091);
xor U12741 (N_12741,N_11042,N_11764);
nor U12742 (N_12742,N_11686,N_11799);
nor U12743 (N_12743,N_11600,N_11470);
nand U12744 (N_12744,N_11601,N_11968);
xnor U12745 (N_12745,N_11378,N_11690);
nor U12746 (N_12746,N_11872,N_11514);
xnor U12747 (N_12747,N_11378,N_11269);
and U12748 (N_12748,N_11158,N_11170);
nor U12749 (N_12749,N_11640,N_11328);
or U12750 (N_12750,N_11816,N_11912);
or U12751 (N_12751,N_11176,N_11272);
nand U12752 (N_12752,N_11101,N_11572);
nand U12753 (N_12753,N_11770,N_11976);
nor U12754 (N_12754,N_11357,N_11957);
or U12755 (N_12755,N_11019,N_11948);
nor U12756 (N_12756,N_11765,N_11946);
nor U12757 (N_12757,N_11570,N_11359);
nand U12758 (N_12758,N_11703,N_11654);
and U12759 (N_12759,N_11152,N_11862);
nor U12760 (N_12760,N_11117,N_11018);
and U12761 (N_12761,N_11463,N_11048);
and U12762 (N_12762,N_11903,N_11701);
and U12763 (N_12763,N_11238,N_11180);
nand U12764 (N_12764,N_11338,N_11696);
nand U12765 (N_12765,N_11469,N_11860);
xnor U12766 (N_12766,N_11888,N_11571);
or U12767 (N_12767,N_11422,N_11392);
nand U12768 (N_12768,N_11960,N_11801);
or U12769 (N_12769,N_11341,N_11599);
xor U12770 (N_12770,N_11510,N_11329);
and U12771 (N_12771,N_11639,N_11380);
xnor U12772 (N_12772,N_11194,N_11976);
xnor U12773 (N_12773,N_11014,N_11274);
nand U12774 (N_12774,N_11323,N_11544);
nand U12775 (N_12775,N_11781,N_11248);
nor U12776 (N_12776,N_11436,N_11765);
nand U12777 (N_12777,N_11107,N_11157);
xnor U12778 (N_12778,N_11944,N_11827);
or U12779 (N_12779,N_11960,N_11961);
xor U12780 (N_12780,N_11933,N_11444);
and U12781 (N_12781,N_11524,N_11072);
nor U12782 (N_12782,N_11767,N_11750);
and U12783 (N_12783,N_11407,N_11672);
nand U12784 (N_12784,N_11313,N_11543);
or U12785 (N_12785,N_11447,N_11928);
xor U12786 (N_12786,N_11583,N_11686);
nand U12787 (N_12787,N_11771,N_11761);
xor U12788 (N_12788,N_11004,N_11714);
xnor U12789 (N_12789,N_11261,N_11090);
or U12790 (N_12790,N_11326,N_11396);
nor U12791 (N_12791,N_11427,N_11268);
or U12792 (N_12792,N_11791,N_11102);
or U12793 (N_12793,N_11997,N_11376);
and U12794 (N_12794,N_11932,N_11805);
nor U12795 (N_12795,N_11745,N_11907);
xor U12796 (N_12796,N_11118,N_11526);
nand U12797 (N_12797,N_11529,N_11337);
nand U12798 (N_12798,N_11708,N_11413);
or U12799 (N_12799,N_11208,N_11104);
xnor U12800 (N_12800,N_11916,N_11423);
and U12801 (N_12801,N_11329,N_11011);
nand U12802 (N_12802,N_11006,N_11847);
and U12803 (N_12803,N_11623,N_11848);
nor U12804 (N_12804,N_11285,N_11539);
nor U12805 (N_12805,N_11007,N_11207);
nand U12806 (N_12806,N_11613,N_11353);
nor U12807 (N_12807,N_11414,N_11794);
nand U12808 (N_12808,N_11049,N_11156);
and U12809 (N_12809,N_11382,N_11187);
xnor U12810 (N_12810,N_11673,N_11233);
nor U12811 (N_12811,N_11735,N_11304);
or U12812 (N_12812,N_11911,N_11330);
or U12813 (N_12813,N_11661,N_11702);
or U12814 (N_12814,N_11748,N_11488);
nand U12815 (N_12815,N_11301,N_11561);
nand U12816 (N_12816,N_11294,N_11604);
nor U12817 (N_12817,N_11667,N_11399);
or U12818 (N_12818,N_11161,N_11430);
or U12819 (N_12819,N_11379,N_11598);
nand U12820 (N_12820,N_11400,N_11824);
nand U12821 (N_12821,N_11877,N_11655);
nand U12822 (N_12822,N_11613,N_11124);
nand U12823 (N_12823,N_11226,N_11065);
or U12824 (N_12824,N_11611,N_11944);
nor U12825 (N_12825,N_11343,N_11057);
or U12826 (N_12826,N_11112,N_11079);
and U12827 (N_12827,N_11109,N_11405);
nor U12828 (N_12828,N_11170,N_11132);
xnor U12829 (N_12829,N_11928,N_11515);
nand U12830 (N_12830,N_11784,N_11630);
or U12831 (N_12831,N_11684,N_11228);
xor U12832 (N_12832,N_11110,N_11359);
xor U12833 (N_12833,N_11090,N_11181);
xnor U12834 (N_12834,N_11783,N_11937);
xnor U12835 (N_12835,N_11071,N_11643);
nand U12836 (N_12836,N_11833,N_11991);
and U12837 (N_12837,N_11493,N_11162);
nor U12838 (N_12838,N_11189,N_11068);
nand U12839 (N_12839,N_11932,N_11006);
xnor U12840 (N_12840,N_11242,N_11582);
and U12841 (N_12841,N_11215,N_11370);
xor U12842 (N_12842,N_11685,N_11664);
nor U12843 (N_12843,N_11151,N_11709);
and U12844 (N_12844,N_11847,N_11698);
or U12845 (N_12845,N_11082,N_11753);
and U12846 (N_12846,N_11135,N_11220);
xnor U12847 (N_12847,N_11915,N_11001);
xor U12848 (N_12848,N_11015,N_11528);
nor U12849 (N_12849,N_11788,N_11046);
or U12850 (N_12850,N_11398,N_11667);
or U12851 (N_12851,N_11959,N_11244);
xnor U12852 (N_12852,N_11410,N_11435);
nand U12853 (N_12853,N_11447,N_11578);
and U12854 (N_12854,N_11862,N_11215);
nor U12855 (N_12855,N_11465,N_11321);
nand U12856 (N_12856,N_11621,N_11302);
nand U12857 (N_12857,N_11835,N_11428);
nand U12858 (N_12858,N_11967,N_11923);
or U12859 (N_12859,N_11230,N_11418);
nor U12860 (N_12860,N_11587,N_11395);
or U12861 (N_12861,N_11407,N_11669);
nor U12862 (N_12862,N_11263,N_11285);
and U12863 (N_12863,N_11331,N_11696);
nor U12864 (N_12864,N_11631,N_11710);
nor U12865 (N_12865,N_11755,N_11359);
nor U12866 (N_12866,N_11397,N_11554);
and U12867 (N_12867,N_11801,N_11895);
nor U12868 (N_12868,N_11290,N_11149);
or U12869 (N_12869,N_11977,N_11119);
xor U12870 (N_12870,N_11212,N_11749);
or U12871 (N_12871,N_11605,N_11847);
nor U12872 (N_12872,N_11989,N_11677);
and U12873 (N_12873,N_11708,N_11182);
nand U12874 (N_12874,N_11714,N_11580);
or U12875 (N_12875,N_11640,N_11291);
nand U12876 (N_12876,N_11498,N_11034);
or U12877 (N_12877,N_11410,N_11056);
nor U12878 (N_12878,N_11010,N_11648);
nor U12879 (N_12879,N_11384,N_11744);
and U12880 (N_12880,N_11606,N_11971);
or U12881 (N_12881,N_11536,N_11107);
xnor U12882 (N_12882,N_11841,N_11414);
and U12883 (N_12883,N_11483,N_11753);
and U12884 (N_12884,N_11914,N_11688);
and U12885 (N_12885,N_11698,N_11719);
or U12886 (N_12886,N_11636,N_11279);
and U12887 (N_12887,N_11185,N_11203);
nand U12888 (N_12888,N_11284,N_11301);
or U12889 (N_12889,N_11783,N_11220);
nand U12890 (N_12890,N_11702,N_11682);
and U12891 (N_12891,N_11569,N_11525);
and U12892 (N_12892,N_11026,N_11915);
nand U12893 (N_12893,N_11861,N_11989);
nand U12894 (N_12894,N_11694,N_11748);
nor U12895 (N_12895,N_11679,N_11563);
nor U12896 (N_12896,N_11536,N_11210);
nand U12897 (N_12897,N_11004,N_11035);
nand U12898 (N_12898,N_11152,N_11650);
and U12899 (N_12899,N_11625,N_11905);
xor U12900 (N_12900,N_11286,N_11555);
nor U12901 (N_12901,N_11180,N_11390);
or U12902 (N_12902,N_11352,N_11426);
nor U12903 (N_12903,N_11617,N_11518);
nor U12904 (N_12904,N_11539,N_11617);
nor U12905 (N_12905,N_11865,N_11711);
nand U12906 (N_12906,N_11481,N_11623);
nor U12907 (N_12907,N_11127,N_11298);
nand U12908 (N_12908,N_11029,N_11208);
xor U12909 (N_12909,N_11714,N_11431);
and U12910 (N_12910,N_11031,N_11867);
xor U12911 (N_12911,N_11812,N_11249);
or U12912 (N_12912,N_11321,N_11874);
and U12913 (N_12913,N_11137,N_11373);
or U12914 (N_12914,N_11569,N_11532);
and U12915 (N_12915,N_11992,N_11993);
xor U12916 (N_12916,N_11437,N_11473);
nand U12917 (N_12917,N_11827,N_11368);
or U12918 (N_12918,N_11591,N_11933);
and U12919 (N_12919,N_11871,N_11787);
or U12920 (N_12920,N_11124,N_11711);
nand U12921 (N_12921,N_11460,N_11391);
or U12922 (N_12922,N_11868,N_11653);
xnor U12923 (N_12923,N_11006,N_11693);
and U12924 (N_12924,N_11948,N_11656);
nand U12925 (N_12925,N_11303,N_11661);
or U12926 (N_12926,N_11122,N_11800);
and U12927 (N_12927,N_11342,N_11510);
xor U12928 (N_12928,N_11937,N_11681);
xor U12929 (N_12929,N_11200,N_11872);
xnor U12930 (N_12930,N_11161,N_11946);
or U12931 (N_12931,N_11560,N_11592);
xnor U12932 (N_12932,N_11029,N_11233);
xnor U12933 (N_12933,N_11649,N_11029);
and U12934 (N_12934,N_11526,N_11244);
nor U12935 (N_12935,N_11553,N_11695);
and U12936 (N_12936,N_11399,N_11282);
nand U12937 (N_12937,N_11686,N_11684);
nor U12938 (N_12938,N_11594,N_11565);
and U12939 (N_12939,N_11540,N_11829);
and U12940 (N_12940,N_11065,N_11911);
and U12941 (N_12941,N_11523,N_11846);
or U12942 (N_12942,N_11577,N_11958);
or U12943 (N_12943,N_11608,N_11727);
nand U12944 (N_12944,N_11340,N_11668);
nor U12945 (N_12945,N_11484,N_11887);
nor U12946 (N_12946,N_11348,N_11414);
nand U12947 (N_12947,N_11613,N_11992);
and U12948 (N_12948,N_11559,N_11838);
and U12949 (N_12949,N_11460,N_11636);
xnor U12950 (N_12950,N_11352,N_11878);
nand U12951 (N_12951,N_11720,N_11116);
xor U12952 (N_12952,N_11715,N_11103);
nand U12953 (N_12953,N_11254,N_11607);
and U12954 (N_12954,N_11302,N_11971);
xor U12955 (N_12955,N_11894,N_11791);
nand U12956 (N_12956,N_11990,N_11156);
xnor U12957 (N_12957,N_11733,N_11873);
or U12958 (N_12958,N_11413,N_11749);
and U12959 (N_12959,N_11614,N_11912);
xor U12960 (N_12960,N_11220,N_11855);
nor U12961 (N_12961,N_11483,N_11578);
nand U12962 (N_12962,N_11020,N_11696);
nand U12963 (N_12963,N_11737,N_11603);
and U12964 (N_12964,N_11933,N_11906);
and U12965 (N_12965,N_11371,N_11179);
nor U12966 (N_12966,N_11967,N_11783);
or U12967 (N_12967,N_11021,N_11175);
nor U12968 (N_12968,N_11343,N_11840);
nand U12969 (N_12969,N_11306,N_11085);
nor U12970 (N_12970,N_11242,N_11576);
nand U12971 (N_12971,N_11358,N_11319);
xor U12972 (N_12972,N_11945,N_11530);
xor U12973 (N_12973,N_11019,N_11096);
nand U12974 (N_12974,N_11070,N_11900);
or U12975 (N_12975,N_11224,N_11591);
nor U12976 (N_12976,N_11176,N_11786);
or U12977 (N_12977,N_11823,N_11873);
or U12978 (N_12978,N_11140,N_11473);
xor U12979 (N_12979,N_11293,N_11797);
xnor U12980 (N_12980,N_11546,N_11215);
and U12981 (N_12981,N_11522,N_11029);
nor U12982 (N_12982,N_11643,N_11494);
nor U12983 (N_12983,N_11215,N_11384);
nor U12984 (N_12984,N_11715,N_11473);
xnor U12985 (N_12985,N_11147,N_11943);
and U12986 (N_12986,N_11927,N_11108);
nand U12987 (N_12987,N_11994,N_11388);
or U12988 (N_12988,N_11434,N_11533);
nor U12989 (N_12989,N_11281,N_11465);
or U12990 (N_12990,N_11178,N_11331);
and U12991 (N_12991,N_11408,N_11851);
nand U12992 (N_12992,N_11295,N_11177);
nor U12993 (N_12993,N_11000,N_11400);
or U12994 (N_12994,N_11941,N_11644);
and U12995 (N_12995,N_11164,N_11627);
nor U12996 (N_12996,N_11117,N_11360);
or U12997 (N_12997,N_11231,N_11238);
and U12998 (N_12998,N_11161,N_11391);
or U12999 (N_12999,N_11498,N_11701);
and U13000 (N_13000,N_12612,N_12794);
and U13001 (N_13001,N_12046,N_12781);
or U13002 (N_13002,N_12658,N_12739);
and U13003 (N_13003,N_12134,N_12171);
nand U13004 (N_13004,N_12244,N_12942);
nor U13005 (N_13005,N_12194,N_12135);
or U13006 (N_13006,N_12029,N_12514);
and U13007 (N_13007,N_12214,N_12912);
xor U13008 (N_13008,N_12614,N_12483);
nor U13009 (N_13009,N_12074,N_12523);
nand U13010 (N_13010,N_12537,N_12247);
and U13011 (N_13011,N_12209,N_12526);
and U13012 (N_13012,N_12619,N_12329);
and U13013 (N_13013,N_12894,N_12227);
and U13014 (N_13014,N_12200,N_12850);
and U13015 (N_13015,N_12138,N_12585);
xnor U13016 (N_13016,N_12718,N_12191);
nand U13017 (N_13017,N_12271,N_12178);
or U13018 (N_13018,N_12277,N_12536);
xor U13019 (N_13019,N_12871,N_12263);
nor U13020 (N_13020,N_12385,N_12500);
nand U13021 (N_13021,N_12701,N_12913);
xor U13022 (N_13022,N_12463,N_12006);
xor U13023 (N_13023,N_12266,N_12529);
xor U13024 (N_13024,N_12787,N_12800);
and U13025 (N_13025,N_12089,N_12717);
or U13026 (N_13026,N_12635,N_12569);
or U13027 (N_13027,N_12328,N_12431);
nand U13028 (N_13028,N_12659,N_12726);
xor U13029 (N_13029,N_12653,N_12770);
and U13030 (N_13030,N_12498,N_12370);
and U13031 (N_13031,N_12306,N_12068);
nor U13032 (N_13032,N_12174,N_12744);
nor U13033 (N_13033,N_12170,N_12272);
or U13034 (N_13034,N_12371,N_12967);
nand U13035 (N_13035,N_12608,N_12821);
and U13036 (N_13036,N_12949,N_12369);
nand U13037 (N_13037,N_12003,N_12777);
nor U13038 (N_13038,N_12384,N_12027);
or U13039 (N_13039,N_12310,N_12522);
or U13040 (N_13040,N_12268,N_12859);
xor U13041 (N_13041,N_12146,N_12270);
nor U13042 (N_13042,N_12565,N_12091);
xor U13043 (N_13043,N_12964,N_12039);
or U13044 (N_13044,N_12466,N_12703);
xor U13045 (N_13045,N_12974,N_12293);
and U13046 (N_13046,N_12583,N_12274);
nand U13047 (N_13047,N_12737,N_12419);
nor U13048 (N_13048,N_12734,N_12405);
nand U13049 (N_13049,N_12389,N_12710);
nand U13050 (N_13050,N_12780,N_12324);
nor U13051 (N_13051,N_12275,N_12305);
or U13052 (N_13052,N_12854,N_12362);
and U13053 (N_13053,N_12096,N_12455);
and U13054 (N_13054,N_12929,N_12311);
and U13055 (N_13055,N_12107,N_12941);
and U13056 (N_13056,N_12136,N_12695);
xnor U13057 (N_13057,N_12985,N_12784);
xor U13058 (N_13058,N_12296,N_12323);
or U13059 (N_13059,N_12811,N_12933);
nor U13060 (N_13060,N_12021,N_12763);
or U13061 (N_13061,N_12613,N_12637);
nand U13062 (N_13062,N_12864,N_12480);
nand U13063 (N_13063,N_12149,N_12461);
or U13064 (N_13064,N_12636,N_12281);
or U13065 (N_13065,N_12278,N_12414);
xor U13066 (N_13066,N_12183,N_12674);
xnor U13067 (N_13067,N_12652,N_12707);
or U13068 (N_13068,N_12660,N_12810);
or U13069 (N_13069,N_12218,N_12140);
or U13070 (N_13070,N_12818,N_12587);
nor U13071 (N_13071,N_12666,N_12350);
xor U13072 (N_13072,N_12258,N_12240);
nor U13073 (N_13073,N_12690,N_12378);
and U13074 (N_13074,N_12457,N_12779);
nor U13075 (N_13075,N_12148,N_12650);
nand U13076 (N_13076,N_12026,N_12465);
nor U13077 (N_13077,N_12827,N_12020);
and U13078 (N_13078,N_12417,N_12482);
nor U13079 (N_13079,N_12077,N_12769);
xor U13080 (N_13080,N_12166,N_12221);
xor U13081 (N_13081,N_12101,N_12682);
nand U13082 (N_13082,N_12072,N_12114);
or U13083 (N_13083,N_12544,N_12713);
nand U13084 (N_13084,N_12848,N_12520);
and U13085 (N_13085,N_12472,N_12868);
or U13086 (N_13086,N_12729,N_12145);
nor U13087 (N_13087,N_12577,N_12447);
nand U13088 (N_13088,N_12299,N_12959);
xor U13089 (N_13089,N_12716,N_12471);
nor U13090 (N_13090,N_12394,N_12357);
or U13091 (N_13091,N_12156,N_12111);
nand U13092 (N_13092,N_12604,N_12273);
or U13093 (N_13093,N_12979,N_12719);
and U13094 (N_13094,N_12343,N_12103);
nand U13095 (N_13095,N_12031,N_12368);
xnor U13096 (N_13096,N_12037,N_12056);
or U13097 (N_13097,N_12566,N_12207);
nand U13098 (N_13098,N_12118,N_12025);
nor U13099 (N_13099,N_12934,N_12918);
and U13100 (N_13100,N_12524,N_12548);
or U13101 (N_13101,N_12632,N_12115);
xor U13102 (N_13102,N_12998,N_12986);
or U13103 (N_13103,N_12880,N_12930);
xor U13104 (N_13104,N_12295,N_12206);
nand U13105 (N_13105,N_12449,N_12014);
xor U13106 (N_13106,N_12494,N_12391);
nor U13107 (N_13107,N_12411,N_12185);
or U13108 (N_13108,N_12751,N_12815);
nand U13109 (N_13109,N_12857,N_12560);
or U13110 (N_13110,N_12944,N_12947);
xnor U13111 (N_13111,N_12144,N_12884);
nor U13112 (N_13112,N_12164,N_12162);
or U13113 (N_13113,N_12973,N_12844);
or U13114 (N_13114,N_12152,N_12557);
and U13115 (N_13115,N_12890,N_12573);
nor U13116 (N_13116,N_12412,N_12182);
nor U13117 (N_13117,N_12983,N_12914);
and U13118 (N_13118,N_12158,N_12749);
and U13119 (N_13119,N_12640,N_12741);
nand U13120 (N_13120,N_12106,N_12697);
and U13121 (N_13121,N_12187,N_12664);
xor U13122 (N_13122,N_12732,N_12831);
nand U13123 (N_13123,N_12216,N_12351);
xor U13124 (N_13124,N_12346,N_12012);
or U13125 (N_13125,N_12321,N_12642);
and U13126 (N_13126,N_12528,N_12755);
nor U13127 (N_13127,N_12793,N_12117);
nor U13128 (N_13128,N_12377,N_12013);
nor U13129 (N_13129,N_12269,N_12338);
nand U13130 (N_13130,N_12341,N_12198);
xnor U13131 (N_13131,N_12990,N_12669);
xor U13132 (N_13132,N_12104,N_12330);
nor U13133 (N_13133,N_12237,N_12497);
or U13134 (N_13134,N_12313,N_12609);
and U13135 (N_13135,N_12980,N_12843);
xor U13136 (N_13136,N_12139,N_12845);
or U13137 (N_13137,N_12647,N_12839);
nor U13138 (N_13138,N_12153,N_12462);
or U13139 (N_13139,N_12775,N_12910);
or U13140 (N_13140,N_12518,N_12813);
xor U13141 (N_13141,N_12379,N_12995);
xnor U13142 (N_13142,N_12167,N_12623);
or U13143 (N_13143,N_12846,N_12870);
nand U13144 (N_13144,N_12927,N_12533);
and U13145 (N_13145,N_12488,N_12802);
nand U13146 (N_13146,N_12965,N_12987);
or U13147 (N_13147,N_12154,N_12331);
xnor U13148 (N_13148,N_12130,N_12893);
and U13149 (N_13149,N_12503,N_12889);
nand U13150 (N_13150,N_12543,N_12515);
and U13151 (N_13151,N_12199,N_12226);
and U13152 (N_13152,N_12219,N_12475);
nor U13153 (N_13153,N_12600,N_12155);
xor U13154 (N_13154,N_12337,N_12646);
and U13155 (N_13155,N_12236,N_12094);
nor U13156 (N_13156,N_12175,N_12806);
nor U13157 (N_13157,N_12651,N_12478);
or U13158 (N_13158,N_12061,N_12804);
nand U13159 (N_13159,N_12381,N_12519);
xnor U13160 (N_13160,N_12142,N_12945);
xnor U13161 (N_13161,N_12648,N_12508);
nor U13162 (N_13162,N_12049,N_12450);
nand U13163 (N_13163,N_12348,N_12264);
and U13164 (N_13164,N_12616,N_12628);
and U13165 (N_13165,N_12017,N_12100);
nor U13166 (N_13166,N_12655,N_12452);
nor U13167 (N_13167,N_12938,N_12639);
or U13168 (N_13168,N_12479,N_12882);
and U13169 (N_13169,N_12773,N_12742);
or U13170 (N_13170,N_12502,N_12113);
and U13171 (N_13171,N_12112,N_12238);
xor U13172 (N_13172,N_12774,N_12783);
nor U13173 (N_13173,N_12066,N_12435);
nor U13174 (N_13174,N_12950,N_12936);
or U13175 (N_13175,N_12960,N_12079);
xor U13176 (N_13176,N_12122,N_12801);
xnor U13177 (N_13177,N_12924,N_12043);
or U13178 (N_13178,N_12454,N_12956);
nor U13179 (N_13179,N_12451,N_12421);
xor U13180 (N_13180,N_12997,N_12428);
or U13181 (N_13181,N_12002,N_12290);
and U13182 (N_13182,N_12649,N_12785);
nor U13183 (N_13183,N_12978,N_12951);
or U13184 (N_13184,N_12193,N_12847);
or U13185 (N_13185,N_12426,N_12404);
nor U13186 (N_13186,N_12285,N_12434);
or U13187 (N_13187,N_12493,N_12119);
or U13188 (N_13188,N_12799,N_12048);
or U13189 (N_13189,N_12791,N_12090);
and U13190 (N_13190,N_12926,N_12991);
or U13191 (N_13191,N_12253,N_12359);
nand U13192 (N_13192,N_12468,N_12334);
nor U13193 (N_13193,N_12764,N_12618);
nand U13194 (N_13194,N_12407,N_12504);
xnor U13195 (N_13195,N_12261,N_12665);
or U13196 (N_13196,N_12023,N_12456);
or U13197 (N_13197,N_12688,N_12365);
or U13198 (N_13198,N_12833,N_12254);
or U13199 (N_13199,N_12474,N_12747);
nand U13200 (N_13200,N_12970,N_12790);
nor U13201 (N_13201,N_12062,N_12469);
nand U13202 (N_13202,N_12491,N_12406);
or U13203 (N_13203,N_12120,N_12436);
and U13204 (N_13204,N_12420,N_12988);
xnor U13205 (N_13205,N_12050,N_12761);
and U13206 (N_13206,N_12069,N_12555);
and U13207 (N_13207,N_12593,N_12205);
and U13208 (N_13208,N_12186,N_12035);
nand U13209 (N_13209,N_12901,N_12953);
and U13210 (N_13210,N_12506,N_12176);
and U13211 (N_13211,N_12302,N_12672);
nand U13212 (N_13212,N_12399,N_12374);
and U13213 (N_13213,N_12731,N_12627);
or U13214 (N_13214,N_12766,N_12347);
xnor U13215 (N_13215,N_12704,N_12257);
and U13216 (N_13216,N_12364,N_12789);
and U13217 (N_13217,N_12634,N_12692);
xor U13218 (N_13218,N_12076,N_12571);
or U13219 (N_13219,N_12395,N_12505);
nand U13220 (N_13220,N_12702,N_12550);
nand U13221 (N_13221,N_12771,N_12955);
nor U13222 (N_13222,N_12099,N_12418);
and U13223 (N_13223,N_12925,N_12181);
nor U13224 (N_13224,N_12909,N_12235);
or U13225 (N_13225,N_12931,N_12098);
nand U13226 (N_13226,N_12291,N_12856);
or U13227 (N_13227,N_12460,N_12935);
nand U13228 (N_13228,N_12429,N_12869);
nor U13229 (N_13229,N_12805,N_12001);
and U13230 (N_13230,N_12629,N_12082);
and U13231 (N_13231,N_12570,N_12724);
nand U13232 (N_13232,N_12999,N_12231);
nand U13233 (N_13233,N_12401,N_12052);
or U13234 (N_13234,N_12150,N_12714);
and U13235 (N_13235,N_12375,N_12427);
or U13236 (N_13236,N_12835,N_12823);
xnor U13237 (N_13237,N_12904,N_12678);
or U13238 (N_13238,N_12592,N_12723);
or U13239 (N_13239,N_12685,N_12891);
nand U13240 (N_13240,N_12750,N_12617);
nand U13241 (N_13241,N_12445,N_12877);
or U13242 (N_13242,N_12189,N_12487);
and U13243 (N_13243,N_12303,N_12591);
nor U13244 (N_13244,N_12495,N_12558);
and U13245 (N_13245,N_12834,N_12301);
xor U13246 (N_13246,N_12849,N_12165);
and U13247 (N_13247,N_12033,N_12952);
nand U13248 (N_13248,N_12215,N_12403);
xor U13249 (N_13249,N_12760,N_12307);
xnor U13250 (N_13250,N_12832,N_12622);
nor U13251 (N_13251,N_12108,N_12073);
xor U13252 (N_13252,N_12318,N_12443);
nor U13253 (N_13253,N_12579,N_12898);
xor U13254 (N_13254,N_12694,N_12851);
xnor U13255 (N_13255,N_12501,N_12525);
or U13256 (N_13256,N_12825,N_12735);
nor U13257 (N_13257,N_12093,N_12123);
and U13258 (N_13258,N_12453,N_12792);
nor U13259 (N_13259,N_12396,N_12433);
and U13260 (N_13260,N_12382,N_12442);
and U13261 (N_13261,N_12315,N_12841);
nor U13262 (N_13262,N_12595,N_12897);
and U13263 (N_13263,N_12996,N_12464);
or U13264 (N_13264,N_12946,N_12060);
and U13265 (N_13265,N_12673,N_12551);
nor U13266 (N_13266,N_12542,N_12065);
and U13267 (N_13267,N_12173,N_12366);
and U13268 (N_13268,N_12441,N_12332);
nor U13269 (N_13269,N_12409,N_12392);
and U13270 (N_13270,N_12981,N_12083);
and U13271 (N_13271,N_12220,N_12905);
or U13272 (N_13272,N_12509,N_12668);
or U13273 (N_13273,N_12872,N_12289);
or U13274 (N_13274,N_12085,N_12473);
and U13275 (N_13275,N_12657,N_12110);
nand U13276 (N_13276,N_12078,N_12222);
xor U13277 (N_13277,N_12019,N_12584);
nor U13278 (N_13278,N_12034,N_12630);
or U13279 (N_13279,N_12080,N_12179);
or U13280 (N_13280,N_12184,N_12853);
nand U13281 (N_13281,N_12758,N_12943);
or U13282 (N_13282,N_12733,N_12873);
nor U13283 (N_13283,N_12625,N_12432);
or U13284 (N_13284,N_12772,N_12992);
xnor U13285 (N_13285,N_12876,N_12410);
nor U13286 (N_13286,N_12481,N_12684);
nand U13287 (N_13287,N_12349,N_12765);
xnor U13288 (N_13288,N_12830,N_12875);
and U13289 (N_13289,N_12358,N_12249);
or U13290 (N_13290,N_12022,N_12024);
nand U13291 (N_13291,N_12000,N_12248);
nand U13292 (N_13292,N_12816,N_12517);
nand U13293 (N_13293,N_12662,N_12393);
nor U13294 (N_13294,N_12958,N_12663);
nor U13295 (N_13295,N_12994,N_12097);
nand U13296 (N_13296,N_12607,N_12372);
or U13297 (N_13297,N_12416,N_12015);
or U13298 (N_13298,N_12881,N_12448);
and U13299 (N_13299,N_12803,N_12671);
xor U13300 (N_13300,N_12667,N_12298);
nand U13301 (N_13301,N_12745,N_12581);
and U13302 (N_13302,N_12109,N_12390);
and U13303 (N_13303,N_12786,N_12353);
nand U13304 (N_13304,N_12210,N_12018);
and U13305 (N_13305,N_12855,N_12458);
or U13306 (N_13306,N_12212,N_12265);
nor U13307 (N_13307,N_12499,N_12916);
xnor U13308 (N_13308,N_12197,N_12243);
and U13309 (N_13309,N_12195,N_12645);
nor U13310 (N_13310,N_12317,N_12711);
nor U13311 (N_13311,N_12388,N_12288);
and U13312 (N_13312,N_12531,N_12356);
nand U13313 (N_13313,N_12796,N_12892);
nor U13314 (N_13314,N_12131,N_12300);
nand U13315 (N_13315,N_12127,N_12975);
nand U13316 (N_13316,N_12010,N_12438);
xnor U13317 (N_13317,N_12923,N_12233);
or U13318 (N_13318,N_12527,N_12538);
and U13319 (N_13319,N_12586,N_12921);
nand U13320 (N_13320,N_12177,N_12865);
or U13321 (N_13321,N_12188,N_12699);
nand U13322 (N_13322,N_12057,N_12255);
nor U13323 (N_13323,N_12599,N_12602);
xnor U13324 (N_13324,N_12788,N_12621);
and U13325 (N_13325,N_12720,N_12376);
xor U13326 (N_13326,N_12256,N_12087);
and U13327 (N_13327,N_12070,N_12322);
or U13328 (N_13328,N_12413,N_12541);
nor U13329 (N_13329,N_12437,N_12888);
and U13330 (N_13330,N_12814,N_12638);
nor U13331 (N_13331,N_12759,N_12670);
xor U13332 (N_13332,N_12721,N_12521);
and U13333 (N_13333,N_12232,N_12032);
nor U13334 (N_13334,N_12116,N_12962);
and U13335 (N_13335,N_12982,N_12675);
xnor U13336 (N_13336,N_12485,N_12677);
or U13337 (N_13337,N_12568,N_12081);
or U13338 (N_13338,N_12819,N_12556);
and U13339 (N_13339,N_12304,N_12597);
or U13340 (N_13340,N_12211,N_12213);
xnor U13341 (N_13341,N_12168,N_12284);
nor U13342 (N_13342,N_12005,N_12467);
and U13343 (N_13343,N_12224,N_12895);
nor U13344 (N_13344,N_12105,N_12228);
or U13345 (N_13345,N_12809,N_12192);
and U13346 (N_13346,N_12267,N_12530);
nor U13347 (N_13347,N_12147,N_12423);
nor U13348 (N_13348,N_12251,N_12545);
xnor U13349 (N_13349,N_12693,N_12425);
or U13350 (N_13350,N_12656,N_12715);
xnor U13351 (N_13351,N_12063,N_12157);
or U13352 (N_13352,N_12092,N_12899);
xnor U13353 (N_13353,N_12601,N_12736);
nand U13354 (N_13354,N_12676,N_12004);
and U13355 (N_13355,N_12594,N_12489);
nand U13356 (N_13356,N_12752,N_12915);
nor U13357 (N_13357,N_12163,N_12308);
nor U13358 (N_13358,N_12572,N_12939);
nand U13359 (N_13359,N_12143,N_12589);
and U13360 (N_13360,N_12795,N_12230);
nor U13361 (N_13361,N_12225,N_12342);
nand U13362 (N_13362,N_12217,N_12606);
xnor U13363 (N_13363,N_12008,N_12680);
and U13364 (N_13364,N_12314,N_12040);
nand U13365 (N_13365,N_12180,N_12798);
xor U13366 (N_13366,N_12561,N_12826);
nand U13367 (N_13367,N_12234,N_12239);
xnor U13368 (N_13368,N_12762,N_12748);
nand U13369 (N_13369,N_12137,N_12753);
xor U13370 (N_13370,N_12546,N_12743);
nor U13371 (N_13371,N_12972,N_12709);
nor U13372 (N_13372,N_12397,N_12576);
xnor U13373 (N_13373,N_12160,N_12387);
nand U13374 (N_13374,N_12047,N_12380);
nand U13375 (N_13375,N_12863,N_12575);
xor U13376 (N_13376,N_12887,N_12287);
and U13377 (N_13377,N_12722,N_12700);
nor U13378 (N_13378,N_12540,N_12917);
xor U13379 (N_13379,N_12820,N_12902);
and U13380 (N_13380,N_12698,N_12446);
xnor U13381 (N_13381,N_12088,N_12730);
xnor U13382 (N_13382,N_12837,N_12776);
xnor U13383 (N_13383,N_12534,N_12202);
nand U13384 (N_13384,N_12125,N_12971);
nand U13385 (N_13385,N_12768,N_12133);
and U13386 (N_13386,N_12679,N_12580);
nand U13387 (N_13387,N_12141,N_12564);
nand U13388 (N_13388,N_12169,N_12554);
and U13389 (N_13389,N_12030,N_12932);
nor U13390 (N_13390,N_12282,N_12363);
xnor U13391 (N_13391,N_12102,N_12828);
nand U13392 (N_13392,N_12782,N_12861);
xor U13393 (N_13393,N_12908,N_12578);
and U13394 (N_13394,N_12883,N_12242);
nor U13395 (N_13395,N_12906,N_12756);
nand U13396 (N_13396,N_12151,N_12687);
and U13397 (N_13397,N_12874,N_12223);
or U13398 (N_13398,N_12757,N_12492);
nor U13399 (N_13399,N_12879,N_12620);
xnor U13400 (N_13400,N_12354,N_12740);
or U13401 (N_13401,N_12340,N_12615);
or U13402 (N_13402,N_12574,N_12294);
or U13403 (N_13403,N_12822,N_12512);
or U13404 (N_13404,N_12262,N_12535);
or U13405 (N_13405,N_12797,N_12778);
nor U13406 (N_13406,N_12496,N_12172);
or U13407 (N_13407,N_12706,N_12402);
nor U13408 (N_13408,N_12327,N_12204);
and U13409 (N_13409,N_12903,N_12028);
nor U13410 (N_13410,N_12336,N_12963);
or U13411 (N_13411,N_12510,N_12132);
nand U13412 (N_13412,N_12058,N_12400);
nor U13413 (N_13413,N_12631,N_12124);
xor U13414 (N_13414,N_12201,N_12922);
xnor U13415 (N_13415,N_12053,N_12245);
or U13416 (N_13416,N_12611,N_12320);
and U13417 (N_13417,N_12588,N_12989);
or U13418 (N_13418,N_12633,N_12563);
xnor U13419 (N_13419,N_12836,N_12807);
or U13420 (N_13420,N_12440,N_12038);
nor U13421 (N_13421,N_12360,N_12691);
and U13422 (N_13422,N_12309,N_12860);
or U13423 (N_13423,N_12486,N_12071);
and U13424 (N_13424,N_12610,N_12075);
xnor U13425 (N_13425,N_12516,N_12067);
and U13426 (N_13426,N_12948,N_12954);
or U13427 (N_13427,N_12367,N_12297);
or U13428 (N_13428,N_12292,N_12817);
nand U13429 (N_13429,N_12016,N_12490);
nor U13430 (N_13430,N_12712,N_12654);
nand U13431 (N_13431,N_12754,N_12373);
xor U13432 (N_13432,N_12009,N_12036);
or U13433 (N_13433,N_12598,N_12624);
xor U13434 (N_13434,N_12626,N_12582);
xnor U13435 (N_13435,N_12829,N_12727);
xor U13436 (N_13436,N_12279,N_12911);
and U13437 (N_13437,N_12852,N_12246);
xnor U13438 (N_13438,N_12547,N_12562);
and U13439 (N_13439,N_12681,N_12661);
nand U13440 (N_13440,N_12689,N_12129);
nand U13441 (N_13441,N_12444,N_12976);
xor U13442 (N_13442,N_12919,N_12885);
and U13443 (N_13443,N_12352,N_12746);
nand U13444 (N_13444,N_12686,N_12567);
xnor U13445 (N_13445,N_12644,N_12126);
and U13446 (N_13446,N_12408,N_12511);
or U13447 (N_13447,N_12459,N_12812);
xor U13448 (N_13448,N_12283,N_12422);
nor U13449 (N_13449,N_12896,N_12552);
and U13450 (N_13450,N_12961,N_12862);
or U13451 (N_13451,N_12241,N_12045);
or U13452 (N_13452,N_12484,N_12229);
nor U13453 (N_13453,N_12333,N_12866);
nor U13454 (N_13454,N_12044,N_12886);
nor U13455 (N_13455,N_12280,N_12312);
or U13456 (N_13456,N_12559,N_12507);
nor U13457 (N_13457,N_12824,N_12250);
or U13458 (N_13458,N_12276,N_12683);
nor U13459 (N_13459,N_12738,N_12553);
nor U13460 (N_13460,N_12054,N_12326);
and U13461 (N_13461,N_12977,N_12470);
nand U13462 (N_13462,N_12252,N_12641);
or U13463 (N_13463,N_12042,N_12513);
and U13464 (N_13464,N_12386,N_12878);
nand U13465 (N_13465,N_12984,N_12842);
and U13466 (N_13466,N_12059,N_12208);
or U13467 (N_13467,N_12957,N_12011);
or U13468 (N_13468,N_12259,N_12603);
nor U13469 (N_13469,N_12708,N_12605);
or U13470 (N_13470,N_12725,N_12383);
or U13471 (N_13471,N_12590,N_12190);
nand U13472 (N_13472,N_12705,N_12339);
xor U13473 (N_13473,N_12361,N_12064);
or U13474 (N_13474,N_12316,N_12335);
nand U13475 (N_13475,N_12532,N_12430);
and U13476 (N_13476,N_12907,N_12398);
or U13477 (N_13477,N_12344,N_12415);
nand U13478 (N_13478,N_12937,N_12767);
xnor U13479 (N_13479,N_12808,N_12286);
and U13480 (N_13480,N_12051,N_12439);
nor U13481 (N_13481,N_12007,N_12095);
and U13482 (N_13482,N_12161,N_12968);
or U13483 (N_13483,N_12728,N_12838);
xnor U13484 (N_13484,N_12055,N_12596);
and U13485 (N_13485,N_12920,N_12858);
and U13486 (N_13486,N_12424,N_12121);
or U13487 (N_13487,N_12928,N_12993);
and U13488 (N_13488,N_12900,N_12966);
or U13489 (N_13489,N_12196,N_12940);
or U13490 (N_13490,N_12696,N_12345);
nor U13491 (N_13491,N_12476,N_12867);
and U13492 (N_13492,N_12477,N_12086);
nor U13493 (N_13493,N_12643,N_12840);
xor U13494 (N_13494,N_12355,N_12084);
nand U13495 (N_13495,N_12325,N_12128);
or U13496 (N_13496,N_12319,N_12041);
nand U13497 (N_13497,N_12260,N_12159);
nand U13498 (N_13498,N_12549,N_12539);
or U13499 (N_13499,N_12969,N_12203);
nor U13500 (N_13500,N_12653,N_12260);
xor U13501 (N_13501,N_12237,N_12731);
or U13502 (N_13502,N_12658,N_12527);
xor U13503 (N_13503,N_12207,N_12336);
nand U13504 (N_13504,N_12016,N_12195);
and U13505 (N_13505,N_12102,N_12384);
xor U13506 (N_13506,N_12990,N_12020);
or U13507 (N_13507,N_12699,N_12298);
or U13508 (N_13508,N_12843,N_12699);
and U13509 (N_13509,N_12263,N_12225);
and U13510 (N_13510,N_12277,N_12713);
or U13511 (N_13511,N_12465,N_12291);
nand U13512 (N_13512,N_12140,N_12913);
nor U13513 (N_13513,N_12106,N_12827);
xnor U13514 (N_13514,N_12263,N_12365);
or U13515 (N_13515,N_12697,N_12098);
xor U13516 (N_13516,N_12624,N_12883);
nand U13517 (N_13517,N_12399,N_12251);
or U13518 (N_13518,N_12488,N_12872);
nor U13519 (N_13519,N_12996,N_12901);
or U13520 (N_13520,N_12387,N_12388);
and U13521 (N_13521,N_12271,N_12839);
nor U13522 (N_13522,N_12423,N_12491);
or U13523 (N_13523,N_12785,N_12705);
xor U13524 (N_13524,N_12391,N_12172);
xnor U13525 (N_13525,N_12291,N_12274);
nand U13526 (N_13526,N_12775,N_12533);
xnor U13527 (N_13527,N_12702,N_12055);
nor U13528 (N_13528,N_12106,N_12559);
xnor U13529 (N_13529,N_12086,N_12940);
or U13530 (N_13530,N_12984,N_12631);
or U13531 (N_13531,N_12198,N_12532);
nor U13532 (N_13532,N_12130,N_12162);
nor U13533 (N_13533,N_12454,N_12980);
nand U13534 (N_13534,N_12869,N_12083);
nor U13535 (N_13535,N_12035,N_12400);
or U13536 (N_13536,N_12662,N_12151);
and U13537 (N_13537,N_12625,N_12108);
nand U13538 (N_13538,N_12896,N_12518);
nor U13539 (N_13539,N_12354,N_12870);
nor U13540 (N_13540,N_12453,N_12817);
or U13541 (N_13541,N_12298,N_12341);
and U13542 (N_13542,N_12513,N_12897);
xor U13543 (N_13543,N_12402,N_12352);
xnor U13544 (N_13544,N_12209,N_12392);
or U13545 (N_13545,N_12201,N_12246);
nand U13546 (N_13546,N_12306,N_12285);
nand U13547 (N_13547,N_12647,N_12080);
or U13548 (N_13548,N_12742,N_12001);
xor U13549 (N_13549,N_12816,N_12276);
nand U13550 (N_13550,N_12581,N_12182);
xor U13551 (N_13551,N_12010,N_12864);
or U13552 (N_13552,N_12570,N_12024);
or U13553 (N_13553,N_12708,N_12975);
or U13554 (N_13554,N_12229,N_12664);
and U13555 (N_13555,N_12368,N_12990);
nand U13556 (N_13556,N_12905,N_12956);
nand U13557 (N_13557,N_12693,N_12151);
xnor U13558 (N_13558,N_12199,N_12768);
xnor U13559 (N_13559,N_12466,N_12865);
and U13560 (N_13560,N_12623,N_12899);
nand U13561 (N_13561,N_12487,N_12683);
nand U13562 (N_13562,N_12690,N_12759);
or U13563 (N_13563,N_12723,N_12542);
nand U13564 (N_13564,N_12558,N_12057);
or U13565 (N_13565,N_12670,N_12569);
nand U13566 (N_13566,N_12953,N_12103);
or U13567 (N_13567,N_12308,N_12471);
nor U13568 (N_13568,N_12954,N_12650);
nand U13569 (N_13569,N_12361,N_12563);
and U13570 (N_13570,N_12791,N_12774);
and U13571 (N_13571,N_12302,N_12190);
nand U13572 (N_13572,N_12766,N_12798);
and U13573 (N_13573,N_12887,N_12097);
nor U13574 (N_13574,N_12225,N_12791);
and U13575 (N_13575,N_12811,N_12706);
nor U13576 (N_13576,N_12345,N_12531);
nand U13577 (N_13577,N_12882,N_12710);
or U13578 (N_13578,N_12008,N_12582);
xor U13579 (N_13579,N_12831,N_12850);
nand U13580 (N_13580,N_12692,N_12780);
nor U13581 (N_13581,N_12884,N_12892);
or U13582 (N_13582,N_12122,N_12243);
nand U13583 (N_13583,N_12833,N_12137);
nand U13584 (N_13584,N_12932,N_12155);
nor U13585 (N_13585,N_12992,N_12552);
nand U13586 (N_13586,N_12930,N_12266);
nor U13587 (N_13587,N_12197,N_12731);
nor U13588 (N_13588,N_12897,N_12444);
nand U13589 (N_13589,N_12692,N_12601);
or U13590 (N_13590,N_12961,N_12017);
xnor U13591 (N_13591,N_12028,N_12935);
and U13592 (N_13592,N_12408,N_12311);
nor U13593 (N_13593,N_12701,N_12537);
or U13594 (N_13594,N_12662,N_12231);
xnor U13595 (N_13595,N_12338,N_12731);
and U13596 (N_13596,N_12126,N_12158);
and U13597 (N_13597,N_12249,N_12996);
and U13598 (N_13598,N_12968,N_12912);
nand U13599 (N_13599,N_12081,N_12900);
nor U13600 (N_13600,N_12879,N_12294);
and U13601 (N_13601,N_12978,N_12461);
nand U13602 (N_13602,N_12979,N_12502);
nor U13603 (N_13603,N_12842,N_12913);
and U13604 (N_13604,N_12294,N_12186);
nand U13605 (N_13605,N_12107,N_12422);
nor U13606 (N_13606,N_12951,N_12071);
nand U13607 (N_13607,N_12538,N_12493);
and U13608 (N_13608,N_12336,N_12441);
and U13609 (N_13609,N_12821,N_12482);
or U13610 (N_13610,N_12373,N_12075);
nand U13611 (N_13611,N_12944,N_12659);
nand U13612 (N_13612,N_12988,N_12186);
and U13613 (N_13613,N_12977,N_12342);
nand U13614 (N_13614,N_12479,N_12235);
or U13615 (N_13615,N_12442,N_12274);
or U13616 (N_13616,N_12423,N_12737);
nand U13617 (N_13617,N_12794,N_12853);
or U13618 (N_13618,N_12375,N_12971);
xnor U13619 (N_13619,N_12386,N_12908);
nand U13620 (N_13620,N_12754,N_12445);
nand U13621 (N_13621,N_12465,N_12303);
or U13622 (N_13622,N_12795,N_12939);
xnor U13623 (N_13623,N_12399,N_12685);
nor U13624 (N_13624,N_12901,N_12863);
and U13625 (N_13625,N_12078,N_12052);
and U13626 (N_13626,N_12460,N_12724);
nand U13627 (N_13627,N_12074,N_12380);
and U13628 (N_13628,N_12139,N_12260);
xor U13629 (N_13629,N_12735,N_12986);
xor U13630 (N_13630,N_12841,N_12063);
xor U13631 (N_13631,N_12843,N_12732);
nor U13632 (N_13632,N_12595,N_12623);
or U13633 (N_13633,N_12455,N_12927);
or U13634 (N_13634,N_12845,N_12164);
and U13635 (N_13635,N_12382,N_12129);
xor U13636 (N_13636,N_12480,N_12208);
nand U13637 (N_13637,N_12282,N_12226);
nand U13638 (N_13638,N_12138,N_12052);
nand U13639 (N_13639,N_12889,N_12600);
nor U13640 (N_13640,N_12393,N_12604);
or U13641 (N_13641,N_12068,N_12275);
nand U13642 (N_13642,N_12184,N_12089);
and U13643 (N_13643,N_12341,N_12224);
or U13644 (N_13644,N_12432,N_12472);
xor U13645 (N_13645,N_12036,N_12214);
or U13646 (N_13646,N_12035,N_12833);
or U13647 (N_13647,N_12763,N_12296);
or U13648 (N_13648,N_12121,N_12308);
xnor U13649 (N_13649,N_12036,N_12028);
xnor U13650 (N_13650,N_12022,N_12369);
xor U13651 (N_13651,N_12333,N_12579);
or U13652 (N_13652,N_12296,N_12442);
or U13653 (N_13653,N_12650,N_12087);
nand U13654 (N_13654,N_12899,N_12687);
nor U13655 (N_13655,N_12915,N_12485);
or U13656 (N_13656,N_12461,N_12121);
xor U13657 (N_13657,N_12574,N_12812);
xnor U13658 (N_13658,N_12524,N_12057);
nor U13659 (N_13659,N_12381,N_12518);
xnor U13660 (N_13660,N_12719,N_12546);
and U13661 (N_13661,N_12008,N_12816);
or U13662 (N_13662,N_12517,N_12808);
and U13663 (N_13663,N_12101,N_12782);
xor U13664 (N_13664,N_12179,N_12746);
and U13665 (N_13665,N_12433,N_12520);
and U13666 (N_13666,N_12049,N_12954);
and U13667 (N_13667,N_12337,N_12586);
nor U13668 (N_13668,N_12411,N_12207);
or U13669 (N_13669,N_12620,N_12108);
nand U13670 (N_13670,N_12993,N_12392);
xnor U13671 (N_13671,N_12256,N_12463);
or U13672 (N_13672,N_12283,N_12367);
and U13673 (N_13673,N_12693,N_12078);
xnor U13674 (N_13674,N_12546,N_12717);
or U13675 (N_13675,N_12261,N_12413);
or U13676 (N_13676,N_12373,N_12701);
xor U13677 (N_13677,N_12824,N_12887);
or U13678 (N_13678,N_12841,N_12785);
nand U13679 (N_13679,N_12127,N_12637);
or U13680 (N_13680,N_12238,N_12893);
nand U13681 (N_13681,N_12735,N_12049);
xor U13682 (N_13682,N_12654,N_12010);
nand U13683 (N_13683,N_12222,N_12995);
or U13684 (N_13684,N_12233,N_12842);
nor U13685 (N_13685,N_12067,N_12786);
xor U13686 (N_13686,N_12354,N_12843);
nor U13687 (N_13687,N_12298,N_12886);
nand U13688 (N_13688,N_12242,N_12095);
nor U13689 (N_13689,N_12851,N_12833);
xnor U13690 (N_13690,N_12767,N_12362);
nor U13691 (N_13691,N_12540,N_12793);
nand U13692 (N_13692,N_12208,N_12751);
xnor U13693 (N_13693,N_12887,N_12013);
or U13694 (N_13694,N_12989,N_12281);
xor U13695 (N_13695,N_12991,N_12770);
nor U13696 (N_13696,N_12793,N_12997);
and U13697 (N_13697,N_12582,N_12949);
nor U13698 (N_13698,N_12512,N_12063);
or U13699 (N_13699,N_12748,N_12343);
or U13700 (N_13700,N_12906,N_12388);
xor U13701 (N_13701,N_12457,N_12768);
nand U13702 (N_13702,N_12475,N_12499);
xor U13703 (N_13703,N_12336,N_12020);
nor U13704 (N_13704,N_12849,N_12060);
xor U13705 (N_13705,N_12371,N_12545);
and U13706 (N_13706,N_12246,N_12988);
nor U13707 (N_13707,N_12069,N_12786);
or U13708 (N_13708,N_12230,N_12201);
nor U13709 (N_13709,N_12250,N_12509);
or U13710 (N_13710,N_12377,N_12030);
nor U13711 (N_13711,N_12333,N_12842);
or U13712 (N_13712,N_12457,N_12064);
xor U13713 (N_13713,N_12677,N_12903);
and U13714 (N_13714,N_12293,N_12084);
or U13715 (N_13715,N_12122,N_12215);
or U13716 (N_13716,N_12768,N_12790);
and U13717 (N_13717,N_12254,N_12516);
or U13718 (N_13718,N_12342,N_12083);
xnor U13719 (N_13719,N_12685,N_12547);
nor U13720 (N_13720,N_12953,N_12719);
nor U13721 (N_13721,N_12130,N_12152);
or U13722 (N_13722,N_12340,N_12091);
or U13723 (N_13723,N_12830,N_12841);
and U13724 (N_13724,N_12072,N_12475);
xor U13725 (N_13725,N_12499,N_12871);
nand U13726 (N_13726,N_12376,N_12398);
nor U13727 (N_13727,N_12396,N_12189);
nand U13728 (N_13728,N_12158,N_12031);
or U13729 (N_13729,N_12595,N_12251);
or U13730 (N_13730,N_12782,N_12086);
nand U13731 (N_13731,N_12876,N_12870);
nand U13732 (N_13732,N_12153,N_12359);
xor U13733 (N_13733,N_12253,N_12643);
nor U13734 (N_13734,N_12827,N_12272);
and U13735 (N_13735,N_12683,N_12041);
nor U13736 (N_13736,N_12986,N_12987);
xor U13737 (N_13737,N_12531,N_12316);
nand U13738 (N_13738,N_12879,N_12196);
or U13739 (N_13739,N_12399,N_12671);
and U13740 (N_13740,N_12716,N_12028);
xor U13741 (N_13741,N_12919,N_12515);
xnor U13742 (N_13742,N_12335,N_12261);
nand U13743 (N_13743,N_12761,N_12070);
nand U13744 (N_13744,N_12170,N_12866);
nand U13745 (N_13745,N_12245,N_12530);
and U13746 (N_13746,N_12897,N_12288);
xnor U13747 (N_13747,N_12576,N_12467);
nand U13748 (N_13748,N_12774,N_12563);
or U13749 (N_13749,N_12667,N_12858);
or U13750 (N_13750,N_12713,N_12591);
and U13751 (N_13751,N_12190,N_12019);
and U13752 (N_13752,N_12969,N_12741);
nand U13753 (N_13753,N_12503,N_12099);
nor U13754 (N_13754,N_12659,N_12963);
xor U13755 (N_13755,N_12519,N_12978);
xor U13756 (N_13756,N_12595,N_12233);
or U13757 (N_13757,N_12540,N_12961);
nor U13758 (N_13758,N_12320,N_12316);
nor U13759 (N_13759,N_12067,N_12827);
nor U13760 (N_13760,N_12845,N_12744);
nor U13761 (N_13761,N_12674,N_12451);
or U13762 (N_13762,N_12057,N_12629);
or U13763 (N_13763,N_12202,N_12189);
nand U13764 (N_13764,N_12338,N_12005);
nor U13765 (N_13765,N_12208,N_12013);
nand U13766 (N_13766,N_12620,N_12658);
xnor U13767 (N_13767,N_12494,N_12722);
and U13768 (N_13768,N_12654,N_12018);
or U13769 (N_13769,N_12629,N_12264);
nand U13770 (N_13770,N_12729,N_12731);
nand U13771 (N_13771,N_12463,N_12738);
xnor U13772 (N_13772,N_12556,N_12414);
or U13773 (N_13773,N_12629,N_12985);
nor U13774 (N_13774,N_12014,N_12203);
and U13775 (N_13775,N_12319,N_12590);
nand U13776 (N_13776,N_12345,N_12546);
nor U13777 (N_13777,N_12352,N_12224);
or U13778 (N_13778,N_12820,N_12620);
or U13779 (N_13779,N_12817,N_12876);
or U13780 (N_13780,N_12538,N_12366);
xnor U13781 (N_13781,N_12752,N_12863);
nor U13782 (N_13782,N_12957,N_12004);
or U13783 (N_13783,N_12665,N_12819);
nand U13784 (N_13784,N_12339,N_12618);
and U13785 (N_13785,N_12699,N_12914);
nand U13786 (N_13786,N_12269,N_12294);
nand U13787 (N_13787,N_12792,N_12488);
and U13788 (N_13788,N_12790,N_12317);
xnor U13789 (N_13789,N_12021,N_12423);
nor U13790 (N_13790,N_12576,N_12523);
nor U13791 (N_13791,N_12596,N_12165);
nor U13792 (N_13792,N_12462,N_12450);
and U13793 (N_13793,N_12680,N_12315);
xnor U13794 (N_13794,N_12719,N_12280);
and U13795 (N_13795,N_12027,N_12551);
nand U13796 (N_13796,N_12405,N_12852);
xnor U13797 (N_13797,N_12329,N_12011);
or U13798 (N_13798,N_12274,N_12771);
and U13799 (N_13799,N_12618,N_12530);
and U13800 (N_13800,N_12300,N_12693);
and U13801 (N_13801,N_12247,N_12014);
nor U13802 (N_13802,N_12211,N_12002);
or U13803 (N_13803,N_12550,N_12797);
and U13804 (N_13804,N_12475,N_12333);
nor U13805 (N_13805,N_12053,N_12803);
nand U13806 (N_13806,N_12196,N_12817);
nand U13807 (N_13807,N_12823,N_12439);
and U13808 (N_13808,N_12399,N_12936);
xnor U13809 (N_13809,N_12777,N_12383);
xnor U13810 (N_13810,N_12633,N_12915);
nand U13811 (N_13811,N_12115,N_12079);
or U13812 (N_13812,N_12760,N_12651);
nor U13813 (N_13813,N_12199,N_12224);
or U13814 (N_13814,N_12752,N_12307);
nor U13815 (N_13815,N_12680,N_12857);
and U13816 (N_13816,N_12277,N_12979);
nand U13817 (N_13817,N_12955,N_12985);
xnor U13818 (N_13818,N_12125,N_12140);
and U13819 (N_13819,N_12104,N_12862);
or U13820 (N_13820,N_12685,N_12048);
nor U13821 (N_13821,N_12354,N_12711);
or U13822 (N_13822,N_12452,N_12490);
or U13823 (N_13823,N_12365,N_12126);
nand U13824 (N_13824,N_12950,N_12293);
and U13825 (N_13825,N_12325,N_12449);
and U13826 (N_13826,N_12187,N_12507);
nand U13827 (N_13827,N_12404,N_12339);
nand U13828 (N_13828,N_12221,N_12923);
and U13829 (N_13829,N_12175,N_12936);
or U13830 (N_13830,N_12497,N_12464);
or U13831 (N_13831,N_12521,N_12749);
xor U13832 (N_13832,N_12629,N_12887);
or U13833 (N_13833,N_12073,N_12888);
and U13834 (N_13834,N_12893,N_12159);
nor U13835 (N_13835,N_12679,N_12253);
xor U13836 (N_13836,N_12005,N_12934);
nand U13837 (N_13837,N_12347,N_12625);
or U13838 (N_13838,N_12616,N_12943);
and U13839 (N_13839,N_12311,N_12454);
xnor U13840 (N_13840,N_12793,N_12557);
nor U13841 (N_13841,N_12427,N_12915);
and U13842 (N_13842,N_12275,N_12206);
or U13843 (N_13843,N_12241,N_12203);
nand U13844 (N_13844,N_12757,N_12811);
nand U13845 (N_13845,N_12847,N_12108);
nand U13846 (N_13846,N_12278,N_12472);
or U13847 (N_13847,N_12399,N_12221);
nand U13848 (N_13848,N_12552,N_12805);
nor U13849 (N_13849,N_12001,N_12558);
and U13850 (N_13850,N_12575,N_12724);
or U13851 (N_13851,N_12453,N_12308);
and U13852 (N_13852,N_12148,N_12550);
nor U13853 (N_13853,N_12255,N_12505);
nor U13854 (N_13854,N_12336,N_12129);
and U13855 (N_13855,N_12270,N_12720);
or U13856 (N_13856,N_12843,N_12434);
nor U13857 (N_13857,N_12222,N_12541);
or U13858 (N_13858,N_12649,N_12921);
nor U13859 (N_13859,N_12034,N_12725);
nor U13860 (N_13860,N_12667,N_12339);
nand U13861 (N_13861,N_12987,N_12348);
nand U13862 (N_13862,N_12209,N_12278);
xnor U13863 (N_13863,N_12287,N_12383);
or U13864 (N_13864,N_12013,N_12080);
and U13865 (N_13865,N_12730,N_12827);
nand U13866 (N_13866,N_12554,N_12556);
nor U13867 (N_13867,N_12073,N_12543);
xnor U13868 (N_13868,N_12091,N_12822);
and U13869 (N_13869,N_12446,N_12684);
xnor U13870 (N_13870,N_12618,N_12973);
and U13871 (N_13871,N_12856,N_12125);
and U13872 (N_13872,N_12480,N_12700);
nand U13873 (N_13873,N_12302,N_12840);
and U13874 (N_13874,N_12533,N_12955);
nor U13875 (N_13875,N_12565,N_12625);
nand U13876 (N_13876,N_12510,N_12206);
xor U13877 (N_13877,N_12851,N_12528);
xnor U13878 (N_13878,N_12065,N_12925);
nor U13879 (N_13879,N_12432,N_12414);
nor U13880 (N_13880,N_12781,N_12972);
nand U13881 (N_13881,N_12698,N_12086);
or U13882 (N_13882,N_12880,N_12527);
and U13883 (N_13883,N_12179,N_12020);
nand U13884 (N_13884,N_12715,N_12088);
and U13885 (N_13885,N_12623,N_12009);
and U13886 (N_13886,N_12370,N_12755);
and U13887 (N_13887,N_12410,N_12147);
or U13888 (N_13888,N_12967,N_12339);
or U13889 (N_13889,N_12329,N_12712);
xnor U13890 (N_13890,N_12932,N_12050);
nor U13891 (N_13891,N_12069,N_12739);
nand U13892 (N_13892,N_12711,N_12573);
nor U13893 (N_13893,N_12905,N_12580);
and U13894 (N_13894,N_12782,N_12663);
xnor U13895 (N_13895,N_12680,N_12707);
or U13896 (N_13896,N_12927,N_12702);
or U13897 (N_13897,N_12043,N_12676);
or U13898 (N_13898,N_12490,N_12546);
nand U13899 (N_13899,N_12935,N_12749);
or U13900 (N_13900,N_12039,N_12740);
nor U13901 (N_13901,N_12971,N_12940);
nor U13902 (N_13902,N_12555,N_12569);
or U13903 (N_13903,N_12843,N_12017);
and U13904 (N_13904,N_12366,N_12540);
or U13905 (N_13905,N_12661,N_12209);
xnor U13906 (N_13906,N_12144,N_12048);
nand U13907 (N_13907,N_12950,N_12122);
xnor U13908 (N_13908,N_12378,N_12654);
nor U13909 (N_13909,N_12732,N_12452);
xnor U13910 (N_13910,N_12322,N_12711);
and U13911 (N_13911,N_12132,N_12642);
and U13912 (N_13912,N_12779,N_12841);
or U13913 (N_13913,N_12058,N_12618);
nor U13914 (N_13914,N_12783,N_12293);
and U13915 (N_13915,N_12139,N_12795);
and U13916 (N_13916,N_12657,N_12861);
nand U13917 (N_13917,N_12866,N_12030);
xor U13918 (N_13918,N_12857,N_12034);
or U13919 (N_13919,N_12107,N_12582);
and U13920 (N_13920,N_12877,N_12126);
and U13921 (N_13921,N_12232,N_12712);
or U13922 (N_13922,N_12072,N_12286);
or U13923 (N_13923,N_12559,N_12901);
nor U13924 (N_13924,N_12609,N_12475);
xnor U13925 (N_13925,N_12323,N_12446);
nor U13926 (N_13926,N_12949,N_12736);
nor U13927 (N_13927,N_12640,N_12784);
nand U13928 (N_13928,N_12768,N_12431);
nor U13929 (N_13929,N_12091,N_12020);
nand U13930 (N_13930,N_12012,N_12130);
or U13931 (N_13931,N_12593,N_12714);
nand U13932 (N_13932,N_12380,N_12350);
or U13933 (N_13933,N_12004,N_12847);
nor U13934 (N_13934,N_12246,N_12790);
and U13935 (N_13935,N_12801,N_12845);
or U13936 (N_13936,N_12652,N_12485);
or U13937 (N_13937,N_12056,N_12918);
nand U13938 (N_13938,N_12552,N_12013);
nand U13939 (N_13939,N_12183,N_12481);
and U13940 (N_13940,N_12755,N_12123);
xnor U13941 (N_13941,N_12840,N_12675);
and U13942 (N_13942,N_12629,N_12231);
nor U13943 (N_13943,N_12321,N_12199);
nand U13944 (N_13944,N_12016,N_12966);
or U13945 (N_13945,N_12021,N_12411);
xor U13946 (N_13946,N_12659,N_12447);
xor U13947 (N_13947,N_12059,N_12578);
nand U13948 (N_13948,N_12257,N_12922);
nor U13949 (N_13949,N_12909,N_12289);
nand U13950 (N_13950,N_12637,N_12108);
nor U13951 (N_13951,N_12433,N_12436);
and U13952 (N_13952,N_12727,N_12497);
or U13953 (N_13953,N_12951,N_12156);
or U13954 (N_13954,N_12506,N_12179);
and U13955 (N_13955,N_12189,N_12344);
and U13956 (N_13956,N_12698,N_12985);
nor U13957 (N_13957,N_12085,N_12883);
and U13958 (N_13958,N_12934,N_12643);
or U13959 (N_13959,N_12626,N_12355);
nand U13960 (N_13960,N_12874,N_12918);
and U13961 (N_13961,N_12275,N_12270);
nand U13962 (N_13962,N_12479,N_12695);
and U13963 (N_13963,N_12252,N_12445);
and U13964 (N_13964,N_12828,N_12825);
nor U13965 (N_13965,N_12184,N_12351);
nor U13966 (N_13966,N_12504,N_12863);
xnor U13967 (N_13967,N_12269,N_12508);
nand U13968 (N_13968,N_12159,N_12872);
xnor U13969 (N_13969,N_12496,N_12627);
and U13970 (N_13970,N_12219,N_12919);
xnor U13971 (N_13971,N_12330,N_12704);
and U13972 (N_13972,N_12288,N_12419);
and U13973 (N_13973,N_12142,N_12542);
or U13974 (N_13974,N_12282,N_12360);
or U13975 (N_13975,N_12577,N_12012);
xor U13976 (N_13976,N_12720,N_12958);
nand U13977 (N_13977,N_12122,N_12031);
nand U13978 (N_13978,N_12376,N_12201);
or U13979 (N_13979,N_12336,N_12113);
nand U13980 (N_13980,N_12093,N_12238);
or U13981 (N_13981,N_12159,N_12768);
or U13982 (N_13982,N_12942,N_12659);
nand U13983 (N_13983,N_12067,N_12525);
nor U13984 (N_13984,N_12640,N_12817);
or U13985 (N_13985,N_12567,N_12604);
nand U13986 (N_13986,N_12329,N_12153);
nand U13987 (N_13987,N_12126,N_12109);
nand U13988 (N_13988,N_12214,N_12281);
nand U13989 (N_13989,N_12979,N_12215);
and U13990 (N_13990,N_12314,N_12916);
and U13991 (N_13991,N_12817,N_12773);
xnor U13992 (N_13992,N_12900,N_12857);
nor U13993 (N_13993,N_12250,N_12482);
and U13994 (N_13994,N_12004,N_12110);
xor U13995 (N_13995,N_12160,N_12203);
nand U13996 (N_13996,N_12971,N_12491);
and U13997 (N_13997,N_12623,N_12665);
or U13998 (N_13998,N_12496,N_12036);
and U13999 (N_13999,N_12845,N_12298);
and U14000 (N_14000,N_13864,N_13402);
xnor U14001 (N_14001,N_13164,N_13742);
nand U14002 (N_14002,N_13494,N_13824);
nor U14003 (N_14003,N_13495,N_13400);
nor U14004 (N_14004,N_13765,N_13027);
nand U14005 (N_14005,N_13235,N_13318);
and U14006 (N_14006,N_13951,N_13143);
nor U14007 (N_14007,N_13776,N_13994);
xor U14008 (N_14008,N_13604,N_13751);
nor U14009 (N_14009,N_13474,N_13024);
nand U14010 (N_14010,N_13968,N_13219);
nand U14011 (N_14011,N_13154,N_13408);
nand U14012 (N_14012,N_13192,N_13735);
or U14013 (N_14013,N_13950,N_13890);
and U14014 (N_14014,N_13882,N_13122);
or U14015 (N_14015,N_13060,N_13306);
xnor U14016 (N_14016,N_13415,N_13443);
nor U14017 (N_14017,N_13791,N_13843);
nor U14018 (N_14018,N_13386,N_13685);
xor U14019 (N_14019,N_13697,N_13709);
or U14020 (N_14020,N_13658,N_13545);
and U14021 (N_14021,N_13194,N_13059);
nor U14022 (N_14022,N_13939,N_13509);
nand U14023 (N_14023,N_13457,N_13915);
nor U14024 (N_14024,N_13207,N_13346);
and U14025 (N_14025,N_13202,N_13562);
and U14026 (N_14026,N_13330,N_13050);
nor U14027 (N_14027,N_13568,N_13260);
or U14028 (N_14028,N_13019,N_13963);
and U14029 (N_14029,N_13577,N_13985);
or U14030 (N_14030,N_13512,N_13584);
xor U14031 (N_14031,N_13233,N_13593);
xnor U14032 (N_14032,N_13838,N_13758);
and U14033 (N_14033,N_13690,N_13480);
nor U14034 (N_14034,N_13935,N_13273);
nand U14035 (N_14035,N_13309,N_13611);
nor U14036 (N_14036,N_13904,N_13669);
xnor U14037 (N_14037,N_13388,N_13392);
xnor U14038 (N_14038,N_13391,N_13767);
or U14039 (N_14039,N_13030,N_13289);
and U14040 (N_14040,N_13799,N_13752);
nand U14041 (N_14041,N_13499,N_13465);
and U14042 (N_14042,N_13720,N_13255);
nor U14043 (N_14043,N_13090,N_13364);
xnor U14044 (N_14044,N_13681,N_13608);
and U14045 (N_14045,N_13874,N_13793);
nand U14046 (N_14046,N_13095,N_13313);
and U14047 (N_14047,N_13597,N_13842);
nand U14048 (N_14048,N_13085,N_13253);
nor U14049 (N_14049,N_13221,N_13769);
nand U14050 (N_14050,N_13013,N_13999);
nor U14051 (N_14051,N_13533,N_13492);
nor U14052 (N_14052,N_13239,N_13215);
nand U14053 (N_14053,N_13600,N_13351);
and U14054 (N_14054,N_13760,N_13020);
xor U14055 (N_14055,N_13908,N_13117);
xor U14056 (N_14056,N_13026,N_13980);
or U14057 (N_14057,N_13648,N_13419);
xor U14058 (N_14058,N_13454,N_13327);
xor U14059 (N_14059,N_13649,N_13097);
or U14060 (N_14060,N_13307,N_13771);
xnor U14061 (N_14061,N_13691,N_13531);
nor U14062 (N_14062,N_13259,N_13815);
nand U14063 (N_14063,N_13749,N_13189);
nor U14064 (N_14064,N_13502,N_13360);
nand U14065 (N_14065,N_13245,N_13755);
nand U14066 (N_14066,N_13088,N_13655);
or U14067 (N_14067,N_13353,N_13661);
nor U14068 (N_14068,N_13078,N_13764);
and U14069 (N_14069,N_13514,N_13437);
nand U14070 (N_14070,N_13871,N_13011);
nor U14071 (N_14071,N_13517,N_13673);
and U14072 (N_14072,N_13038,N_13425);
xnor U14073 (N_14073,N_13003,N_13031);
xor U14074 (N_14074,N_13879,N_13010);
nand U14075 (N_14075,N_13505,N_13487);
xor U14076 (N_14076,N_13863,N_13200);
xnor U14077 (N_14077,N_13894,N_13250);
and U14078 (N_14078,N_13845,N_13814);
xor U14079 (N_14079,N_13158,N_13797);
or U14080 (N_14080,N_13766,N_13537);
nand U14081 (N_14081,N_13867,N_13712);
nand U14082 (N_14082,N_13989,N_13555);
and U14083 (N_14083,N_13988,N_13801);
nand U14084 (N_14084,N_13466,N_13970);
or U14085 (N_14085,N_13785,N_13302);
nand U14086 (N_14086,N_13380,N_13934);
and U14087 (N_14087,N_13439,N_13852);
or U14088 (N_14088,N_13528,N_13228);
and U14089 (N_14089,N_13226,N_13706);
xor U14090 (N_14090,N_13264,N_13204);
and U14091 (N_14091,N_13075,N_13998);
and U14092 (N_14092,N_13639,N_13628);
nand U14093 (N_14093,N_13096,N_13780);
xnor U14094 (N_14094,N_13813,N_13564);
and U14095 (N_14095,N_13556,N_13162);
nor U14096 (N_14096,N_13073,N_13042);
or U14097 (N_14097,N_13525,N_13111);
or U14098 (N_14098,N_13405,N_13535);
and U14099 (N_14099,N_13906,N_13914);
and U14100 (N_14100,N_13884,N_13184);
and U14101 (N_14101,N_13945,N_13316);
nor U14102 (N_14102,N_13576,N_13949);
xnor U14103 (N_14103,N_13279,N_13188);
nor U14104 (N_14104,N_13686,N_13272);
or U14105 (N_14105,N_13147,N_13034);
or U14106 (N_14106,N_13682,N_13716);
nand U14107 (N_14107,N_13243,N_13479);
or U14108 (N_14108,N_13047,N_13839);
nor U14109 (N_14109,N_13298,N_13917);
nand U14110 (N_14110,N_13549,N_13293);
nor U14111 (N_14111,N_13782,N_13654);
and U14112 (N_14112,N_13249,N_13621);
and U14113 (N_14113,N_13507,N_13984);
or U14114 (N_14114,N_13009,N_13893);
nor U14115 (N_14115,N_13952,N_13727);
or U14116 (N_14116,N_13053,N_13996);
or U14117 (N_14117,N_13394,N_13198);
nor U14118 (N_14118,N_13961,N_13421);
or U14119 (N_14119,N_13041,N_13777);
nand U14120 (N_14120,N_13510,N_13598);
or U14121 (N_14121,N_13878,N_13211);
or U14122 (N_14122,N_13678,N_13521);
and U14123 (N_14123,N_13870,N_13213);
and U14124 (N_14124,N_13627,N_13885);
nand U14125 (N_14125,N_13633,N_13331);
nand U14126 (N_14126,N_13396,N_13435);
and U14127 (N_14127,N_13978,N_13444);
and U14128 (N_14128,N_13106,N_13163);
and U14129 (N_14129,N_13569,N_13848);
nand U14130 (N_14130,N_13017,N_13729);
and U14131 (N_14131,N_13612,N_13965);
nor U14132 (N_14132,N_13734,N_13288);
nand U14133 (N_14133,N_13744,N_13028);
and U14134 (N_14134,N_13553,N_13183);
and U14135 (N_14135,N_13857,N_13937);
nor U14136 (N_14136,N_13354,N_13077);
or U14137 (N_14137,N_13614,N_13543);
or U14138 (N_14138,N_13818,N_13508);
nand U14139 (N_14139,N_13299,N_13315);
nand U14140 (N_14140,N_13365,N_13643);
nor U14141 (N_14141,N_13370,N_13770);
xor U14142 (N_14142,N_13805,N_13208);
and U14143 (N_14143,N_13640,N_13150);
or U14144 (N_14144,N_13087,N_13976);
xnor U14145 (N_14145,N_13625,N_13240);
nor U14146 (N_14146,N_13109,N_13779);
xor U14147 (N_14147,N_13825,N_13483);
nor U14148 (N_14148,N_13647,N_13303);
xnor U14149 (N_14149,N_13763,N_13702);
xnor U14150 (N_14150,N_13110,N_13039);
or U14151 (N_14151,N_13834,N_13317);
or U14152 (N_14152,N_13114,N_13218);
nor U14153 (N_14153,N_13574,N_13982);
nor U14154 (N_14154,N_13276,N_13187);
xnor U14155 (N_14155,N_13237,N_13775);
xor U14156 (N_14156,N_13103,N_13458);
nor U14157 (N_14157,N_13137,N_13389);
xor U14158 (N_14158,N_13591,N_13589);
nand U14159 (N_14159,N_13877,N_13212);
xor U14160 (N_14160,N_13100,N_13349);
or U14161 (N_14161,N_13638,N_13489);
or U14162 (N_14162,N_13446,N_13520);
xnor U14163 (N_14163,N_13918,N_13025);
nor U14164 (N_14164,N_13049,N_13714);
nor U14165 (N_14165,N_13384,N_13282);
nand U14166 (N_14166,N_13196,N_13107);
and U14167 (N_14167,N_13021,N_13862);
xor U14168 (N_14168,N_13821,N_13367);
and U14169 (N_14169,N_13660,N_13515);
nand U14170 (N_14170,N_13693,N_13227);
or U14171 (N_14171,N_13179,N_13504);
or U14172 (N_14172,N_13886,N_13448);
xor U14173 (N_14173,N_13414,N_13539);
xnor U14174 (N_14174,N_13800,N_13610);
nor U14175 (N_14175,N_13708,N_13888);
nand U14176 (N_14176,N_13420,N_13944);
nor U14177 (N_14177,N_13571,N_13062);
xnor U14178 (N_14178,N_13832,N_13692);
or U14179 (N_14179,N_13687,N_13773);
and U14180 (N_14180,N_13244,N_13133);
and U14181 (N_14181,N_13417,N_13881);
nor U14182 (N_14182,N_13067,N_13456);
nor U14183 (N_14183,N_13153,N_13513);
and U14184 (N_14184,N_13830,N_13728);
nor U14185 (N_14185,N_13375,N_13296);
or U14186 (N_14186,N_13201,N_13322);
and U14187 (N_14187,N_13694,N_13928);
xor U14188 (N_14188,N_13004,N_13563);
xnor U14189 (N_14189,N_13339,N_13946);
and U14190 (N_14190,N_13646,N_13450);
nor U14191 (N_14191,N_13018,N_13971);
xor U14192 (N_14192,N_13256,N_13230);
or U14193 (N_14193,N_13721,N_13740);
or U14194 (N_14194,N_13193,N_13962);
or U14195 (N_14195,N_13441,N_13461);
and U14196 (N_14196,N_13623,N_13774);
nor U14197 (N_14197,N_13008,N_13328);
nand U14198 (N_14198,N_13223,N_13398);
nand U14199 (N_14199,N_13580,N_13558);
nor U14200 (N_14200,N_13873,N_13599);
and U14201 (N_14201,N_13592,N_13897);
nand U14202 (N_14202,N_13467,N_13300);
nor U14203 (N_14203,N_13206,N_13642);
or U14204 (N_14204,N_13175,N_13772);
nand U14205 (N_14205,N_13098,N_13145);
or U14206 (N_14206,N_13975,N_13231);
or U14207 (N_14207,N_13781,N_13203);
nand U14208 (N_14208,N_13899,N_13040);
nor U14209 (N_14209,N_13858,N_13176);
nor U14210 (N_14210,N_13002,N_13093);
or U14211 (N_14211,N_13822,N_13632);
nor U14212 (N_14212,N_13058,N_13674);
nor U14213 (N_14213,N_13872,N_13254);
and U14214 (N_14214,N_13321,N_13333);
nand U14215 (N_14215,N_13529,N_13631);
and U14216 (N_14216,N_13565,N_13941);
or U14217 (N_14217,N_13753,N_13526);
or U14218 (N_14218,N_13068,N_13156);
and U14219 (N_14219,N_13451,N_13338);
xor U14220 (N_14220,N_13119,N_13554);
xor U14221 (N_14221,N_13719,N_13836);
and U14222 (N_14222,N_13178,N_13329);
and U14223 (N_14223,N_13074,N_13341);
xnor U14224 (N_14224,N_13345,N_13622);
nor U14225 (N_14225,N_13807,N_13966);
and U14226 (N_14226,N_13585,N_13356);
xnor U14227 (N_14227,N_13596,N_13146);
and U14228 (N_14228,N_13159,N_13748);
or U14229 (N_14229,N_13485,N_13662);
or U14230 (N_14230,N_13995,N_13355);
xor U14231 (N_14231,N_13573,N_13875);
nand U14232 (N_14232,N_13866,N_13155);
nand U14233 (N_14233,N_13594,N_13536);
nand U14234 (N_14234,N_13173,N_13301);
and U14235 (N_14235,N_13091,N_13855);
and U14236 (N_14236,N_13972,N_13348);
nand U14237 (N_14237,N_13992,N_13718);
and U14238 (N_14238,N_13261,N_13581);
xnor U14239 (N_14239,N_13374,N_13715);
nand U14240 (N_14240,N_13506,N_13583);
or U14241 (N_14241,N_13029,N_13248);
nand U14242 (N_14242,N_13251,N_13079);
xnor U14243 (N_14243,N_13567,N_13524);
xor U14244 (N_14244,N_13634,N_13007);
and U14245 (N_14245,N_13683,N_13063);
and U14246 (N_14246,N_13490,N_13698);
nor U14247 (N_14247,N_13116,N_13786);
xnor U14248 (N_14248,N_13501,N_13166);
nor U14249 (N_14249,N_13932,N_13387);
xor U14250 (N_14250,N_13579,N_13666);
xor U14251 (N_14251,N_13741,N_13991);
xnor U14252 (N_14252,N_13667,N_13217);
or U14253 (N_14253,N_13500,N_13071);
and U14254 (N_14254,N_13768,N_13268);
and U14255 (N_14255,N_13787,N_13267);
nand U14256 (N_14256,N_13413,N_13933);
nor U14257 (N_14257,N_13403,N_13738);
nor U14258 (N_14258,N_13656,N_13689);
nor U14259 (N_14259,N_13283,N_13121);
nand U14260 (N_14260,N_13829,N_13802);
xnor U14261 (N_14261,N_13120,N_13817);
nor U14262 (N_14262,N_13503,N_13379);
xnor U14263 (N_14263,N_13497,N_13925);
and U14264 (N_14264,N_13828,N_13523);
nand U14265 (N_14265,N_13860,N_13827);
nand U14266 (N_14266,N_13544,N_13588);
nor U14267 (N_14267,N_13312,N_13703);
nor U14268 (N_14268,N_13089,N_13901);
nor U14269 (N_14269,N_13723,N_13618);
or U14270 (N_14270,N_13141,N_13232);
nor U14271 (N_14271,N_13916,N_13725);
nand U14272 (N_14272,N_13134,N_13280);
and U14273 (N_14273,N_13603,N_13923);
or U14274 (N_14274,N_13366,N_13803);
or U14275 (N_14275,N_13900,N_13205);
and U14276 (N_14276,N_13960,N_13488);
nor U14277 (N_14277,N_13587,N_13859);
nand U14278 (N_14278,N_13129,N_13304);
or U14279 (N_14279,N_13938,N_13373);
xor U14280 (N_14280,N_13459,N_13149);
or U14281 (N_14281,N_13650,N_13064);
and U14282 (N_14282,N_13383,N_13411);
xor U14283 (N_14283,N_13516,N_13433);
nand U14284 (N_14284,N_13144,N_13710);
xor U14285 (N_14285,N_13665,N_13644);
nand U14286 (N_14286,N_13796,N_13378);
xor U14287 (N_14287,N_13167,N_13455);
and U14288 (N_14288,N_13498,N_13371);
or U14289 (N_14289,N_13854,N_13376);
or U14290 (N_14290,N_13462,N_13086);
nand U14291 (N_14291,N_13595,N_13438);
nand U14292 (N_14292,N_13065,N_13668);
nor U14293 (N_14293,N_13344,N_13547);
nand U14294 (N_14294,N_13534,N_13808);
xor U14295 (N_14295,N_13546,N_13810);
nor U14296 (N_14296,N_13056,N_13615);
nor U14297 (N_14297,N_13473,N_13757);
or U14298 (N_14298,N_13132,N_13586);
nand U14299 (N_14299,N_13138,N_13055);
or U14300 (N_14300,N_13139,N_13182);
nor U14301 (N_14301,N_13442,N_13731);
or U14302 (N_14302,N_13334,N_13426);
nand U14303 (N_14303,N_13191,N_13675);
nor U14304 (N_14304,N_13983,N_13907);
xnor U14305 (N_14305,N_13696,N_13127);
or U14306 (N_14306,N_13266,N_13432);
or U14307 (N_14307,N_13294,N_13036);
and U14308 (N_14308,N_13607,N_13912);
and U14309 (N_14309,N_13561,N_13151);
nand U14310 (N_14310,N_13477,N_13436);
or U14311 (N_14311,N_13157,N_13820);
nor U14312 (N_14312,N_13620,N_13072);
or U14313 (N_14313,N_13393,N_13320);
or U14314 (N_14314,N_13726,N_13560);
or U14315 (N_14315,N_13286,N_13883);
nand U14316 (N_14316,N_13680,N_13125);
xor U14317 (N_14317,N_13229,N_13979);
and U14318 (N_14318,N_13676,N_13406);
nor U14319 (N_14319,N_13493,N_13342);
or U14320 (N_14320,N_13238,N_13126);
nor U14321 (N_14321,N_13833,N_13168);
nor U14322 (N_14322,N_13572,N_13804);
or U14323 (N_14323,N_13352,N_13084);
or U14324 (N_14324,N_13737,N_13269);
or U14325 (N_14325,N_13453,N_13128);
or U14326 (N_14326,N_13142,N_13395);
and U14327 (N_14327,N_13789,N_13958);
xor U14328 (N_14328,N_13242,N_13246);
or U14329 (N_14329,N_13214,N_13275);
nor U14330 (N_14330,N_13340,N_13409);
and U14331 (N_14331,N_13012,N_13898);
nor U14332 (N_14332,N_13762,N_13337);
xnor U14333 (N_14333,N_13362,N_13861);
nor U14334 (N_14334,N_13434,N_13684);
and U14335 (N_14335,N_13548,N_13241);
nand U14336 (N_14336,N_13051,N_13806);
and U14337 (N_14337,N_13407,N_13739);
nand U14338 (N_14338,N_13278,N_13343);
or U14339 (N_14339,N_13636,N_13974);
and U14340 (N_14340,N_13990,N_13177);
nor U14341 (N_14341,N_13291,N_13478);
nor U14342 (N_14342,N_13000,N_13940);
xor U14343 (N_14343,N_13118,N_13936);
nand U14344 (N_14344,N_13284,N_13629);
nand U14345 (N_14345,N_13601,N_13794);
nor U14346 (N_14346,N_13688,N_13981);
and U14347 (N_14347,N_13037,N_13993);
nor U14348 (N_14348,N_13997,N_13837);
nor U14349 (N_14349,N_13161,N_13181);
xor U14350 (N_14350,N_13148,N_13043);
nor U14351 (N_14351,N_13209,N_13428);
xor U14352 (N_14352,N_13530,N_13606);
or U14353 (N_14353,N_13846,N_13713);
or U14354 (N_14354,N_13361,N_13609);
and U14355 (N_14355,N_13277,N_13310);
nand U14356 (N_14356,N_13171,N_13657);
nand U14357 (N_14357,N_13613,N_13112);
and U14358 (N_14358,N_13224,N_13423);
nor U14359 (N_14359,N_13750,N_13197);
nand U14360 (N_14360,N_13397,N_13174);
or U14361 (N_14361,N_13195,N_13672);
nand U14362 (N_14362,N_13566,N_13977);
nand U14363 (N_14363,N_13105,N_13115);
xor U14364 (N_14364,N_13108,N_13853);
xor U14365 (N_14365,N_13736,N_13390);
nor U14366 (N_14366,N_13418,N_13880);
and U14367 (N_14367,N_13677,N_13323);
and U14368 (N_14368,N_13826,N_13022);
or U14369 (N_14369,N_13236,N_13430);
or U14370 (N_14370,N_13840,N_13066);
and U14371 (N_14371,N_13987,N_13258);
and U14372 (N_14372,N_13033,N_13169);
and U14373 (N_14373,N_13788,N_13947);
xor U14374 (N_14374,N_13369,N_13519);
nor U14375 (N_14375,N_13257,N_13557);
or U14376 (N_14376,N_13054,N_13730);
and U14377 (N_14377,N_13185,N_13052);
or U14378 (N_14378,N_13921,N_13092);
and U14379 (N_14379,N_13372,N_13460);
xnor U14380 (N_14380,N_13124,N_13332);
nor U14381 (N_14381,N_13954,N_13522);
nor U14382 (N_14382,N_13160,N_13216);
or U14383 (N_14383,N_13659,N_13496);
and U14384 (N_14384,N_13297,N_13913);
nor U14385 (N_14385,N_13305,N_13717);
xnor U14386 (N_14386,N_13180,N_13541);
or U14387 (N_14387,N_13252,N_13001);
nor U14388 (N_14388,N_13819,N_13445);
and U14389 (N_14389,N_13210,N_13699);
nor U14390 (N_14390,N_13399,N_13724);
and U14391 (N_14391,N_13247,N_13057);
and U14392 (N_14392,N_13582,N_13412);
and U14393 (N_14393,N_13926,N_13876);
or U14394 (N_14394,N_13271,N_13889);
and U14395 (N_14395,N_13263,N_13358);
xnor U14396 (N_14396,N_13104,N_13722);
xnor U14397 (N_14397,N_13401,N_13754);
nand U14398 (N_14398,N_13005,N_13746);
nor U14399 (N_14399,N_13705,N_13792);
or U14400 (N_14400,N_13551,N_13835);
and U14401 (N_14401,N_13790,N_13641);
nor U14402 (N_14402,N_13082,N_13903);
and U14403 (N_14403,N_13319,N_13747);
nor U14404 (N_14404,N_13955,N_13578);
xnor U14405 (N_14405,N_13942,N_13482);
nand U14406 (N_14406,N_13759,N_13905);
nand U14407 (N_14407,N_13652,N_13637);
nor U14408 (N_14408,N_13070,N_13131);
nor U14409 (N_14409,N_13326,N_13484);
xnor U14410 (N_14410,N_13416,N_13491);
xor U14411 (N_14411,N_13651,N_13045);
nor U14412 (N_14412,N_13140,N_13927);
and U14413 (N_14413,N_13948,N_13919);
nand U14414 (N_14414,N_13325,N_13469);
nand U14415 (N_14415,N_13812,N_13559);
nand U14416 (N_14416,N_13920,N_13048);
or U14417 (N_14417,N_13404,N_13518);
nor U14418 (N_14418,N_13743,N_13381);
nor U14419 (N_14419,N_13552,N_13895);
and U14420 (N_14420,N_13700,N_13670);
nand U14421 (N_14421,N_13102,N_13130);
nand U14422 (N_14422,N_13964,N_13679);
xor U14423 (N_14423,N_13671,N_13849);
and U14424 (N_14424,N_13816,N_13841);
nor U14425 (N_14425,N_13382,N_13851);
nor U14426 (N_14426,N_13101,N_13570);
xnor U14427 (N_14427,N_13464,N_13014);
nor U14428 (N_14428,N_13527,N_13135);
or U14429 (N_14429,N_13290,N_13220);
nor U14430 (N_14430,N_13626,N_13347);
and U14431 (N_14431,N_13959,N_13429);
or U14432 (N_14432,N_13733,N_13083);
nor U14433 (N_14433,N_13784,N_13186);
and U14434 (N_14434,N_13909,N_13069);
nand U14435 (N_14435,N_13481,N_13969);
nor U14436 (N_14436,N_13080,N_13165);
and U14437 (N_14437,N_13645,N_13359);
nor U14438 (N_14438,N_13778,N_13540);
or U14439 (N_14439,N_13311,N_13590);
and U14440 (N_14440,N_13427,N_13287);
nor U14441 (N_14441,N_13061,N_13424);
and U14442 (N_14442,N_13225,N_13016);
xnor U14443 (N_14443,N_13973,N_13447);
xnor U14444 (N_14444,N_13471,N_13314);
nor U14445 (N_14445,N_13123,N_13511);
and U14446 (N_14446,N_13046,N_13274);
nand U14447 (N_14447,N_13199,N_13930);
and U14448 (N_14448,N_13486,N_13619);
xor U14449 (N_14449,N_13902,N_13023);
xor U14450 (N_14450,N_13422,N_13953);
nor U14451 (N_14451,N_13265,N_13711);
xnor U14452 (N_14452,N_13811,N_13887);
or U14453 (N_14453,N_13136,N_13865);
xnor U14454 (N_14454,N_13911,N_13295);
or U14455 (N_14455,N_13368,N_13663);
and U14456 (N_14456,N_13431,N_13234);
or U14457 (N_14457,N_13152,N_13281);
and U14458 (N_14458,N_13015,N_13336);
nand U14459 (N_14459,N_13463,N_13761);
or U14460 (N_14460,N_13910,N_13099);
and U14461 (N_14461,N_13308,N_13172);
and U14462 (N_14462,N_13868,N_13844);
xor U14463 (N_14463,N_13831,N_13896);
or U14464 (N_14464,N_13170,N_13624);
xor U14465 (N_14465,N_13350,N_13285);
or U14466 (N_14466,N_13410,N_13470);
or U14467 (N_14467,N_13850,N_13542);
xnor U14468 (N_14468,N_13924,N_13575);
or U14469 (N_14469,N_13449,N_13892);
nor U14470 (N_14470,N_13094,N_13856);
nand U14471 (N_14471,N_13967,N_13695);
nor U14472 (N_14472,N_13076,N_13704);
nand U14473 (N_14473,N_13756,N_13986);
or U14474 (N_14474,N_13292,N_13809);
and U14475 (N_14475,N_13616,N_13032);
nor U14476 (N_14476,N_13081,N_13222);
nand U14477 (N_14477,N_13617,N_13190);
nand U14478 (N_14478,N_13476,N_13452);
nand U14479 (N_14479,N_13943,N_13957);
or U14480 (N_14480,N_13798,N_13113);
or U14481 (N_14481,N_13783,N_13602);
nand U14482 (N_14482,N_13044,N_13035);
nand U14483 (N_14483,N_13891,N_13385);
xor U14484 (N_14484,N_13468,N_13630);
xor U14485 (N_14485,N_13532,N_13270);
xor U14486 (N_14486,N_13440,N_13931);
and U14487 (N_14487,N_13922,N_13745);
nand U14488 (N_14488,N_13707,N_13869);
and U14489 (N_14489,N_13363,N_13472);
nor U14490 (N_14490,N_13823,N_13475);
nor U14491 (N_14491,N_13550,N_13653);
and U14492 (N_14492,N_13377,N_13795);
or U14493 (N_14493,N_13605,N_13538);
and U14494 (N_14494,N_13929,N_13956);
and U14495 (N_14495,N_13664,N_13357);
nand U14496 (N_14496,N_13324,N_13847);
or U14497 (N_14497,N_13262,N_13635);
xor U14498 (N_14498,N_13335,N_13701);
nand U14499 (N_14499,N_13006,N_13732);
and U14500 (N_14500,N_13626,N_13608);
nand U14501 (N_14501,N_13110,N_13623);
nor U14502 (N_14502,N_13539,N_13425);
or U14503 (N_14503,N_13773,N_13919);
nor U14504 (N_14504,N_13658,N_13149);
or U14505 (N_14505,N_13778,N_13075);
and U14506 (N_14506,N_13358,N_13968);
xnor U14507 (N_14507,N_13384,N_13488);
xnor U14508 (N_14508,N_13716,N_13440);
xor U14509 (N_14509,N_13128,N_13351);
nand U14510 (N_14510,N_13305,N_13430);
xor U14511 (N_14511,N_13375,N_13526);
and U14512 (N_14512,N_13840,N_13280);
nor U14513 (N_14513,N_13940,N_13666);
xnor U14514 (N_14514,N_13137,N_13440);
and U14515 (N_14515,N_13004,N_13392);
and U14516 (N_14516,N_13101,N_13373);
nor U14517 (N_14517,N_13120,N_13213);
and U14518 (N_14518,N_13254,N_13507);
or U14519 (N_14519,N_13758,N_13411);
nor U14520 (N_14520,N_13045,N_13641);
nand U14521 (N_14521,N_13923,N_13520);
and U14522 (N_14522,N_13027,N_13527);
xor U14523 (N_14523,N_13117,N_13137);
and U14524 (N_14524,N_13013,N_13083);
nor U14525 (N_14525,N_13510,N_13151);
nor U14526 (N_14526,N_13246,N_13743);
xnor U14527 (N_14527,N_13061,N_13894);
and U14528 (N_14528,N_13457,N_13603);
nand U14529 (N_14529,N_13446,N_13648);
or U14530 (N_14530,N_13920,N_13288);
xor U14531 (N_14531,N_13866,N_13114);
nor U14532 (N_14532,N_13803,N_13787);
nand U14533 (N_14533,N_13617,N_13028);
or U14534 (N_14534,N_13027,N_13385);
xnor U14535 (N_14535,N_13027,N_13468);
nor U14536 (N_14536,N_13780,N_13144);
nand U14537 (N_14537,N_13755,N_13945);
nor U14538 (N_14538,N_13549,N_13292);
xor U14539 (N_14539,N_13848,N_13498);
nor U14540 (N_14540,N_13517,N_13550);
and U14541 (N_14541,N_13568,N_13038);
or U14542 (N_14542,N_13211,N_13812);
xnor U14543 (N_14543,N_13111,N_13554);
nand U14544 (N_14544,N_13764,N_13519);
nand U14545 (N_14545,N_13249,N_13518);
nand U14546 (N_14546,N_13782,N_13212);
or U14547 (N_14547,N_13692,N_13525);
and U14548 (N_14548,N_13747,N_13127);
and U14549 (N_14549,N_13375,N_13341);
and U14550 (N_14550,N_13575,N_13170);
nor U14551 (N_14551,N_13597,N_13550);
and U14552 (N_14552,N_13597,N_13152);
and U14553 (N_14553,N_13737,N_13319);
xor U14554 (N_14554,N_13868,N_13939);
and U14555 (N_14555,N_13833,N_13005);
and U14556 (N_14556,N_13087,N_13962);
nor U14557 (N_14557,N_13877,N_13692);
xnor U14558 (N_14558,N_13974,N_13470);
or U14559 (N_14559,N_13126,N_13301);
nor U14560 (N_14560,N_13092,N_13304);
xor U14561 (N_14561,N_13772,N_13682);
or U14562 (N_14562,N_13183,N_13109);
nor U14563 (N_14563,N_13823,N_13747);
nor U14564 (N_14564,N_13968,N_13759);
nor U14565 (N_14565,N_13413,N_13587);
nor U14566 (N_14566,N_13152,N_13364);
and U14567 (N_14567,N_13918,N_13178);
nand U14568 (N_14568,N_13736,N_13212);
and U14569 (N_14569,N_13753,N_13120);
nand U14570 (N_14570,N_13202,N_13482);
or U14571 (N_14571,N_13672,N_13733);
or U14572 (N_14572,N_13460,N_13771);
and U14573 (N_14573,N_13810,N_13596);
or U14574 (N_14574,N_13619,N_13150);
xor U14575 (N_14575,N_13519,N_13979);
or U14576 (N_14576,N_13885,N_13975);
or U14577 (N_14577,N_13907,N_13754);
or U14578 (N_14578,N_13845,N_13173);
nor U14579 (N_14579,N_13285,N_13822);
xnor U14580 (N_14580,N_13328,N_13264);
nor U14581 (N_14581,N_13592,N_13167);
nor U14582 (N_14582,N_13749,N_13338);
nand U14583 (N_14583,N_13072,N_13924);
or U14584 (N_14584,N_13030,N_13596);
and U14585 (N_14585,N_13737,N_13209);
and U14586 (N_14586,N_13926,N_13136);
and U14587 (N_14587,N_13975,N_13003);
xor U14588 (N_14588,N_13519,N_13060);
nand U14589 (N_14589,N_13243,N_13639);
nor U14590 (N_14590,N_13810,N_13993);
xnor U14591 (N_14591,N_13735,N_13449);
xor U14592 (N_14592,N_13496,N_13584);
nand U14593 (N_14593,N_13628,N_13763);
nor U14594 (N_14594,N_13917,N_13824);
nand U14595 (N_14595,N_13993,N_13406);
and U14596 (N_14596,N_13950,N_13953);
or U14597 (N_14597,N_13151,N_13354);
nor U14598 (N_14598,N_13911,N_13617);
or U14599 (N_14599,N_13099,N_13025);
nand U14600 (N_14600,N_13114,N_13488);
nor U14601 (N_14601,N_13714,N_13435);
xnor U14602 (N_14602,N_13552,N_13939);
xor U14603 (N_14603,N_13476,N_13892);
xnor U14604 (N_14604,N_13737,N_13188);
and U14605 (N_14605,N_13982,N_13525);
or U14606 (N_14606,N_13475,N_13957);
nand U14607 (N_14607,N_13740,N_13873);
nand U14608 (N_14608,N_13362,N_13504);
and U14609 (N_14609,N_13599,N_13089);
and U14610 (N_14610,N_13466,N_13395);
nor U14611 (N_14611,N_13570,N_13287);
xnor U14612 (N_14612,N_13641,N_13301);
nand U14613 (N_14613,N_13898,N_13787);
nand U14614 (N_14614,N_13509,N_13210);
xnor U14615 (N_14615,N_13215,N_13294);
nor U14616 (N_14616,N_13140,N_13856);
or U14617 (N_14617,N_13343,N_13357);
nor U14618 (N_14618,N_13746,N_13145);
nand U14619 (N_14619,N_13591,N_13726);
and U14620 (N_14620,N_13395,N_13886);
or U14621 (N_14621,N_13188,N_13714);
nand U14622 (N_14622,N_13553,N_13056);
nor U14623 (N_14623,N_13212,N_13977);
or U14624 (N_14624,N_13580,N_13667);
nor U14625 (N_14625,N_13401,N_13797);
nand U14626 (N_14626,N_13632,N_13932);
or U14627 (N_14627,N_13465,N_13981);
xor U14628 (N_14628,N_13270,N_13010);
nand U14629 (N_14629,N_13662,N_13699);
xor U14630 (N_14630,N_13716,N_13733);
or U14631 (N_14631,N_13813,N_13701);
nor U14632 (N_14632,N_13495,N_13628);
nor U14633 (N_14633,N_13828,N_13619);
nor U14634 (N_14634,N_13700,N_13160);
nor U14635 (N_14635,N_13173,N_13148);
nor U14636 (N_14636,N_13890,N_13255);
or U14637 (N_14637,N_13180,N_13344);
xor U14638 (N_14638,N_13846,N_13630);
and U14639 (N_14639,N_13637,N_13466);
and U14640 (N_14640,N_13228,N_13147);
nor U14641 (N_14641,N_13102,N_13394);
and U14642 (N_14642,N_13732,N_13363);
nor U14643 (N_14643,N_13857,N_13993);
nand U14644 (N_14644,N_13115,N_13130);
or U14645 (N_14645,N_13278,N_13557);
xnor U14646 (N_14646,N_13737,N_13283);
and U14647 (N_14647,N_13419,N_13003);
and U14648 (N_14648,N_13444,N_13903);
or U14649 (N_14649,N_13209,N_13597);
xnor U14650 (N_14650,N_13478,N_13018);
xnor U14651 (N_14651,N_13009,N_13555);
and U14652 (N_14652,N_13888,N_13330);
nand U14653 (N_14653,N_13814,N_13371);
nand U14654 (N_14654,N_13124,N_13893);
xor U14655 (N_14655,N_13263,N_13122);
or U14656 (N_14656,N_13206,N_13432);
nand U14657 (N_14657,N_13506,N_13049);
nand U14658 (N_14658,N_13267,N_13133);
and U14659 (N_14659,N_13429,N_13210);
xnor U14660 (N_14660,N_13546,N_13605);
nor U14661 (N_14661,N_13367,N_13923);
and U14662 (N_14662,N_13395,N_13966);
nand U14663 (N_14663,N_13330,N_13871);
or U14664 (N_14664,N_13747,N_13157);
nor U14665 (N_14665,N_13208,N_13067);
and U14666 (N_14666,N_13420,N_13720);
and U14667 (N_14667,N_13648,N_13426);
xnor U14668 (N_14668,N_13728,N_13987);
nand U14669 (N_14669,N_13289,N_13396);
or U14670 (N_14670,N_13686,N_13976);
xnor U14671 (N_14671,N_13124,N_13460);
nor U14672 (N_14672,N_13317,N_13723);
xnor U14673 (N_14673,N_13152,N_13227);
or U14674 (N_14674,N_13265,N_13745);
or U14675 (N_14675,N_13647,N_13214);
xnor U14676 (N_14676,N_13192,N_13786);
and U14677 (N_14677,N_13615,N_13070);
nor U14678 (N_14678,N_13820,N_13199);
xnor U14679 (N_14679,N_13329,N_13935);
xnor U14680 (N_14680,N_13097,N_13376);
xnor U14681 (N_14681,N_13499,N_13334);
xor U14682 (N_14682,N_13731,N_13607);
or U14683 (N_14683,N_13742,N_13501);
xnor U14684 (N_14684,N_13564,N_13124);
or U14685 (N_14685,N_13365,N_13881);
or U14686 (N_14686,N_13000,N_13665);
or U14687 (N_14687,N_13856,N_13311);
nand U14688 (N_14688,N_13897,N_13851);
nor U14689 (N_14689,N_13265,N_13528);
xnor U14690 (N_14690,N_13975,N_13655);
and U14691 (N_14691,N_13413,N_13321);
nor U14692 (N_14692,N_13849,N_13061);
nand U14693 (N_14693,N_13100,N_13484);
nor U14694 (N_14694,N_13785,N_13819);
or U14695 (N_14695,N_13198,N_13105);
nor U14696 (N_14696,N_13964,N_13998);
nor U14697 (N_14697,N_13828,N_13068);
nor U14698 (N_14698,N_13645,N_13320);
nor U14699 (N_14699,N_13115,N_13569);
nor U14700 (N_14700,N_13820,N_13934);
and U14701 (N_14701,N_13160,N_13401);
or U14702 (N_14702,N_13999,N_13878);
nand U14703 (N_14703,N_13991,N_13631);
and U14704 (N_14704,N_13834,N_13348);
or U14705 (N_14705,N_13753,N_13269);
or U14706 (N_14706,N_13149,N_13723);
xor U14707 (N_14707,N_13039,N_13231);
nor U14708 (N_14708,N_13824,N_13638);
xnor U14709 (N_14709,N_13269,N_13086);
nor U14710 (N_14710,N_13772,N_13149);
and U14711 (N_14711,N_13241,N_13682);
nor U14712 (N_14712,N_13508,N_13591);
and U14713 (N_14713,N_13025,N_13961);
and U14714 (N_14714,N_13857,N_13226);
or U14715 (N_14715,N_13888,N_13731);
xor U14716 (N_14716,N_13732,N_13688);
xor U14717 (N_14717,N_13801,N_13907);
or U14718 (N_14718,N_13660,N_13781);
nor U14719 (N_14719,N_13497,N_13511);
xnor U14720 (N_14720,N_13000,N_13620);
xnor U14721 (N_14721,N_13015,N_13600);
nor U14722 (N_14722,N_13946,N_13401);
nand U14723 (N_14723,N_13349,N_13172);
or U14724 (N_14724,N_13267,N_13922);
and U14725 (N_14725,N_13075,N_13472);
or U14726 (N_14726,N_13135,N_13788);
and U14727 (N_14727,N_13135,N_13011);
and U14728 (N_14728,N_13217,N_13619);
and U14729 (N_14729,N_13900,N_13814);
nor U14730 (N_14730,N_13062,N_13157);
or U14731 (N_14731,N_13110,N_13409);
and U14732 (N_14732,N_13384,N_13672);
nor U14733 (N_14733,N_13346,N_13713);
nand U14734 (N_14734,N_13573,N_13164);
nor U14735 (N_14735,N_13705,N_13433);
nand U14736 (N_14736,N_13126,N_13269);
nor U14737 (N_14737,N_13522,N_13704);
nor U14738 (N_14738,N_13236,N_13820);
xnor U14739 (N_14739,N_13147,N_13789);
xnor U14740 (N_14740,N_13967,N_13183);
xor U14741 (N_14741,N_13999,N_13183);
or U14742 (N_14742,N_13552,N_13831);
xnor U14743 (N_14743,N_13803,N_13815);
or U14744 (N_14744,N_13047,N_13141);
or U14745 (N_14745,N_13924,N_13558);
xor U14746 (N_14746,N_13039,N_13592);
or U14747 (N_14747,N_13454,N_13734);
and U14748 (N_14748,N_13628,N_13672);
and U14749 (N_14749,N_13100,N_13910);
xnor U14750 (N_14750,N_13856,N_13167);
or U14751 (N_14751,N_13981,N_13597);
and U14752 (N_14752,N_13393,N_13098);
nand U14753 (N_14753,N_13320,N_13751);
and U14754 (N_14754,N_13705,N_13132);
nand U14755 (N_14755,N_13982,N_13875);
nor U14756 (N_14756,N_13223,N_13789);
xor U14757 (N_14757,N_13932,N_13928);
nand U14758 (N_14758,N_13906,N_13895);
and U14759 (N_14759,N_13897,N_13827);
xnor U14760 (N_14760,N_13863,N_13664);
and U14761 (N_14761,N_13180,N_13538);
and U14762 (N_14762,N_13795,N_13331);
nor U14763 (N_14763,N_13209,N_13667);
nand U14764 (N_14764,N_13063,N_13226);
nand U14765 (N_14765,N_13004,N_13415);
xor U14766 (N_14766,N_13687,N_13134);
nor U14767 (N_14767,N_13442,N_13315);
nor U14768 (N_14768,N_13897,N_13591);
xor U14769 (N_14769,N_13833,N_13504);
xnor U14770 (N_14770,N_13357,N_13129);
and U14771 (N_14771,N_13232,N_13305);
or U14772 (N_14772,N_13958,N_13506);
nor U14773 (N_14773,N_13050,N_13860);
xnor U14774 (N_14774,N_13509,N_13414);
nor U14775 (N_14775,N_13931,N_13138);
and U14776 (N_14776,N_13483,N_13869);
or U14777 (N_14777,N_13873,N_13886);
xor U14778 (N_14778,N_13804,N_13566);
nand U14779 (N_14779,N_13015,N_13192);
or U14780 (N_14780,N_13474,N_13559);
xnor U14781 (N_14781,N_13274,N_13341);
and U14782 (N_14782,N_13930,N_13510);
xnor U14783 (N_14783,N_13136,N_13535);
and U14784 (N_14784,N_13916,N_13460);
or U14785 (N_14785,N_13285,N_13940);
xor U14786 (N_14786,N_13112,N_13131);
nor U14787 (N_14787,N_13377,N_13767);
and U14788 (N_14788,N_13145,N_13390);
xnor U14789 (N_14789,N_13376,N_13629);
nor U14790 (N_14790,N_13232,N_13206);
xor U14791 (N_14791,N_13827,N_13494);
or U14792 (N_14792,N_13052,N_13899);
xnor U14793 (N_14793,N_13192,N_13592);
nor U14794 (N_14794,N_13931,N_13585);
and U14795 (N_14795,N_13307,N_13976);
xor U14796 (N_14796,N_13133,N_13138);
xnor U14797 (N_14797,N_13633,N_13681);
nand U14798 (N_14798,N_13349,N_13263);
nor U14799 (N_14799,N_13638,N_13528);
nor U14800 (N_14800,N_13366,N_13956);
nand U14801 (N_14801,N_13552,N_13568);
nand U14802 (N_14802,N_13638,N_13094);
nor U14803 (N_14803,N_13525,N_13996);
nand U14804 (N_14804,N_13870,N_13167);
nor U14805 (N_14805,N_13749,N_13421);
and U14806 (N_14806,N_13004,N_13487);
and U14807 (N_14807,N_13042,N_13402);
nor U14808 (N_14808,N_13129,N_13376);
nor U14809 (N_14809,N_13140,N_13855);
xnor U14810 (N_14810,N_13208,N_13827);
nor U14811 (N_14811,N_13706,N_13419);
nor U14812 (N_14812,N_13779,N_13008);
or U14813 (N_14813,N_13769,N_13448);
or U14814 (N_14814,N_13967,N_13502);
nor U14815 (N_14815,N_13510,N_13612);
nor U14816 (N_14816,N_13165,N_13843);
or U14817 (N_14817,N_13791,N_13778);
nor U14818 (N_14818,N_13770,N_13804);
nand U14819 (N_14819,N_13089,N_13137);
or U14820 (N_14820,N_13645,N_13618);
nand U14821 (N_14821,N_13173,N_13537);
and U14822 (N_14822,N_13967,N_13442);
nand U14823 (N_14823,N_13024,N_13727);
and U14824 (N_14824,N_13315,N_13945);
xor U14825 (N_14825,N_13847,N_13077);
nor U14826 (N_14826,N_13350,N_13717);
nand U14827 (N_14827,N_13114,N_13884);
xnor U14828 (N_14828,N_13993,N_13564);
or U14829 (N_14829,N_13070,N_13308);
nor U14830 (N_14830,N_13077,N_13136);
nor U14831 (N_14831,N_13046,N_13735);
and U14832 (N_14832,N_13711,N_13442);
nand U14833 (N_14833,N_13990,N_13314);
xnor U14834 (N_14834,N_13528,N_13724);
and U14835 (N_14835,N_13446,N_13247);
and U14836 (N_14836,N_13326,N_13075);
nand U14837 (N_14837,N_13525,N_13020);
nor U14838 (N_14838,N_13158,N_13095);
and U14839 (N_14839,N_13352,N_13661);
nand U14840 (N_14840,N_13751,N_13133);
nor U14841 (N_14841,N_13426,N_13675);
or U14842 (N_14842,N_13301,N_13282);
or U14843 (N_14843,N_13211,N_13772);
xnor U14844 (N_14844,N_13944,N_13857);
xnor U14845 (N_14845,N_13767,N_13902);
nor U14846 (N_14846,N_13674,N_13947);
nor U14847 (N_14847,N_13966,N_13398);
nor U14848 (N_14848,N_13660,N_13446);
or U14849 (N_14849,N_13302,N_13548);
nand U14850 (N_14850,N_13332,N_13354);
or U14851 (N_14851,N_13023,N_13337);
nand U14852 (N_14852,N_13680,N_13113);
or U14853 (N_14853,N_13615,N_13074);
and U14854 (N_14854,N_13858,N_13155);
and U14855 (N_14855,N_13123,N_13121);
nand U14856 (N_14856,N_13765,N_13857);
nand U14857 (N_14857,N_13705,N_13524);
or U14858 (N_14858,N_13337,N_13671);
or U14859 (N_14859,N_13792,N_13230);
and U14860 (N_14860,N_13335,N_13018);
xor U14861 (N_14861,N_13466,N_13381);
nand U14862 (N_14862,N_13804,N_13570);
xor U14863 (N_14863,N_13387,N_13205);
nand U14864 (N_14864,N_13832,N_13728);
or U14865 (N_14865,N_13170,N_13100);
and U14866 (N_14866,N_13869,N_13046);
nand U14867 (N_14867,N_13682,N_13728);
or U14868 (N_14868,N_13680,N_13273);
nor U14869 (N_14869,N_13356,N_13226);
nand U14870 (N_14870,N_13883,N_13726);
nor U14871 (N_14871,N_13080,N_13936);
or U14872 (N_14872,N_13939,N_13726);
nand U14873 (N_14873,N_13523,N_13656);
and U14874 (N_14874,N_13176,N_13052);
xor U14875 (N_14875,N_13584,N_13463);
nor U14876 (N_14876,N_13458,N_13572);
xnor U14877 (N_14877,N_13843,N_13274);
and U14878 (N_14878,N_13989,N_13724);
and U14879 (N_14879,N_13180,N_13728);
nor U14880 (N_14880,N_13871,N_13947);
nand U14881 (N_14881,N_13462,N_13678);
xor U14882 (N_14882,N_13379,N_13949);
nand U14883 (N_14883,N_13958,N_13837);
and U14884 (N_14884,N_13278,N_13400);
nand U14885 (N_14885,N_13826,N_13456);
and U14886 (N_14886,N_13075,N_13779);
xnor U14887 (N_14887,N_13122,N_13657);
and U14888 (N_14888,N_13973,N_13098);
or U14889 (N_14889,N_13400,N_13630);
and U14890 (N_14890,N_13101,N_13077);
xnor U14891 (N_14891,N_13856,N_13973);
nand U14892 (N_14892,N_13771,N_13547);
nand U14893 (N_14893,N_13961,N_13153);
xor U14894 (N_14894,N_13992,N_13923);
and U14895 (N_14895,N_13144,N_13782);
and U14896 (N_14896,N_13266,N_13955);
or U14897 (N_14897,N_13179,N_13043);
nand U14898 (N_14898,N_13392,N_13681);
nor U14899 (N_14899,N_13423,N_13307);
nor U14900 (N_14900,N_13053,N_13375);
or U14901 (N_14901,N_13183,N_13023);
nand U14902 (N_14902,N_13156,N_13721);
nand U14903 (N_14903,N_13447,N_13539);
nor U14904 (N_14904,N_13057,N_13804);
xor U14905 (N_14905,N_13512,N_13910);
nand U14906 (N_14906,N_13646,N_13811);
and U14907 (N_14907,N_13648,N_13296);
and U14908 (N_14908,N_13415,N_13156);
nand U14909 (N_14909,N_13247,N_13595);
or U14910 (N_14910,N_13719,N_13401);
nor U14911 (N_14911,N_13883,N_13894);
or U14912 (N_14912,N_13733,N_13276);
nor U14913 (N_14913,N_13922,N_13886);
nor U14914 (N_14914,N_13637,N_13005);
xor U14915 (N_14915,N_13367,N_13347);
nor U14916 (N_14916,N_13262,N_13055);
and U14917 (N_14917,N_13809,N_13264);
xnor U14918 (N_14918,N_13354,N_13404);
nor U14919 (N_14919,N_13286,N_13685);
and U14920 (N_14920,N_13915,N_13446);
or U14921 (N_14921,N_13532,N_13613);
nand U14922 (N_14922,N_13746,N_13834);
nand U14923 (N_14923,N_13976,N_13032);
nand U14924 (N_14924,N_13145,N_13014);
and U14925 (N_14925,N_13146,N_13278);
nand U14926 (N_14926,N_13567,N_13182);
or U14927 (N_14927,N_13335,N_13545);
xnor U14928 (N_14928,N_13699,N_13951);
and U14929 (N_14929,N_13677,N_13577);
xor U14930 (N_14930,N_13535,N_13183);
nand U14931 (N_14931,N_13267,N_13695);
and U14932 (N_14932,N_13787,N_13741);
nor U14933 (N_14933,N_13280,N_13260);
nand U14934 (N_14934,N_13337,N_13626);
nand U14935 (N_14935,N_13970,N_13877);
and U14936 (N_14936,N_13665,N_13284);
or U14937 (N_14937,N_13055,N_13957);
nand U14938 (N_14938,N_13533,N_13040);
or U14939 (N_14939,N_13983,N_13332);
and U14940 (N_14940,N_13395,N_13457);
nand U14941 (N_14941,N_13398,N_13730);
nor U14942 (N_14942,N_13900,N_13625);
xnor U14943 (N_14943,N_13582,N_13783);
xnor U14944 (N_14944,N_13357,N_13062);
and U14945 (N_14945,N_13145,N_13462);
nand U14946 (N_14946,N_13135,N_13512);
nor U14947 (N_14947,N_13451,N_13719);
xor U14948 (N_14948,N_13316,N_13379);
or U14949 (N_14949,N_13717,N_13973);
nor U14950 (N_14950,N_13719,N_13437);
xnor U14951 (N_14951,N_13191,N_13413);
and U14952 (N_14952,N_13844,N_13568);
nor U14953 (N_14953,N_13407,N_13588);
nor U14954 (N_14954,N_13395,N_13866);
nor U14955 (N_14955,N_13984,N_13358);
and U14956 (N_14956,N_13975,N_13601);
and U14957 (N_14957,N_13129,N_13190);
or U14958 (N_14958,N_13820,N_13139);
or U14959 (N_14959,N_13747,N_13803);
or U14960 (N_14960,N_13070,N_13044);
nand U14961 (N_14961,N_13314,N_13367);
and U14962 (N_14962,N_13346,N_13187);
nand U14963 (N_14963,N_13945,N_13775);
or U14964 (N_14964,N_13470,N_13932);
nand U14965 (N_14965,N_13479,N_13163);
nand U14966 (N_14966,N_13346,N_13011);
nand U14967 (N_14967,N_13865,N_13751);
xnor U14968 (N_14968,N_13666,N_13200);
nor U14969 (N_14969,N_13381,N_13063);
nor U14970 (N_14970,N_13870,N_13039);
nand U14971 (N_14971,N_13641,N_13227);
nor U14972 (N_14972,N_13289,N_13640);
xnor U14973 (N_14973,N_13029,N_13950);
nor U14974 (N_14974,N_13461,N_13377);
xnor U14975 (N_14975,N_13628,N_13303);
or U14976 (N_14976,N_13636,N_13564);
xnor U14977 (N_14977,N_13597,N_13540);
nand U14978 (N_14978,N_13858,N_13692);
or U14979 (N_14979,N_13318,N_13641);
nor U14980 (N_14980,N_13511,N_13896);
nor U14981 (N_14981,N_13992,N_13464);
xor U14982 (N_14982,N_13116,N_13495);
nand U14983 (N_14983,N_13644,N_13411);
nand U14984 (N_14984,N_13091,N_13265);
nand U14985 (N_14985,N_13091,N_13006);
nor U14986 (N_14986,N_13940,N_13039);
and U14987 (N_14987,N_13551,N_13774);
nor U14988 (N_14988,N_13197,N_13443);
xnor U14989 (N_14989,N_13312,N_13904);
or U14990 (N_14990,N_13565,N_13662);
and U14991 (N_14991,N_13737,N_13652);
nand U14992 (N_14992,N_13947,N_13465);
and U14993 (N_14993,N_13622,N_13679);
or U14994 (N_14994,N_13396,N_13262);
xnor U14995 (N_14995,N_13467,N_13960);
nor U14996 (N_14996,N_13587,N_13940);
xor U14997 (N_14997,N_13027,N_13925);
xnor U14998 (N_14998,N_13895,N_13311);
and U14999 (N_14999,N_13206,N_13810);
xnor U15000 (N_15000,N_14577,N_14763);
or U15001 (N_15001,N_14775,N_14150);
xnor U15002 (N_15002,N_14981,N_14537);
and U15003 (N_15003,N_14183,N_14691);
nand U15004 (N_15004,N_14166,N_14969);
nor U15005 (N_15005,N_14097,N_14890);
and U15006 (N_15006,N_14787,N_14870);
xor U15007 (N_15007,N_14606,N_14370);
xnor U15008 (N_15008,N_14622,N_14340);
nand U15009 (N_15009,N_14324,N_14955);
and U15010 (N_15010,N_14589,N_14611);
nand U15011 (N_15011,N_14125,N_14842);
and U15012 (N_15012,N_14313,N_14274);
xor U15013 (N_15013,N_14235,N_14396);
or U15014 (N_15014,N_14701,N_14090);
or U15015 (N_15015,N_14619,N_14655);
nand U15016 (N_15016,N_14908,N_14957);
nand U15017 (N_15017,N_14586,N_14584);
nand U15018 (N_15018,N_14251,N_14751);
xnor U15019 (N_15019,N_14364,N_14839);
nand U15020 (N_15020,N_14989,N_14788);
or U15021 (N_15021,N_14774,N_14224);
or U15022 (N_15022,N_14412,N_14781);
nor U15023 (N_15023,N_14757,N_14769);
and U15024 (N_15024,N_14050,N_14399);
and U15025 (N_15025,N_14026,N_14209);
nor U15026 (N_15026,N_14003,N_14398);
or U15027 (N_15027,N_14850,N_14108);
nor U15028 (N_15028,N_14938,N_14545);
or U15029 (N_15029,N_14871,N_14880);
and U15030 (N_15030,N_14185,N_14151);
or U15031 (N_15031,N_14401,N_14335);
or U15032 (N_15032,N_14178,N_14266);
and U15033 (N_15033,N_14264,N_14698);
nor U15034 (N_15034,N_14749,N_14427);
or U15035 (N_15035,N_14591,N_14991);
nand U15036 (N_15036,N_14466,N_14675);
xor U15037 (N_15037,N_14269,N_14136);
nor U15038 (N_15038,N_14789,N_14400);
nor U15039 (N_15039,N_14948,N_14336);
nor U15040 (N_15040,N_14806,N_14208);
xnor U15041 (N_15041,N_14230,N_14270);
and U15042 (N_15042,N_14629,N_14404);
xnor U15043 (N_15043,N_14359,N_14999);
or U15044 (N_15044,N_14276,N_14565);
and U15045 (N_15045,N_14343,N_14099);
xor U15046 (N_15046,N_14403,N_14608);
nand U15047 (N_15047,N_14295,N_14685);
nor U15048 (N_15048,N_14961,N_14258);
xor U15049 (N_15049,N_14283,N_14570);
xor U15050 (N_15050,N_14993,N_14538);
nand U15051 (N_15051,N_14587,N_14502);
or U15052 (N_15052,N_14816,N_14501);
and U15053 (N_15053,N_14539,N_14883);
and U15054 (N_15054,N_14508,N_14817);
nand U15055 (N_15055,N_14992,N_14031);
xor U15056 (N_15056,N_14020,N_14238);
nor U15057 (N_15057,N_14059,N_14953);
and U15058 (N_15058,N_14014,N_14366);
and U15059 (N_15059,N_14225,N_14511);
or U15060 (N_15060,N_14024,N_14673);
or U15061 (N_15061,N_14793,N_14437);
xnor U15062 (N_15062,N_14474,N_14909);
and U15063 (N_15063,N_14686,N_14068);
nand U15064 (N_15064,N_14895,N_14277);
and U15065 (N_15065,N_14557,N_14203);
nand U15066 (N_15066,N_14206,N_14833);
nor U15067 (N_15067,N_14598,N_14709);
or U15068 (N_15068,N_14055,N_14137);
nand U15069 (N_15069,N_14845,N_14947);
and U15070 (N_15070,N_14113,N_14245);
xor U15071 (N_15071,N_14844,N_14350);
and U15072 (N_15072,N_14797,N_14296);
and U15073 (N_15073,N_14504,N_14541);
nand U15074 (N_15074,N_14796,N_14865);
xnor U15075 (N_15075,N_14741,N_14637);
or U15076 (N_15076,N_14906,N_14426);
or U15077 (N_15077,N_14188,N_14920);
xor U15078 (N_15078,N_14728,N_14980);
and U15079 (N_15079,N_14123,N_14771);
and U15080 (N_15080,N_14243,N_14919);
nand U15081 (N_15081,N_14424,N_14913);
nor U15082 (N_15082,N_14451,N_14391);
or U15083 (N_15083,N_14814,N_14857);
nor U15084 (N_15084,N_14580,N_14450);
or U15085 (N_15085,N_14627,N_14832);
nand U15086 (N_15086,N_14928,N_14661);
xor U15087 (N_15087,N_14569,N_14975);
nand U15088 (N_15088,N_14599,N_14660);
xor U15089 (N_15089,N_14516,N_14896);
nand U15090 (N_15090,N_14601,N_14885);
and U15091 (N_15091,N_14902,N_14439);
or U15092 (N_15092,N_14776,N_14218);
nand U15093 (N_15093,N_14679,N_14231);
or U15094 (N_15094,N_14745,N_14233);
xor U15095 (N_15095,N_14915,N_14659);
nand U15096 (N_15096,N_14965,N_14668);
nor U15097 (N_15097,N_14051,N_14517);
nand U15098 (N_15098,N_14272,N_14509);
nand U15099 (N_15099,N_14176,N_14593);
nor U15100 (N_15100,N_14316,N_14973);
and U15101 (N_15101,N_14874,N_14070);
and U15102 (N_15102,N_14917,N_14220);
and U15103 (N_15103,N_14344,N_14049);
or U15104 (N_15104,N_14597,N_14294);
nor U15105 (N_15105,N_14899,N_14469);
or U15106 (N_15106,N_14669,N_14664);
nor U15107 (N_15107,N_14574,N_14280);
xor U15108 (N_15108,N_14066,N_14760);
xnor U15109 (N_15109,N_14872,N_14009);
or U15110 (N_15110,N_14595,N_14354);
or U15111 (N_15111,N_14889,N_14513);
nand U15112 (N_15112,N_14162,N_14618);
nor U15113 (N_15113,N_14607,N_14782);
nand U15114 (N_15114,N_14950,N_14645);
xnor U15115 (N_15115,N_14397,N_14860);
and U15116 (N_15116,N_14080,N_14624);
or U15117 (N_15117,N_14374,N_14442);
xor U15118 (N_15118,N_14304,N_14954);
or U15119 (N_15119,N_14575,N_14143);
nor U15120 (N_15120,N_14652,N_14468);
or U15121 (N_15121,N_14930,N_14657);
nand U15122 (N_15122,N_14293,N_14485);
nand U15123 (N_15123,N_14968,N_14402);
nand U15124 (N_15124,N_14520,N_14353);
and U15125 (N_15125,N_14951,N_14002);
and U15126 (N_15126,N_14138,N_14772);
xnor U15127 (N_15127,N_14376,N_14383);
nand U15128 (N_15128,N_14356,N_14102);
and U15129 (N_15129,N_14228,N_14423);
nor U15130 (N_15130,N_14484,N_14388);
nor U15131 (N_15131,N_14467,N_14907);
xor U15132 (N_15132,N_14351,N_14210);
and U15133 (N_15133,N_14363,N_14854);
xnor U15134 (N_15134,N_14255,N_14482);
and U15135 (N_15135,N_14445,N_14674);
and U15136 (N_15136,N_14145,N_14934);
nor U15137 (N_15137,N_14931,N_14180);
xor U15138 (N_15138,N_14711,N_14916);
nand U15139 (N_15139,N_14804,N_14984);
and U15140 (N_15140,N_14253,N_14381);
or U15141 (N_15141,N_14834,N_14933);
and U15142 (N_15142,N_14358,N_14382);
nor U15143 (N_15143,N_14091,N_14963);
or U15144 (N_15144,N_14721,N_14654);
nor U15145 (N_15145,N_14229,N_14643);
xnor U15146 (N_15146,N_14519,N_14135);
or U15147 (N_15147,N_14415,N_14084);
xor U15148 (N_15148,N_14670,N_14753);
or U15149 (N_15149,N_14128,N_14744);
xor U15150 (N_15150,N_14488,N_14186);
xnor U15151 (N_15151,N_14572,N_14446);
and U15152 (N_15152,N_14073,N_14853);
nand U15153 (N_15153,N_14472,N_14811);
nor U15154 (N_15154,N_14800,N_14329);
and U15155 (N_15155,N_14495,N_14406);
or U15156 (N_15156,N_14801,N_14241);
nand U15157 (N_15157,N_14115,N_14704);
xor U15158 (N_15158,N_14805,N_14822);
nand U15159 (N_15159,N_14200,N_14820);
xnor U15160 (N_15160,N_14785,N_14886);
and U15161 (N_15161,N_14368,N_14418);
or U15162 (N_15162,N_14809,N_14723);
and U15163 (N_15163,N_14286,N_14944);
or U15164 (N_15164,N_14199,N_14167);
or U15165 (N_15165,N_14856,N_14473);
or U15166 (N_15166,N_14430,N_14148);
nor U15167 (N_15167,N_14677,N_14434);
nand U15168 (N_15168,N_14958,N_14144);
and U15169 (N_15169,N_14579,N_14734);
xnor U15170 (N_15170,N_14616,N_14935);
nor U15171 (N_15171,N_14288,N_14433);
nor U15172 (N_15172,N_14553,N_14825);
nor U15173 (N_15173,N_14332,N_14682);
nor U15174 (N_15174,N_14267,N_14551);
xor U15175 (N_15175,N_14710,N_14464);
nand U15176 (N_15176,N_14048,N_14175);
and U15177 (N_15177,N_14492,N_14649);
and U15178 (N_15178,N_14232,N_14821);
or U15179 (N_15179,N_14985,N_14526);
nor U15180 (N_15180,N_14481,N_14337);
or U15181 (N_15181,N_14559,N_14858);
nand U15182 (N_15182,N_14515,N_14561);
nor U15183 (N_15183,N_14360,N_14006);
or U15184 (N_15184,N_14912,N_14667);
nor U15185 (N_15185,N_14592,N_14945);
nor U15186 (N_15186,N_14892,N_14375);
xor U15187 (N_15187,N_14695,N_14982);
xnor U15188 (N_15188,N_14927,N_14847);
and U15189 (N_15189,N_14217,N_14072);
or U15190 (N_15190,N_14191,N_14187);
xnor U15191 (N_15191,N_14813,N_14583);
xnor U15192 (N_15192,N_14325,N_14555);
and U15193 (N_15193,N_14321,N_14155);
or U15194 (N_15194,N_14803,N_14349);
xnor U15195 (N_15195,N_14019,N_14285);
nor U15196 (N_15196,N_14204,N_14315);
nand U15197 (N_15197,N_14271,N_14477);
nand U15198 (N_15198,N_14452,N_14635);
nand U15199 (N_15199,N_14065,N_14490);
nand U15200 (N_15200,N_14621,N_14921);
or U15201 (N_15201,N_14234,N_14071);
nand U15202 (N_15202,N_14112,N_14052);
nand U15203 (N_15203,N_14612,N_14389);
nor U15204 (N_15204,N_14139,N_14491);
nor U15205 (N_15205,N_14518,N_14613);
or U15206 (N_15206,N_14314,N_14904);
and U15207 (N_15207,N_14680,N_14303);
and U15208 (N_15208,N_14829,N_14761);
or U15209 (N_15209,N_14505,N_14609);
or U15210 (N_15210,N_14159,N_14998);
and U15211 (N_15211,N_14897,N_14205);
nor U15212 (N_15212,N_14197,N_14465);
xnor U15213 (N_15213,N_14893,N_14960);
and U15214 (N_15214,N_14265,N_14838);
and U15215 (N_15215,N_14222,N_14348);
and U15216 (N_15216,N_14798,N_14039);
nor U15217 (N_15217,N_14639,N_14733);
nor U15218 (N_15218,N_14170,N_14507);
and U15219 (N_15219,N_14700,N_14417);
nor U15220 (N_15220,N_14578,N_14207);
or U15221 (N_15221,N_14731,N_14770);
and U15222 (N_15222,N_14367,N_14715);
nand U15223 (N_15223,N_14300,N_14929);
and U15224 (N_15224,N_14305,N_14021);
nand U15225 (N_15225,N_14863,N_14964);
nand U15226 (N_15226,N_14281,N_14489);
xor U15227 (N_15227,N_14076,N_14263);
and U15228 (N_15228,N_14740,N_14487);
nand U15229 (N_15229,N_14808,N_14617);
and U15230 (N_15230,N_14932,N_14610);
and U15231 (N_15231,N_14441,N_14540);
and U15232 (N_15232,N_14497,N_14543);
xnor U15233 (N_15233,N_14848,N_14646);
or U15234 (N_15234,N_14626,N_14096);
nor U15235 (N_15235,N_14550,N_14792);
nor U15236 (N_15236,N_14330,N_14837);
and U15237 (N_15237,N_14869,N_14802);
and U15238 (N_15238,N_14810,N_14385);
nor U15239 (N_15239,N_14878,N_14328);
and U15240 (N_15240,N_14596,N_14449);
xnor U15241 (N_15241,N_14082,N_14949);
or U15242 (N_15242,N_14987,N_14133);
xor U15243 (N_15243,N_14086,N_14498);
nor U15244 (N_15244,N_14160,N_14239);
and U15245 (N_15245,N_14215,N_14393);
and U15246 (N_15246,N_14877,N_14289);
or U15247 (N_15247,N_14131,N_14098);
nor U15248 (N_15248,N_14005,N_14118);
nor U15249 (N_15249,N_14346,N_14812);
nand U15250 (N_15250,N_14712,N_14830);
and U15251 (N_15251,N_14693,N_14983);
or U15252 (N_15252,N_14739,N_14996);
nand U15253 (N_15253,N_14341,N_14632);
and U15254 (N_15254,N_14422,N_14292);
and U15255 (N_15255,N_14764,N_14807);
or U15256 (N_15256,N_14369,N_14355);
or U15257 (N_15257,N_14320,N_14053);
or U15258 (N_15258,N_14758,N_14500);
nand U15259 (N_15259,N_14784,N_14372);
or U15260 (N_15260,N_14824,N_14081);
xor U15261 (N_15261,N_14476,N_14903);
and U15262 (N_15262,N_14549,N_14891);
xor U15263 (N_15263,N_14408,N_14684);
and U15264 (N_15264,N_14202,N_14773);
nand U15265 (N_15265,N_14212,N_14478);
nand U15266 (N_15266,N_14994,N_14568);
nand U15267 (N_15267,N_14132,N_14022);
and U15268 (N_15268,N_14158,N_14729);
and U15269 (N_15269,N_14326,N_14563);
nor U15270 (N_15270,N_14730,N_14881);
nand U15271 (N_15271,N_14706,N_14377);
xnor U15272 (N_15272,N_14530,N_14640);
nor U15273 (N_15273,N_14547,N_14861);
and U15274 (N_15274,N_14614,N_14479);
and U15275 (N_15275,N_14995,N_14588);
nor U15276 (N_15276,N_14074,N_14117);
or U15277 (N_15277,N_14783,N_14017);
xnor U15278 (N_15278,N_14297,N_14259);
or U15279 (N_15279,N_14536,N_14552);
or U15280 (N_15280,N_14748,N_14566);
nor U15281 (N_15281,N_14436,N_14528);
and U15282 (N_15282,N_14767,N_14378);
or U15283 (N_15283,N_14154,N_14088);
xnor U15284 (N_15284,N_14105,N_14153);
or U15285 (N_15285,N_14110,N_14725);
nand U15286 (N_15286,N_14103,N_14647);
nand U15287 (N_15287,N_14717,N_14008);
nor U15288 (N_15288,N_14826,N_14615);
or U15289 (N_15289,N_14959,N_14460);
xor U15290 (N_15290,N_14683,N_14431);
and U15291 (N_15291,N_14699,N_14855);
nand U15292 (N_15292,N_14004,N_14339);
nor U15293 (N_15293,N_14361,N_14390);
xor U15294 (N_15294,N_14195,N_14425);
xor U15295 (N_15295,N_14936,N_14713);
xnor U15296 (N_15296,N_14278,N_14282);
xor U15297 (N_15297,N_14054,N_14171);
or U15298 (N_15298,N_14828,N_14970);
nand U15299 (N_15299,N_14688,N_14768);
nand U15300 (N_15300,N_14815,N_14001);
and U15301 (N_15301,N_14556,N_14142);
nand U15302 (N_15302,N_14317,N_14835);
nand U15303 (N_15303,N_14689,N_14444);
nand U15304 (N_15304,N_14237,N_14496);
nand U15305 (N_15305,N_14571,N_14514);
nor U15306 (N_15306,N_14666,N_14100);
nand U15307 (N_15307,N_14058,N_14213);
nand U15308 (N_15308,N_14190,N_14978);
and U15309 (N_15309,N_14236,N_14122);
nand U15310 (N_15310,N_14146,N_14535);
nand U15311 (N_15311,N_14750,N_14106);
and U15312 (N_15312,N_14040,N_14141);
nand U15313 (N_15313,N_14067,N_14119);
nand U15314 (N_15314,N_14057,N_14095);
xnor U15315 (N_15315,N_14419,N_14777);
or U15316 (N_15316,N_14077,N_14345);
or U15317 (N_15317,N_14905,N_14174);
xor U15318 (N_15318,N_14562,N_14576);
or U15319 (N_15319,N_14172,N_14311);
nor U15320 (N_15320,N_14720,N_14416);
nand U15321 (N_15321,N_14494,N_14193);
nand U15322 (N_15322,N_14028,N_14475);
nor U15323 (N_15323,N_14018,N_14448);
and U15324 (N_15324,N_14653,N_14988);
or U15325 (N_15325,N_14087,N_14184);
and U15326 (N_15326,N_14503,N_14823);
nand U15327 (N_15327,N_14116,N_14911);
xnor U15328 (N_15328,N_14631,N_14149);
xor U15329 (N_15329,N_14273,N_14602);
nand U15330 (N_15330,N_14457,N_14062);
nor U15331 (N_15331,N_14083,N_14884);
or U15332 (N_15332,N_14638,N_14323);
nor U15333 (N_15333,N_14221,N_14510);
nand U15334 (N_15334,N_14037,N_14275);
nor U15335 (N_15335,N_14879,N_14795);
nand U15336 (N_15336,N_14952,N_14512);
xor U15337 (N_15337,N_14990,N_14290);
and U15338 (N_15338,N_14025,N_14279);
or U15339 (N_15339,N_14859,N_14333);
xor U15340 (N_15340,N_14976,N_14651);
and U15341 (N_15341,N_14152,N_14681);
nor U15342 (N_15342,N_14078,N_14016);
nand U15343 (N_15343,N_14027,N_14214);
and U15344 (N_15344,N_14979,N_14094);
xor U15345 (N_15345,N_14521,N_14093);
and U15346 (N_15346,N_14582,N_14898);
xnor U15347 (N_15347,N_14762,N_14522);
and U15348 (N_15348,N_14173,N_14227);
and U15349 (N_15349,N_14943,N_14240);
or U15350 (N_15350,N_14922,N_14414);
and U15351 (N_15351,N_14506,N_14244);
nor U15352 (N_15352,N_14157,N_14379);
xor U15353 (N_15353,N_14179,N_14705);
nor U15354 (N_15354,N_14127,N_14558);
nand U15355 (N_15355,N_14888,N_14453);
nor U15356 (N_15356,N_14261,N_14941);
and U15357 (N_15357,N_14529,N_14900);
or U15358 (N_15358,N_14322,N_14676);
nor U15359 (N_15359,N_14046,N_14605);
xor U15360 (N_15360,N_14129,N_14696);
or U15361 (N_15361,N_14818,N_14420);
nor U15362 (N_15362,N_14851,N_14038);
and U15363 (N_15363,N_14428,N_14334);
nor U15364 (N_15364,N_14169,N_14780);
nand U15365 (N_15365,N_14407,N_14480);
and U15366 (N_15366,N_14738,N_14254);
xor U15367 (N_15367,N_14962,N_14924);
or U15368 (N_15368,N_14534,N_14268);
xor U15369 (N_15369,N_14023,N_14940);
nand U15370 (N_15370,N_14779,N_14794);
nor U15371 (N_15371,N_14752,N_14971);
and U15372 (N_15372,N_14918,N_14035);
and U15373 (N_15373,N_14581,N_14743);
or U15374 (N_15374,N_14849,N_14386);
nand U15375 (N_15375,N_14542,N_14164);
nor U15376 (N_15376,N_14216,N_14318);
nor U15377 (N_15377,N_14926,N_14628);
nor U15378 (N_15378,N_14168,N_14189);
xor U15379 (N_15379,N_14047,N_14650);
nor U15380 (N_15380,N_14470,N_14876);
nor U15381 (N_15381,N_14032,N_14260);
nand U15382 (N_15382,N_14124,N_14778);
or U15383 (N_15383,N_14548,N_14015);
nand U15384 (N_15384,N_14567,N_14085);
nand U15385 (N_15385,N_14942,N_14755);
and U15386 (N_15386,N_14732,N_14302);
nand U15387 (N_15387,N_14625,N_14182);
xor U15388 (N_15388,N_14636,N_14373);
and U15389 (N_15389,N_14714,N_14063);
xnor U15390 (N_15390,N_14012,N_14013);
nor U15391 (N_15391,N_14707,N_14246);
nor U15392 (N_15392,N_14658,N_14690);
nor U15393 (N_15393,N_14045,N_14923);
and U15394 (N_15394,N_14347,N_14827);
nand U15395 (N_15395,N_14410,N_14447);
and U15396 (N_15396,N_14946,N_14440);
and U15397 (N_15397,N_14306,N_14413);
xor U15398 (N_15398,N_14527,N_14977);
nor U15399 (N_15399,N_14868,N_14737);
and U15400 (N_15400,N_14836,N_14546);
nor U15401 (N_15401,N_14463,N_14533);
and U15402 (N_15402,N_14034,N_14791);
xor U15403 (N_15403,N_14287,N_14121);
or U15404 (N_15404,N_14727,N_14443);
nor U15405 (N_15405,N_14831,N_14043);
nand U15406 (N_15406,N_14064,N_14252);
xnor U15407 (N_15407,N_14130,N_14365);
and U15408 (N_15408,N_14724,N_14882);
xnor U15409 (N_15409,N_14114,N_14662);
or U15410 (N_15410,N_14307,N_14310);
or U15411 (N_15411,N_14722,N_14411);
nor U15412 (N_15412,N_14493,N_14641);
or U15413 (N_15413,N_14697,N_14873);
nand U15414 (N_15414,N_14846,N_14703);
nand U15415 (N_15415,N_14060,N_14387);
and U15416 (N_15416,N_14937,N_14248);
or U15417 (N_15417,N_14716,N_14692);
nor U15418 (N_15418,N_14041,N_14997);
nand U15419 (N_15419,N_14371,N_14841);
xor U15420 (N_15420,N_14455,N_14967);
xnor U15421 (N_15421,N_14181,N_14765);
nand U15422 (N_15422,N_14069,N_14630);
xnor U15423 (N_15423,N_14986,N_14875);
and U15424 (N_15424,N_14454,N_14177);
nor U15425 (N_15425,N_14198,N_14623);
nor U15426 (N_15426,N_14421,N_14790);
nor U15427 (N_15427,N_14438,N_14042);
or U15428 (N_15428,N_14107,N_14291);
and U15429 (N_15429,N_14362,N_14432);
nand U15430 (N_15430,N_14862,N_14678);
xor U15431 (N_15431,N_14554,N_14840);
nor U15432 (N_15432,N_14380,N_14766);
nor U15433 (N_15433,N_14726,N_14544);
or U15434 (N_15434,N_14201,N_14901);
and U15435 (N_15435,N_14395,N_14357);
nor U15436 (N_15436,N_14120,N_14799);
xor U15437 (N_15437,N_14910,N_14165);
xor U15438 (N_15438,N_14163,N_14392);
nand U15439 (N_15439,N_14192,N_14011);
xor U15440 (N_15440,N_14458,N_14089);
and U15441 (N_15441,N_14298,N_14687);
or U15442 (N_15442,N_14161,N_14914);
and U15443 (N_15443,N_14754,N_14342);
or U15444 (N_15444,N_14648,N_14247);
nand U15445 (N_15445,N_14079,N_14663);
nand U15446 (N_15446,N_14759,N_14887);
and U15447 (N_15447,N_14603,N_14974);
or U15448 (N_15448,N_14718,N_14532);
nor U15449 (N_15449,N_14429,N_14249);
nor U15450 (N_15450,N_14708,N_14327);
nor U15451 (N_15451,N_14262,N_14044);
nor U15452 (N_15452,N_14308,N_14746);
nor U15453 (N_15453,N_14620,N_14459);
nor U15454 (N_15454,N_14109,N_14742);
and U15455 (N_15455,N_14409,N_14384);
nand U15456 (N_15456,N_14223,N_14633);
or U15457 (N_15457,N_14819,N_14672);
xnor U15458 (N_15458,N_14736,N_14564);
nand U15459 (N_15459,N_14756,N_14256);
nor U15460 (N_15460,N_14257,N_14007);
nor U15461 (N_15461,N_14140,N_14925);
nor U15462 (N_15462,N_14101,N_14644);
nor U15463 (N_15463,N_14242,N_14331);
and U15464 (N_15464,N_14211,N_14523);
or U15465 (N_15465,N_14634,N_14594);
nor U15466 (N_15466,N_14694,N_14104);
or U15467 (N_15467,N_14000,N_14156);
or U15468 (N_15468,N_14604,N_14435);
xnor U15469 (N_15469,N_14461,N_14894);
or U15470 (N_15470,N_14033,N_14219);
nor U15471 (N_15471,N_14600,N_14147);
nand U15472 (N_15472,N_14299,N_14309);
xnor U15473 (N_15473,N_14312,N_14111);
nand U15474 (N_15474,N_14056,N_14573);
or U15475 (N_15475,N_14560,N_14656);
or U15476 (N_15476,N_14499,N_14671);
and U15477 (N_15477,N_14665,N_14524);
nor U15478 (N_15478,N_14735,N_14531);
nand U15479 (N_15479,N_14483,N_14867);
or U15480 (N_15480,N_14702,N_14405);
nor U15481 (N_15481,N_14843,N_14866);
nand U15482 (N_15482,N_14036,N_14126);
and U15483 (N_15483,N_14338,N_14972);
nand U15484 (N_15484,N_14486,N_14456);
and U15485 (N_15485,N_14194,N_14284);
nor U15486 (N_15486,N_14642,N_14585);
nor U15487 (N_15487,N_14075,N_14226);
or U15488 (N_15488,N_14061,N_14134);
xor U15489 (N_15489,N_14747,N_14010);
nand U15490 (N_15490,N_14939,N_14525);
nor U15491 (N_15491,N_14250,N_14956);
or U15492 (N_15492,N_14966,N_14030);
nand U15493 (N_15493,N_14786,N_14590);
or U15494 (N_15494,N_14029,N_14319);
nand U15495 (N_15495,N_14864,N_14352);
nand U15496 (N_15496,N_14196,N_14471);
xor U15497 (N_15497,N_14719,N_14462);
xor U15498 (N_15498,N_14301,N_14394);
nand U15499 (N_15499,N_14092,N_14852);
xor U15500 (N_15500,N_14120,N_14719);
nor U15501 (N_15501,N_14915,N_14133);
or U15502 (N_15502,N_14898,N_14979);
and U15503 (N_15503,N_14782,N_14339);
nand U15504 (N_15504,N_14637,N_14311);
nand U15505 (N_15505,N_14058,N_14136);
nand U15506 (N_15506,N_14718,N_14445);
xnor U15507 (N_15507,N_14534,N_14936);
nor U15508 (N_15508,N_14831,N_14562);
xor U15509 (N_15509,N_14253,N_14467);
and U15510 (N_15510,N_14534,N_14058);
xor U15511 (N_15511,N_14813,N_14848);
nand U15512 (N_15512,N_14991,N_14172);
xor U15513 (N_15513,N_14429,N_14577);
and U15514 (N_15514,N_14860,N_14366);
xor U15515 (N_15515,N_14703,N_14983);
xnor U15516 (N_15516,N_14717,N_14404);
xor U15517 (N_15517,N_14304,N_14660);
nor U15518 (N_15518,N_14822,N_14727);
and U15519 (N_15519,N_14459,N_14503);
nor U15520 (N_15520,N_14249,N_14243);
nand U15521 (N_15521,N_14190,N_14720);
xnor U15522 (N_15522,N_14938,N_14039);
and U15523 (N_15523,N_14106,N_14340);
xor U15524 (N_15524,N_14799,N_14413);
or U15525 (N_15525,N_14452,N_14584);
or U15526 (N_15526,N_14932,N_14111);
or U15527 (N_15527,N_14635,N_14476);
or U15528 (N_15528,N_14898,N_14388);
or U15529 (N_15529,N_14040,N_14903);
and U15530 (N_15530,N_14199,N_14916);
xor U15531 (N_15531,N_14190,N_14071);
xnor U15532 (N_15532,N_14830,N_14746);
or U15533 (N_15533,N_14153,N_14961);
xnor U15534 (N_15534,N_14763,N_14908);
and U15535 (N_15535,N_14064,N_14608);
nand U15536 (N_15536,N_14819,N_14640);
nand U15537 (N_15537,N_14884,N_14008);
nor U15538 (N_15538,N_14673,N_14235);
nand U15539 (N_15539,N_14958,N_14334);
nand U15540 (N_15540,N_14178,N_14646);
xor U15541 (N_15541,N_14880,N_14291);
nand U15542 (N_15542,N_14624,N_14744);
and U15543 (N_15543,N_14672,N_14423);
or U15544 (N_15544,N_14332,N_14145);
nor U15545 (N_15545,N_14383,N_14776);
and U15546 (N_15546,N_14325,N_14150);
nor U15547 (N_15547,N_14810,N_14996);
nand U15548 (N_15548,N_14933,N_14417);
or U15549 (N_15549,N_14674,N_14679);
xor U15550 (N_15550,N_14528,N_14631);
xor U15551 (N_15551,N_14945,N_14559);
nand U15552 (N_15552,N_14959,N_14348);
xnor U15553 (N_15553,N_14897,N_14669);
nand U15554 (N_15554,N_14749,N_14459);
nand U15555 (N_15555,N_14448,N_14841);
xor U15556 (N_15556,N_14072,N_14938);
nor U15557 (N_15557,N_14046,N_14623);
xor U15558 (N_15558,N_14608,N_14316);
nand U15559 (N_15559,N_14898,N_14316);
nand U15560 (N_15560,N_14133,N_14093);
xor U15561 (N_15561,N_14725,N_14423);
or U15562 (N_15562,N_14217,N_14859);
nor U15563 (N_15563,N_14017,N_14436);
nor U15564 (N_15564,N_14904,N_14739);
nor U15565 (N_15565,N_14904,N_14658);
xor U15566 (N_15566,N_14101,N_14914);
nor U15567 (N_15567,N_14591,N_14613);
nor U15568 (N_15568,N_14472,N_14195);
nand U15569 (N_15569,N_14935,N_14535);
xor U15570 (N_15570,N_14109,N_14985);
xor U15571 (N_15571,N_14874,N_14868);
or U15572 (N_15572,N_14562,N_14333);
xor U15573 (N_15573,N_14010,N_14165);
nor U15574 (N_15574,N_14459,N_14319);
nand U15575 (N_15575,N_14577,N_14693);
and U15576 (N_15576,N_14085,N_14439);
and U15577 (N_15577,N_14074,N_14312);
nor U15578 (N_15578,N_14807,N_14125);
nand U15579 (N_15579,N_14565,N_14340);
nor U15580 (N_15580,N_14377,N_14956);
nand U15581 (N_15581,N_14706,N_14399);
nor U15582 (N_15582,N_14686,N_14225);
nor U15583 (N_15583,N_14616,N_14605);
nand U15584 (N_15584,N_14580,N_14797);
nor U15585 (N_15585,N_14652,N_14770);
or U15586 (N_15586,N_14560,N_14385);
or U15587 (N_15587,N_14401,N_14426);
or U15588 (N_15588,N_14231,N_14057);
nand U15589 (N_15589,N_14616,N_14869);
nand U15590 (N_15590,N_14309,N_14581);
nand U15591 (N_15591,N_14277,N_14063);
or U15592 (N_15592,N_14923,N_14787);
nor U15593 (N_15593,N_14432,N_14478);
and U15594 (N_15594,N_14829,N_14131);
xor U15595 (N_15595,N_14838,N_14776);
or U15596 (N_15596,N_14864,N_14949);
nor U15597 (N_15597,N_14611,N_14714);
or U15598 (N_15598,N_14867,N_14815);
and U15599 (N_15599,N_14625,N_14049);
nand U15600 (N_15600,N_14992,N_14900);
xor U15601 (N_15601,N_14387,N_14962);
and U15602 (N_15602,N_14752,N_14983);
xnor U15603 (N_15603,N_14174,N_14117);
or U15604 (N_15604,N_14009,N_14759);
nand U15605 (N_15605,N_14955,N_14218);
nor U15606 (N_15606,N_14212,N_14147);
and U15607 (N_15607,N_14134,N_14202);
nand U15608 (N_15608,N_14422,N_14914);
or U15609 (N_15609,N_14469,N_14380);
and U15610 (N_15610,N_14817,N_14707);
xor U15611 (N_15611,N_14586,N_14858);
and U15612 (N_15612,N_14735,N_14676);
or U15613 (N_15613,N_14878,N_14372);
nor U15614 (N_15614,N_14185,N_14855);
and U15615 (N_15615,N_14143,N_14553);
xnor U15616 (N_15616,N_14157,N_14296);
or U15617 (N_15617,N_14875,N_14752);
nand U15618 (N_15618,N_14498,N_14219);
nand U15619 (N_15619,N_14343,N_14600);
xor U15620 (N_15620,N_14940,N_14657);
xor U15621 (N_15621,N_14429,N_14939);
and U15622 (N_15622,N_14112,N_14179);
nand U15623 (N_15623,N_14640,N_14537);
and U15624 (N_15624,N_14569,N_14220);
and U15625 (N_15625,N_14662,N_14808);
or U15626 (N_15626,N_14408,N_14042);
xor U15627 (N_15627,N_14319,N_14475);
nand U15628 (N_15628,N_14023,N_14036);
or U15629 (N_15629,N_14615,N_14164);
nand U15630 (N_15630,N_14195,N_14221);
nand U15631 (N_15631,N_14269,N_14307);
nand U15632 (N_15632,N_14423,N_14253);
xor U15633 (N_15633,N_14938,N_14954);
and U15634 (N_15634,N_14426,N_14836);
nand U15635 (N_15635,N_14939,N_14087);
xor U15636 (N_15636,N_14647,N_14335);
nand U15637 (N_15637,N_14371,N_14197);
nand U15638 (N_15638,N_14307,N_14455);
and U15639 (N_15639,N_14643,N_14587);
nor U15640 (N_15640,N_14528,N_14032);
nor U15641 (N_15641,N_14443,N_14431);
xor U15642 (N_15642,N_14319,N_14180);
or U15643 (N_15643,N_14082,N_14906);
or U15644 (N_15644,N_14995,N_14974);
xnor U15645 (N_15645,N_14909,N_14409);
nand U15646 (N_15646,N_14655,N_14475);
nand U15647 (N_15647,N_14977,N_14681);
or U15648 (N_15648,N_14111,N_14711);
nor U15649 (N_15649,N_14237,N_14220);
nor U15650 (N_15650,N_14144,N_14935);
nor U15651 (N_15651,N_14752,N_14117);
nor U15652 (N_15652,N_14726,N_14154);
nand U15653 (N_15653,N_14561,N_14308);
and U15654 (N_15654,N_14619,N_14735);
nand U15655 (N_15655,N_14169,N_14712);
nor U15656 (N_15656,N_14316,N_14629);
or U15657 (N_15657,N_14779,N_14142);
nor U15658 (N_15658,N_14880,N_14211);
and U15659 (N_15659,N_14399,N_14865);
and U15660 (N_15660,N_14812,N_14694);
xor U15661 (N_15661,N_14677,N_14034);
and U15662 (N_15662,N_14757,N_14856);
xor U15663 (N_15663,N_14603,N_14582);
nor U15664 (N_15664,N_14057,N_14221);
xnor U15665 (N_15665,N_14556,N_14495);
nor U15666 (N_15666,N_14790,N_14369);
nand U15667 (N_15667,N_14165,N_14815);
nand U15668 (N_15668,N_14318,N_14029);
nand U15669 (N_15669,N_14566,N_14998);
and U15670 (N_15670,N_14529,N_14742);
xnor U15671 (N_15671,N_14179,N_14113);
or U15672 (N_15672,N_14842,N_14654);
nand U15673 (N_15673,N_14249,N_14718);
nor U15674 (N_15674,N_14056,N_14433);
nand U15675 (N_15675,N_14324,N_14696);
nor U15676 (N_15676,N_14565,N_14503);
nand U15677 (N_15677,N_14258,N_14191);
nor U15678 (N_15678,N_14494,N_14932);
or U15679 (N_15679,N_14759,N_14056);
xnor U15680 (N_15680,N_14160,N_14459);
nor U15681 (N_15681,N_14667,N_14122);
xor U15682 (N_15682,N_14357,N_14745);
nand U15683 (N_15683,N_14415,N_14752);
nor U15684 (N_15684,N_14323,N_14514);
xor U15685 (N_15685,N_14830,N_14587);
xor U15686 (N_15686,N_14450,N_14014);
and U15687 (N_15687,N_14724,N_14270);
and U15688 (N_15688,N_14242,N_14993);
and U15689 (N_15689,N_14156,N_14397);
and U15690 (N_15690,N_14132,N_14406);
or U15691 (N_15691,N_14966,N_14408);
nand U15692 (N_15692,N_14186,N_14838);
nor U15693 (N_15693,N_14735,N_14617);
and U15694 (N_15694,N_14234,N_14022);
xnor U15695 (N_15695,N_14604,N_14362);
xor U15696 (N_15696,N_14374,N_14897);
and U15697 (N_15697,N_14983,N_14451);
xor U15698 (N_15698,N_14438,N_14709);
xnor U15699 (N_15699,N_14108,N_14599);
xor U15700 (N_15700,N_14872,N_14116);
or U15701 (N_15701,N_14037,N_14183);
nor U15702 (N_15702,N_14795,N_14990);
and U15703 (N_15703,N_14706,N_14245);
nor U15704 (N_15704,N_14795,N_14160);
nor U15705 (N_15705,N_14350,N_14303);
or U15706 (N_15706,N_14147,N_14601);
nand U15707 (N_15707,N_14440,N_14302);
and U15708 (N_15708,N_14062,N_14714);
xnor U15709 (N_15709,N_14523,N_14632);
or U15710 (N_15710,N_14798,N_14145);
xor U15711 (N_15711,N_14594,N_14153);
nor U15712 (N_15712,N_14833,N_14345);
nand U15713 (N_15713,N_14280,N_14062);
nand U15714 (N_15714,N_14267,N_14563);
and U15715 (N_15715,N_14897,N_14421);
nand U15716 (N_15716,N_14467,N_14869);
nand U15717 (N_15717,N_14557,N_14066);
xnor U15718 (N_15718,N_14956,N_14995);
xnor U15719 (N_15719,N_14187,N_14233);
or U15720 (N_15720,N_14383,N_14780);
xor U15721 (N_15721,N_14319,N_14400);
nor U15722 (N_15722,N_14878,N_14853);
nor U15723 (N_15723,N_14375,N_14522);
and U15724 (N_15724,N_14475,N_14817);
nor U15725 (N_15725,N_14872,N_14960);
nand U15726 (N_15726,N_14941,N_14746);
xor U15727 (N_15727,N_14189,N_14852);
xor U15728 (N_15728,N_14803,N_14004);
nand U15729 (N_15729,N_14257,N_14718);
xnor U15730 (N_15730,N_14972,N_14421);
nor U15731 (N_15731,N_14739,N_14347);
or U15732 (N_15732,N_14140,N_14152);
xor U15733 (N_15733,N_14764,N_14331);
or U15734 (N_15734,N_14261,N_14324);
nor U15735 (N_15735,N_14468,N_14159);
nand U15736 (N_15736,N_14397,N_14823);
or U15737 (N_15737,N_14439,N_14575);
or U15738 (N_15738,N_14432,N_14831);
and U15739 (N_15739,N_14878,N_14816);
or U15740 (N_15740,N_14355,N_14435);
or U15741 (N_15741,N_14092,N_14989);
xor U15742 (N_15742,N_14551,N_14863);
nand U15743 (N_15743,N_14274,N_14734);
or U15744 (N_15744,N_14231,N_14535);
xnor U15745 (N_15745,N_14602,N_14416);
or U15746 (N_15746,N_14683,N_14216);
or U15747 (N_15747,N_14077,N_14834);
nor U15748 (N_15748,N_14740,N_14175);
and U15749 (N_15749,N_14905,N_14928);
nor U15750 (N_15750,N_14725,N_14775);
or U15751 (N_15751,N_14681,N_14127);
nor U15752 (N_15752,N_14180,N_14344);
nor U15753 (N_15753,N_14778,N_14794);
nor U15754 (N_15754,N_14446,N_14342);
nor U15755 (N_15755,N_14421,N_14110);
nor U15756 (N_15756,N_14014,N_14855);
and U15757 (N_15757,N_14631,N_14968);
and U15758 (N_15758,N_14222,N_14448);
and U15759 (N_15759,N_14706,N_14835);
nor U15760 (N_15760,N_14524,N_14452);
nand U15761 (N_15761,N_14591,N_14103);
and U15762 (N_15762,N_14680,N_14715);
or U15763 (N_15763,N_14681,N_14139);
xnor U15764 (N_15764,N_14256,N_14731);
xor U15765 (N_15765,N_14470,N_14363);
nor U15766 (N_15766,N_14770,N_14581);
and U15767 (N_15767,N_14097,N_14896);
xor U15768 (N_15768,N_14018,N_14469);
xor U15769 (N_15769,N_14445,N_14462);
xnor U15770 (N_15770,N_14055,N_14025);
or U15771 (N_15771,N_14317,N_14399);
nand U15772 (N_15772,N_14229,N_14913);
nand U15773 (N_15773,N_14147,N_14348);
or U15774 (N_15774,N_14783,N_14794);
and U15775 (N_15775,N_14871,N_14748);
xor U15776 (N_15776,N_14417,N_14113);
and U15777 (N_15777,N_14605,N_14778);
and U15778 (N_15778,N_14111,N_14521);
nor U15779 (N_15779,N_14849,N_14671);
xnor U15780 (N_15780,N_14163,N_14288);
nor U15781 (N_15781,N_14140,N_14344);
nor U15782 (N_15782,N_14741,N_14414);
nor U15783 (N_15783,N_14114,N_14082);
and U15784 (N_15784,N_14053,N_14204);
nand U15785 (N_15785,N_14829,N_14973);
and U15786 (N_15786,N_14143,N_14011);
nor U15787 (N_15787,N_14456,N_14904);
and U15788 (N_15788,N_14837,N_14508);
nand U15789 (N_15789,N_14289,N_14910);
and U15790 (N_15790,N_14999,N_14863);
xor U15791 (N_15791,N_14279,N_14421);
and U15792 (N_15792,N_14226,N_14504);
xor U15793 (N_15793,N_14102,N_14419);
or U15794 (N_15794,N_14475,N_14163);
xor U15795 (N_15795,N_14887,N_14946);
nand U15796 (N_15796,N_14425,N_14199);
or U15797 (N_15797,N_14102,N_14571);
nand U15798 (N_15798,N_14262,N_14002);
nand U15799 (N_15799,N_14486,N_14241);
or U15800 (N_15800,N_14701,N_14648);
nor U15801 (N_15801,N_14166,N_14818);
xor U15802 (N_15802,N_14851,N_14675);
or U15803 (N_15803,N_14566,N_14984);
or U15804 (N_15804,N_14937,N_14720);
or U15805 (N_15805,N_14144,N_14128);
nand U15806 (N_15806,N_14083,N_14455);
nand U15807 (N_15807,N_14470,N_14656);
nand U15808 (N_15808,N_14716,N_14837);
nor U15809 (N_15809,N_14967,N_14299);
nand U15810 (N_15810,N_14908,N_14528);
nand U15811 (N_15811,N_14976,N_14901);
or U15812 (N_15812,N_14263,N_14964);
or U15813 (N_15813,N_14227,N_14930);
nand U15814 (N_15814,N_14481,N_14058);
nor U15815 (N_15815,N_14476,N_14320);
nor U15816 (N_15816,N_14537,N_14016);
and U15817 (N_15817,N_14083,N_14364);
nor U15818 (N_15818,N_14945,N_14492);
nand U15819 (N_15819,N_14262,N_14342);
xor U15820 (N_15820,N_14938,N_14034);
nand U15821 (N_15821,N_14196,N_14694);
nor U15822 (N_15822,N_14093,N_14404);
and U15823 (N_15823,N_14465,N_14716);
and U15824 (N_15824,N_14166,N_14305);
nand U15825 (N_15825,N_14241,N_14655);
or U15826 (N_15826,N_14867,N_14446);
nor U15827 (N_15827,N_14790,N_14798);
and U15828 (N_15828,N_14073,N_14002);
xnor U15829 (N_15829,N_14891,N_14092);
or U15830 (N_15830,N_14943,N_14065);
or U15831 (N_15831,N_14441,N_14757);
nor U15832 (N_15832,N_14597,N_14975);
xnor U15833 (N_15833,N_14283,N_14192);
nand U15834 (N_15834,N_14381,N_14742);
nand U15835 (N_15835,N_14779,N_14181);
nor U15836 (N_15836,N_14202,N_14135);
nor U15837 (N_15837,N_14194,N_14744);
or U15838 (N_15838,N_14756,N_14492);
and U15839 (N_15839,N_14924,N_14646);
nand U15840 (N_15840,N_14232,N_14962);
nor U15841 (N_15841,N_14900,N_14017);
nand U15842 (N_15842,N_14142,N_14638);
or U15843 (N_15843,N_14534,N_14873);
and U15844 (N_15844,N_14641,N_14190);
nor U15845 (N_15845,N_14719,N_14908);
or U15846 (N_15846,N_14769,N_14187);
nand U15847 (N_15847,N_14480,N_14972);
nand U15848 (N_15848,N_14852,N_14254);
nand U15849 (N_15849,N_14609,N_14566);
and U15850 (N_15850,N_14285,N_14400);
nor U15851 (N_15851,N_14960,N_14545);
nand U15852 (N_15852,N_14731,N_14468);
xor U15853 (N_15853,N_14586,N_14943);
nor U15854 (N_15854,N_14882,N_14701);
nand U15855 (N_15855,N_14058,N_14490);
or U15856 (N_15856,N_14182,N_14122);
nor U15857 (N_15857,N_14612,N_14697);
nand U15858 (N_15858,N_14627,N_14665);
or U15859 (N_15859,N_14992,N_14863);
nand U15860 (N_15860,N_14999,N_14170);
nand U15861 (N_15861,N_14828,N_14029);
nor U15862 (N_15862,N_14695,N_14398);
xnor U15863 (N_15863,N_14066,N_14861);
or U15864 (N_15864,N_14011,N_14043);
or U15865 (N_15865,N_14945,N_14878);
xnor U15866 (N_15866,N_14600,N_14028);
nor U15867 (N_15867,N_14443,N_14894);
and U15868 (N_15868,N_14696,N_14613);
nand U15869 (N_15869,N_14333,N_14700);
nor U15870 (N_15870,N_14446,N_14901);
xor U15871 (N_15871,N_14047,N_14009);
nand U15872 (N_15872,N_14721,N_14568);
or U15873 (N_15873,N_14597,N_14915);
nand U15874 (N_15874,N_14677,N_14830);
nand U15875 (N_15875,N_14845,N_14584);
nor U15876 (N_15876,N_14949,N_14621);
xnor U15877 (N_15877,N_14311,N_14316);
nand U15878 (N_15878,N_14238,N_14779);
nand U15879 (N_15879,N_14758,N_14502);
and U15880 (N_15880,N_14153,N_14823);
or U15881 (N_15881,N_14239,N_14541);
xor U15882 (N_15882,N_14279,N_14024);
nor U15883 (N_15883,N_14439,N_14966);
or U15884 (N_15884,N_14130,N_14266);
and U15885 (N_15885,N_14442,N_14015);
or U15886 (N_15886,N_14643,N_14983);
nor U15887 (N_15887,N_14494,N_14997);
nor U15888 (N_15888,N_14534,N_14708);
xor U15889 (N_15889,N_14122,N_14044);
or U15890 (N_15890,N_14506,N_14561);
and U15891 (N_15891,N_14794,N_14796);
nand U15892 (N_15892,N_14208,N_14758);
nand U15893 (N_15893,N_14481,N_14003);
nor U15894 (N_15894,N_14701,N_14188);
nor U15895 (N_15895,N_14150,N_14674);
nor U15896 (N_15896,N_14873,N_14612);
and U15897 (N_15897,N_14906,N_14468);
and U15898 (N_15898,N_14903,N_14637);
xor U15899 (N_15899,N_14077,N_14854);
nor U15900 (N_15900,N_14285,N_14426);
or U15901 (N_15901,N_14565,N_14576);
xor U15902 (N_15902,N_14908,N_14235);
nor U15903 (N_15903,N_14610,N_14187);
nand U15904 (N_15904,N_14335,N_14455);
or U15905 (N_15905,N_14419,N_14615);
and U15906 (N_15906,N_14372,N_14246);
and U15907 (N_15907,N_14556,N_14565);
xnor U15908 (N_15908,N_14204,N_14246);
nand U15909 (N_15909,N_14978,N_14797);
xnor U15910 (N_15910,N_14162,N_14463);
nand U15911 (N_15911,N_14679,N_14040);
nor U15912 (N_15912,N_14603,N_14861);
or U15913 (N_15913,N_14488,N_14006);
nand U15914 (N_15914,N_14127,N_14329);
nand U15915 (N_15915,N_14927,N_14667);
xor U15916 (N_15916,N_14407,N_14022);
and U15917 (N_15917,N_14263,N_14422);
nor U15918 (N_15918,N_14374,N_14697);
xor U15919 (N_15919,N_14251,N_14396);
nor U15920 (N_15920,N_14190,N_14751);
xnor U15921 (N_15921,N_14261,N_14166);
and U15922 (N_15922,N_14294,N_14579);
or U15923 (N_15923,N_14551,N_14245);
nor U15924 (N_15924,N_14812,N_14663);
or U15925 (N_15925,N_14713,N_14106);
nor U15926 (N_15926,N_14692,N_14047);
nand U15927 (N_15927,N_14886,N_14216);
and U15928 (N_15928,N_14125,N_14179);
nor U15929 (N_15929,N_14272,N_14109);
nor U15930 (N_15930,N_14652,N_14293);
and U15931 (N_15931,N_14919,N_14136);
or U15932 (N_15932,N_14334,N_14339);
xor U15933 (N_15933,N_14647,N_14998);
and U15934 (N_15934,N_14159,N_14296);
xor U15935 (N_15935,N_14523,N_14241);
xor U15936 (N_15936,N_14664,N_14320);
nand U15937 (N_15937,N_14316,N_14140);
nand U15938 (N_15938,N_14957,N_14891);
or U15939 (N_15939,N_14156,N_14727);
or U15940 (N_15940,N_14952,N_14799);
and U15941 (N_15941,N_14330,N_14426);
nor U15942 (N_15942,N_14407,N_14540);
nor U15943 (N_15943,N_14706,N_14357);
xor U15944 (N_15944,N_14426,N_14750);
nor U15945 (N_15945,N_14642,N_14975);
or U15946 (N_15946,N_14258,N_14132);
nor U15947 (N_15947,N_14431,N_14098);
or U15948 (N_15948,N_14871,N_14575);
nand U15949 (N_15949,N_14358,N_14529);
nand U15950 (N_15950,N_14595,N_14781);
nor U15951 (N_15951,N_14265,N_14400);
nor U15952 (N_15952,N_14014,N_14865);
and U15953 (N_15953,N_14048,N_14059);
and U15954 (N_15954,N_14130,N_14612);
nand U15955 (N_15955,N_14906,N_14238);
or U15956 (N_15956,N_14109,N_14118);
nor U15957 (N_15957,N_14443,N_14928);
nand U15958 (N_15958,N_14510,N_14110);
xnor U15959 (N_15959,N_14199,N_14594);
xor U15960 (N_15960,N_14300,N_14735);
and U15961 (N_15961,N_14051,N_14006);
and U15962 (N_15962,N_14218,N_14309);
or U15963 (N_15963,N_14012,N_14744);
or U15964 (N_15964,N_14119,N_14210);
xor U15965 (N_15965,N_14014,N_14035);
nand U15966 (N_15966,N_14798,N_14911);
nand U15967 (N_15967,N_14925,N_14266);
xor U15968 (N_15968,N_14330,N_14961);
xnor U15969 (N_15969,N_14749,N_14171);
nand U15970 (N_15970,N_14491,N_14512);
nor U15971 (N_15971,N_14074,N_14054);
nor U15972 (N_15972,N_14351,N_14063);
or U15973 (N_15973,N_14618,N_14890);
and U15974 (N_15974,N_14225,N_14523);
and U15975 (N_15975,N_14198,N_14365);
nor U15976 (N_15976,N_14347,N_14250);
and U15977 (N_15977,N_14755,N_14981);
xnor U15978 (N_15978,N_14289,N_14856);
and U15979 (N_15979,N_14987,N_14068);
nand U15980 (N_15980,N_14359,N_14629);
and U15981 (N_15981,N_14465,N_14479);
nand U15982 (N_15982,N_14608,N_14443);
xnor U15983 (N_15983,N_14780,N_14630);
nand U15984 (N_15984,N_14642,N_14444);
and U15985 (N_15985,N_14744,N_14927);
nor U15986 (N_15986,N_14882,N_14044);
or U15987 (N_15987,N_14841,N_14886);
and U15988 (N_15988,N_14538,N_14866);
and U15989 (N_15989,N_14522,N_14686);
and U15990 (N_15990,N_14677,N_14992);
and U15991 (N_15991,N_14499,N_14750);
xor U15992 (N_15992,N_14720,N_14550);
nor U15993 (N_15993,N_14623,N_14436);
or U15994 (N_15994,N_14099,N_14904);
xnor U15995 (N_15995,N_14220,N_14533);
xor U15996 (N_15996,N_14167,N_14055);
nand U15997 (N_15997,N_14948,N_14731);
xnor U15998 (N_15998,N_14107,N_14428);
xor U15999 (N_15999,N_14470,N_14066);
nand U16000 (N_16000,N_15169,N_15145);
and U16001 (N_16001,N_15049,N_15783);
nand U16002 (N_16002,N_15286,N_15102);
nor U16003 (N_16003,N_15067,N_15668);
nor U16004 (N_16004,N_15302,N_15309);
nand U16005 (N_16005,N_15831,N_15106);
xor U16006 (N_16006,N_15517,N_15187);
nor U16007 (N_16007,N_15122,N_15873);
or U16008 (N_16008,N_15489,N_15841);
nor U16009 (N_16009,N_15919,N_15300);
nor U16010 (N_16010,N_15260,N_15340);
nand U16011 (N_16011,N_15764,N_15289);
nand U16012 (N_16012,N_15775,N_15405);
and U16013 (N_16013,N_15147,N_15570);
and U16014 (N_16014,N_15768,N_15709);
or U16015 (N_16015,N_15110,N_15786);
xor U16016 (N_16016,N_15227,N_15165);
nand U16017 (N_16017,N_15151,N_15513);
or U16018 (N_16018,N_15735,N_15663);
nand U16019 (N_16019,N_15058,N_15642);
xor U16020 (N_16020,N_15705,N_15141);
xor U16021 (N_16021,N_15238,N_15393);
and U16022 (N_16022,N_15987,N_15878);
nor U16023 (N_16023,N_15906,N_15082);
nor U16024 (N_16024,N_15785,N_15745);
nor U16025 (N_16025,N_15686,N_15799);
xnor U16026 (N_16026,N_15299,N_15031);
xor U16027 (N_16027,N_15379,N_15247);
nand U16028 (N_16028,N_15407,N_15641);
nor U16029 (N_16029,N_15531,N_15898);
or U16030 (N_16030,N_15751,N_15885);
or U16031 (N_16031,N_15943,N_15884);
and U16032 (N_16032,N_15046,N_15606);
or U16033 (N_16033,N_15318,N_15837);
and U16034 (N_16034,N_15638,N_15723);
xnor U16035 (N_16035,N_15479,N_15500);
or U16036 (N_16036,N_15903,N_15211);
or U16037 (N_16037,N_15365,N_15436);
nand U16038 (N_16038,N_15478,N_15864);
and U16039 (N_16039,N_15331,N_15862);
xor U16040 (N_16040,N_15076,N_15139);
nand U16041 (N_16041,N_15372,N_15054);
nand U16042 (N_16042,N_15448,N_15839);
nor U16043 (N_16043,N_15215,N_15875);
xor U16044 (N_16044,N_15652,N_15883);
and U16045 (N_16045,N_15213,N_15869);
nor U16046 (N_16046,N_15132,N_15959);
xnor U16047 (N_16047,N_15524,N_15616);
nand U16048 (N_16048,N_15635,N_15874);
nor U16049 (N_16049,N_15386,N_15565);
nand U16050 (N_16050,N_15738,N_15251);
or U16051 (N_16051,N_15353,N_15858);
xnor U16052 (N_16052,N_15265,N_15782);
nand U16053 (N_16053,N_15576,N_15117);
xnor U16054 (N_16054,N_15792,N_15441);
nor U16055 (N_16055,N_15167,N_15494);
xor U16056 (N_16056,N_15722,N_15254);
nand U16057 (N_16057,N_15469,N_15274);
or U16058 (N_16058,N_15264,N_15714);
and U16059 (N_16059,N_15654,N_15623);
or U16060 (N_16060,N_15776,N_15276);
xnor U16061 (N_16061,N_15281,N_15672);
xor U16062 (N_16062,N_15596,N_15371);
nand U16063 (N_16063,N_15356,N_15221);
and U16064 (N_16064,N_15970,N_15643);
nor U16065 (N_16065,N_15320,N_15438);
xor U16066 (N_16066,N_15189,N_15475);
nor U16067 (N_16067,N_15508,N_15470);
and U16068 (N_16068,N_15428,N_15892);
and U16069 (N_16069,N_15501,N_15505);
or U16070 (N_16070,N_15346,N_15385);
nor U16071 (N_16071,N_15061,N_15902);
or U16072 (N_16072,N_15112,N_15933);
or U16073 (N_16073,N_15198,N_15509);
and U16074 (N_16074,N_15760,N_15806);
nand U16075 (N_16075,N_15460,N_15486);
nand U16076 (N_16076,N_15521,N_15242);
xnor U16077 (N_16077,N_15421,N_15612);
xor U16078 (N_16078,N_15868,N_15120);
and U16079 (N_16079,N_15793,N_15588);
nor U16080 (N_16080,N_15975,N_15537);
xor U16081 (N_16081,N_15182,N_15996);
nand U16082 (N_16082,N_15894,N_15599);
and U16083 (N_16083,N_15010,N_15856);
nor U16084 (N_16084,N_15375,N_15832);
or U16085 (N_16085,N_15396,N_15064);
nor U16086 (N_16086,N_15288,N_15284);
nor U16087 (N_16087,N_15569,N_15457);
and U16088 (N_16088,N_15133,N_15471);
xnor U16089 (N_16089,N_15940,N_15810);
xor U16090 (N_16090,N_15794,N_15620);
or U16091 (N_16091,N_15949,N_15997);
xnor U16092 (N_16092,N_15495,N_15155);
and U16093 (N_16093,N_15752,N_15945);
and U16094 (N_16094,N_15081,N_15192);
and U16095 (N_16095,N_15631,N_15637);
xnor U16096 (N_16096,N_15740,N_15941);
nor U16097 (N_16097,N_15473,N_15684);
and U16098 (N_16098,N_15472,N_15159);
and U16099 (N_16099,N_15548,N_15149);
xor U16100 (N_16100,N_15555,N_15851);
nand U16101 (N_16101,N_15844,N_15582);
and U16102 (N_16102,N_15339,N_15886);
or U16103 (N_16103,N_15063,N_15560);
nor U16104 (N_16104,N_15235,N_15414);
and U16105 (N_16105,N_15158,N_15127);
xor U16106 (N_16106,N_15437,N_15540);
xnor U16107 (N_16107,N_15821,N_15131);
xor U16108 (N_16108,N_15050,N_15079);
or U16109 (N_16109,N_15335,N_15271);
xnor U16110 (N_16110,N_15001,N_15921);
and U16111 (N_16111,N_15715,N_15329);
and U16112 (N_16112,N_15880,N_15912);
nand U16113 (N_16113,N_15754,N_15241);
xor U16114 (N_16114,N_15700,N_15711);
xnor U16115 (N_16115,N_15930,N_15237);
nand U16116 (N_16116,N_15412,N_15310);
or U16117 (N_16117,N_15963,N_15577);
and U16118 (N_16118,N_15729,N_15293);
nor U16119 (N_16119,N_15915,N_15815);
nand U16120 (N_16120,N_15662,N_15180);
nor U16121 (N_16121,N_15511,N_15474);
and U16122 (N_16122,N_15246,N_15009);
nor U16123 (N_16123,N_15233,N_15163);
or U16124 (N_16124,N_15273,N_15721);
or U16125 (N_16125,N_15748,N_15143);
and U16126 (N_16126,N_15332,N_15173);
or U16127 (N_16127,N_15649,N_15602);
nand U16128 (N_16128,N_15998,N_15944);
nor U16129 (N_16129,N_15953,N_15590);
or U16130 (N_16130,N_15529,N_15258);
or U16131 (N_16131,N_15086,N_15157);
xor U16132 (N_16132,N_15653,N_15974);
xnor U16133 (N_16133,N_15384,N_15275);
nand U16134 (N_16134,N_15267,N_15303);
nor U16135 (N_16135,N_15931,N_15435);
or U16136 (N_16136,N_15466,N_15349);
or U16137 (N_16137,N_15950,N_15717);
xnor U16138 (N_16138,N_15680,N_15694);
nor U16139 (N_16139,N_15695,N_15593);
and U16140 (N_16140,N_15036,N_15160);
nand U16141 (N_16141,N_15223,N_15727);
nand U16142 (N_16142,N_15399,N_15222);
or U16143 (N_16143,N_15625,N_15034);
or U16144 (N_16144,N_15481,N_15947);
nand U16145 (N_16145,N_15546,N_15003);
or U16146 (N_16146,N_15601,N_15055);
or U16147 (N_16147,N_15614,N_15467);
xnor U16148 (N_16148,N_15195,N_15913);
xnor U16149 (N_16149,N_15011,N_15609);
or U16150 (N_16150,N_15762,N_15536);
nor U16151 (N_16151,N_15772,N_15589);
xnor U16152 (N_16152,N_15644,N_15820);
and U16153 (N_16153,N_15871,N_15390);
nand U16154 (N_16154,N_15788,N_15659);
or U16155 (N_16155,N_15315,N_15454);
or U16156 (N_16156,N_15453,N_15938);
and U16157 (N_16157,N_15655,N_15295);
and U16158 (N_16158,N_15716,N_15564);
nand U16159 (N_16159,N_15370,N_15013);
nor U16160 (N_16160,N_15171,N_15351);
or U16161 (N_16161,N_15743,N_15713);
xnor U16162 (N_16162,N_15100,N_15243);
and U16163 (N_16163,N_15140,N_15733);
or U16164 (N_16164,N_15592,N_15850);
nand U16165 (N_16165,N_15480,N_15763);
nand U16166 (N_16166,N_15965,N_15447);
or U16167 (N_16167,N_15545,N_15861);
nand U16168 (N_16168,N_15982,N_15515);
and U16169 (N_16169,N_15089,N_15019);
or U16170 (N_16170,N_15683,N_15865);
and U16171 (N_16171,N_15035,N_15988);
xnor U16172 (N_16172,N_15336,N_15119);
nand U16173 (N_16173,N_15566,N_15897);
and U16174 (N_16174,N_15773,N_15877);
xnor U16175 (N_16175,N_15825,N_15424);
and U16176 (N_16176,N_15226,N_15634);
and U16177 (N_16177,N_15301,N_15319);
nand U16178 (N_16178,N_15551,N_15607);
xnor U16179 (N_16179,N_15113,N_15224);
or U16180 (N_16180,N_15430,N_15840);
nor U16181 (N_16181,N_15528,N_15125);
or U16182 (N_16182,N_15463,N_15855);
or U16183 (N_16183,N_15981,N_15502);
and U16184 (N_16184,N_15419,N_15870);
nand U16185 (N_16185,N_15842,N_15976);
and U16186 (N_16186,N_15362,N_15829);
or U16187 (N_16187,N_15962,N_15395);
nor U16188 (N_16188,N_15583,N_15377);
xnor U16189 (N_16189,N_15193,N_15893);
nand U16190 (N_16190,N_15206,N_15854);
nand U16191 (N_16191,N_15742,N_15306);
nor U16192 (N_16192,N_15044,N_15039);
xor U16193 (N_16193,N_15542,N_15890);
xor U16194 (N_16194,N_15758,N_15809);
nand U16195 (N_16195,N_15461,N_15613);
and U16196 (N_16196,N_15325,N_15423);
and U16197 (N_16197,N_15016,N_15344);
or U16198 (N_16198,N_15692,N_15863);
xor U16199 (N_16199,N_15527,N_15484);
or U16200 (N_16200,N_15843,N_15532);
nand U16201 (N_16201,N_15148,N_15170);
xnor U16202 (N_16202,N_15357,N_15123);
and U16203 (N_16203,N_15969,N_15400);
xor U16204 (N_16204,N_15739,N_15465);
xor U16205 (N_16205,N_15455,N_15350);
nand U16206 (N_16206,N_15369,N_15647);
or U16207 (N_16207,N_15209,N_15701);
xnor U16208 (N_16208,N_15784,N_15543);
or U16209 (N_16209,N_15578,N_15420);
nand U16210 (N_16210,N_15980,N_15923);
xnor U16211 (N_16211,N_15628,N_15699);
nor U16212 (N_16212,N_15935,N_15955);
nand U16213 (N_16213,N_15586,N_15707);
nor U16214 (N_16214,N_15905,N_15728);
and U16215 (N_16215,N_15026,N_15525);
nor U16216 (N_16216,N_15427,N_15909);
nor U16217 (N_16217,N_15972,N_15622);
and U16218 (N_16218,N_15138,N_15093);
and U16219 (N_16219,N_15126,N_15805);
or U16220 (N_16220,N_15376,N_15107);
nand U16221 (N_16221,N_15136,N_15746);
nor U16222 (N_16222,N_15388,N_15040);
xnor U16223 (N_16223,N_15826,N_15166);
nand U16224 (N_16224,N_15450,N_15835);
and U16225 (N_16225,N_15533,N_15355);
xnor U16226 (N_16226,N_15304,N_15585);
nor U16227 (N_16227,N_15757,N_15676);
nand U16228 (N_16228,N_15364,N_15324);
xor U16229 (N_16229,N_15530,N_15939);
nor U16230 (N_16230,N_15552,N_15904);
or U16231 (N_16231,N_15047,N_15704);
nand U16232 (N_16232,N_15462,N_15814);
nand U16233 (N_16233,N_15538,N_15587);
nor U16234 (N_16234,N_15108,N_15492);
xnor U16235 (N_16235,N_15404,N_15121);
and U16236 (N_16236,N_15337,N_15024);
nand U16237 (N_16237,N_15358,N_15808);
xor U16238 (N_16238,N_15852,N_15681);
xnor U16239 (N_16239,N_15190,N_15703);
xor U16240 (N_16240,N_15732,N_15907);
and U16241 (N_16241,N_15270,N_15071);
nor U16242 (N_16242,N_15347,N_15266);
or U16243 (N_16243,N_15656,N_15651);
xnor U16244 (N_16244,N_15261,N_15203);
nand U16245 (N_16245,N_15901,N_15429);
nor U16246 (N_16246,N_15150,N_15401);
nand U16247 (N_16247,N_15640,N_15137);
or U16248 (N_16248,N_15510,N_15617);
or U16249 (N_16249,N_15294,N_15797);
and U16250 (N_16250,N_15368,N_15824);
or U16251 (N_16251,N_15848,N_15128);
xnor U16252 (N_16252,N_15181,N_15177);
xnor U16253 (N_16253,N_15927,N_15403);
or U16254 (N_16254,N_15697,N_15766);
nor U16255 (N_16255,N_15553,N_15971);
nor U16256 (N_16256,N_15750,N_15657);
or U16257 (N_16257,N_15954,N_15426);
nand U16258 (N_16258,N_15391,N_15452);
xnor U16259 (N_16259,N_15204,N_15269);
or U16260 (N_16260,N_15085,N_15398);
and U16261 (N_16261,N_15658,N_15250);
nor U16262 (N_16262,N_15410,N_15216);
nand U16263 (N_16263,N_15519,N_15896);
nor U16264 (N_16264,N_15146,N_15522);
xor U16265 (N_16265,N_15575,N_15926);
and U16266 (N_16266,N_15632,N_15803);
nand U16267 (N_16267,N_15708,N_15178);
nand U16268 (N_16268,N_15661,N_15456);
and U16269 (N_16269,N_15020,N_15790);
nor U16270 (N_16270,N_15446,N_15174);
and U16271 (N_16271,N_15175,N_15394);
and U16272 (N_16272,N_15556,N_15065);
nand U16273 (N_16273,N_15090,N_15853);
nand U16274 (N_16274,N_15374,N_15753);
xnor U16275 (N_16275,N_15696,N_15413);
or U16276 (N_16276,N_15099,N_15443);
nand U16277 (N_16277,N_15262,N_15296);
xnor U16278 (N_16278,N_15240,N_15033);
nor U16279 (N_16279,N_15539,N_15664);
and U16280 (N_16280,N_15879,N_15341);
nand U16281 (N_16281,N_15859,N_15581);
nor U16282 (N_16282,N_15053,N_15778);
and U16283 (N_16283,N_15605,N_15411);
and U16284 (N_16284,N_15951,N_15691);
nand U16285 (N_16285,N_15352,N_15279);
and U16286 (N_16286,N_15978,N_15818);
nor U16287 (N_16287,N_15381,N_15078);
nor U16288 (N_16288,N_15201,N_15208);
xnor U16289 (N_16289,N_15719,N_15630);
nor U16290 (N_16290,N_15493,N_15343);
nand U16291 (N_16291,N_15629,N_15194);
nand U16292 (N_16292,N_15600,N_15779);
xor U16293 (N_16293,N_15857,N_15562);
and U16294 (N_16294,N_15698,N_15777);
nor U16295 (N_16295,N_15268,N_15115);
or U16296 (N_16296,N_15162,N_15451);
nand U16297 (N_16297,N_15021,N_15042);
nor U16298 (N_16298,N_15256,N_15060);
xor U16299 (N_16299,N_15311,N_15769);
and U16300 (N_16300,N_15406,N_15029);
and U16301 (N_16301,N_15671,N_15520);
nor U16302 (N_16302,N_15409,N_15490);
nor U16303 (N_16303,N_15670,N_15449);
nor U16304 (N_16304,N_15008,N_15477);
nand U16305 (N_16305,N_15229,N_15822);
and U16306 (N_16306,N_15800,N_15022);
or U16307 (N_16307,N_15482,N_15734);
xor U16308 (N_16308,N_15559,N_15230);
or U16309 (N_16309,N_15544,N_15487);
xor U16310 (N_16310,N_15297,N_15253);
xor U16311 (N_16311,N_15780,N_15690);
xor U16312 (N_16312,N_15847,N_15366);
nor U16313 (N_16313,N_15184,N_15702);
nor U16314 (N_16314,N_15819,N_15983);
nand U16315 (N_16315,N_15767,N_15259);
or U16316 (N_16316,N_15077,N_15756);
nand U16317 (N_16317,N_15737,N_15041);
and U16318 (N_16318,N_15402,N_15882);
or U16319 (N_16319,N_15387,N_15730);
nand U16320 (N_16320,N_15706,N_15354);
xor U16321 (N_16321,N_15849,N_15316);
nand U16322 (N_16322,N_15574,N_15660);
xnor U16323 (N_16323,N_15114,N_15636);
nor U16324 (N_16324,N_15291,N_15639);
and U16325 (N_16325,N_15973,N_15669);
and U16326 (N_16326,N_15891,N_15827);
nor U16327 (N_16327,N_15367,N_15550);
nor U16328 (N_16328,N_15693,N_15389);
nand U16329 (N_16329,N_15549,N_15594);
or U16330 (N_16330,N_15334,N_15363);
nand U16331 (N_16331,N_15307,N_15097);
nand U16332 (N_16332,N_15277,N_15263);
nor U16333 (N_16333,N_15504,N_15791);
and U16334 (N_16334,N_15345,N_15084);
nand U16335 (N_16335,N_15666,N_15018);
nor U16336 (N_16336,N_15313,N_15872);
xnor U16337 (N_16337,N_15360,N_15272);
nand U16338 (N_16338,N_15129,N_15506);
and U16339 (N_16339,N_15098,N_15507);
nor U16340 (N_16340,N_15012,N_15887);
nor U16341 (N_16341,N_15993,N_15744);
nor U16342 (N_16342,N_15104,N_15995);
nor U16343 (N_16343,N_15967,N_15069);
nor U16344 (N_16344,N_15817,N_15212);
xor U16345 (N_16345,N_15028,N_15860);
nand U16346 (N_16346,N_15535,N_15244);
xor U16347 (N_16347,N_15228,N_15483);
and U16348 (N_16348,N_15239,N_15152);
nor U16349 (N_16349,N_15154,N_15074);
or U16350 (N_16350,N_15442,N_15322);
nor U16351 (N_16351,N_15936,N_15679);
nor U16352 (N_16352,N_15218,N_15185);
nor U16353 (N_16353,N_15673,N_15781);
nor U16354 (N_16354,N_15397,N_15846);
and U16355 (N_16355,N_15172,N_15283);
and U16356 (N_16356,N_15627,N_15795);
nor U16357 (N_16357,N_15937,N_15312);
xor U16358 (N_16358,N_15674,N_15801);
nor U16359 (N_16359,N_15045,N_15444);
nor U16360 (N_16360,N_15603,N_15186);
xnor U16361 (N_16361,N_15798,N_15914);
and U16362 (N_16362,N_15488,N_15207);
or U16363 (N_16363,N_15497,N_15979);
nor U16364 (N_16364,N_15986,N_15095);
xnor U16365 (N_16365,N_15677,N_15205);
and U16366 (N_16366,N_15485,N_15000);
xnor U16367 (N_16367,N_15881,N_15498);
nor U16368 (N_16368,N_15416,N_15116);
nand U16369 (N_16369,N_15408,N_15580);
xor U16370 (N_16370,N_15816,N_15070);
nor U16371 (N_16371,N_15749,N_15561);
xnor U16372 (N_16372,N_15889,N_15828);
nand U16373 (N_16373,N_15968,N_15179);
xor U16374 (N_16374,N_15161,N_15468);
and U16375 (N_16375,N_15232,N_15910);
xnor U16376 (N_16376,N_15811,N_15595);
and U16377 (N_16377,N_15014,N_15929);
nor U16378 (N_16378,N_15499,N_15491);
xor U16379 (N_16379,N_15526,N_15459);
or U16380 (N_16380,N_15415,N_15431);
nand U16381 (N_16381,N_15091,N_15168);
nand U16382 (N_16382,N_15619,N_15802);
xnor U16383 (N_16383,N_15323,N_15432);
nor U16384 (N_16384,N_15961,N_15087);
xnor U16385 (N_16385,N_15004,N_15867);
and U16386 (N_16386,N_15056,N_15964);
nor U16387 (N_16387,N_15571,N_15188);
xnor U16388 (N_16388,N_15200,N_15958);
nor U16389 (N_16389,N_15002,N_15759);
xnor U16390 (N_16390,N_15573,N_15217);
nor U16391 (N_16391,N_15458,N_15027);
and U16392 (N_16392,N_15895,N_15496);
and U16393 (N_16393,N_15048,N_15567);
nor U16394 (N_16394,N_15135,N_15920);
xor U16395 (N_16395,N_15285,N_15199);
and U16396 (N_16396,N_15900,N_15298);
or U16397 (N_16397,N_15557,N_15946);
nand U16398 (N_16398,N_15023,N_15665);
nand U16399 (N_16399,N_15876,N_15830);
and U16400 (N_16400,N_15621,N_15183);
or U16401 (N_16401,N_15476,N_15908);
and U16402 (N_16402,N_15984,N_15292);
nand U16403 (N_16403,N_15770,N_15057);
or U16404 (N_16404,N_15142,N_15675);
and U16405 (N_16405,N_15037,N_15888);
nand U16406 (N_16406,N_15833,N_15418);
nor U16407 (N_16407,N_15796,N_15092);
xnor U16408 (N_16408,N_15164,N_15032);
nand U16409 (N_16409,N_15989,N_15667);
and U16410 (N_16410,N_15966,N_15597);
or U16411 (N_16411,N_15080,N_15234);
nor U16412 (N_16412,N_15718,N_15321);
or U16413 (N_16413,N_15030,N_15836);
or U16414 (N_16414,N_15006,N_15382);
nor U16415 (N_16415,N_15682,N_15096);
xor U16416 (N_16416,N_15922,N_15725);
nand U16417 (N_16417,N_15823,N_15248);
nor U16418 (N_16418,N_15236,N_15807);
or U16419 (N_16419,N_15918,N_15305);
xnor U16420 (N_16420,N_15615,N_15417);
nor U16421 (N_16421,N_15604,N_15066);
nor U16422 (N_16422,N_15225,N_15584);
nor U16423 (N_16423,N_15308,N_15361);
and U16424 (N_16424,N_15156,N_15153);
xnor U16425 (N_16425,N_15977,N_15608);
xnor U16426 (N_16426,N_15917,N_15523);
or U16427 (N_16427,N_15747,N_15838);
nand U16428 (N_16428,N_15678,N_15359);
or U16429 (N_16429,N_15942,N_15202);
and U16430 (N_16430,N_15755,N_15257);
or U16431 (N_16431,N_15025,N_15934);
nand U16432 (N_16432,N_15547,N_15518);
nand U16433 (N_16433,N_15072,N_15924);
nor U16434 (N_16434,N_15541,N_15124);
or U16435 (N_16435,N_15990,N_15591);
and U16436 (N_16436,N_15327,N_15813);
nor U16437 (N_16437,N_15383,N_15255);
and U16438 (N_16438,N_15991,N_15911);
or U16439 (N_16439,N_15088,N_15646);
nand U16440 (N_16440,N_15017,N_15439);
xor U16441 (N_16441,N_15985,N_15252);
and U16442 (N_16442,N_15598,N_15710);
and U16443 (N_16443,N_15111,N_15220);
and U16444 (N_16444,N_15464,N_15994);
nand U16445 (N_16445,N_15068,N_15130);
nor U16446 (N_16446,N_15568,N_15342);
nor U16447 (N_16447,N_15380,N_15624);
and U16448 (N_16448,N_15689,N_15774);
or U16449 (N_16449,N_15916,N_15197);
xnor U16450 (N_16450,N_15043,N_15348);
or U16451 (N_16451,N_15957,N_15433);
and U16452 (N_16452,N_15075,N_15059);
xor U16453 (N_16453,N_15960,N_15720);
nand U16454 (N_16454,N_15512,N_15736);
nand U16455 (N_16455,N_15196,N_15290);
and U16456 (N_16456,N_15952,N_15118);
nor U16457 (N_16457,N_15326,N_15245);
nor U16458 (N_16458,N_15038,N_15214);
nand U16459 (N_16459,N_15534,N_15176);
and U16460 (N_16460,N_15094,N_15378);
or U16461 (N_16461,N_15134,N_15191);
xor U16462 (N_16462,N_15109,N_15650);
nor U16463 (N_16463,N_15330,N_15333);
or U16464 (N_16464,N_15611,N_15563);
nor U16465 (N_16465,N_15278,N_15249);
xor U16466 (N_16466,N_15688,N_15282);
nand U16467 (N_16467,N_15062,N_15645);
and U16468 (N_16468,N_15899,N_15610);
nand U16469 (N_16469,N_15516,N_15834);
xnor U16470 (N_16470,N_15434,N_15626);
and U16471 (N_16471,N_15787,N_15932);
nor U16472 (N_16472,N_15948,N_15314);
nand U16473 (N_16473,N_15724,N_15579);
and U16474 (N_16474,N_15812,N_15726);
xnor U16475 (N_16475,N_15992,N_15445);
or U16476 (N_16476,N_15633,N_15103);
or U16477 (N_16477,N_15144,N_15845);
nor U16478 (N_16478,N_15514,N_15572);
or U16479 (N_16479,N_15928,N_15373);
and U16480 (N_16480,N_15083,N_15422);
and U16481 (N_16481,N_15956,N_15005);
xnor U16482 (N_16482,N_15712,N_15231);
or U16483 (N_16483,N_15999,N_15771);
xnor U16484 (N_16484,N_15741,N_15051);
nor U16485 (N_16485,N_15052,N_15618);
xor U16486 (N_16486,N_15425,N_15338);
nor U16487 (N_16487,N_15101,N_15925);
xor U16488 (N_16488,N_15328,N_15804);
or U16489 (N_16489,N_15554,N_15392);
nor U16490 (N_16490,N_15685,N_15219);
and U16491 (N_16491,N_15015,N_15866);
nand U16492 (N_16492,N_15558,N_15210);
or U16493 (N_16493,N_15503,N_15280);
nand U16494 (N_16494,N_15761,N_15007);
and U16495 (N_16495,N_15687,N_15105);
xor U16496 (N_16496,N_15440,N_15765);
nand U16497 (N_16497,N_15073,N_15287);
or U16498 (N_16498,N_15731,N_15789);
xor U16499 (N_16499,N_15317,N_15648);
nand U16500 (N_16500,N_15883,N_15893);
nand U16501 (N_16501,N_15236,N_15148);
and U16502 (N_16502,N_15068,N_15835);
or U16503 (N_16503,N_15209,N_15327);
nor U16504 (N_16504,N_15738,N_15298);
xor U16505 (N_16505,N_15538,N_15744);
xnor U16506 (N_16506,N_15963,N_15558);
and U16507 (N_16507,N_15122,N_15954);
nand U16508 (N_16508,N_15783,N_15787);
xnor U16509 (N_16509,N_15464,N_15083);
nand U16510 (N_16510,N_15802,N_15035);
or U16511 (N_16511,N_15456,N_15995);
nor U16512 (N_16512,N_15065,N_15186);
xnor U16513 (N_16513,N_15459,N_15333);
or U16514 (N_16514,N_15270,N_15349);
or U16515 (N_16515,N_15051,N_15356);
or U16516 (N_16516,N_15339,N_15469);
xnor U16517 (N_16517,N_15297,N_15375);
nor U16518 (N_16518,N_15029,N_15010);
xnor U16519 (N_16519,N_15499,N_15406);
or U16520 (N_16520,N_15138,N_15614);
or U16521 (N_16521,N_15146,N_15865);
xnor U16522 (N_16522,N_15609,N_15111);
xor U16523 (N_16523,N_15524,N_15370);
xnor U16524 (N_16524,N_15792,N_15842);
or U16525 (N_16525,N_15520,N_15236);
nand U16526 (N_16526,N_15816,N_15394);
nor U16527 (N_16527,N_15806,N_15702);
nor U16528 (N_16528,N_15095,N_15862);
xnor U16529 (N_16529,N_15165,N_15540);
xnor U16530 (N_16530,N_15340,N_15212);
nand U16531 (N_16531,N_15940,N_15452);
nand U16532 (N_16532,N_15013,N_15623);
nor U16533 (N_16533,N_15602,N_15505);
and U16534 (N_16534,N_15212,N_15242);
and U16535 (N_16535,N_15043,N_15878);
or U16536 (N_16536,N_15847,N_15518);
or U16537 (N_16537,N_15650,N_15337);
nand U16538 (N_16538,N_15679,N_15784);
nor U16539 (N_16539,N_15177,N_15462);
or U16540 (N_16540,N_15100,N_15017);
and U16541 (N_16541,N_15148,N_15584);
and U16542 (N_16542,N_15659,N_15979);
nand U16543 (N_16543,N_15699,N_15192);
nor U16544 (N_16544,N_15819,N_15086);
nor U16545 (N_16545,N_15979,N_15418);
nand U16546 (N_16546,N_15598,N_15014);
and U16547 (N_16547,N_15583,N_15829);
nand U16548 (N_16548,N_15753,N_15583);
nor U16549 (N_16549,N_15378,N_15095);
or U16550 (N_16550,N_15759,N_15932);
nand U16551 (N_16551,N_15167,N_15048);
and U16552 (N_16552,N_15767,N_15084);
nand U16553 (N_16553,N_15189,N_15950);
and U16554 (N_16554,N_15296,N_15155);
xnor U16555 (N_16555,N_15615,N_15107);
nor U16556 (N_16556,N_15562,N_15498);
and U16557 (N_16557,N_15052,N_15915);
or U16558 (N_16558,N_15229,N_15648);
xor U16559 (N_16559,N_15228,N_15498);
or U16560 (N_16560,N_15796,N_15111);
and U16561 (N_16561,N_15922,N_15710);
or U16562 (N_16562,N_15422,N_15328);
or U16563 (N_16563,N_15122,N_15988);
or U16564 (N_16564,N_15295,N_15152);
nor U16565 (N_16565,N_15430,N_15244);
nand U16566 (N_16566,N_15429,N_15405);
nand U16567 (N_16567,N_15460,N_15615);
or U16568 (N_16568,N_15685,N_15106);
xnor U16569 (N_16569,N_15049,N_15344);
or U16570 (N_16570,N_15114,N_15495);
and U16571 (N_16571,N_15262,N_15241);
nor U16572 (N_16572,N_15004,N_15752);
nor U16573 (N_16573,N_15591,N_15348);
and U16574 (N_16574,N_15541,N_15594);
xnor U16575 (N_16575,N_15417,N_15169);
and U16576 (N_16576,N_15795,N_15075);
xor U16577 (N_16577,N_15263,N_15472);
nor U16578 (N_16578,N_15980,N_15939);
nand U16579 (N_16579,N_15606,N_15421);
nand U16580 (N_16580,N_15521,N_15524);
xnor U16581 (N_16581,N_15343,N_15952);
or U16582 (N_16582,N_15200,N_15181);
nand U16583 (N_16583,N_15702,N_15213);
nand U16584 (N_16584,N_15492,N_15450);
xnor U16585 (N_16585,N_15077,N_15708);
nand U16586 (N_16586,N_15913,N_15817);
and U16587 (N_16587,N_15725,N_15356);
nand U16588 (N_16588,N_15497,N_15378);
nor U16589 (N_16589,N_15493,N_15803);
nand U16590 (N_16590,N_15390,N_15062);
xor U16591 (N_16591,N_15697,N_15357);
or U16592 (N_16592,N_15969,N_15291);
and U16593 (N_16593,N_15072,N_15604);
nor U16594 (N_16594,N_15078,N_15415);
or U16595 (N_16595,N_15240,N_15744);
nor U16596 (N_16596,N_15096,N_15273);
or U16597 (N_16597,N_15317,N_15820);
xor U16598 (N_16598,N_15073,N_15729);
or U16599 (N_16599,N_15336,N_15357);
and U16600 (N_16600,N_15890,N_15173);
nor U16601 (N_16601,N_15567,N_15755);
and U16602 (N_16602,N_15648,N_15875);
or U16603 (N_16603,N_15381,N_15893);
or U16604 (N_16604,N_15120,N_15245);
or U16605 (N_16605,N_15918,N_15591);
nand U16606 (N_16606,N_15675,N_15957);
or U16607 (N_16607,N_15567,N_15634);
or U16608 (N_16608,N_15750,N_15927);
xnor U16609 (N_16609,N_15464,N_15084);
or U16610 (N_16610,N_15782,N_15711);
xnor U16611 (N_16611,N_15371,N_15867);
and U16612 (N_16612,N_15762,N_15670);
nor U16613 (N_16613,N_15583,N_15028);
or U16614 (N_16614,N_15546,N_15517);
xnor U16615 (N_16615,N_15690,N_15016);
or U16616 (N_16616,N_15211,N_15974);
nand U16617 (N_16617,N_15021,N_15731);
nor U16618 (N_16618,N_15135,N_15013);
and U16619 (N_16619,N_15585,N_15042);
xnor U16620 (N_16620,N_15063,N_15043);
xnor U16621 (N_16621,N_15829,N_15572);
or U16622 (N_16622,N_15253,N_15489);
nand U16623 (N_16623,N_15415,N_15741);
xor U16624 (N_16624,N_15958,N_15455);
nor U16625 (N_16625,N_15662,N_15072);
nand U16626 (N_16626,N_15746,N_15789);
nor U16627 (N_16627,N_15393,N_15235);
and U16628 (N_16628,N_15364,N_15331);
nand U16629 (N_16629,N_15372,N_15736);
nor U16630 (N_16630,N_15514,N_15578);
or U16631 (N_16631,N_15404,N_15732);
xor U16632 (N_16632,N_15711,N_15455);
or U16633 (N_16633,N_15395,N_15635);
nor U16634 (N_16634,N_15178,N_15188);
and U16635 (N_16635,N_15014,N_15077);
nor U16636 (N_16636,N_15545,N_15999);
and U16637 (N_16637,N_15387,N_15756);
or U16638 (N_16638,N_15351,N_15923);
nand U16639 (N_16639,N_15196,N_15119);
and U16640 (N_16640,N_15707,N_15309);
xnor U16641 (N_16641,N_15629,N_15384);
nor U16642 (N_16642,N_15568,N_15654);
and U16643 (N_16643,N_15249,N_15525);
nor U16644 (N_16644,N_15067,N_15269);
xnor U16645 (N_16645,N_15836,N_15845);
or U16646 (N_16646,N_15477,N_15206);
xnor U16647 (N_16647,N_15855,N_15698);
nor U16648 (N_16648,N_15195,N_15428);
nor U16649 (N_16649,N_15790,N_15074);
or U16650 (N_16650,N_15265,N_15450);
nor U16651 (N_16651,N_15541,N_15102);
xor U16652 (N_16652,N_15409,N_15460);
or U16653 (N_16653,N_15448,N_15381);
and U16654 (N_16654,N_15285,N_15400);
nand U16655 (N_16655,N_15312,N_15463);
or U16656 (N_16656,N_15468,N_15948);
and U16657 (N_16657,N_15980,N_15168);
nand U16658 (N_16658,N_15886,N_15969);
or U16659 (N_16659,N_15790,N_15471);
nand U16660 (N_16660,N_15008,N_15192);
nor U16661 (N_16661,N_15423,N_15508);
nor U16662 (N_16662,N_15837,N_15111);
and U16663 (N_16663,N_15475,N_15253);
and U16664 (N_16664,N_15443,N_15043);
and U16665 (N_16665,N_15054,N_15438);
xor U16666 (N_16666,N_15113,N_15774);
or U16667 (N_16667,N_15910,N_15003);
and U16668 (N_16668,N_15112,N_15809);
and U16669 (N_16669,N_15206,N_15394);
or U16670 (N_16670,N_15395,N_15416);
and U16671 (N_16671,N_15678,N_15516);
nand U16672 (N_16672,N_15265,N_15849);
or U16673 (N_16673,N_15068,N_15637);
nor U16674 (N_16674,N_15833,N_15839);
and U16675 (N_16675,N_15156,N_15792);
and U16676 (N_16676,N_15705,N_15792);
or U16677 (N_16677,N_15303,N_15774);
or U16678 (N_16678,N_15381,N_15706);
or U16679 (N_16679,N_15489,N_15433);
or U16680 (N_16680,N_15765,N_15501);
or U16681 (N_16681,N_15012,N_15178);
or U16682 (N_16682,N_15533,N_15847);
or U16683 (N_16683,N_15117,N_15459);
or U16684 (N_16684,N_15734,N_15882);
nand U16685 (N_16685,N_15316,N_15201);
or U16686 (N_16686,N_15996,N_15098);
or U16687 (N_16687,N_15121,N_15220);
nor U16688 (N_16688,N_15345,N_15942);
nand U16689 (N_16689,N_15821,N_15910);
nand U16690 (N_16690,N_15555,N_15781);
nor U16691 (N_16691,N_15237,N_15455);
xor U16692 (N_16692,N_15013,N_15151);
nand U16693 (N_16693,N_15230,N_15936);
nor U16694 (N_16694,N_15276,N_15814);
nand U16695 (N_16695,N_15727,N_15659);
or U16696 (N_16696,N_15757,N_15063);
nand U16697 (N_16697,N_15914,N_15852);
nand U16698 (N_16698,N_15947,N_15398);
xnor U16699 (N_16699,N_15959,N_15649);
nor U16700 (N_16700,N_15612,N_15276);
nand U16701 (N_16701,N_15410,N_15536);
xor U16702 (N_16702,N_15147,N_15233);
nand U16703 (N_16703,N_15348,N_15027);
or U16704 (N_16704,N_15830,N_15680);
nand U16705 (N_16705,N_15447,N_15314);
or U16706 (N_16706,N_15052,N_15178);
nor U16707 (N_16707,N_15755,N_15762);
and U16708 (N_16708,N_15711,N_15428);
nor U16709 (N_16709,N_15261,N_15495);
and U16710 (N_16710,N_15729,N_15375);
xnor U16711 (N_16711,N_15744,N_15059);
nor U16712 (N_16712,N_15036,N_15189);
nand U16713 (N_16713,N_15041,N_15526);
nor U16714 (N_16714,N_15419,N_15214);
nor U16715 (N_16715,N_15961,N_15380);
and U16716 (N_16716,N_15222,N_15795);
xnor U16717 (N_16717,N_15643,N_15332);
and U16718 (N_16718,N_15256,N_15902);
or U16719 (N_16719,N_15535,N_15705);
and U16720 (N_16720,N_15057,N_15157);
or U16721 (N_16721,N_15619,N_15326);
nand U16722 (N_16722,N_15898,N_15117);
xor U16723 (N_16723,N_15792,N_15599);
or U16724 (N_16724,N_15550,N_15818);
xnor U16725 (N_16725,N_15035,N_15322);
nand U16726 (N_16726,N_15847,N_15190);
nand U16727 (N_16727,N_15468,N_15374);
xnor U16728 (N_16728,N_15238,N_15326);
nand U16729 (N_16729,N_15560,N_15940);
nor U16730 (N_16730,N_15370,N_15418);
xnor U16731 (N_16731,N_15210,N_15289);
or U16732 (N_16732,N_15135,N_15402);
and U16733 (N_16733,N_15220,N_15842);
nand U16734 (N_16734,N_15756,N_15007);
and U16735 (N_16735,N_15805,N_15760);
xnor U16736 (N_16736,N_15821,N_15782);
or U16737 (N_16737,N_15703,N_15431);
nor U16738 (N_16738,N_15429,N_15238);
and U16739 (N_16739,N_15708,N_15257);
xnor U16740 (N_16740,N_15801,N_15053);
nand U16741 (N_16741,N_15672,N_15724);
nand U16742 (N_16742,N_15896,N_15682);
xor U16743 (N_16743,N_15517,N_15962);
or U16744 (N_16744,N_15922,N_15300);
nand U16745 (N_16745,N_15269,N_15046);
nor U16746 (N_16746,N_15691,N_15365);
xnor U16747 (N_16747,N_15752,N_15891);
or U16748 (N_16748,N_15261,N_15284);
xnor U16749 (N_16749,N_15658,N_15771);
and U16750 (N_16750,N_15643,N_15302);
or U16751 (N_16751,N_15008,N_15406);
nand U16752 (N_16752,N_15644,N_15846);
and U16753 (N_16753,N_15305,N_15101);
or U16754 (N_16754,N_15714,N_15555);
xnor U16755 (N_16755,N_15154,N_15853);
or U16756 (N_16756,N_15530,N_15409);
and U16757 (N_16757,N_15093,N_15024);
and U16758 (N_16758,N_15516,N_15276);
xnor U16759 (N_16759,N_15739,N_15781);
nor U16760 (N_16760,N_15552,N_15263);
nor U16761 (N_16761,N_15957,N_15429);
xnor U16762 (N_16762,N_15631,N_15484);
nor U16763 (N_16763,N_15893,N_15691);
nand U16764 (N_16764,N_15783,N_15884);
nand U16765 (N_16765,N_15510,N_15060);
xor U16766 (N_16766,N_15242,N_15762);
and U16767 (N_16767,N_15590,N_15177);
and U16768 (N_16768,N_15526,N_15982);
and U16769 (N_16769,N_15886,N_15417);
nor U16770 (N_16770,N_15928,N_15521);
nand U16771 (N_16771,N_15609,N_15804);
xor U16772 (N_16772,N_15092,N_15986);
nand U16773 (N_16773,N_15215,N_15621);
or U16774 (N_16774,N_15553,N_15061);
nand U16775 (N_16775,N_15675,N_15578);
and U16776 (N_16776,N_15925,N_15747);
nand U16777 (N_16777,N_15926,N_15459);
nand U16778 (N_16778,N_15044,N_15284);
nand U16779 (N_16779,N_15515,N_15071);
nand U16780 (N_16780,N_15535,N_15037);
and U16781 (N_16781,N_15367,N_15521);
nand U16782 (N_16782,N_15269,N_15648);
nor U16783 (N_16783,N_15721,N_15713);
nand U16784 (N_16784,N_15360,N_15286);
nand U16785 (N_16785,N_15464,N_15302);
nand U16786 (N_16786,N_15566,N_15151);
nor U16787 (N_16787,N_15921,N_15491);
nand U16788 (N_16788,N_15281,N_15532);
xnor U16789 (N_16789,N_15774,N_15741);
and U16790 (N_16790,N_15695,N_15592);
xnor U16791 (N_16791,N_15330,N_15733);
and U16792 (N_16792,N_15371,N_15853);
or U16793 (N_16793,N_15960,N_15426);
nor U16794 (N_16794,N_15348,N_15274);
nor U16795 (N_16795,N_15471,N_15845);
xor U16796 (N_16796,N_15635,N_15188);
and U16797 (N_16797,N_15675,N_15822);
nand U16798 (N_16798,N_15835,N_15244);
nor U16799 (N_16799,N_15739,N_15038);
nor U16800 (N_16800,N_15902,N_15159);
nand U16801 (N_16801,N_15673,N_15455);
nand U16802 (N_16802,N_15642,N_15497);
or U16803 (N_16803,N_15785,N_15850);
nor U16804 (N_16804,N_15947,N_15083);
nand U16805 (N_16805,N_15933,N_15066);
nand U16806 (N_16806,N_15441,N_15753);
xnor U16807 (N_16807,N_15616,N_15474);
or U16808 (N_16808,N_15463,N_15691);
nor U16809 (N_16809,N_15184,N_15497);
nor U16810 (N_16810,N_15124,N_15978);
nor U16811 (N_16811,N_15514,N_15880);
nor U16812 (N_16812,N_15160,N_15524);
or U16813 (N_16813,N_15353,N_15420);
nand U16814 (N_16814,N_15586,N_15493);
and U16815 (N_16815,N_15755,N_15025);
xnor U16816 (N_16816,N_15841,N_15920);
and U16817 (N_16817,N_15711,N_15469);
nor U16818 (N_16818,N_15526,N_15236);
xnor U16819 (N_16819,N_15446,N_15881);
nor U16820 (N_16820,N_15335,N_15314);
nand U16821 (N_16821,N_15433,N_15184);
nand U16822 (N_16822,N_15217,N_15212);
nand U16823 (N_16823,N_15540,N_15434);
or U16824 (N_16824,N_15549,N_15744);
nand U16825 (N_16825,N_15878,N_15889);
xor U16826 (N_16826,N_15812,N_15002);
or U16827 (N_16827,N_15451,N_15823);
nand U16828 (N_16828,N_15515,N_15978);
nor U16829 (N_16829,N_15427,N_15895);
nor U16830 (N_16830,N_15431,N_15272);
nor U16831 (N_16831,N_15722,N_15125);
or U16832 (N_16832,N_15422,N_15600);
nand U16833 (N_16833,N_15282,N_15783);
nand U16834 (N_16834,N_15905,N_15278);
nor U16835 (N_16835,N_15847,N_15099);
nand U16836 (N_16836,N_15655,N_15501);
and U16837 (N_16837,N_15067,N_15153);
or U16838 (N_16838,N_15045,N_15290);
or U16839 (N_16839,N_15678,N_15082);
and U16840 (N_16840,N_15093,N_15931);
nor U16841 (N_16841,N_15471,N_15111);
nand U16842 (N_16842,N_15360,N_15172);
nand U16843 (N_16843,N_15251,N_15668);
xnor U16844 (N_16844,N_15837,N_15997);
and U16845 (N_16845,N_15836,N_15866);
xor U16846 (N_16846,N_15368,N_15045);
nor U16847 (N_16847,N_15116,N_15673);
or U16848 (N_16848,N_15091,N_15546);
and U16849 (N_16849,N_15541,N_15821);
nand U16850 (N_16850,N_15078,N_15318);
and U16851 (N_16851,N_15222,N_15636);
xor U16852 (N_16852,N_15156,N_15535);
or U16853 (N_16853,N_15155,N_15803);
and U16854 (N_16854,N_15509,N_15361);
nand U16855 (N_16855,N_15571,N_15421);
or U16856 (N_16856,N_15381,N_15394);
nand U16857 (N_16857,N_15548,N_15201);
nor U16858 (N_16858,N_15534,N_15934);
nor U16859 (N_16859,N_15738,N_15203);
or U16860 (N_16860,N_15082,N_15526);
or U16861 (N_16861,N_15331,N_15272);
and U16862 (N_16862,N_15627,N_15198);
nand U16863 (N_16863,N_15722,N_15296);
and U16864 (N_16864,N_15972,N_15508);
nor U16865 (N_16865,N_15081,N_15851);
xnor U16866 (N_16866,N_15363,N_15083);
nor U16867 (N_16867,N_15617,N_15610);
or U16868 (N_16868,N_15540,N_15583);
or U16869 (N_16869,N_15691,N_15174);
and U16870 (N_16870,N_15009,N_15344);
or U16871 (N_16871,N_15185,N_15083);
or U16872 (N_16872,N_15601,N_15547);
or U16873 (N_16873,N_15336,N_15455);
nor U16874 (N_16874,N_15904,N_15886);
and U16875 (N_16875,N_15563,N_15419);
or U16876 (N_16876,N_15050,N_15504);
nor U16877 (N_16877,N_15823,N_15516);
nand U16878 (N_16878,N_15667,N_15137);
xor U16879 (N_16879,N_15070,N_15543);
and U16880 (N_16880,N_15387,N_15919);
and U16881 (N_16881,N_15336,N_15206);
and U16882 (N_16882,N_15798,N_15633);
nand U16883 (N_16883,N_15007,N_15378);
or U16884 (N_16884,N_15673,N_15585);
nand U16885 (N_16885,N_15303,N_15799);
nand U16886 (N_16886,N_15773,N_15916);
nand U16887 (N_16887,N_15993,N_15896);
nor U16888 (N_16888,N_15094,N_15326);
xor U16889 (N_16889,N_15458,N_15140);
nor U16890 (N_16890,N_15794,N_15701);
xor U16891 (N_16891,N_15892,N_15942);
or U16892 (N_16892,N_15144,N_15060);
and U16893 (N_16893,N_15727,N_15354);
xor U16894 (N_16894,N_15649,N_15850);
and U16895 (N_16895,N_15008,N_15772);
nor U16896 (N_16896,N_15874,N_15817);
or U16897 (N_16897,N_15544,N_15172);
nand U16898 (N_16898,N_15132,N_15862);
nand U16899 (N_16899,N_15536,N_15900);
nand U16900 (N_16900,N_15321,N_15635);
xor U16901 (N_16901,N_15582,N_15223);
or U16902 (N_16902,N_15409,N_15370);
or U16903 (N_16903,N_15909,N_15251);
or U16904 (N_16904,N_15986,N_15585);
or U16905 (N_16905,N_15586,N_15598);
nand U16906 (N_16906,N_15155,N_15701);
nand U16907 (N_16907,N_15500,N_15255);
nor U16908 (N_16908,N_15655,N_15029);
or U16909 (N_16909,N_15589,N_15842);
or U16910 (N_16910,N_15122,N_15007);
or U16911 (N_16911,N_15045,N_15548);
xnor U16912 (N_16912,N_15701,N_15649);
xor U16913 (N_16913,N_15523,N_15822);
nand U16914 (N_16914,N_15311,N_15661);
or U16915 (N_16915,N_15668,N_15988);
xor U16916 (N_16916,N_15795,N_15655);
or U16917 (N_16917,N_15773,N_15377);
and U16918 (N_16918,N_15921,N_15623);
nor U16919 (N_16919,N_15499,N_15578);
nor U16920 (N_16920,N_15039,N_15685);
xor U16921 (N_16921,N_15344,N_15834);
and U16922 (N_16922,N_15179,N_15063);
nor U16923 (N_16923,N_15055,N_15717);
or U16924 (N_16924,N_15291,N_15887);
and U16925 (N_16925,N_15283,N_15533);
xnor U16926 (N_16926,N_15230,N_15709);
and U16927 (N_16927,N_15829,N_15481);
or U16928 (N_16928,N_15784,N_15793);
nand U16929 (N_16929,N_15521,N_15011);
xnor U16930 (N_16930,N_15423,N_15990);
and U16931 (N_16931,N_15749,N_15200);
or U16932 (N_16932,N_15735,N_15533);
nand U16933 (N_16933,N_15697,N_15316);
xor U16934 (N_16934,N_15458,N_15259);
xor U16935 (N_16935,N_15181,N_15938);
and U16936 (N_16936,N_15601,N_15203);
and U16937 (N_16937,N_15466,N_15012);
nor U16938 (N_16938,N_15099,N_15983);
xnor U16939 (N_16939,N_15133,N_15886);
nor U16940 (N_16940,N_15961,N_15247);
nor U16941 (N_16941,N_15144,N_15023);
nand U16942 (N_16942,N_15689,N_15786);
or U16943 (N_16943,N_15717,N_15911);
nor U16944 (N_16944,N_15050,N_15326);
xor U16945 (N_16945,N_15492,N_15409);
nand U16946 (N_16946,N_15211,N_15495);
and U16947 (N_16947,N_15487,N_15519);
or U16948 (N_16948,N_15733,N_15923);
xnor U16949 (N_16949,N_15284,N_15112);
or U16950 (N_16950,N_15904,N_15926);
nand U16951 (N_16951,N_15793,N_15477);
xor U16952 (N_16952,N_15807,N_15659);
nand U16953 (N_16953,N_15364,N_15519);
or U16954 (N_16954,N_15767,N_15470);
or U16955 (N_16955,N_15032,N_15109);
or U16956 (N_16956,N_15113,N_15294);
or U16957 (N_16957,N_15922,N_15782);
nor U16958 (N_16958,N_15603,N_15363);
or U16959 (N_16959,N_15569,N_15182);
nand U16960 (N_16960,N_15941,N_15273);
nand U16961 (N_16961,N_15040,N_15742);
xnor U16962 (N_16962,N_15762,N_15144);
and U16963 (N_16963,N_15265,N_15982);
xnor U16964 (N_16964,N_15416,N_15998);
nor U16965 (N_16965,N_15546,N_15378);
nand U16966 (N_16966,N_15448,N_15505);
or U16967 (N_16967,N_15362,N_15148);
nand U16968 (N_16968,N_15313,N_15815);
or U16969 (N_16969,N_15090,N_15624);
and U16970 (N_16970,N_15767,N_15903);
or U16971 (N_16971,N_15471,N_15855);
nor U16972 (N_16972,N_15140,N_15766);
and U16973 (N_16973,N_15620,N_15210);
nand U16974 (N_16974,N_15152,N_15724);
or U16975 (N_16975,N_15009,N_15928);
xnor U16976 (N_16976,N_15942,N_15778);
or U16977 (N_16977,N_15771,N_15679);
xnor U16978 (N_16978,N_15884,N_15904);
nor U16979 (N_16979,N_15715,N_15152);
and U16980 (N_16980,N_15585,N_15071);
and U16981 (N_16981,N_15963,N_15044);
or U16982 (N_16982,N_15677,N_15068);
xnor U16983 (N_16983,N_15698,N_15466);
or U16984 (N_16984,N_15956,N_15509);
and U16985 (N_16985,N_15874,N_15243);
and U16986 (N_16986,N_15657,N_15866);
xnor U16987 (N_16987,N_15828,N_15143);
or U16988 (N_16988,N_15174,N_15557);
xnor U16989 (N_16989,N_15731,N_15594);
nand U16990 (N_16990,N_15678,N_15352);
nand U16991 (N_16991,N_15174,N_15157);
and U16992 (N_16992,N_15804,N_15564);
nand U16993 (N_16993,N_15440,N_15046);
nand U16994 (N_16994,N_15371,N_15631);
xnor U16995 (N_16995,N_15498,N_15026);
or U16996 (N_16996,N_15791,N_15382);
or U16997 (N_16997,N_15924,N_15066);
xor U16998 (N_16998,N_15461,N_15992);
and U16999 (N_16999,N_15060,N_15859);
or U17000 (N_17000,N_16982,N_16957);
nor U17001 (N_17001,N_16429,N_16016);
and U17002 (N_17002,N_16195,N_16824);
and U17003 (N_17003,N_16585,N_16618);
nor U17004 (N_17004,N_16104,N_16326);
nor U17005 (N_17005,N_16673,N_16591);
nand U17006 (N_17006,N_16480,N_16811);
nor U17007 (N_17007,N_16004,N_16595);
nand U17008 (N_17008,N_16122,N_16170);
or U17009 (N_17009,N_16850,N_16518);
nor U17010 (N_17010,N_16972,N_16665);
or U17011 (N_17011,N_16049,N_16523);
xnor U17012 (N_17012,N_16501,N_16137);
and U17013 (N_17013,N_16302,N_16428);
xnor U17014 (N_17014,N_16040,N_16263);
or U17015 (N_17015,N_16332,N_16319);
nand U17016 (N_17016,N_16756,N_16861);
and U17017 (N_17017,N_16228,N_16866);
or U17018 (N_17018,N_16366,N_16583);
and U17019 (N_17019,N_16990,N_16022);
nand U17020 (N_17020,N_16478,N_16590);
nor U17021 (N_17021,N_16145,N_16808);
or U17022 (N_17022,N_16785,N_16610);
or U17023 (N_17023,N_16368,N_16928);
nand U17024 (N_17024,N_16453,N_16183);
and U17025 (N_17025,N_16846,N_16419);
or U17026 (N_17026,N_16098,N_16210);
and U17027 (N_17027,N_16830,N_16679);
xnor U17028 (N_17028,N_16773,N_16044);
nor U17029 (N_17029,N_16031,N_16181);
nor U17030 (N_17030,N_16248,N_16669);
or U17031 (N_17031,N_16742,N_16331);
nand U17032 (N_17032,N_16985,N_16015);
or U17033 (N_17033,N_16639,N_16500);
xor U17034 (N_17034,N_16382,N_16338);
xnor U17035 (N_17035,N_16176,N_16576);
nor U17036 (N_17036,N_16127,N_16254);
and U17037 (N_17037,N_16447,N_16130);
or U17038 (N_17038,N_16000,N_16281);
and U17039 (N_17039,N_16617,N_16086);
or U17040 (N_17040,N_16198,N_16173);
xor U17041 (N_17041,N_16117,N_16153);
and U17042 (N_17042,N_16735,N_16242);
or U17043 (N_17043,N_16490,N_16370);
or U17044 (N_17044,N_16530,N_16247);
xor U17045 (N_17045,N_16476,N_16746);
xnor U17046 (N_17046,N_16213,N_16816);
nand U17047 (N_17047,N_16645,N_16788);
nand U17048 (N_17048,N_16479,N_16201);
nand U17049 (N_17049,N_16291,N_16712);
xor U17050 (N_17050,N_16792,N_16837);
xnor U17051 (N_17051,N_16027,N_16601);
or U17052 (N_17052,N_16282,N_16457);
nand U17053 (N_17053,N_16165,N_16743);
or U17054 (N_17054,N_16007,N_16573);
or U17055 (N_17055,N_16339,N_16769);
nor U17056 (N_17056,N_16310,N_16449);
nand U17057 (N_17057,N_16536,N_16632);
nand U17058 (N_17058,N_16731,N_16580);
or U17059 (N_17059,N_16111,N_16971);
or U17060 (N_17060,N_16316,N_16094);
and U17061 (N_17061,N_16693,N_16290);
nor U17062 (N_17062,N_16570,N_16634);
and U17063 (N_17063,N_16546,N_16134);
or U17064 (N_17064,N_16096,N_16726);
or U17065 (N_17065,N_16912,N_16556);
xor U17066 (N_17066,N_16287,N_16073);
or U17067 (N_17067,N_16562,N_16091);
xnor U17068 (N_17068,N_16032,N_16880);
nor U17069 (N_17069,N_16361,N_16904);
nor U17070 (N_17070,N_16818,N_16256);
and U17071 (N_17071,N_16289,N_16897);
xor U17072 (N_17072,N_16118,N_16847);
nand U17073 (N_17073,N_16891,N_16531);
or U17074 (N_17074,N_16283,N_16421);
and U17075 (N_17075,N_16009,N_16789);
nand U17076 (N_17076,N_16780,N_16638);
xor U17077 (N_17077,N_16119,N_16061);
xor U17078 (N_17078,N_16822,N_16615);
nor U17079 (N_17079,N_16411,N_16517);
nor U17080 (N_17080,N_16948,N_16875);
or U17081 (N_17081,N_16935,N_16285);
xor U17082 (N_17082,N_16143,N_16910);
or U17083 (N_17083,N_16343,N_16803);
xor U17084 (N_17084,N_16486,N_16755);
xor U17085 (N_17085,N_16724,N_16744);
nor U17086 (N_17086,N_16065,N_16710);
nor U17087 (N_17087,N_16322,N_16495);
or U17088 (N_17088,N_16359,N_16342);
or U17089 (N_17089,N_16661,N_16124);
or U17090 (N_17090,N_16223,N_16823);
and U17091 (N_17091,N_16688,N_16074);
or U17092 (N_17092,N_16162,N_16771);
nand U17093 (N_17093,N_16271,N_16221);
or U17094 (N_17094,N_16001,N_16510);
nand U17095 (N_17095,N_16083,N_16732);
and U17096 (N_17096,N_16494,N_16676);
xnor U17097 (N_17097,N_16574,N_16164);
and U17098 (N_17098,N_16055,N_16471);
nor U17099 (N_17099,N_16779,N_16078);
and U17100 (N_17100,N_16514,N_16709);
nand U17101 (N_17101,N_16047,N_16862);
xnor U17102 (N_17102,N_16983,N_16072);
nor U17103 (N_17103,N_16774,N_16696);
nand U17104 (N_17104,N_16140,N_16565);
or U17105 (N_17105,N_16468,N_16087);
or U17106 (N_17106,N_16413,N_16068);
or U17107 (N_17107,N_16253,N_16733);
xnor U17108 (N_17108,N_16351,N_16416);
and U17109 (N_17109,N_16033,N_16795);
nand U17110 (N_17110,N_16986,N_16019);
nand U17111 (N_17111,N_16970,N_16876);
and U17112 (N_17112,N_16113,N_16269);
and U17113 (N_17113,N_16108,N_16937);
and U17114 (N_17114,N_16608,N_16435);
xor U17115 (N_17115,N_16809,N_16105);
nand U17116 (N_17116,N_16489,N_16660);
and U17117 (N_17117,N_16511,N_16587);
and U17118 (N_17118,N_16672,N_16540);
or U17119 (N_17119,N_16558,N_16666);
nand U17120 (N_17120,N_16923,N_16241);
or U17121 (N_17121,N_16272,N_16424);
or U17122 (N_17122,N_16978,N_16778);
nand U17123 (N_17123,N_16103,N_16488);
nor U17124 (N_17124,N_16062,N_16526);
nand U17125 (N_17125,N_16635,N_16456);
and U17126 (N_17126,N_16594,N_16155);
nand U17127 (N_17127,N_16944,N_16147);
nand U17128 (N_17128,N_16474,N_16005);
xnor U17129 (N_17129,N_16920,N_16825);
xnor U17130 (N_17130,N_16030,N_16237);
or U17131 (N_17131,N_16954,N_16029);
nand U17132 (N_17132,N_16403,N_16204);
or U17133 (N_17133,N_16884,N_16790);
nor U17134 (N_17134,N_16492,N_16350);
nor U17135 (N_17135,N_16649,N_16292);
or U17136 (N_17136,N_16782,N_16497);
nor U17137 (N_17137,N_16801,N_16431);
or U17138 (N_17138,N_16462,N_16849);
nor U17139 (N_17139,N_16303,N_16512);
nand U17140 (N_17140,N_16056,N_16740);
and U17141 (N_17141,N_16569,N_16642);
and U17142 (N_17142,N_16123,N_16998);
and U17143 (N_17143,N_16442,N_16171);
nand U17144 (N_17144,N_16674,N_16685);
nor U17145 (N_17145,N_16467,N_16960);
nor U17146 (N_17146,N_16966,N_16539);
xor U17147 (N_17147,N_16426,N_16956);
nor U17148 (N_17148,N_16994,N_16037);
and U17149 (N_17149,N_16232,N_16973);
and U17150 (N_17150,N_16355,N_16715);
and U17151 (N_17151,N_16596,N_16804);
nor U17152 (N_17152,N_16295,N_16358);
or U17153 (N_17153,N_16433,N_16243);
xor U17154 (N_17154,N_16329,N_16592);
nor U17155 (N_17155,N_16036,N_16304);
nand U17156 (N_17156,N_16927,N_16132);
nand U17157 (N_17157,N_16485,N_16727);
nor U17158 (N_17158,N_16088,N_16257);
nand U17159 (N_17159,N_16692,N_16373);
or U17160 (N_17160,N_16741,N_16440);
or U17161 (N_17161,N_16600,N_16643);
and U17162 (N_17162,N_16187,N_16258);
or U17163 (N_17163,N_16131,N_16318);
xnor U17164 (N_17164,N_16084,N_16878);
nor U17165 (N_17165,N_16947,N_16992);
xnor U17166 (N_17166,N_16964,N_16991);
nand U17167 (N_17167,N_16315,N_16425);
xor U17168 (N_17168,N_16621,N_16858);
and U17169 (N_17169,N_16656,N_16081);
nand U17170 (N_17170,N_16690,N_16519);
or U17171 (N_17171,N_16936,N_16838);
xnor U17172 (N_17172,N_16603,N_16444);
nor U17173 (N_17173,N_16612,N_16196);
nand U17174 (N_17174,N_16921,N_16739);
xor U17175 (N_17175,N_16265,N_16197);
xor U17176 (N_17176,N_16959,N_16231);
nand U17177 (N_17177,N_16079,N_16899);
xor U17178 (N_17178,N_16598,N_16346);
nand U17179 (N_17179,N_16648,N_16568);
nor U17180 (N_17180,N_16244,N_16763);
or U17181 (N_17181,N_16586,N_16611);
nand U17182 (N_17182,N_16507,N_16535);
nand U17183 (N_17183,N_16521,N_16160);
xnor U17184 (N_17184,N_16252,N_16699);
and U17185 (N_17185,N_16802,N_16234);
xnor U17186 (N_17186,N_16736,N_16503);
xor U17187 (N_17187,N_16002,N_16890);
nand U17188 (N_17188,N_16260,N_16943);
and U17189 (N_17189,N_16924,N_16867);
nand U17190 (N_17190,N_16174,N_16833);
or U17191 (N_17191,N_16023,N_16455);
xnor U17192 (N_17192,N_16085,N_16344);
xor U17193 (N_17193,N_16534,N_16212);
or U17194 (N_17194,N_16892,N_16797);
nand U17195 (N_17195,N_16422,N_16848);
and U17196 (N_17196,N_16602,N_16567);
nor U17197 (N_17197,N_16820,N_16463);
xor U17198 (N_17198,N_16868,N_16336);
nor U17199 (N_17199,N_16386,N_16057);
and U17200 (N_17200,N_16473,N_16718);
and U17201 (N_17201,N_16932,N_16175);
xnor U17202 (N_17202,N_16734,N_16894);
and U17203 (N_17203,N_16538,N_16925);
or U17204 (N_17204,N_16375,N_16719);
or U17205 (N_17205,N_16067,N_16919);
xor U17206 (N_17206,N_16136,N_16750);
nand U17207 (N_17207,N_16063,N_16167);
nor U17208 (N_17208,N_16048,N_16312);
nor U17209 (N_17209,N_16843,N_16264);
nor U17210 (N_17210,N_16657,N_16819);
nand U17211 (N_17211,N_16321,N_16465);
nor U17212 (N_17212,N_16458,N_16853);
nor U17213 (N_17213,N_16139,N_16787);
xor U17214 (N_17214,N_16909,N_16786);
nand U17215 (N_17215,N_16548,N_16933);
xnor U17216 (N_17216,N_16039,N_16099);
and U17217 (N_17217,N_16466,N_16730);
nand U17218 (N_17218,N_16683,N_16385);
and U17219 (N_17219,N_16371,N_16410);
xor U17220 (N_17220,N_16409,N_16522);
or U17221 (N_17221,N_16186,N_16220);
xnor U17222 (N_17222,N_16070,N_16356);
nor U17223 (N_17223,N_16148,N_16387);
xor U17224 (N_17224,N_16578,N_16012);
xnor U17225 (N_17225,N_16481,N_16713);
nand U17226 (N_17226,N_16156,N_16362);
nor U17227 (N_17227,N_16266,N_16747);
and U17228 (N_17228,N_16214,N_16914);
xor U17229 (N_17229,N_16775,N_16193);
nor U17230 (N_17230,N_16681,N_16758);
nor U17231 (N_17231,N_16008,N_16549);
nor U17232 (N_17232,N_16093,N_16589);
and U17233 (N_17233,N_16374,N_16398);
xor U17234 (N_17234,N_16369,N_16934);
nor U17235 (N_17235,N_16844,N_16760);
or U17236 (N_17236,N_16584,N_16161);
and U17237 (N_17237,N_16581,N_16793);
and U17238 (N_17238,N_16505,N_16547);
and U17239 (N_17239,N_16702,N_16508);
or U17240 (N_17240,N_16624,N_16146);
xnor U17241 (N_17241,N_16185,N_16179);
nand U17242 (N_17242,N_16560,N_16622);
nand U17243 (N_17243,N_16939,N_16407);
or U17244 (N_17244,N_16593,N_16427);
nand U17245 (N_17245,N_16895,N_16544);
nand U17246 (N_17246,N_16951,N_16834);
nand U17247 (N_17247,N_16013,N_16296);
nand U17248 (N_17248,N_16141,N_16053);
or U17249 (N_17249,N_16046,N_16306);
nand U17250 (N_17250,N_16883,N_16286);
nor U17251 (N_17251,N_16450,N_16906);
xnor U17252 (N_17252,N_16764,N_16077);
nor U17253 (N_17253,N_16977,N_16828);
nor U17254 (N_17254,N_16695,N_16700);
and U17255 (N_17255,N_16377,N_16694);
nor U17256 (N_17256,N_16034,N_16353);
or U17257 (N_17257,N_16807,N_16969);
nor U17258 (N_17258,N_16184,N_16121);
or U17259 (N_17259,N_16206,N_16776);
and U17260 (N_17260,N_16020,N_16794);
xnor U17261 (N_17261,N_16445,N_16235);
or U17262 (N_17262,N_16138,N_16394);
xor U17263 (N_17263,N_16813,N_16869);
or U17264 (N_17264,N_16873,N_16506);
xnor U17265 (N_17265,N_16294,N_16224);
nor U17266 (N_17266,N_16995,N_16475);
xor U17267 (N_17267,N_16064,N_16227);
xnor U17268 (N_17268,N_16831,N_16110);
nor U17269 (N_17269,N_16472,N_16835);
nor U17270 (N_17270,N_16434,N_16491);
and U17271 (N_17271,N_16588,N_16630);
xor U17272 (N_17272,N_16126,N_16177);
nand U17273 (N_17273,N_16262,N_16115);
or U17274 (N_17274,N_16940,N_16832);
and U17275 (N_17275,N_16738,N_16682);
or U17276 (N_17276,N_16107,N_16708);
nor U17277 (N_17277,N_16192,N_16106);
nor U17278 (N_17278,N_16655,N_16035);
nand U17279 (N_17279,N_16571,N_16041);
and U17280 (N_17280,N_16381,N_16840);
nor U17281 (N_17281,N_16211,N_16650);
or U17282 (N_17282,N_16404,N_16348);
and U17283 (N_17283,N_16406,N_16483);
and U17284 (N_17284,N_16273,N_16753);
nor U17285 (N_17285,N_16857,N_16144);
xor U17286 (N_17286,N_16089,N_16652);
or U17287 (N_17287,N_16199,N_16783);
or U17288 (N_17288,N_16222,N_16900);
or U17289 (N_17289,N_16737,N_16052);
or U17290 (N_17290,N_16018,N_16327);
nand U17291 (N_17291,N_16524,N_16380);
xnor U17292 (N_17292,N_16142,N_16997);
xor U17293 (N_17293,N_16284,N_16553);
xnor U17294 (N_17294,N_16393,N_16529);
and U17295 (N_17295,N_16552,N_16050);
nand U17296 (N_17296,N_16090,N_16974);
xnor U17297 (N_17297,N_16852,N_16414);
and U17298 (N_17298,N_16979,N_16885);
and U17299 (N_17299,N_16097,N_16791);
nand U17300 (N_17300,N_16563,N_16918);
nand U17301 (N_17301,N_16662,N_16270);
or U17302 (N_17302,N_16114,N_16651);
nand U17303 (N_17303,N_16365,N_16239);
nand U17304 (N_17304,N_16668,N_16839);
and U17305 (N_17305,N_16278,N_16360);
and U17306 (N_17306,N_16765,N_16976);
or U17307 (N_17307,N_16705,N_16941);
xnor U17308 (N_17308,N_16942,N_16109);
or U17309 (N_17309,N_16915,N_16766);
nor U17310 (N_17310,N_16207,N_16543);
or U17311 (N_17311,N_16597,N_16328);
nand U17312 (N_17312,N_16300,N_16806);
or U17313 (N_17313,N_16417,N_16245);
and U17314 (N_17314,N_16439,N_16686);
nor U17315 (N_17315,N_16101,N_16180);
and U17316 (N_17316,N_16233,N_16397);
and U17317 (N_17317,N_16745,N_16125);
xnor U17318 (N_17318,N_16372,N_16477);
or U17319 (N_17319,N_16929,N_16172);
xor U17320 (N_17320,N_16922,N_16953);
xor U17321 (N_17321,N_16996,N_16827);
and U17322 (N_17322,N_16582,N_16768);
xnor U17323 (N_17323,N_16579,N_16268);
nand U17324 (N_17324,N_16572,N_16341);
xnor U17325 (N_17325,N_16017,N_16217);
and U17326 (N_17326,N_16874,N_16812);
or U17327 (N_17327,N_16190,N_16059);
nor U17328 (N_17328,N_16376,N_16149);
nor U17329 (N_17329,N_16527,N_16150);
and U17330 (N_17330,N_16958,N_16208);
or U17331 (N_17331,N_16337,N_16357);
and U17332 (N_17332,N_16605,N_16886);
or U17333 (N_17333,N_16205,N_16469);
nand U17334 (N_17334,N_16946,N_16432);
and U17335 (N_17335,N_16965,N_16902);
or U17336 (N_17336,N_16395,N_16664);
or U17337 (N_17337,N_16716,N_16420);
and U17338 (N_17338,N_16408,N_16949);
xnor U17339 (N_17339,N_16200,N_16043);
or U17340 (N_17340,N_16644,N_16261);
or U17341 (N_17341,N_16152,N_16178);
nand U17342 (N_17342,N_16333,N_16051);
and U17343 (N_17343,N_16810,N_16100);
nand U17344 (N_17344,N_16276,N_16250);
or U17345 (N_17345,N_16637,N_16498);
nand U17346 (N_17346,N_16721,N_16952);
nand U17347 (N_17347,N_16903,N_16717);
and U17348 (N_17348,N_16038,N_16392);
nor U17349 (N_17349,N_16749,N_16631);
nor U17350 (N_17350,N_16202,N_16267);
and U17351 (N_17351,N_16461,N_16026);
or U17352 (N_17352,N_16288,N_16159);
xnor U17353 (N_17353,N_16158,N_16279);
nand U17354 (N_17354,N_16045,N_16767);
and U17355 (N_17355,N_16646,N_16451);
and U17356 (N_17356,N_16378,N_16859);
nand U17357 (N_17357,N_16907,N_16961);
xor U17358 (N_17358,N_16759,N_16251);
xor U17359 (N_17359,N_16725,N_16663);
nand U17360 (N_17360,N_16135,N_16226);
nand U17361 (N_17361,N_16550,N_16218);
xnor U17362 (N_17362,N_16545,N_16363);
and U17363 (N_17363,N_16128,N_16757);
nand U17364 (N_17364,N_16120,N_16805);
or U17365 (N_17365,N_16075,N_16826);
nand U17366 (N_17366,N_16945,N_16566);
or U17367 (N_17367,N_16887,N_16402);
xnor U17368 (N_17368,N_16396,N_16905);
and U17369 (N_17369,N_16423,N_16599);
or U17370 (N_17370,N_16352,N_16515);
and U17371 (N_17371,N_16754,N_16893);
xnor U17372 (N_17372,N_16877,N_16784);
nand U17373 (N_17373,N_16799,N_16854);
and U17374 (N_17374,N_16219,N_16698);
or U17375 (N_17375,N_16559,N_16470);
nor U17376 (N_17376,N_16317,N_16537);
and U17377 (N_17377,N_16908,N_16418);
xnor U17378 (N_17378,N_16459,N_16028);
and U17379 (N_17379,N_16667,N_16334);
nand U17380 (N_17380,N_16707,N_16274);
xnor U17381 (N_17381,N_16723,N_16703);
and U17382 (N_17382,N_16313,N_16653);
and U17383 (N_17383,N_16349,N_16354);
nor U17384 (N_17384,N_16323,N_16714);
or U17385 (N_17385,N_16401,N_16391);
nand U17386 (N_17386,N_16555,N_16781);
and U17387 (N_17387,N_16704,N_16627);
or U17388 (N_17388,N_16129,N_16330);
xnor U17389 (N_17389,N_16870,N_16364);
and U17390 (N_17390,N_16389,N_16541);
nor U17391 (N_17391,N_16379,N_16275);
nor U17392 (N_17392,N_16796,N_16441);
nand U17393 (N_17393,N_16772,N_16728);
and U17394 (N_17394,N_16215,N_16298);
and U17395 (N_17395,N_16194,N_16060);
nand U17396 (N_17396,N_16169,N_16412);
nor U17397 (N_17397,N_16388,N_16102);
and U17398 (N_17398,N_16438,N_16430);
nor U17399 (N_17399,N_16821,N_16623);
and U17400 (N_17400,N_16770,N_16926);
or U17401 (N_17401,N_16151,N_16443);
or U17402 (N_17402,N_16855,N_16080);
nor U17403 (N_17403,N_16836,N_16249);
nor U17404 (N_17404,N_16320,N_16236);
xor U17405 (N_17405,N_16367,N_16962);
and U17406 (N_17406,N_16689,N_16325);
and U17407 (N_17407,N_16066,N_16814);
nand U17408 (N_17408,N_16482,N_16533);
nor U17409 (N_17409,N_16641,N_16701);
or U17410 (N_17410,N_16845,N_16095);
nor U17411 (N_17411,N_16647,N_16720);
or U17412 (N_17412,N_16864,N_16841);
nand U17413 (N_17413,N_16554,N_16499);
and U17414 (N_17414,N_16116,N_16452);
xor U17415 (N_17415,N_16684,N_16577);
or U17416 (N_17416,N_16188,N_16729);
and U17417 (N_17417,N_16889,N_16238);
and U17418 (N_17418,N_16896,N_16751);
nor U17419 (N_17419,N_16575,N_16860);
and U17420 (N_17420,N_16680,N_16993);
nor U17421 (N_17421,N_16340,N_16777);
nor U17422 (N_17422,N_16464,N_16629);
and U17423 (N_17423,N_16454,N_16335);
nand U17424 (N_17424,N_16950,N_16293);
and U17425 (N_17425,N_16011,N_16988);
or U17426 (N_17426,N_16888,N_16301);
and U17427 (N_17427,N_16092,N_16913);
nand U17428 (N_17428,N_16259,N_16619);
nand U17429 (N_17429,N_16609,N_16405);
or U17430 (N_17430,N_16021,N_16625);
nor U17431 (N_17431,N_16532,N_16561);
nand U17432 (N_17432,N_16484,N_16182);
nor U17433 (N_17433,N_16604,N_16916);
xor U17434 (N_17434,N_16390,N_16042);
nand U17435 (N_17435,N_16670,N_16157);
nand U17436 (N_17436,N_16678,N_16437);
nand U17437 (N_17437,N_16297,N_16606);
nand U17438 (N_17438,N_16071,N_16311);
and U17439 (N_17439,N_16014,N_16383);
nand U17440 (N_17440,N_16626,N_16133);
xnor U17441 (N_17441,N_16054,N_16968);
xnor U17442 (N_17442,N_16614,N_16240);
or U17443 (N_17443,N_16930,N_16076);
nor U17444 (N_17444,N_16898,N_16659);
or U17445 (N_17445,N_16671,N_16460);
xor U17446 (N_17446,N_16516,N_16931);
xnor U17447 (N_17447,N_16938,N_16980);
and U17448 (N_17448,N_16069,N_16865);
or U17449 (N_17449,N_16347,N_16761);
nand U17450 (N_17450,N_16955,N_16520);
and U17451 (N_17451,N_16191,N_16706);
xor U17452 (N_17452,N_16748,N_16687);
nor U17453 (N_17453,N_16166,N_16871);
nand U17454 (N_17454,N_16879,N_16299);
nand U17455 (N_17455,N_16163,N_16168);
nand U17456 (N_17456,N_16345,N_16399);
nand U17457 (N_17457,N_16872,N_16246);
xor U17458 (N_17458,N_16446,N_16654);
and U17459 (N_17459,N_16255,N_16024);
nand U17460 (N_17460,N_16752,N_16628);
nor U17461 (N_17461,N_16496,N_16798);
or U17462 (N_17462,N_16082,N_16967);
nor U17463 (N_17463,N_16448,N_16006);
xnor U17464 (N_17464,N_16963,N_16722);
or U17465 (N_17465,N_16984,N_16436);
nor U17466 (N_17466,N_16842,N_16691);
nor U17467 (N_17467,N_16711,N_16384);
or U17468 (N_17468,N_16415,N_16502);
nand U17469 (N_17469,N_16229,N_16154);
or U17470 (N_17470,N_16917,N_16975);
and U17471 (N_17471,N_16209,N_16230);
nand U17472 (N_17472,N_16987,N_16989);
xnor U17473 (N_17473,N_16277,N_16493);
or U17474 (N_17474,N_16487,N_16307);
xor U17475 (N_17475,N_16658,N_16856);
nor U17476 (N_17476,N_16981,N_16677);
or U17477 (N_17477,N_16528,N_16216);
nor U17478 (N_17478,N_16633,N_16607);
or U17479 (N_17479,N_16509,N_16400);
nor U17480 (N_17480,N_16851,N_16829);
or U17481 (N_17481,N_16557,N_16620);
or U17482 (N_17482,N_16305,N_16636);
nand U17483 (N_17483,N_16504,N_16640);
nand U17484 (N_17484,N_16525,N_16675);
and U17485 (N_17485,N_16616,N_16911);
and U17486 (N_17486,N_16817,N_16513);
xor U17487 (N_17487,N_16189,N_16863);
and U17488 (N_17488,N_16112,N_16025);
nor U17489 (N_17489,N_16613,N_16010);
nand U17490 (N_17490,N_16697,N_16901);
xor U17491 (N_17491,N_16308,N_16314);
nor U17492 (N_17492,N_16800,N_16815);
and U17493 (N_17493,N_16882,N_16881);
or U17494 (N_17494,N_16542,N_16551);
or U17495 (N_17495,N_16762,N_16309);
nor U17496 (N_17496,N_16058,N_16280);
nor U17497 (N_17497,N_16564,N_16225);
or U17498 (N_17498,N_16999,N_16324);
xnor U17499 (N_17499,N_16003,N_16203);
or U17500 (N_17500,N_16553,N_16326);
nand U17501 (N_17501,N_16017,N_16231);
or U17502 (N_17502,N_16160,N_16112);
xor U17503 (N_17503,N_16513,N_16780);
nand U17504 (N_17504,N_16169,N_16652);
nand U17505 (N_17505,N_16546,N_16357);
nand U17506 (N_17506,N_16120,N_16784);
nand U17507 (N_17507,N_16053,N_16492);
and U17508 (N_17508,N_16604,N_16304);
and U17509 (N_17509,N_16560,N_16555);
nand U17510 (N_17510,N_16256,N_16351);
or U17511 (N_17511,N_16540,N_16423);
xor U17512 (N_17512,N_16348,N_16762);
or U17513 (N_17513,N_16377,N_16552);
xnor U17514 (N_17514,N_16584,N_16383);
or U17515 (N_17515,N_16121,N_16873);
nor U17516 (N_17516,N_16857,N_16487);
or U17517 (N_17517,N_16222,N_16286);
and U17518 (N_17518,N_16718,N_16879);
and U17519 (N_17519,N_16131,N_16632);
nor U17520 (N_17520,N_16540,N_16851);
and U17521 (N_17521,N_16853,N_16299);
and U17522 (N_17522,N_16329,N_16456);
and U17523 (N_17523,N_16814,N_16272);
xnor U17524 (N_17524,N_16706,N_16599);
xnor U17525 (N_17525,N_16510,N_16688);
nand U17526 (N_17526,N_16984,N_16835);
nor U17527 (N_17527,N_16378,N_16438);
or U17528 (N_17528,N_16070,N_16169);
xor U17529 (N_17529,N_16592,N_16131);
or U17530 (N_17530,N_16412,N_16086);
or U17531 (N_17531,N_16748,N_16202);
xor U17532 (N_17532,N_16547,N_16461);
nand U17533 (N_17533,N_16405,N_16942);
nor U17534 (N_17534,N_16710,N_16929);
nand U17535 (N_17535,N_16838,N_16466);
nand U17536 (N_17536,N_16516,N_16548);
and U17537 (N_17537,N_16181,N_16375);
or U17538 (N_17538,N_16851,N_16603);
nor U17539 (N_17539,N_16127,N_16195);
nor U17540 (N_17540,N_16652,N_16425);
and U17541 (N_17541,N_16497,N_16857);
or U17542 (N_17542,N_16854,N_16520);
nor U17543 (N_17543,N_16301,N_16527);
or U17544 (N_17544,N_16729,N_16069);
nor U17545 (N_17545,N_16449,N_16513);
or U17546 (N_17546,N_16482,N_16736);
or U17547 (N_17547,N_16241,N_16553);
and U17548 (N_17548,N_16128,N_16405);
nor U17549 (N_17549,N_16843,N_16524);
or U17550 (N_17550,N_16085,N_16668);
or U17551 (N_17551,N_16317,N_16380);
nand U17552 (N_17552,N_16645,N_16202);
nand U17553 (N_17553,N_16482,N_16692);
nor U17554 (N_17554,N_16907,N_16292);
xor U17555 (N_17555,N_16278,N_16922);
nand U17556 (N_17556,N_16342,N_16479);
or U17557 (N_17557,N_16385,N_16512);
or U17558 (N_17558,N_16849,N_16274);
nand U17559 (N_17559,N_16960,N_16690);
or U17560 (N_17560,N_16731,N_16576);
and U17561 (N_17561,N_16340,N_16239);
nor U17562 (N_17562,N_16587,N_16921);
and U17563 (N_17563,N_16464,N_16146);
or U17564 (N_17564,N_16536,N_16484);
and U17565 (N_17565,N_16685,N_16429);
xor U17566 (N_17566,N_16287,N_16440);
xor U17567 (N_17567,N_16106,N_16928);
xnor U17568 (N_17568,N_16311,N_16770);
or U17569 (N_17569,N_16991,N_16957);
or U17570 (N_17570,N_16905,N_16256);
or U17571 (N_17571,N_16941,N_16604);
xnor U17572 (N_17572,N_16628,N_16896);
and U17573 (N_17573,N_16283,N_16709);
nor U17574 (N_17574,N_16135,N_16332);
xor U17575 (N_17575,N_16612,N_16368);
xor U17576 (N_17576,N_16733,N_16099);
and U17577 (N_17577,N_16901,N_16612);
nand U17578 (N_17578,N_16033,N_16109);
nor U17579 (N_17579,N_16827,N_16176);
xor U17580 (N_17580,N_16676,N_16663);
xnor U17581 (N_17581,N_16860,N_16414);
and U17582 (N_17582,N_16142,N_16350);
nor U17583 (N_17583,N_16274,N_16598);
xnor U17584 (N_17584,N_16036,N_16804);
and U17585 (N_17585,N_16221,N_16544);
or U17586 (N_17586,N_16805,N_16554);
nand U17587 (N_17587,N_16355,N_16607);
nand U17588 (N_17588,N_16858,N_16809);
nor U17589 (N_17589,N_16185,N_16592);
or U17590 (N_17590,N_16129,N_16056);
nand U17591 (N_17591,N_16293,N_16599);
nand U17592 (N_17592,N_16507,N_16945);
or U17593 (N_17593,N_16568,N_16369);
nor U17594 (N_17594,N_16695,N_16739);
or U17595 (N_17595,N_16033,N_16500);
nand U17596 (N_17596,N_16021,N_16714);
nor U17597 (N_17597,N_16887,N_16406);
and U17598 (N_17598,N_16816,N_16759);
nand U17599 (N_17599,N_16389,N_16919);
and U17600 (N_17600,N_16174,N_16245);
or U17601 (N_17601,N_16111,N_16772);
nand U17602 (N_17602,N_16374,N_16682);
nand U17603 (N_17603,N_16013,N_16265);
and U17604 (N_17604,N_16284,N_16679);
and U17605 (N_17605,N_16622,N_16134);
nand U17606 (N_17606,N_16390,N_16905);
nor U17607 (N_17607,N_16166,N_16690);
or U17608 (N_17608,N_16986,N_16313);
xor U17609 (N_17609,N_16576,N_16162);
nor U17610 (N_17610,N_16147,N_16519);
xor U17611 (N_17611,N_16232,N_16655);
xor U17612 (N_17612,N_16756,N_16921);
and U17613 (N_17613,N_16697,N_16885);
xnor U17614 (N_17614,N_16889,N_16025);
nor U17615 (N_17615,N_16673,N_16330);
nand U17616 (N_17616,N_16409,N_16850);
or U17617 (N_17617,N_16291,N_16178);
xor U17618 (N_17618,N_16914,N_16389);
xnor U17619 (N_17619,N_16068,N_16834);
nand U17620 (N_17620,N_16778,N_16648);
and U17621 (N_17621,N_16529,N_16017);
and U17622 (N_17622,N_16537,N_16212);
nand U17623 (N_17623,N_16075,N_16445);
and U17624 (N_17624,N_16718,N_16184);
nor U17625 (N_17625,N_16913,N_16918);
nand U17626 (N_17626,N_16264,N_16536);
nor U17627 (N_17627,N_16041,N_16238);
xor U17628 (N_17628,N_16281,N_16052);
nor U17629 (N_17629,N_16253,N_16474);
nor U17630 (N_17630,N_16363,N_16458);
xor U17631 (N_17631,N_16980,N_16338);
and U17632 (N_17632,N_16328,N_16163);
and U17633 (N_17633,N_16770,N_16121);
xor U17634 (N_17634,N_16478,N_16234);
or U17635 (N_17635,N_16079,N_16924);
and U17636 (N_17636,N_16407,N_16581);
nor U17637 (N_17637,N_16961,N_16158);
nand U17638 (N_17638,N_16709,N_16838);
nand U17639 (N_17639,N_16361,N_16117);
xnor U17640 (N_17640,N_16137,N_16507);
or U17641 (N_17641,N_16500,N_16090);
nand U17642 (N_17642,N_16689,N_16573);
nor U17643 (N_17643,N_16756,N_16850);
nor U17644 (N_17644,N_16450,N_16989);
and U17645 (N_17645,N_16618,N_16555);
nor U17646 (N_17646,N_16156,N_16002);
or U17647 (N_17647,N_16015,N_16669);
nor U17648 (N_17648,N_16354,N_16899);
nand U17649 (N_17649,N_16213,N_16957);
xnor U17650 (N_17650,N_16703,N_16338);
nand U17651 (N_17651,N_16358,N_16293);
xor U17652 (N_17652,N_16285,N_16918);
or U17653 (N_17653,N_16012,N_16483);
and U17654 (N_17654,N_16185,N_16277);
or U17655 (N_17655,N_16652,N_16135);
xor U17656 (N_17656,N_16539,N_16527);
xnor U17657 (N_17657,N_16727,N_16889);
or U17658 (N_17658,N_16312,N_16332);
nor U17659 (N_17659,N_16759,N_16091);
or U17660 (N_17660,N_16212,N_16913);
and U17661 (N_17661,N_16494,N_16026);
nand U17662 (N_17662,N_16126,N_16590);
or U17663 (N_17663,N_16156,N_16323);
xnor U17664 (N_17664,N_16909,N_16891);
or U17665 (N_17665,N_16018,N_16767);
xnor U17666 (N_17666,N_16239,N_16476);
or U17667 (N_17667,N_16643,N_16859);
nand U17668 (N_17668,N_16512,N_16602);
xor U17669 (N_17669,N_16641,N_16271);
or U17670 (N_17670,N_16306,N_16814);
and U17671 (N_17671,N_16431,N_16507);
nand U17672 (N_17672,N_16984,N_16407);
nand U17673 (N_17673,N_16129,N_16335);
or U17674 (N_17674,N_16282,N_16342);
or U17675 (N_17675,N_16560,N_16201);
nand U17676 (N_17676,N_16251,N_16984);
or U17677 (N_17677,N_16252,N_16865);
or U17678 (N_17678,N_16028,N_16653);
nand U17679 (N_17679,N_16803,N_16377);
and U17680 (N_17680,N_16845,N_16318);
and U17681 (N_17681,N_16486,N_16297);
nor U17682 (N_17682,N_16565,N_16906);
and U17683 (N_17683,N_16539,N_16389);
xor U17684 (N_17684,N_16471,N_16791);
nand U17685 (N_17685,N_16415,N_16340);
nor U17686 (N_17686,N_16066,N_16905);
nor U17687 (N_17687,N_16499,N_16841);
nor U17688 (N_17688,N_16388,N_16908);
and U17689 (N_17689,N_16405,N_16740);
and U17690 (N_17690,N_16198,N_16066);
and U17691 (N_17691,N_16745,N_16806);
and U17692 (N_17692,N_16702,N_16185);
nand U17693 (N_17693,N_16022,N_16303);
and U17694 (N_17694,N_16620,N_16477);
xnor U17695 (N_17695,N_16098,N_16228);
and U17696 (N_17696,N_16708,N_16672);
xnor U17697 (N_17697,N_16271,N_16984);
or U17698 (N_17698,N_16373,N_16785);
nand U17699 (N_17699,N_16154,N_16383);
nor U17700 (N_17700,N_16885,N_16859);
nand U17701 (N_17701,N_16405,N_16017);
or U17702 (N_17702,N_16074,N_16017);
or U17703 (N_17703,N_16969,N_16317);
xor U17704 (N_17704,N_16459,N_16744);
nor U17705 (N_17705,N_16581,N_16300);
xor U17706 (N_17706,N_16617,N_16192);
xnor U17707 (N_17707,N_16627,N_16053);
nand U17708 (N_17708,N_16781,N_16108);
nor U17709 (N_17709,N_16463,N_16254);
nor U17710 (N_17710,N_16123,N_16656);
nand U17711 (N_17711,N_16961,N_16489);
and U17712 (N_17712,N_16269,N_16794);
xor U17713 (N_17713,N_16250,N_16569);
or U17714 (N_17714,N_16127,N_16784);
nand U17715 (N_17715,N_16278,N_16952);
and U17716 (N_17716,N_16014,N_16941);
xor U17717 (N_17717,N_16304,N_16079);
nor U17718 (N_17718,N_16707,N_16498);
and U17719 (N_17719,N_16272,N_16173);
xor U17720 (N_17720,N_16624,N_16140);
nand U17721 (N_17721,N_16371,N_16038);
xnor U17722 (N_17722,N_16480,N_16538);
and U17723 (N_17723,N_16913,N_16988);
or U17724 (N_17724,N_16968,N_16766);
xnor U17725 (N_17725,N_16220,N_16580);
or U17726 (N_17726,N_16435,N_16790);
nor U17727 (N_17727,N_16413,N_16999);
nor U17728 (N_17728,N_16008,N_16276);
xnor U17729 (N_17729,N_16640,N_16850);
or U17730 (N_17730,N_16231,N_16462);
nor U17731 (N_17731,N_16282,N_16796);
nand U17732 (N_17732,N_16535,N_16889);
nor U17733 (N_17733,N_16315,N_16002);
and U17734 (N_17734,N_16056,N_16154);
nor U17735 (N_17735,N_16749,N_16712);
and U17736 (N_17736,N_16492,N_16983);
xor U17737 (N_17737,N_16807,N_16442);
or U17738 (N_17738,N_16940,N_16301);
nand U17739 (N_17739,N_16907,N_16781);
and U17740 (N_17740,N_16420,N_16534);
nand U17741 (N_17741,N_16290,N_16551);
nand U17742 (N_17742,N_16363,N_16512);
nor U17743 (N_17743,N_16798,N_16203);
xnor U17744 (N_17744,N_16768,N_16396);
nor U17745 (N_17745,N_16184,N_16509);
nand U17746 (N_17746,N_16413,N_16512);
xor U17747 (N_17747,N_16670,N_16843);
nand U17748 (N_17748,N_16261,N_16457);
and U17749 (N_17749,N_16768,N_16061);
nor U17750 (N_17750,N_16397,N_16469);
and U17751 (N_17751,N_16688,N_16917);
xnor U17752 (N_17752,N_16343,N_16025);
and U17753 (N_17753,N_16740,N_16297);
and U17754 (N_17754,N_16631,N_16473);
or U17755 (N_17755,N_16023,N_16395);
xor U17756 (N_17756,N_16368,N_16660);
nand U17757 (N_17757,N_16629,N_16120);
and U17758 (N_17758,N_16796,N_16183);
and U17759 (N_17759,N_16832,N_16689);
and U17760 (N_17760,N_16938,N_16072);
nand U17761 (N_17761,N_16892,N_16331);
or U17762 (N_17762,N_16933,N_16209);
xor U17763 (N_17763,N_16029,N_16783);
nor U17764 (N_17764,N_16456,N_16757);
or U17765 (N_17765,N_16954,N_16281);
xnor U17766 (N_17766,N_16329,N_16773);
or U17767 (N_17767,N_16448,N_16286);
xor U17768 (N_17768,N_16465,N_16224);
xor U17769 (N_17769,N_16281,N_16612);
or U17770 (N_17770,N_16983,N_16521);
xnor U17771 (N_17771,N_16026,N_16056);
nor U17772 (N_17772,N_16777,N_16936);
xor U17773 (N_17773,N_16459,N_16470);
or U17774 (N_17774,N_16197,N_16534);
xnor U17775 (N_17775,N_16237,N_16821);
or U17776 (N_17776,N_16523,N_16946);
or U17777 (N_17777,N_16975,N_16737);
or U17778 (N_17778,N_16509,N_16467);
nor U17779 (N_17779,N_16921,N_16133);
xnor U17780 (N_17780,N_16150,N_16665);
nand U17781 (N_17781,N_16676,N_16762);
nand U17782 (N_17782,N_16085,N_16664);
nor U17783 (N_17783,N_16984,N_16772);
and U17784 (N_17784,N_16354,N_16287);
or U17785 (N_17785,N_16392,N_16295);
xnor U17786 (N_17786,N_16059,N_16116);
nor U17787 (N_17787,N_16252,N_16431);
xor U17788 (N_17788,N_16986,N_16835);
nand U17789 (N_17789,N_16247,N_16581);
and U17790 (N_17790,N_16199,N_16291);
and U17791 (N_17791,N_16080,N_16366);
nor U17792 (N_17792,N_16050,N_16338);
nor U17793 (N_17793,N_16449,N_16212);
xor U17794 (N_17794,N_16499,N_16647);
or U17795 (N_17795,N_16754,N_16816);
or U17796 (N_17796,N_16580,N_16918);
xnor U17797 (N_17797,N_16751,N_16063);
and U17798 (N_17798,N_16356,N_16254);
and U17799 (N_17799,N_16888,N_16165);
nor U17800 (N_17800,N_16192,N_16052);
xnor U17801 (N_17801,N_16297,N_16689);
xor U17802 (N_17802,N_16375,N_16775);
nor U17803 (N_17803,N_16471,N_16474);
and U17804 (N_17804,N_16131,N_16975);
xor U17805 (N_17805,N_16881,N_16230);
xor U17806 (N_17806,N_16242,N_16221);
nand U17807 (N_17807,N_16440,N_16395);
xnor U17808 (N_17808,N_16580,N_16845);
xnor U17809 (N_17809,N_16262,N_16763);
nand U17810 (N_17810,N_16669,N_16437);
or U17811 (N_17811,N_16748,N_16575);
or U17812 (N_17812,N_16474,N_16066);
nand U17813 (N_17813,N_16009,N_16930);
xnor U17814 (N_17814,N_16675,N_16145);
xnor U17815 (N_17815,N_16723,N_16059);
nor U17816 (N_17816,N_16434,N_16142);
nor U17817 (N_17817,N_16012,N_16526);
xor U17818 (N_17818,N_16023,N_16147);
nor U17819 (N_17819,N_16084,N_16294);
or U17820 (N_17820,N_16625,N_16188);
and U17821 (N_17821,N_16476,N_16437);
nor U17822 (N_17822,N_16929,N_16222);
nand U17823 (N_17823,N_16846,N_16962);
nor U17824 (N_17824,N_16205,N_16321);
nand U17825 (N_17825,N_16469,N_16353);
and U17826 (N_17826,N_16214,N_16172);
or U17827 (N_17827,N_16180,N_16338);
and U17828 (N_17828,N_16006,N_16659);
nor U17829 (N_17829,N_16607,N_16869);
nand U17830 (N_17830,N_16291,N_16701);
nor U17831 (N_17831,N_16958,N_16786);
nand U17832 (N_17832,N_16114,N_16685);
or U17833 (N_17833,N_16966,N_16623);
xor U17834 (N_17834,N_16124,N_16070);
or U17835 (N_17835,N_16697,N_16788);
nor U17836 (N_17836,N_16554,N_16465);
and U17837 (N_17837,N_16513,N_16336);
nand U17838 (N_17838,N_16628,N_16652);
or U17839 (N_17839,N_16854,N_16213);
and U17840 (N_17840,N_16754,N_16328);
and U17841 (N_17841,N_16511,N_16647);
and U17842 (N_17842,N_16851,N_16418);
and U17843 (N_17843,N_16202,N_16219);
nand U17844 (N_17844,N_16208,N_16731);
and U17845 (N_17845,N_16823,N_16484);
xor U17846 (N_17846,N_16839,N_16389);
xor U17847 (N_17847,N_16087,N_16682);
or U17848 (N_17848,N_16469,N_16383);
xnor U17849 (N_17849,N_16497,N_16134);
and U17850 (N_17850,N_16617,N_16204);
xor U17851 (N_17851,N_16915,N_16567);
nand U17852 (N_17852,N_16156,N_16854);
and U17853 (N_17853,N_16835,N_16037);
nand U17854 (N_17854,N_16389,N_16110);
and U17855 (N_17855,N_16917,N_16235);
or U17856 (N_17856,N_16395,N_16000);
xor U17857 (N_17857,N_16595,N_16982);
and U17858 (N_17858,N_16939,N_16594);
xor U17859 (N_17859,N_16096,N_16665);
and U17860 (N_17860,N_16838,N_16524);
nand U17861 (N_17861,N_16745,N_16566);
nor U17862 (N_17862,N_16933,N_16215);
nor U17863 (N_17863,N_16575,N_16423);
nand U17864 (N_17864,N_16041,N_16878);
nand U17865 (N_17865,N_16454,N_16443);
and U17866 (N_17866,N_16263,N_16081);
and U17867 (N_17867,N_16646,N_16896);
xnor U17868 (N_17868,N_16856,N_16919);
nand U17869 (N_17869,N_16365,N_16597);
or U17870 (N_17870,N_16547,N_16031);
xor U17871 (N_17871,N_16748,N_16625);
and U17872 (N_17872,N_16531,N_16563);
or U17873 (N_17873,N_16485,N_16174);
or U17874 (N_17874,N_16138,N_16806);
or U17875 (N_17875,N_16383,N_16145);
nor U17876 (N_17876,N_16248,N_16093);
and U17877 (N_17877,N_16098,N_16040);
nor U17878 (N_17878,N_16295,N_16551);
and U17879 (N_17879,N_16429,N_16399);
xnor U17880 (N_17880,N_16452,N_16137);
nor U17881 (N_17881,N_16765,N_16961);
nor U17882 (N_17882,N_16204,N_16777);
nand U17883 (N_17883,N_16051,N_16515);
and U17884 (N_17884,N_16554,N_16080);
xor U17885 (N_17885,N_16401,N_16296);
xnor U17886 (N_17886,N_16182,N_16921);
xor U17887 (N_17887,N_16207,N_16164);
nand U17888 (N_17888,N_16396,N_16215);
nor U17889 (N_17889,N_16420,N_16189);
xnor U17890 (N_17890,N_16233,N_16055);
xor U17891 (N_17891,N_16738,N_16455);
and U17892 (N_17892,N_16258,N_16022);
xnor U17893 (N_17893,N_16504,N_16460);
and U17894 (N_17894,N_16536,N_16415);
and U17895 (N_17895,N_16217,N_16562);
nor U17896 (N_17896,N_16038,N_16053);
nand U17897 (N_17897,N_16690,N_16937);
and U17898 (N_17898,N_16321,N_16620);
nand U17899 (N_17899,N_16265,N_16740);
nor U17900 (N_17900,N_16124,N_16302);
or U17901 (N_17901,N_16762,N_16197);
and U17902 (N_17902,N_16423,N_16133);
or U17903 (N_17903,N_16083,N_16777);
or U17904 (N_17904,N_16396,N_16174);
nand U17905 (N_17905,N_16348,N_16158);
or U17906 (N_17906,N_16112,N_16117);
or U17907 (N_17907,N_16690,N_16432);
xor U17908 (N_17908,N_16616,N_16145);
nor U17909 (N_17909,N_16666,N_16361);
or U17910 (N_17910,N_16799,N_16043);
xnor U17911 (N_17911,N_16127,N_16242);
xor U17912 (N_17912,N_16979,N_16857);
or U17913 (N_17913,N_16308,N_16812);
nor U17914 (N_17914,N_16550,N_16446);
and U17915 (N_17915,N_16082,N_16402);
nand U17916 (N_17916,N_16194,N_16833);
nor U17917 (N_17917,N_16924,N_16778);
nand U17918 (N_17918,N_16586,N_16076);
nor U17919 (N_17919,N_16262,N_16652);
and U17920 (N_17920,N_16218,N_16180);
or U17921 (N_17921,N_16891,N_16020);
or U17922 (N_17922,N_16220,N_16764);
xor U17923 (N_17923,N_16305,N_16218);
or U17924 (N_17924,N_16291,N_16883);
nor U17925 (N_17925,N_16611,N_16781);
and U17926 (N_17926,N_16693,N_16423);
nor U17927 (N_17927,N_16709,N_16387);
or U17928 (N_17928,N_16826,N_16879);
xor U17929 (N_17929,N_16228,N_16377);
xor U17930 (N_17930,N_16296,N_16076);
xnor U17931 (N_17931,N_16347,N_16198);
nand U17932 (N_17932,N_16436,N_16171);
nor U17933 (N_17933,N_16843,N_16961);
nor U17934 (N_17934,N_16868,N_16809);
xor U17935 (N_17935,N_16305,N_16826);
xnor U17936 (N_17936,N_16796,N_16701);
and U17937 (N_17937,N_16934,N_16810);
or U17938 (N_17938,N_16050,N_16520);
or U17939 (N_17939,N_16185,N_16187);
nand U17940 (N_17940,N_16276,N_16157);
nand U17941 (N_17941,N_16969,N_16131);
or U17942 (N_17942,N_16238,N_16622);
and U17943 (N_17943,N_16664,N_16723);
xnor U17944 (N_17944,N_16340,N_16701);
nor U17945 (N_17945,N_16311,N_16666);
and U17946 (N_17946,N_16867,N_16249);
nand U17947 (N_17947,N_16897,N_16158);
and U17948 (N_17948,N_16809,N_16207);
xor U17949 (N_17949,N_16948,N_16326);
xnor U17950 (N_17950,N_16603,N_16803);
nor U17951 (N_17951,N_16870,N_16447);
and U17952 (N_17952,N_16417,N_16009);
or U17953 (N_17953,N_16087,N_16906);
nor U17954 (N_17954,N_16788,N_16388);
and U17955 (N_17955,N_16563,N_16633);
xnor U17956 (N_17956,N_16974,N_16860);
nor U17957 (N_17957,N_16105,N_16304);
nor U17958 (N_17958,N_16134,N_16873);
nand U17959 (N_17959,N_16679,N_16164);
or U17960 (N_17960,N_16034,N_16009);
nand U17961 (N_17961,N_16361,N_16933);
and U17962 (N_17962,N_16843,N_16284);
or U17963 (N_17963,N_16693,N_16015);
nand U17964 (N_17964,N_16678,N_16821);
xnor U17965 (N_17965,N_16091,N_16575);
xor U17966 (N_17966,N_16158,N_16054);
xor U17967 (N_17967,N_16667,N_16674);
and U17968 (N_17968,N_16144,N_16979);
and U17969 (N_17969,N_16709,N_16115);
nor U17970 (N_17970,N_16802,N_16698);
xor U17971 (N_17971,N_16506,N_16440);
or U17972 (N_17972,N_16424,N_16775);
nand U17973 (N_17973,N_16893,N_16352);
xnor U17974 (N_17974,N_16893,N_16158);
nand U17975 (N_17975,N_16987,N_16397);
nor U17976 (N_17976,N_16702,N_16385);
or U17977 (N_17977,N_16841,N_16606);
nand U17978 (N_17978,N_16890,N_16546);
xor U17979 (N_17979,N_16761,N_16887);
and U17980 (N_17980,N_16463,N_16175);
xnor U17981 (N_17981,N_16276,N_16913);
xor U17982 (N_17982,N_16210,N_16481);
nor U17983 (N_17983,N_16629,N_16391);
xnor U17984 (N_17984,N_16843,N_16746);
xor U17985 (N_17985,N_16377,N_16988);
nand U17986 (N_17986,N_16740,N_16206);
nand U17987 (N_17987,N_16375,N_16594);
and U17988 (N_17988,N_16801,N_16628);
or U17989 (N_17989,N_16317,N_16410);
nand U17990 (N_17990,N_16392,N_16260);
nor U17991 (N_17991,N_16531,N_16166);
nor U17992 (N_17992,N_16572,N_16069);
nor U17993 (N_17993,N_16791,N_16531);
nand U17994 (N_17994,N_16460,N_16500);
xor U17995 (N_17995,N_16702,N_16032);
or U17996 (N_17996,N_16598,N_16575);
nand U17997 (N_17997,N_16926,N_16363);
nor U17998 (N_17998,N_16440,N_16611);
nand U17999 (N_17999,N_16479,N_16556);
and U18000 (N_18000,N_17370,N_17755);
xor U18001 (N_18001,N_17657,N_17814);
nor U18002 (N_18002,N_17598,N_17284);
nand U18003 (N_18003,N_17086,N_17422);
xor U18004 (N_18004,N_17184,N_17476);
or U18005 (N_18005,N_17860,N_17804);
nand U18006 (N_18006,N_17368,N_17308);
or U18007 (N_18007,N_17128,N_17219);
and U18008 (N_18008,N_17993,N_17637);
nand U18009 (N_18009,N_17578,N_17207);
and U18010 (N_18010,N_17734,N_17831);
xnor U18011 (N_18011,N_17615,N_17844);
nand U18012 (N_18012,N_17066,N_17316);
nor U18013 (N_18013,N_17740,N_17566);
or U18014 (N_18014,N_17882,N_17433);
nor U18015 (N_18015,N_17732,N_17796);
xor U18016 (N_18016,N_17183,N_17388);
and U18017 (N_18017,N_17247,N_17298);
nor U18018 (N_18018,N_17406,N_17214);
and U18019 (N_18019,N_17843,N_17285);
and U18020 (N_18020,N_17603,N_17681);
nand U18021 (N_18021,N_17594,N_17399);
or U18022 (N_18022,N_17835,N_17992);
and U18023 (N_18023,N_17961,N_17957);
nand U18024 (N_18024,N_17038,N_17596);
nand U18025 (N_18025,N_17450,N_17274);
and U18026 (N_18026,N_17828,N_17773);
xor U18027 (N_18027,N_17717,N_17980);
and U18028 (N_18028,N_17339,N_17515);
xor U18029 (N_18029,N_17726,N_17213);
xor U18030 (N_18030,N_17712,N_17911);
or U18031 (N_18031,N_17210,N_17565);
and U18032 (N_18032,N_17341,N_17574);
nor U18033 (N_18033,N_17281,N_17628);
nand U18034 (N_18034,N_17558,N_17150);
xnor U18035 (N_18035,N_17462,N_17355);
or U18036 (N_18036,N_17968,N_17039);
nand U18037 (N_18037,N_17060,N_17514);
nor U18038 (N_18038,N_17738,N_17364);
nor U18039 (N_18039,N_17189,N_17556);
xor U18040 (N_18040,N_17386,N_17700);
nor U18041 (N_18041,N_17375,N_17995);
nand U18042 (N_18042,N_17280,N_17588);
nand U18043 (N_18043,N_17496,N_17401);
nand U18044 (N_18044,N_17173,N_17176);
xor U18045 (N_18045,N_17982,N_17591);
nor U18046 (N_18046,N_17627,N_17157);
nand U18047 (N_18047,N_17049,N_17265);
nand U18048 (N_18048,N_17387,N_17249);
xor U18049 (N_18049,N_17886,N_17235);
and U18050 (N_18050,N_17609,N_17632);
or U18051 (N_18051,N_17013,N_17393);
or U18052 (N_18052,N_17942,N_17221);
xor U18053 (N_18053,N_17120,N_17233);
nand U18054 (N_18054,N_17534,N_17822);
nor U18055 (N_18055,N_17690,N_17267);
and U18056 (N_18056,N_17789,N_17010);
nor U18057 (N_18057,N_17569,N_17344);
or U18058 (N_18058,N_17254,N_17939);
and U18059 (N_18059,N_17015,N_17731);
nor U18060 (N_18060,N_17916,N_17996);
xor U18061 (N_18061,N_17290,N_17354);
xor U18062 (N_18062,N_17849,N_17977);
nand U18063 (N_18063,N_17779,N_17643);
nand U18064 (N_18064,N_17226,N_17990);
nor U18065 (N_18065,N_17635,N_17498);
xnor U18066 (N_18066,N_17915,N_17276);
and U18067 (N_18067,N_17914,N_17570);
and U18068 (N_18068,N_17115,N_17062);
xor U18069 (N_18069,N_17042,N_17746);
or U18070 (N_18070,N_17193,N_17516);
nor U18071 (N_18071,N_17252,N_17701);
nor U18072 (N_18072,N_17061,N_17946);
xor U18073 (N_18073,N_17492,N_17521);
nor U18074 (N_18074,N_17381,N_17453);
nor U18075 (N_18075,N_17620,N_17715);
or U18076 (N_18076,N_17582,N_17662);
nand U18077 (N_18077,N_17294,N_17812);
or U18078 (N_18078,N_17847,N_17885);
and U18079 (N_18079,N_17474,N_17117);
nand U18080 (N_18080,N_17763,N_17478);
xnor U18081 (N_18081,N_17456,N_17325);
nor U18082 (N_18082,N_17180,N_17411);
nand U18083 (N_18083,N_17610,N_17500);
and U18084 (N_18084,N_17818,N_17649);
xor U18085 (N_18085,N_17630,N_17084);
nor U18086 (N_18086,N_17146,N_17211);
xnor U18087 (N_18087,N_17958,N_17768);
xnor U18088 (N_18088,N_17182,N_17658);
nor U18089 (N_18089,N_17848,N_17862);
or U18090 (N_18090,N_17664,N_17338);
nand U18091 (N_18091,N_17722,N_17633);
nor U18092 (N_18092,N_17340,N_17937);
xnor U18093 (N_18093,N_17728,N_17602);
and U18094 (N_18094,N_17676,N_17932);
or U18095 (N_18095,N_17349,N_17047);
nand U18096 (N_18096,N_17251,N_17268);
nor U18097 (N_18097,N_17537,N_17951);
xnor U18098 (N_18098,N_17177,N_17971);
and U18099 (N_18099,N_17218,N_17287);
or U18100 (N_18100,N_17997,N_17679);
nand U18101 (N_18101,N_17156,N_17924);
or U18102 (N_18102,N_17321,N_17170);
xor U18103 (N_18103,N_17994,N_17810);
or U18104 (N_18104,N_17873,N_17979);
nor U18105 (N_18105,N_17684,N_17947);
nor U18106 (N_18106,N_17402,N_17391);
and U18107 (N_18107,N_17612,N_17032);
or U18108 (N_18108,N_17694,N_17890);
xnor U18109 (N_18109,N_17833,N_17148);
nor U18110 (N_18110,N_17766,N_17646);
nor U18111 (N_18111,N_17459,N_17445);
nand U18112 (N_18112,N_17052,N_17113);
nand U18113 (N_18113,N_17102,N_17634);
nor U18114 (N_18114,N_17371,N_17020);
or U18115 (N_18115,N_17056,N_17877);
nor U18116 (N_18116,N_17442,N_17236);
xnor U18117 (N_18117,N_17794,N_17353);
nor U18118 (N_18118,N_17449,N_17346);
and U18119 (N_18119,N_17699,N_17665);
nor U18120 (N_18120,N_17366,N_17545);
nand U18121 (N_18121,N_17095,N_17686);
or U18122 (N_18122,N_17929,N_17969);
and U18123 (N_18123,N_17432,N_17716);
xor U18124 (N_18124,N_17670,N_17229);
or U18125 (N_18125,N_17495,N_17583);
or U18126 (N_18126,N_17261,N_17892);
nand U18127 (N_18127,N_17225,N_17908);
and U18128 (N_18128,N_17174,N_17467);
xor U18129 (N_18129,N_17869,N_17222);
or U18130 (N_18130,N_17295,N_17300);
and U18131 (N_18131,N_17764,N_17175);
nor U18132 (N_18132,N_17255,N_17641);
or U18133 (N_18133,N_17902,N_17741);
xnor U18134 (N_18134,N_17923,N_17934);
nor U18135 (N_18135,N_17035,N_17104);
nor U18136 (N_18136,N_17579,N_17553);
and U18137 (N_18137,N_17105,N_17837);
nand U18138 (N_18138,N_17648,N_17473);
nor U18139 (N_18139,N_17520,N_17082);
and U18140 (N_18140,N_17145,N_17262);
and U18141 (N_18141,N_17457,N_17607);
or U18142 (N_18142,N_17487,N_17959);
and U18143 (N_18143,N_17337,N_17484);
nand U18144 (N_18144,N_17392,N_17040);
and U18145 (N_18145,N_17412,N_17116);
or U18146 (N_18146,N_17654,N_17667);
nor U18147 (N_18147,N_17577,N_17382);
xor U18148 (N_18148,N_17573,N_17031);
and U18149 (N_18149,N_17400,N_17505);
nand U18150 (N_18150,N_17303,N_17024);
xnor U18151 (N_18151,N_17824,N_17048);
nor U18152 (N_18152,N_17385,N_17147);
xor U18153 (N_18153,N_17164,N_17504);
xor U18154 (N_18154,N_17533,N_17782);
nor U18155 (N_18155,N_17350,N_17983);
nand U18156 (N_18156,N_17736,N_17608);
and U18157 (N_18157,N_17752,N_17754);
and U18158 (N_18158,N_17016,N_17852);
nor U18159 (N_18159,N_17542,N_17378);
nand U18160 (N_18160,N_17875,N_17253);
and U18161 (N_18161,N_17129,N_17054);
and U18162 (N_18162,N_17239,N_17441);
or U18163 (N_18163,N_17687,N_17380);
or U18164 (N_18164,N_17486,N_17282);
xnor U18165 (N_18165,N_17688,N_17819);
xor U18166 (N_18166,N_17889,N_17224);
and U18167 (N_18167,N_17403,N_17037);
xnor U18168 (N_18168,N_17377,N_17933);
nand U18169 (N_18169,N_17352,N_17851);
nor U18170 (N_18170,N_17685,N_17530);
or U18171 (N_18171,N_17394,N_17012);
nor U18172 (N_18172,N_17523,N_17518);
and U18173 (N_18173,N_17151,N_17975);
nand U18174 (N_18174,N_17872,N_17335);
nand U18175 (N_18175,N_17970,N_17571);
nor U18176 (N_18176,N_17167,N_17479);
or U18177 (N_18177,N_17238,N_17072);
and U18178 (N_18178,N_17597,N_17705);
or U18179 (N_18179,N_17692,N_17109);
or U18180 (N_18180,N_17493,N_17540);
or U18181 (N_18181,N_17126,N_17470);
xor U18182 (N_18182,N_17960,N_17414);
or U18183 (N_18183,N_17477,N_17522);
nand U18184 (N_18184,N_17784,N_17348);
or U18185 (N_18185,N_17605,N_17407);
and U18186 (N_18186,N_17075,N_17083);
nand U18187 (N_18187,N_17695,N_17333);
xor U18188 (N_18188,N_17244,N_17372);
nor U18189 (N_18189,N_17159,N_17033);
nand U18190 (N_18190,N_17972,N_17390);
nor U18191 (N_18191,N_17880,N_17606);
and U18192 (N_18192,N_17743,N_17861);
and U18193 (N_18193,N_17625,N_17733);
nand U18194 (N_18194,N_17645,N_17409);
xor U18195 (N_18195,N_17132,N_17927);
nand U18196 (N_18196,N_17698,N_17724);
and U18197 (N_18197,N_17737,N_17904);
nor U18198 (N_18198,N_17134,N_17876);
xor U18199 (N_18199,N_17554,N_17976);
nor U18200 (N_18200,N_17271,N_17144);
nand U18201 (N_18201,N_17895,N_17771);
nor U18202 (N_18202,N_17878,N_17543);
or U18203 (N_18203,N_17466,N_17136);
xor U18204 (N_18204,N_17948,N_17623);
and U18205 (N_18205,N_17720,N_17240);
and U18206 (N_18206,N_17342,N_17998);
nor U18207 (N_18207,N_17027,N_17601);
xor U18208 (N_18208,N_17191,N_17863);
and U18209 (N_18209,N_17272,N_17074);
nor U18210 (N_18210,N_17008,N_17906);
and U18211 (N_18211,N_17059,N_17689);
or U18212 (N_18212,N_17650,N_17455);
or U18213 (N_18213,N_17963,N_17389);
xnor U18214 (N_18214,N_17044,N_17317);
nor U18215 (N_18215,N_17204,N_17891);
nand U18216 (N_18216,N_17775,N_17110);
nor U18217 (N_18217,N_17107,N_17702);
and U18218 (N_18218,N_17791,N_17119);
and U18219 (N_18219,N_17666,N_17919);
or U18220 (N_18220,N_17660,N_17435);
and U18221 (N_18221,N_17071,N_17944);
nor U18222 (N_18222,N_17021,N_17858);
and U18223 (N_18223,N_17838,N_17723);
xnor U18224 (N_18224,N_17057,N_17727);
nor U18225 (N_18225,N_17396,N_17683);
or U18226 (N_18226,N_17100,N_17376);
or U18227 (N_18227,N_17912,N_17900);
xor U18228 (N_18228,N_17626,N_17131);
xor U18229 (N_18229,N_17550,N_17857);
or U18230 (N_18230,N_17536,N_17677);
xnor U18231 (N_18231,N_17673,N_17328);
nand U18232 (N_18232,N_17011,N_17094);
or U18233 (N_18233,N_17792,N_17940);
and U18234 (N_18234,N_17510,N_17546);
and U18235 (N_18235,N_17142,N_17326);
or U18236 (N_18236,N_17758,N_17899);
xor U18237 (N_18237,N_17809,N_17721);
xnor U18238 (N_18238,N_17043,N_17549);
nor U18239 (N_18239,N_17888,N_17133);
nor U18240 (N_18240,N_17894,N_17616);
or U18241 (N_18241,N_17121,N_17513);
xor U18242 (N_18242,N_17245,N_17202);
and U18243 (N_18243,N_17587,N_17089);
or U18244 (N_18244,N_17777,N_17710);
nor U18245 (N_18245,N_17840,N_17436);
nor U18246 (N_18246,N_17030,N_17647);
xor U18247 (N_18247,N_17519,N_17216);
xor U18248 (N_18248,N_17561,N_17171);
nand U18249 (N_18249,N_17122,N_17706);
and U18250 (N_18250,N_17362,N_17163);
nor U18251 (N_18251,N_17839,N_17471);
nor U18252 (N_18252,N_17258,N_17767);
nor U18253 (N_18253,N_17999,N_17604);
and U18254 (N_18254,N_17301,N_17770);
or U18255 (N_18255,N_17331,N_17805);
nor U18256 (N_18256,N_17621,N_17966);
nand U18257 (N_18257,N_17329,N_17172);
nand U18258 (N_18258,N_17434,N_17774);
nand U18259 (N_18259,N_17855,N_17859);
xnor U18260 (N_18260,N_17611,N_17475);
xnor U18261 (N_18261,N_17160,N_17334);
nand U18262 (N_18262,N_17953,N_17697);
xor U18263 (N_18263,N_17709,N_17526);
or U18264 (N_18264,N_17811,N_17090);
xor U18265 (N_18265,N_17696,N_17600);
and U18266 (N_18266,N_17181,N_17114);
nor U18267 (N_18267,N_17324,N_17237);
and U18268 (N_18268,N_17884,N_17155);
nand U18269 (N_18269,N_17599,N_17283);
nand U18270 (N_18270,N_17555,N_17964);
nand U18271 (N_18271,N_17096,N_17575);
nand U18272 (N_18272,N_17420,N_17832);
nor U18273 (N_18273,N_17419,N_17581);
or U18274 (N_18274,N_17425,N_17950);
nor U18275 (N_18275,N_17985,N_17395);
xor U18276 (N_18276,N_17524,N_17101);
nor U18277 (N_18277,N_17788,N_17800);
nor U18278 (N_18278,N_17817,N_17759);
nand U18279 (N_18279,N_17140,N_17750);
xnor U18280 (N_18280,N_17987,N_17935);
nor U18281 (N_18281,N_17661,N_17231);
nor U18282 (N_18282,N_17437,N_17489);
or U18283 (N_18283,N_17444,N_17488);
and U18284 (N_18284,N_17356,N_17671);
and U18285 (N_18285,N_17644,N_17201);
xnor U18286 (N_18286,N_17921,N_17846);
xnor U18287 (N_18287,N_17808,N_17619);
and U18288 (N_18288,N_17988,N_17397);
or U18289 (N_18289,N_17305,N_17564);
or U18290 (N_18290,N_17154,N_17512);
xor U18291 (N_18291,N_17803,N_17106);
or U18292 (N_18292,N_17413,N_17866);
xnor U18293 (N_18293,N_17622,N_17454);
nor U18294 (N_18294,N_17659,N_17139);
or U18295 (N_18295,N_17336,N_17879);
and U18296 (N_18296,N_17208,N_17464);
xnor U18297 (N_18297,N_17351,N_17118);
or U18298 (N_18298,N_17802,N_17404);
and U18299 (N_18299,N_17497,N_17299);
nor U18300 (N_18300,N_17028,N_17168);
or U18301 (N_18301,N_17242,N_17507);
xnor U18302 (N_18302,N_17651,N_17593);
and U18303 (N_18303,N_17408,N_17922);
xor U18304 (N_18304,N_17166,N_17112);
nand U18305 (N_18305,N_17557,N_17003);
or U18306 (N_18306,N_17785,N_17568);
and U18307 (N_18307,N_17141,N_17769);
or U18308 (N_18308,N_17297,N_17410);
nand U18309 (N_18309,N_17672,N_17631);
and U18310 (N_18310,N_17091,N_17069);
nand U18311 (N_18311,N_17135,N_17078);
xnor U18312 (N_18312,N_17874,N_17482);
nor U18313 (N_18313,N_17509,N_17077);
nor U18314 (N_18314,N_17322,N_17552);
and U18315 (N_18315,N_17358,N_17468);
or U18316 (N_18316,N_17765,N_17956);
or U18317 (N_18317,N_17315,N_17374);
nor U18318 (N_18318,N_17535,N_17451);
and U18319 (N_18319,N_17506,N_17430);
nand U18320 (N_18320,N_17029,N_17674);
and U18321 (N_18321,N_17006,N_17795);
nand U18322 (N_18322,N_17901,N_17359);
nand U18323 (N_18323,N_17241,N_17820);
xor U18324 (N_18324,N_17757,N_17002);
nor U18325 (N_18325,N_17458,N_17097);
or U18326 (N_18326,N_17865,N_17429);
xor U18327 (N_18327,N_17707,N_17823);
xnor U18328 (N_18328,N_17580,N_17761);
and U18329 (N_18329,N_17563,N_17169);
xnor U18330 (N_18330,N_17292,N_17469);
xor U18331 (N_18331,N_17682,N_17936);
nor U18332 (N_18332,N_17826,N_17289);
and U18333 (N_18333,N_17311,N_17978);
nand U18334 (N_18334,N_17544,N_17250);
nand U18335 (N_18335,N_17192,N_17248);
or U18336 (N_18336,N_17228,N_17323);
xnor U18337 (N_18337,N_17439,N_17896);
nor U18338 (N_18338,N_17909,N_17827);
nand U18339 (N_18339,N_17065,N_17918);
nand U18340 (N_18340,N_17137,N_17952);
nor U18341 (N_18341,N_17871,N_17318);
and U18342 (N_18342,N_17360,N_17187);
and U18343 (N_18343,N_17125,N_17864);
nand U18344 (N_18344,N_17053,N_17127);
and U18345 (N_18345,N_17188,N_17491);
or U18346 (N_18346,N_17307,N_17655);
xnor U18347 (N_18347,N_17798,N_17320);
nand U18348 (N_18348,N_17357,N_17185);
nor U18349 (N_18349,N_17275,N_17001);
xnor U18350 (N_18350,N_17025,N_17103);
nand U18351 (N_18351,N_17306,N_17165);
nand U18352 (N_18352,N_17989,N_17675);
and U18353 (N_18353,N_17910,N_17829);
nor U18354 (N_18354,N_17428,N_17232);
nand U18355 (N_18355,N_17678,N_17636);
nand U18356 (N_18356,N_17017,N_17215);
or U18357 (N_18357,N_17585,N_17373);
or U18358 (N_18358,N_17220,N_17034);
or U18359 (N_18359,N_17617,N_17898);
xor U18360 (N_18360,N_17286,N_17304);
nand U18361 (N_18361,N_17527,N_17799);
xnor U18362 (N_18362,N_17614,N_17931);
and U18363 (N_18363,N_17551,N_17205);
nor U18364 (N_18364,N_17092,N_17541);
nor U18365 (N_18365,N_17050,N_17529);
nor U18366 (N_18366,N_17807,N_17856);
nor U18367 (N_18367,N_17780,N_17263);
xor U18368 (N_18368,N_17893,N_17938);
and U18369 (N_18369,N_17361,N_17567);
nand U18370 (N_18370,N_17797,N_17485);
and U18371 (N_18371,N_17423,N_17009);
or U18372 (N_18372,N_17343,N_17532);
nor U18373 (N_18373,N_17196,N_17854);
nand U18374 (N_18374,N_17981,N_17273);
nand U18375 (N_18375,N_17076,N_17022);
xor U18376 (N_18376,N_17446,N_17162);
nor U18377 (N_18377,N_17088,N_17517);
or U18378 (N_18378,N_17230,N_17045);
or U18379 (N_18379,N_17153,N_17085);
or U18380 (N_18380,N_17055,N_17149);
or U18381 (N_18381,N_17748,N_17111);
xor U18382 (N_18382,N_17881,N_17772);
xnor U18383 (N_18383,N_17227,N_17161);
nor U18384 (N_18384,N_17190,N_17954);
nor U18385 (N_18385,N_17036,N_17786);
or U18386 (N_18386,N_17461,N_17842);
nand U18387 (N_18387,N_17714,N_17447);
xnor U18388 (N_18388,N_17443,N_17576);
and U18389 (N_18389,N_17490,N_17018);
or U18390 (N_18390,N_17023,N_17920);
nand U18391 (N_18391,N_17680,N_17955);
xor U18392 (N_18392,N_17613,N_17749);
and U18393 (N_18393,N_17051,N_17595);
xnor U18394 (N_18394,N_17691,N_17815);
nand U18395 (N_18395,N_17291,N_17525);
and U18396 (N_18396,N_17730,N_17783);
and U18397 (N_18397,N_17246,N_17440);
xor U18398 (N_18398,N_17431,N_17897);
and U18399 (N_18399,N_17004,N_17278);
and U18400 (N_18400,N_17309,N_17448);
nor U18401 (N_18401,N_17124,N_17365);
xnor U18402 (N_18402,N_17415,N_17590);
xnor U18403 (N_18403,N_17000,N_17269);
or U18404 (N_18404,N_17367,N_17158);
or U18405 (N_18405,N_17776,N_17624);
or U18406 (N_18406,N_17531,N_17312);
or U18407 (N_18407,N_17821,N_17511);
nor U18408 (N_18408,N_17508,N_17868);
or U18409 (N_18409,N_17825,N_17778);
nor U18410 (N_18410,N_17186,N_17058);
or U18411 (N_18411,N_17926,N_17747);
nor U18412 (N_18412,N_17539,N_17907);
or U18413 (N_18413,N_17538,N_17418);
nor U18414 (N_18414,N_17480,N_17756);
or U18415 (N_18415,N_17481,N_17925);
xor U18416 (N_18416,N_17398,N_17943);
and U18417 (N_18417,N_17203,N_17967);
or U18418 (N_18418,N_17369,N_17383);
xor U18419 (N_18419,N_17787,N_17266);
xnor U18420 (N_18420,N_17903,N_17194);
and U18421 (N_18421,N_17499,N_17417);
and U18422 (N_18422,N_17426,N_17427);
or U18423 (N_18423,N_17302,N_17656);
and U18424 (N_18424,N_17087,N_17589);
and U18425 (N_18425,N_17974,N_17629);
and U18426 (N_18426,N_17347,N_17363);
or U18427 (N_18427,N_17494,N_17870);
xor U18428 (N_18428,N_17640,N_17288);
nand U18429 (N_18429,N_17206,N_17345);
and U18430 (N_18430,N_17693,N_17729);
nand U18431 (N_18431,N_17279,N_17501);
or U18432 (N_18432,N_17836,N_17930);
xnor U18433 (N_18433,N_17212,N_17708);
xor U18434 (N_18434,N_17080,N_17424);
nand U18435 (N_18435,N_17123,N_17296);
nand U18436 (N_18436,N_17079,N_17421);
and U18437 (N_18437,N_17019,N_17713);
or U18438 (N_18438,N_17949,N_17928);
nand U18439 (N_18439,N_17070,N_17270);
xor U18440 (N_18440,N_17548,N_17562);
nand U18441 (N_18441,N_17379,N_17790);
nor U18442 (N_18442,N_17744,N_17572);
and U18443 (N_18443,N_17760,N_17735);
and U18444 (N_18444,N_17256,N_17405);
xnor U18445 (N_18445,N_17547,N_17319);
xnor U18446 (N_18446,N_17867,N_17669);
and U18447 (N_18447,N_17668,N_17098);
nand U18448 (N_18448,N_17941,N_17719);
nand U18449 (N_18449,N_17130,N_17753);
xor U18450 (N_18450,N_17986,N_17064);
and U18451 (N_18451,N_17465,N_17711);
or U18452 (N_18452,N_17108,N_17200);
xnor U18453 (N_18453,N_17416,N_17138);
nor U18454 (N_18454,N_17093,N_17483);
nand U18455 (N_18455,N_17472,N_17143);
and U18456 (N_18456,N_17830,N_17528);
or U18457 (N_18457,N_17041,N_17816);
xor U18458 (N_18458,N_17806,N_17652);
nand U18459 (N_18459,N_17327,N_17739);
or U18460 (N_18460,N_17330,N_17850);
nand U18461 (N_18461,N_17046,N_17560);
xor U18462 (N_18462,N_17007,N_17917);
and U18463 (N_18463,N_17310,N_17197);
nor U18464 (N_18464,N_17463,N_17293);
or U18465 (N_18465,N_17217,N_17452);
nor U18466 (N_18466,N_17026,N_17973);
xnor U18467 (N_18467,N_17099,N_17887);
nand U18468 (N_18468,N_17703,N_17068);
nor U18469 (N_18469,N_17781,N_17984);
nand U18470 (N_18470,N_17991,N_17801);
and U18471 (N_18471,N_17313,N_17314);
or U18472 (N_18472,N_17243,N_17259);
nor U18473 (N_18473,N_17586,N_17725);
or U18474 (N_18474,N_17618,N_17751);
and U18475 (N_18475,N_17178,N_17592);
and U18476 (N_18476,N_17718,N_17841);
and U18477 (N_18477,N_17502,N_17845);
xnor U18478 (N_18478,N_17179,N_17198);
xnor U18479 (N_18479,N_17063,N_17209);
nor U18480 (N_18480,N_17260,N_17199);
and U18481 (N_18481,N_17742,N_17913);
and U18482 (N_18482,N_17073,N_17195);
and U18483 (N_18483,N_17081,N_17460);
xnor U18484 (N_18484,N_17223,N_17384);
xor U18485 (N_18485,N_17793,N_17067);
xnor U18486 (N_18486,N_17853,N_17642);
xnor U18487 (N_18487,N_17503,N_17653);
and U18488 (N_18488,N_17584,N_17834);
or U18489 (N_18489,N_17438,N_17704);
xor U18490 (N_18490,N_17883,N_17264);
or U18491 (N_18491,N_17014,N_17965);
and U18492 (N_18492,N_17257,N_17745);
nor U18493 (N_18493,N_17332,N_17234);
nor U18494 (N_18494,N_17813,N_17663);
or U18495 (N_18495,N_17005,N_17559);
xnor U18496 (N_18496,N_17152,N_17639);
nand U18497 (N_18497,N_17945,N_17277);
nand U18498 (N_18498,N_17638,N_17905);
xnor U18499 (N_18499,N_17962,N_17762);
nand U18500 (N_18500,N_17031,N_17541);
nand U18501 (N_18501,N_17249,N_17046);
and U18502 (N_18502,N_17915,N_17602);
and U18503 (N_18503,N_17666,N_17810);
and U18504 (N_18504,N_17029,N_17960);
nor U18505 (N_18505,N_17024,N_17040);
or U18506 (N_18506,N_17255,N_17006);
or U18507 (N_18507,N_17416,N_17716);
nand U18508 (N_18508,N_17420,N_17607);
or U18509 (N_18509,N_17605,N_17055);
nor U18510 (N_18510,N_17971,N_17531);
or U18511 (N_18511,N_17004,N_17470);
and U18512 (N_18512,N_17753,N_17059);
and U18513 (N_18513,N_17896,N_17727);
nor U18514 (N_18514,N_17036,N_17970);
or U18515 (N_18515,N_17372,N_17935);
nor U18516 (N_18516,N_17951,N_17755);
nand U18517 (N_18517,N_17355,N_17949);
nand U18518 (N_18518,N_17048,N_17542);
or U18519 (N_18519,N_17536,N_17207);
and U18520 (N_18520,N_17143,N_17260);
or U18521 (N_18521,N_17170,N_17382);
or U18522 (N_18522,N_17523,N_17026);
nand U18523 (N_18523,N_17506,N_17865);
or U18524 (N_18524,N_17678,N_17459);
nand U18525 (N_18525,N_17105,N_17352);
xor U18526 (N_18526,N_17062,N_17360);
or U18527 (N_18527,N_17949,N_17457);
or U18528 (N_18528,N_17863,N_17414);
nor U18529 (N_18529,N_17342,N_17346);
and U18530 (N_18530,N_17192,N_17879);
nand U18531 (N_18531,N_17332,N_17027);
xnor U18532 (N_18532,N_17939,N_17634);
xor U18533 (N_18533,N_17241,N_17628);
nand U18534 (N_18534,N_17083,N_17930);
or U18535 (N_18535,N_17948,N_17366);
nand U18536 (N_18536,N_17163,N_17453);
nand U18537 (N_18537,N_17101,N_17004);
and U18538 (N_18538,N_17341,N_17749);
xor U18539 (N_18539,N_17921,N_17989);
nand U18540 (N_18540,N_17850,N_17778);
nand U18541 (N_18541,N_17062,N_17848);
nor U18542 (N_18542,N_17365,N_17441);
xnor U18543 (N_18543,N_17069,N_17867);
nand U18544 (N_18544,N_17540,N_17788);
or U18545 (N_18545,N_17830,N_17185);
nand U18546 (N_18546,N_17809,N_17723);
and U18547 (N_18547,N_17877,N_17197);
nand U18548 (N_18548,N_17849,N_17518);
and U18549 (N_18549,N_17993,N_17980);
and U18550 (N_18550,N_17753,N_17662);
nor U18551 (N_18551,N_17410,N_17454);
and U18552 (N_18552,N_17231,N_17094);
or U18553 (N_18553,N_17838,N_17696);
nand U18554 (N_18554,N_17804,N_17806);
and U18555 (N_18555,N_17938,N_17632);
nand U18556 (N_18556,N_17445,N_17685);
and U18557 (N_18557,N_17856,N_17668);
and U18558 (N_18558,N_17232,N_17999);
and U18559 (N_18559,N_17110,N_17740);
and U18560 (N_18560,N_17924,N_17413);
nor U18561 (N_18561,N_17214,N_17292);
and U18562 (N_18562,N_17549,N_17147);
nor U18563 (N_18563,N_17815,N_17388);
and U18564 (N_18564,N_17922,N_17495);
nor U18565 (N_18565,N_17954,N_17288);
and U18566 (N_18566,N_17273,N_17856);
or U18567 (N_18567,N_17149,N_17410);
xor U18568 (N_18568,N_17719,N_17050);
and U18569 (N_18569,N_17098,N_17465);
xor U18570 (N_18570,N_17456,N_17438);
or U18571 (N_18571,N_17527,N_17645);
and U18572 (N_18572,N_17760,N_17876);
xor U18573 (N_18573,N_17081,N_17526);
or U18574 (N_18574,N_17741,N_17012);
xor U18575 (N_18575,N_17417,N_17581);
or U18576 (N_18576,N_17576,N_17857);
xor U18577 (N_18577,N_17821,N_17783);
or U18578 (N_18578,N_17852,N_17295);
nand U18579 (N_18579,N_17830,N_17315);
nor U18580 (N_18580,N_17521,N_17276);
and U18581 (N_18581,N_17708,N_17559);
nand U18582 (N_18582,N_17070,N_17893);
and U18583 (N_18583,N_17203,N_17745);
xor U18584 (N_18584,N_17883,N_17803);
nand U18585 (N_18585,N_17321,N_17977);
nor U18586 (N_18586,N_17313,N_17158);
nand U18587 (N_18587,N_17478,N_17363);
nor U18588 (N_18588,N_17805,N_17722);
and U18589 (N_18589,N_17402,N_17296);
and U18590 (N_18590,N_17743,N_17153);
or U18591 (N_18591,N_17288,N_17285);
xor U18592 (N_18592,N_17835,N_17108);
or U18593 (N_18593,N_17809,N_17473);
or U18594 (N_18594,N_17084,N_17856);
or U18595 (N_18595,N_17859,N_17160);
nand U18596 (N_18596,N_17512,N_17374);
nand U18597 (N_18597,N_17538,N_17216);
nand U18598 (N_18598,N_17629,N_17950);
nor U18599 (N_18599,N_17164,N_17379);
nand U18600 (N_18600,N_17789,N_17575);
or U18601 (N_18601,N_17592,N_17729);
nand U18602 (N_18602,N_17737,N_17231);
and U18603 (N_18603,N_17679,N_17047);
xor U18604 (N_18604,N_17260,N_17196);
or U18605 (N_18605,N_17185,N_17074);
and U18606 (N_18606,N_17555,N_17250);
and U18607 (N_18607,N_17927,N_17586);
nor U18608 (N_18608,N_17904,N_17919);
xnor U18609 (N_18609,N_17977,N_17170);
nand U18610 (N_18610,N_17597,N_17386);
and U18611 (N_18611,N_17357,N_17607);
xnor U18612 (N_18612,N_17094,N_17781);
and U18613 (N_18613,N_17005,N_17887);
xnor U18614 (N_18614,N_17557,N_17233);
or U18615 (N_18615,N_17711,N_17978);
xor U18616 (N_18616,N_17772,N_17572);
xnor U18617 (N_18617,N_17639,N_17800);
nor U18618 (N_18618,N_17657,N_17563);
or U18619 (N_18619,N_17877,N_17639);
nor U18620 (N_18620,N_17976,N_17233);
xnor U18621 (N_18621,N_17794,N_17594);
nor U18622 (N_18622,N_17944,N_17183);
nor U18623 (N_18623,N_17650,N_17925);
nor U18624 (N_18624,N_17164,N_17532);
and U18625 (N_18625,N_17245,N_17256);
and U18626 (N_18626,N_17776,N_17691);
xnor U18627 (N_18627,N_17396,N_17736);
and U18628 (N_18628,N_17768,N_17759);
and U18629 (N_18629,N_17219,N_17012);
xor U18630 (N_18630,N_17279,N_17637);
nor U18631 (N_18631,N_17225,N_17162);
nor U18632 (N_18632,N_17336,N_17721);
nand U18633 (N_18633,N_17515,N_17384);
and U18634 (N_18634,N_17608,N_17697);
or U18635 (N_18635,N_17242,N_17807);
nor U18636 (N_18636,N_17334,N_17133);
nor U18637 (N_18637,N_17691,N_17421);
and U18638 (N_18638,N_17833,N_17814);
and U18639 (N_18639,N_17894,N_17611);
or U18640 (N_18640,N_17412,N_17394);
or U18641 (N_18641,N_17592,N_17104);
and U18642 (N_18642,N_17989,N_17384);
nor U18643 (N_18643,N_17968,N_17261);
nand U18644 (N_18644,N_17454,N_17055);
and U18645 (N_18645,N_17767,N_17145);
or U18646 (N_18646,N_17208,N_17147);
and U18647 (N_18647,N_17853,N_17495);
nor U18648 (N_18648,N_17573,N_17960);
and U18649 (N_18649,N_17843,N_17775);
and U18650 (N_18650,N_17403,N_17476);
nor U18651 (N_18651,N_17090,N_17097);
xnor U18652 (N_18652,N_17654,N_17348);
or U18653 (N_18653,N_17417,N_17307);
nor U18654 (N_18654,N_17010,N_17537);
nor U18655 (N_18655,N_17665,N_17055);
xor U18656 (N_18656,N_17567,N_17052);
or U18657 (N_18657,N_17856,N_17058);
or U18658 (N_18658,N_17497,N_17133);
nand U18659 (N_18659,N_17382,N_17311);
xor U18660 (N_18660,N_17181,N_17459);
nor U18661 (N_18661,N_17222,N_17511);
xor U18662 (N_18662,N_17242,N_17026);
nand U18663 (N_18663,N_17254,N_17084);
nor U18664 (N_18664,N_17191,N_17271);
and U18665 (N_18665,N_17948,N_17293);
nand U18666 (N_18666,N_17627,N_17120);
and U18667 (N_18667,N_17057,N_17278);
nand U18668 (N_18668,N_17540,N_17299);
or U18669 (N_18669,N_17095,N_17866);
nor U18670 (N_18670,N_17019,N_17189);
or U18671 (N_18671,N_17208,N_17128);
nor U18672 (N_18672,N_17401,N_17421);
xor U18673 (N_18673,N_17205,N_17856);
or U18674 (N_18674,N_17840,N_17459);
nor U18675 (N_18675,N_17028,N_17899);
nor U18676 (N_18676,N_17436,N_17621);
and U18677 (N_18677,N_17945,N_17949);
and U18678 (N_18678,N_17324,N_17721);
or U18679 (N_18679,N_17116,N_17108);
xor U18680 (N_18680,N_17951,N_17753);
and U18681 (N_18681,N_17354,N_17507);
and U18682 (N_18682,N_17073,N_17228);
nand U18683 (N_18683,N_17563,N_17157);
nor U18684 (N_18684,N_17455,N_17033);
xor U18685 (N_18685,N_17438,N_17403);
and U18686 (N_18686,N_17240,N_17225);
nor U18687 (N_18687,N_17228,N_17065);
xor U18688 (N_18688,N_17880,N_17167);
and U18689 (N_18689,N_17350,N_17850);
nor U18690 (N_18690,N_17311,N_17306);
nand U18691 (N_18691,N_17355,N_17936);
or U18692 (N_18692,N_17445,N_17109);
nand U18693 (N_18693,N_17435,N_17230);
nor U18694 (N_18694,N_17395,N_17341);
nor U18695 (N_18695,N_17021,N_17723);
or U18696 (N_18696,N_17861,N_17735);
nand U18697 (N_18697,N_17546,N_17864);
and U18698 (N_18698,N_17477,N_17419);
nor U18699 (N_18699,N_17926,N_17070);
and U18700 (N_18700,N_17943,N_17376);
nor U18701 (N_18701,N_17426,N_17819);
and U18702 (N_18702,N_17046,N_17346);
nand U18703 (N_18703,N_17914,N_17670);
xor U18704 (N_18704,N_17315,N_17154);
and U18705 (N_18705,N_17205,N_17352);
and U18706 (N_18706,N_17122,N_17357);
or U18707 (N_18707,N_17755,N_17245);
nor U18708 (N_18708,N_17807,N_17028);
xnor U18709 (N_18709,N_17983,N_17945);
xnor U18710 (N_18710,N_17252,N_17383);
xnor U18711 (N_18711,N_17905,N_17092);
xor U18712 (N_18712,N_17885,N_17180);
nor U18713 (N_18713,N_17831,N_17523);
nand U18714 (N_18714,N_17290,N_17610);
or U18715 (N_18715,N_17002,N_17186);
xor U18716 (N_18716,N_17321,N_17481);
or U18717 (N_18717,N_17896,N_17282);
and U18718 (N_18718,N_17618,N_17607);
xor U18719 (N_18719,N_17551,N_17925);
xnor U18720 (N_18720,N_17145,N_17221);
nand U18721 (N_18721,N_17314,N_17366);
nor U18722 (N_18722,N_17102,N_17995);
or U18723 (N_18723,N_17563,N_17405);
or U18724 (N_18724,N_17799,N_17261);
xnor U18725 (N_18725,N_17569,N_17610);
xnor U18726 (N_18726,N_17590,N_17666);
xor U18727 (N_18727,N_17456,N_17853);
or U18728 (N_18728,N_17303,N_17651);
xnor U18729 (N_18729,N_17335,N_17229);
xnor U18730 (N_18730,N_17484,N_17376);
nand U18731 (N_18731,N_17233,N_17076);
nor U18732 (N_18732,N_17008,N_17010);
or U18733 (N_18733,N_17160,N_17028);
nand U18734 (N_18734,N_17519,N_17668);
and U18735 (N_18735,N_17134,N_17635);
and U18736 (N_18736,N_17936,N_17216);
or U18737 (N_18737,N_17584,N_17992);
nor U18738 (N_18738,N_17121,N_17986);
nand U18739 (N_18739,N_17521,N_17264);
nand U18740 (N_18740,N_17016,N_17499);
xor U18741 (N_18741,N_17505,N_17064);
nor U18742 (N_18742,N_17497,N_17910);
nand U18743 (N_18743,N_17090,N_17013);
xor U18744 (N_18744,N_17093,N_17123);
or U18745 (N_18745,N_17464,N_17490);
and U18746 (N_18746,N_17709,N_17550);
xnor U18747 (N_18747,N_17609,N_17593);
nand U18748 (N_18748,N_17138,N_17903);
nand U18749 (N_18749,N_17816,N_17930);
nand U18750 (N_18750,N_17828,N_17222);
nor U18751 (N_18751,N_17475,N_17109);
or U18752 (N_18752,N_17642,N_17036);
and U18753 (N_18753,N_17269,N_17945);
or U18754 (N_18754,N_17604,N_17457);
and U18755 (N_18755,N_17275,N_17698);
nand U18756 (N_18756,N_17364,N_17300);
or U18757 (N_18757,N_17803,N_17947);
xnor U18758 (N_18758,N_17748,N_17774);
nand U18759 (N_18759,N_17671,N_17723);
xnor U18760 (N_18760,N_17082,N_17672);
nor U18761 (N_18761,N_17537,N_17267);
xor U18762 (N_18762,N_17409,N_17186);
and U18763 (N_18763,N_17820,N_17907);
xnor U18764 (N_18764,N_17204,N_17449);
nand U18765 (N_18765,N_17537,N_17719);
nand U18766 (N_18766,N_17179,N_17917);
and U18767 (N_18767,N_17269,N_17417);
xnor U18768 (N_18768,N_17114,N_17205);
or U18769 (N_18769,N_17681,N_17438);
and U18770 (N_18770,N_17331,N_17258);
or U18771 (N_18771,N_17008,N_17872);
and U18772 (N_18772,N_17824,N_17280);
xor U18773 (N_18773,N_17219,N_17826);
or U18774 (N_18774,N_17367,N_17535);
nand U18775 (N_18775,N_17220,N_17854);
and U18776 (N_18776,N_17620,N_17571);
xor U18777 (N_18777,N_17339,N_17722);
or U18778 (N_18778,N_17522,N_17303);
nor U18779 (N_18779,N_17344,N_17261);
xor U18780 (N_18780,N_17169,N_17896);
and U18781 (N_18781,N_17252,N_17852);
nor U18782 (N_18782,N_17722,N_17999);
nor U18783 (N_18783,N_17834,N_17836);
or U18784 (N_18784,N_17594,N_17065);
xnor U18785 (N_18785,N_17989,N_17467);
and U18786 (N_18786,N_17734,N_17321);
or U18787 (N_18787,N_17788,N_17655);
nor U18788 (N_18788,N_17047,N_17528);
nand U18789 (N_18789,N_17397,N_17930);
or U18790 (N_18790,N_17289,N_17117);
nor U18791 (N_18791,N_17243,N_17785);
nor U18792 (N_18792,N_17856,N_17735);
and U18793 (N_18793,N_17072,N_17215);
nand U18794 (N_18794,N_17717,N_17197);
xor U18795 (N_18795,N_17496,N_17475);
or U18796 (N_18796,N_17831,N_17391);
xor U18797 (N_18797,N_17102,N_17393);
nor U18798 (N_18798,N_17882,N_17074);
and U18799 (N_18799,N_17743,N_17457);
and U18800 (N_18800,N_17063,N_17374);
xor U18801 (N_18801,N_17443,N_17437);
and U18802 (N_18802,N_17480,N_17079);
nand U18803 (N_18803,N_17838,N_17033);
nor U18804 (N_18804,N_17725,N_17031);
xor U18805 (N_18805,N_17743,N_17310);
and U18806 (N_18806,N_17896,N_17987);
xor U18807 (N_18807,N_17621,N_17431);
nor U18808 (N_18808,N_17910,N_17127);
or U18809 (N_18809,N_17096,N_17103);
and U18810 (N_18810,N_17382,N_17221);
xor U18811 (N_18811,N_17256,N_17014);
nor U18812 (N_18812,N_17136,N_17109);
or U18813 (N_18813,N_17339,N_17543);
and U18814 (N_18814,N_17691,N_17052);
nand U18815 (N_18815,N_17989,N_17943);
nand U18816 (N_18816,N_17998,N_17693);
and U18817 (N_18817,N_17437,N_17468);
xnor U18818 (N_18818,N_17213,N_17580);
nor U18819 (N_18819,N_17263,N_17397);
and U18820 (N_18820,N_17911,N_17778);
nand U18821 (N_18821,N_17741,N_17027);
xnor U18822 (N_18822,N_17781,N_17449);
xnor U18823 (N_18823,N_17294,N_17968);
or U18824 (N_18824,N_17550,N_17524);
xnor U18825 (N_18825,N_17832,N_17547);
and U18826 (N_18826,N_17604,N_17998);
or U18827 (N_18827,N_17967,N_17694);
xor U18828 (N_18828,N_17471,N_17005);
or U18829 (N_18829,N_17510,N_17499);
xor U18830 (N_18830,N_17288,N_17208);
and U18831 (N_18831,N_17890,N_17452);
xnor U18832 (N_18832,N_17182,N_17056);
and U18833 (N_18833,N_17307,N_17735);
and U18834 (N_18834,N_17937,N_17288);
xor U18835 (N_18835,N_17545,N_17070);
or U18836 (N_18836,N_17426,N_17381);
nand U18837 (N_18837,N_17396,N_17343);
and U18838 (N_18838,N_17064,N_17494);
xor U18839 (N_18839,N_17014,N_17312);
xnor U18840 (N_18840,N_17803,N_17921);
xor U18841 (N_18841,N_17824,N_17503);
nand U18842 (N_18842,N_17139,N_17649);
nor U18843 (N_18843,N_17841,N_17292);
or U18844 (N_18844,N_17731,N_17394);
and U18845 (N_18845,N_17935,N_17871);
xnor U18846 (N_18846,N_17884,N_17621);
xor U18847 (N_18847,N_17936,N_17087);
and U18848 (N_18848,N_17146,N_17291);
and U18849 (N_18849,N_17901,N_17994);
nor U18850 (N_18850,N_17045,N_17760);
xnor U18851 (N_18851,N_17596,N_17811);
nor U18852 (N_18852,N_17315,N_17077);
nand U18853 (N_18853,N_17364,N_17956);
xnor U18854 (N_18854,N_17942,N_17289);
nor U18855 (N_18855,N_17722,N_17835);
nand U18856 (N_18856,N_17514,N_17530);
nor U18857 (N_18857,N_17996,N_17233);
nor U18858 (N_18858,N_17391,N_17255);
nand U18859 (N_18859,N_17976,N_17306);
xnor U18860 (N_18860,N_17451,N_17635);
nor U18861 (N_18861,N_17366,N_17535);
nor U18862 (N_18862,N_17206,N_17718);
or U18863 (N_18863,N_17641,N_17460);
and U18864 (N_18864,N_17876,N_17747);
and U18865 (N_18865,N_17659,N_17392);
xor U18866 (N_18866,N_17105,N_17713);
nand U18867 (N_18867,N_17777,N_17493);
nand U18868 (N_18868,N_17009,N_17581);
xnor U18869 (N_18869,N_17846,N_17750);
nand U18870 (N_18870,N_17427,N_17555);
nand U18871 (N_18871,N_17408,N_17574);
nand U18872 (N_18872,N_17016,N_17038);
nor U18873 (N_18873,N_17977,N_17810);
nor U18874 (N_18874,N_17501,N_17586);
xnor U18875 (N_18875,N_17902,N_17287);
and U18876 (N_18876,N_17858,N_17432);
or U18877 (N_18877,N_17440,N_17612);
xnor U18878 (N_18878,N_17252,N_17787);
nor U18879 (N_18879,N_17262,N_17609);
nand U18880 (N_18880,N_17684,N_17637);
and U18881 (N_18881,N_17985,N_17281);
xor U18882 (N_18882,N_17327,N_17377);
and U18883 (N_18883,N_17066,N_17123);
nor U18884 (N_18884,N_17413,N_17827);
nor U18885 (N_18885,N_17161,N_17577);
nand U18886 (N_18886,N_17173,N_17717);
and U18887 (N_18887,N_17821,N_17276);
and U18888 (N_18888,N_17228,N_17883);
nand U18889 (N_18889,N_17038,N_17828);
nor U18890 (N_18890,N_17789,N_17193);
nand U18891 (N_18891,N_17614,N_17016);
nor U18892 (N_18892,N_17635,N_17670);
and U18893 (N_18893,N_17938,N_17929);
nor U18894 (N_18894,N_17598,N_17541);
xor U18895 (N_18895,N_17538,N_17987);
nor U18896 (N_18896,N_17418,N_17059);
xor U18897 (N_18897,N_17296,N_17991);
nand U18898 (N_18898,N_17648,N_17031);
and U18899 (N_18899,N_17971,N_17656);
nand U18900 (N_18900,N_17901,N_17482);
nor U18901 (N_18901,N_17700,N_17067);
nor U18902 (N_18902,N_17729,N_17361);
nand U18903 (N_18903,N_17955,N_17816);
xor U18904 (N_18904,N_17138,N_17411);
nand U18905 (N_18905,N_17747,N_17872);
xnor U18906 (N_18906,N_17551,N_17629);
nor U18907 (N_18907,N_17373,N_17217);
or U18908 (N_18908,N_17637,N_17673);
or U18909 (N_18909,N_17535,N_17726);
xnor U18910 (N_18910,N_17364,N_17955);
xor U18911 (N_18911,N_17909,N_17239);
xor U18912 (N_18912,N_17836,N_17753);
xor U18913 (N_18913,N_17600,N_17812);
nor U18914 (N_18914,N_17928,N_17435);
xnor U18915 (N_18915,N_17798,N_17129);
or U18916 (N_18916,N_17413,N_17314);
nand U18917 (N_18917,N_17744,N_17512);
nor U18918 (N_18918,N_17303,N_17071);
nor U18919 (N_18919,N_17598,N_17454);
nor U18920 (N_18920,N_17435,N_17995);
or U18921 (N_18921,N_17308,N_17677);
and U18922 (N_18922,N_17478,N_17093);
and U18923 (N_18923,N_17687,N_17819);
nor U18924 (N_18924,N_17783,N_17241);
or U18925 (N_18925,N_17623,N_17467);
and U18926 (N_18926,N_17282,N_17828);
nor U18927 (N_18927,N_17089,N_17103);
or U18928 (N_18928,N_17385,N_17728);
nand U18929 (N_18929,N_17931,N_17997);
nor U18930 (N_18930,N_17678,N_17027);
nor U18931 (N_18931,N_17084,N_17128);
nor U18932 (N_18932,N_17570,N_17502);
nor U18933 (N_18933,N_17341,N_17075);
nor U18934 (N_18934,N_17265,N_17922);
nand U18935 (N_18935,N_17473,N_17967);
and U18936 (N_18936,N_17810,N_17017);
or U18937 (N_18937,N_17723,N_17914);
xnor U18938 (N_18938,N_17902,N_17627);
and U18939 (N_18939,N_17203,N_17803);
or U18940 (N_18940,N_17030,N_17638);
xnor U18941 (N_18941,N_17965,N_17106);
nor U18942 (N_18942,N_17448,N_17605);
nand U18943 (N_18943,N_17317,N_17100);
or U18944 (N_18944,N_17414,N_17814);
nor U18945 (N_18945,N_17336,N_17943);
and U18946 (N_18946,N_17722,N_17616);
or U18947 (N_18947,N_17414,N_17815);
nor U18948 (N_18948,N_17199,N_17442);
nor U18949 (N_18949,N_17314,N_17753);
or U18950 (N_18950,N_17297,N_17449);
nand U18951 (N_18951,N_17630,N_17733);
nor U18952 (N_18952,N_17320,N_17862);
nor U18953 (N_18953,N_17529,N_17203);
nor U18954 (N_18954,N_17991,N_17895);
nor U18955 (N_18955,N_17496,N_17859);
nor U18956 (N_18956,N_17763,N_17006);
or U18957 (N_18957,N_17985,N_17264);
and U18958 (N_18958,N_17111,N_17482);
nor U18959 (N_18959,N_17855,N_17526);
or U18960 (N_18960,N_17733,N_17964);
nand U18961 (N_18961,N_17790,N_17611);
or U18962 (N_18962,N_17979,N_17157);
or U18963 (N_18963,N_17685,N_17894);
nor U18964 (N_18964,N_17108,N_17433);
xnor U18965 (N_18965,N_17206,N_17278);
or U18966 (N_18966,N_17774,N_17481);
xnor U18967 (N_18967,N_17040,N_17321);
nor U18968 (N_18968,N_17667,N_17404);
xor U18969 (N_18969,N_17753,N_17697);
nand U18970 (N_18970,N_17403,N_17694);
and U18971 (N_18971,N_17974,N_17436);
and U18972 (N_18972,N_17366,N_17380);
or U18973 (N_18973,N_17662,N_17902);
nand U18974 (N_18974,N_17779,N_17649);
xor U18975 (N_18975,N_17563,N_17397);
or U18976 (N_18976,N_17329,N_17472);
nor U18977 (N_18977,N_17541,N_17922);
and U18978 (N_18978,N_17702,N_17962);
nand U18979 (N_18979,N_17113,N_17871);
or U18980 (N_18980,N_17196,N_17731);
or U18981 (N_18981,N_17666,N_17893);
and U18982 (N_18982,N_17830,N_17618);
or U18983 (N_18983,N_17986,N_17618);
and U18984 (N_18984,N_17566,N_17595);
nor U18985 (N_18985,N_17317,N_17153);
nor U18986 (N_18986,N_17482,N_17425);
nor U18987 (N_18987,N_17021,N_17866);
or U18988 (N_18988,N_17874,N_17400);
or U18989 (N_18989,N_17401,N_17622);
nand U18990 (N_18990,N_17329,N_17070);
and U18991 (N_18991,N_17861,N_17051);
nand U18992 (N_18992,N_17616,N_17884);
and U18993 (N_18993,N_17057,N_17852);
xnor U18994 (N_18994,N_17739,N_17956);
nor U18995 (N_18995,N_17814,N_17183);
xor U18996 (N_18996,N_17836,N_17224);
nand U18997 (N_18997,N_17594,N_17074);
and U18998 (N_18998,N_17626,N_17762);
and U18999 (N_18999,N_17252,N_17833);
or U19000 (N_19000,N_18009,N_18305);
and U19001 (N_19001,N_18197,N_18394);
nor U19002 (N_19002,N_18904,N_18911);
or U19003 (N_19003,N_18857,N_18443);
nor U19004 (N_19004,N_18730,N_18528);
or U19005 (N_19005,N_18574,N_18117);
xnor U19006 (N_19006,N_18993,N_18057);
nand U19007 (N_19007,N_18508,N_18504);
xor U19008 (N_19008,N_18994,N_18845);
nor U19009 (N_19009,N_18489,N_18400);
nand U19010 (N_19010,N_18273,N_18841);
and U19011 (N_19011,N_18014,N_18580);
and U19012 (N_19012,N_18427,N_18720);
or U19013 (N_19013,N_18541,N_18870);
and U19014 (N_19014,N_18654,N_18352);
and U19015 (N_19015,N_18091,N_18538);
nand U19016 (N_19016,N_18038,N_18656);
xor U19017 (N_19017,N_18045,N_18444);
nor U19018 (N_19018,N_18258,N_18061);
or U19019 (N_19019,N_18991,N_18207);
or U19020 (N_19020,N_18692,N_18025);
xnor U19021 (N_19021,N_18526,N_18493);
xnor U19022 (N_19022,N_18088,N_18058);
nor U19023 (N_19023,N_18124,N_18941);
nor U19024 (N_19024,N_18502,N_18474);
nor U19025 (N_19025,N_18155,N_18228);
nand U19026 (N_19026,N_18587,N_18497);
nor U19027 (N_19027,N_18436,N_18896);
nand U19028 (N_19028,N_18562,N_18787);
and U19029 (N_19029,N_18825,N_18962);
nor U19030 (N_19030,N_18871,N_18487);
nor U19031 (N_19031,N_18147,N_18894);
nor U19032 (N_19032,N_18143,N_18711);
nand U19033 (N_19033,N_18529,N_18432);
xnor U19034 (N_19034,N_18568,N_18681);
nand U19035 (N_19035,N_18165,N_18012);
nand U19036 (N_19036,N_18630,N_18341);
nand U19037 (N_19037,N_18843,N_18007);
nand U19038 (N_19038,N_18086,N_18334);
and U19039 (N_19039,N_18733,N_18388);
nor U19040 (N_19040,N_18861,N_18839);
or U19041 (N_19041,N_18326,N_18652);
and U19042 (N_19042,N_18216,N_18028);
xnor U19043 (N_19043,N_18187,N_18132);
or U19044 (N_19044,N_18914,N_18488);
and U19045 (N_19045,N_18530,N_18224);
and U19046 (N_19046,N_18189,N_18913);
or U19047 (N_19047,N_18675,N_18726);
nor U19048 (N_19048,N_18328,N_18174);
and U19049 (N_19049,N_18697,N_18545);
xor U19050 (N_19050,N_18442,N_18840);
nor U19051 (N_19051,N_18389,N_18679);
nor U19052 (N_19052,N_18982,N_18073);
nor U19053 (N_19053,N_18002,N_18929);
xnor U19054 (N_19054,N_18880,N_18138);
xnor U19055 (N_19055,N_18186,N_18721);
and U19056 (N_19056,N_18875,N_18828);
xor U19057 (N_19057,N_18585,N_18844);
xor U19058 (N_19058,N_18668,N_18931);
and U19059 (N_19059,N_18837,N_18008);
xnor U19060 (N_19060,N_18616,N_18856);
or U19061 (N_19061,N_18010,N_18121);
xor U19062 (N_19062,N_18715,N_18410);
nand U19063 (N_19063,N_18859,N_18280);
xnor U19064 (N_19064,N_18286,N_18027);
or U19065 (N_19065,N_18683,N_18324);
and U19066 (N_19066,N_18098,N_18114);
nand U19067 (N_19067,N_18246,N_18808);
nand U19068 (N_19068,N_18811,N_18851);
nand U19069 (N_19069,N_18229,N_18212);
nand U19070 (N_19070,N_18393,N_18603);
xor U19071 (N_19071,N_18325,N_18357);
and U19072 (N_19072,N_18135,N_18524);
xor U19073 (N_19073,N_18672,N_18621);
xnor U19074 (N_19074,N_18759,N_18312);
xor U19075 (N_19075,N_18635,N_18832);
xnor U19076 (N_19076,N_18315,N_18815);
xor U19077 (N_19077,N_18707,N_18582);
or U19078 (N_19078,N_18985,N_18492);
nor U19079 (N_19079,N_18951,N_18932);
and U19080 (N_19080,N_18773,N_18997);
or U19081 (N_19081,N_18686,N_18744);
nand U19082 (N_19082,N_18862,N_18006);
xnor U19083 (N_19083,N_18860,N_18042);
or U19084 (N_19084,N_18299,N_18657);
xnor U19085 (N_19085,N_18163,N_18314);
or U19086 (N_19086,N_18421,N_18570);
or U19087 (N_19087,N_18351,N_18694);
or U19088 (N_19088,N_18849,N_18483);
xor U19089 (N_19089,N_18999,N_18550);
or U19090 (N_19090,N_18321,N_18477);
nor U19091 (N_19091,N_18531,N_18262);
nand U19092 (N_19092,N_18522,N_18283);
and U19093 (N_19093,N_18847,N_18642);
and U19094 (N_19094,N_18395,N_18544);
nand U19095 (N_19095,N_18131,N_18573);
xor U19096 (N_19096,N_18969,N_18942);
and U19097 (N_19097,N_18031,N_18247);
and U19098 (N_19098,N_18542,N_18727);
or U19099 (N_19099,N_18986,N_18592);
and U19100 (N_19100,N_18591,N_18925);
nand U19101 (N_19101,N_18636,N_18223);
and U19102 (N_19102,N_18895,N_18500);
and U19103 (N_19103,N_18157,N_18863);
xor U19104 (N_19104,N_18846,N_18375);
xnor U19105 (N_19105,N_18786,N_18797);
and U19106 (N_19106,N_18893,N_18300);
or U19107 (N_19107,N_18429,N_18596);
nand U19108 (N_19108,N_18584,N_18149);
nor U19109 (N_19109,N_18739,N_18118);
and U19110 (N_19110,N_18891,N_18037);
and U19111 (N_19111,N_18505,N_18298);
xor U19112 (N_19112,N_18885,N_18762);
xnor U19113 (N_19113,N_18938,N_18619);
nor U19114 (N_19114,N_18434,N_18793);
or U19115 (N_19115,N_18276,N_18818);
xnor U19116 (N_19116,N_18688,N_18192);
xnor U19117 (N_19117,N_18651,N_18018);
and U19118 (N_19118,N_18778,N_18052);
nand U19119 (N_19119,N_18598,N_18318);
nor U19120 (N_19120,N_18139,N_18816);
or U19121 (N_19121,N_18869,N_18235);
and U19122 (N_19122,N_18983,N_18764);
nor U19123 (N_19123,N_18170,N_18961);
and U19124 (N_19124,N_18742,N_18771);
nand U19125 (N_19125,N_18198,N_18693);
and U19126 (N_19126,N_18466,N_18700);
nor U19127 (N_19127,N_18438,N_18958);
nand U19128 (N_19128,N_18096,N_18467);
and U19129 (N_19129,N_18250,N_18704);
nand U19130 (N_19130,N_18070,N_18168);
and U19131 (N_19131,N_18960,N_18490);
and U19132 (N_19132,N_18349,N_18971);
xnor U19133 (N_19133,N_18777,N_18785);
or U19134 (N_19134,N_18220,N_18144);
and U19135 (N_19135,N_18689,N_18026);
nand U19136 (N_19136,N_18113,N_18459);
xor U19137 (N_19137,N_18678,N_18639);
nor U19138 (N_19138,N_18676,N_18158);
and U19139 (N_19139,N_18680,N_18552);
nor U19140 (N_19140,N_18032,N_18838);
nor U19141 (N_19141,N_18485,N_18213);
nand U19142 (N_19142,N_18368,N_18384);
nor U19143 (N_19143,N_18747,N_18106);
xor U19144 (N_19144,N_18080,N_18369);
and U19145 (N_19145,N_18980,N_18017);
or U19146 (N_19146,N_18476,N_18669);
and U19147 (N_19147,N_18077,N_18399);
nor U19148 (N_19148,N_18004,N_18362);
and U19149 (N_19149,N_18067,N_18184);
xor U19150 (N_19150,N_18370,N_18236);
xor U19151 (N_19151,N_18270,N_18978);
nor U19152 (N_19152,N_18852,N_18374);
nor U19153 (N_19153,N_18154,N_18548);
nand U19154 (N_19154,N_18699,N_18059);
xor U19155 (N_19155,N_18036,N_18906);
and U19156 (N_19156,N_18511,N_18064);
or U19157 (N_19157,N_18202,N_18243);
and U19158 (N_19158,N_18191,N_18926);
xor U19159 (N_19159,N_18850,N_18858);
nand U19160 (N_19160,N_18551,N_18332);
and U19161 (N_19161,N_18687,N_18446);
or U19162 (N_19162,N_18946,N_18418);
nor U19163 (N_19163,N_18322,N_18167);
xor U19164 (N_19164,N_18617,N_18901);
nor U19165 (N_19165,N_18970,N_18746);
xnor U19166 (N_19166,N_18741,N_18354);
or U19167 (N_19167,N_18610,N_18520);
and U19168 (N_19168,N_18897,N_18166);
or U19169 (N_19169,N_18296,N_18110);
nor U19170 (N_19170,N_18525,N_18761);
and U19171 (N_19171,N_18792,N_18956);
nor U19172 (N_19172,N_18209,N_18082);
or U19173 (N_19173,N_18356,N_18160);
nor U19174 (N_19174,N_18478,N_18363);
and U19175 (N_19175,N_18930,N_18431);
xor U19176 (N_19176,N_18396,N_18968);
and U19177 (N_19177,N_18966,N_18087);
or U19178 (N_19178,N_18921,N_18285);
xor U19179 (N_19179,N_18378,N_18104);
xor U19180 (N_19180,N_18424,N_18953);
xor U19181 (N_19181,N_18109,N_18809);
and U19182 (N_19182,N_18648,N_18724);
nor U19183 (N_19183,N_18084,N_18078);
nor U19184 (N_19184,N_18575,N_18013);
and U19185 (N_19185,N_18164,N_18075);
or U19186 (N_19186,N_18597,N_18658);
xnor U19187 (N_19187,N_18241,N_18887);
or U19188 (N_19188,N_18812,N_18376);
and U19189 (N_19189,N_18288,N_18682);
nor U19190 (N_19190,N_18646,N_18173);
or U19191 (N_19191,N_18965,N_18107);
xor U19192 (N_19192,N_18563,N_18874);
xnor U19193 (N_19193,N_18532,N_18267);
nor U19194 (N_19194,N_18799,N_18567);
or U19195 (N_19195,N_18348,N_18453);
nor U19196 (N_19196,N_18264,N_18898);
nor U19197 (N_19197,N_18623,N_18074);
or U19198 (N_19198,N_18397,N_18450);
and U19199 (N_19199,N_18364,N_18632);
and U19200 (N_19200,N_18503,N_18625);
or U19201 (N_19201,N_18171,N_18448);
and U19202 (N_19202,N_18051,N_18779);
or U19203 (N_19203,N_18804,N_18757);
and U19204 (N_19204,N_18222,N_18948);
xor U19205 (N_19205,N_18736,N_18304);
nand U19206 (N_19206,N_18095,N_18302);
xnor U19207 (N_19207,N_18054,N_18172);
nand U19208 (N_19208,N_18536,N_18398);
or U19209 (N_19209,N_18272,N_18415);
or U19210 (N_19210,N_18631,N_18461);
nor U19211 (N_19211,N_18872,N_18089);
and U19212 (N_19212,N_18440,N_18310);
xor U19213 (N_19213,N_18830,N_18937);
or U19214 (N_19214,N_18001,N_18784);
or U19215 (N_19215,N_18756,N_18760);
xor U19216 (N_19216,N_18578,N_18411);
nor U19217 (N_19217,N_18482,N_18122);
xnor U19218 (N_19218,N_18782,N_18385);
and U19219 (N_19219,N_18182,N_18260);
nand U19220 (N_19220,N_18136,N_18607);
xnor U19221 (N_19221,N_18293,N_18557);
nor U19222 (N_19222,N_18691,N_18053);
nand U19223 (N_19223,N_18734,N_18180);
or U19224 (N_19224,N_18126,N_18454);
and U19225 (N_19225,N_18769,N_18056);
xor U19226 (N_19226,N_18589,N_18824);
nand U19227 (N_19227,N_18281,N_18663);
xor U19228 (N_19228,N_18350,N_18881);
or U19229 (N_19229,N_18346,N_18046);
xor U19230 (N_19230,N_18430,N_18748);
nand U19231 (N_19231,N_18392,N_18817);
or U19232 (N_19232,N_18470,N_18237);
nand U19233 (N_19233,N_18671,N_18102);
or U19234 (N_19234,N_18065,N_18827);
nor U19235 (N_19235,N_18199,N_18156);
or U19236 (N_19236,N_18445,N_18565);
nor U19237 (N_19237,N_18789,N_18920);
or U19238 (N_19238,N_18535,N_18826);
and U19239 (N_19239,N_18219,N_18422);
or U19240 (N_19240,N_18781,N_18030);
or U19241 (N_19241,N_18405,N_18447);
xor U19242 (N_19242,N_18716,N_18390);
xnor U19243 (N_19243,N_18566,N_18383);
nor U19244 (N_19244,N_18115,N_18755);
and U19245 (N_19245,N_18643,N_18848);
or U19246 (N_19246,N_18605,N_18303);
or U19247 (N_19247,N_18068,N_18402);
xnor U19248 (N_19248,N_18945,N_18463);
or U19249 (N_19249,N_18516,N_18586);
nor U19250 (N_19250,N_18420,N_18540);
nor U19251 (N_19251,N_18079,N_18944);
or U19252 (N_19252,N_18279,N_18361);
nor U19253 (N_19253,N_18003,N_18788);
and U19254 (N_19254,N_18048,N_18269);
xor U19255 (N_19255,N_18776,N_18329);
and U19256 (N_19256,N_18853,N_18278);
xor U19257 (N_19257,N_18918,N_18015);
nand U19258 (N_19258,N_18206,N_18622);
and U19259 (N_19259,N_18758,N_18878);
nor U19260 (N_19260,N_18338,N_18204);
nor U19261 (N_19261,N_18468,N_18255);
or U19262 (N_19262,N_18287,N_18103);
and U19263 (N_19263,N_18290,N_18670);
nand U19264 (N_19264,N_18798,N_18701);
nand U19265 (N_19265,N_18801,N_18127);
nand U19266 (N_19266,N_18768,N_18995);
nand U19267 (N_19267,N_18256,N_18695);
xnor U19268 (N_19268,N_18604,N_18481);
nand U19269 (N_19269,N_18822,N_18647);
nand U19270 (N_19270,N_18577,N_18150);
or U19271 (N_19271,N_18458,N_18169);
nand U19272 (N_19272,N_18595,N_18049);
nor U19273 (N_19273,N_18641,N_18090);
nand U19274 (N_19274,N_18738,N_18033);
nand U19275 (N_19275,N_18553,N_18130);
xor U19276 (N_19276,N_18309,N_18765);
xor U19277 (N_19277,N_18772,N_18441);
xor U19278 (N_19278,N_18791,N_18706);
and U19279 (N_19279,N_18200,N_18608);
or U19280 (N_19280,N_18729,N_18336);
nor U19281 (N_19281,N_18218,N_18928);
nor U19282 (N_19282,N_18062,N_18882);
or U19283 (N_19283,N_18713,N_18101);
or U19284 (N_19284,N_18659,N_18455);
or U19285 (N_19285,N_18534,N_18569);
and U19286 (N_19286,N_18094,N_18677);
nand U19287 (N_19287,N_18696,N_18217);
xnor U19288 (N_19288,N_18909,N_18099);
xnor U19289 (N_19289,N_18673,N_18473);
and U19290 (N_19290,N_18274,N_18890);
xnor U19291 (N_19291,N_18559,N_18833);
and U19292 (N_19292,N_18634,N_18905);
and U19293 (N_19293,N_18611,N_18649);
xor U19294 (N_19294,N_18423,N_18989);
or U19295 (N_19295,N_18666,N_18590);
nor U19296 (N_19296,N_18251,N_18041);
nand U19297 (N_19297,N_18203,N_18231);
xor U19298 (N_19298,N_18992,N_18100);
nor U19299 (N_19299,N_18479,N_18813);
xor U19300 (N_19300,N_18208,N_18069);
or U19301 (N_19301,N_18108,N_18594);
or U19302 (N_19302,N_18021,N_18717);
and U19303 (N_19303,N_18831,N_18185);
nand U19304 (N_19304,N_18959,N_18564);
xnor U19305 (N_19305,N_18365,N_18855);
and U19306 (N_19306,N_18775,N_18645);
and U19307 (N_19307,N_18234,N_18740);
nand U19308 (N_19308,N_18723,N_18360);
and U19309 (N_19309,N_18934,N_18076);
nand U19310 (N_19310,N_18915,N_18205);
nor U19311 (N_19311,N_18266,N_18661);
nand U19312 (N_19312,N_18371,N_18387);
xor U19313 (N_19313,N_18331,N_18404);
and U19314 (N_19314,N_18097,N_18519);
or U19315 (N_19315,N_18381,N_18974);
xor U19316 (N_19316,N_18233,N_18380);
xnor U19317 (N_19317,N_18879,N_18320);
nand U19318 (N_19318,N_18521,N_18665);
nand U19319 (N_19319,N_18496,N_18176);
xor U19320 (N_19320,N_18876,N_18214);
nand U19321 (N_19321,N_18494,N_18549);
nor U19322 (N_19322,N_18282,N_18957);
or U19323 (N_19323,N_18092,N_18821);
and U19324 (N_19324,N_18763,N_18177);
and U19325 (N_19325,N_18311,N_18916);
and U19326 (N_19326,N_18152,N_18924);
or U19327 (N_19327,N_18674,N_18967);
nor U19328 (N_19328,N_18638,N_18343);
xnor U19329 (N_19329,N_18047,N_18181);
nor U19330 (N_19330,N_18615,N_18066);
xnor U19331 (N_19331,N_18766,N_18612);
nand U19332 (N_19332,N_18195,N_18588);
or U19333 (N_19333,N_18864,N_18019);
nor U19334 (N_19334,N_18579,N_18936);
nor U19335 (N_19335,N_18624,N_18698);
or U19336 (N_19336,N_18419,N_18752);
and U19337 (N_19337,N_18248,N_18367);
or U19338 (N_19338,N_18000,N_18345);
and U19339 (N_19339,N_18323,N_18745);
nand U19340 (N_19340,N_18307,N_18884);
nor U19341 (N_19341,N_18133,N_18501);
and U19342 (N_19342,N_18178,N_18249);
nand U19343 (N_19343,N_18333,N_18710);
and U19344 (N_19344,N_18335,N_18317);
nor U19345 (N_19345,N_18795,N_18907);
xor U19346 (N_19346,N_18128,N_18509);
nor U19347 (N_19347,N_18690,N_18964);
xnor U19348 (N_19348,N_18919,N_18794);
or U19349 (N_19349,N_18796,N_18460);
nor U19350 (N_19350,N_18819,N_18451);
or U19351 (N_19351,N_18471,N_18024);
nor U19352 (N_19352,N_18653,N_18543);
nor U19353 (N_19353,N_18391,N_18016);
or U19354 (N_19354,N_18313,N_18063);
nand U19355 (N_19355,N_18977,N_18774);
nor U19356 (N_19356,N_18599,N_18407);
or U19357 (N_19357,N_18120,N_18908);
nor U19358 (N_19358,N_18606,N_18245);
xnor U19359 (N_19359,N_18252,N_18339);
or U19360 (N_19360,N_18877,N_18265);
xnor U19361 (N_19361,N_18437,N_18227);
or U19362 (N_19362,N_18083,N_18572);
xor U19363 (N_19363,N_18259,N_18963);
xor U19364 (N_19364,N_18188,N_18226);
nand U19365 (N_19365,N_18515,N_18655);
or U19366 (N_19366,N_18297,N_18593);
nor U19367 (N_19367,N_18221,N_18523);
nor U19368 (N_19368,N_18836,N_18193);
or U19369 (N_19369,N_18854,N_18040);
and U19370 (N_19370,N_18112,N_18952);
and U19371 (N_19371,N_18238,N_18190);
nand U19372 (N_19372,N_18292,N_18725);
nor U19373 (N_19373,N_18988,N_18556);
xnor U19374 (N_19374,N_18412,N_18947);
or U19375 (N_19375,N_18435,N_18950);
nand U19376 (N_19376,N_18034,N_18533);
nand U19377 (N_19377,N_18277,N_18372);
or U19378 (N_19378,N_18512,N_18949);
nor U19379 (N_19379,N_18814,N_18240);
nor U19380 (N_19380,N_18413,N_18685);
xor U19381 (N_19381,N_18660,N_18601);
xor U19382 (N_19382,N_18119,N_18306);
or U19383 (N_19383,N_18513,N_18990);
nor U19384 (N_19384,N_18142,N_18011);
and U19385 (N_19385,N_18626,N_18770);
xnor U19386 (N_19386,N_18749,N_18495);
nor U19387 (N_19387,N_18475,N_18976);
and U19388 (N_19388,N_18137,N_18708);
and U19389 (N_19389,N_18480,N_18330);
nor U19390 (N_19390,N_18537,N_18629);
and U19391 (N_19391,N_18873,N_18469);
xor U19392 (N_19392,N_18464,N_18294);
and U19393 (N_19393,N_18401,N_18116);
nand U19394 (N_19394,N_18344,N_18291);
and U19395 (N_19395,N_18123,N_18600);
xor U19396 (N_19396,N_18506,N_18927);
or U19397 (N_19397,N_18664,N_18633);
nor U19398 (N_19398,N_18620,N_18714);
nand U19399 (N_19399,N_18886,N_18614);
and U19400 (N_19400,N_18984,N_18428);
and U19401 (N_19401,N_18373,N_18790);
nor U19402 (N_19402,N_18050,N_18868);
nor U19403 (N_19403,N_18379,N_18308);
or U19404 (N_19404,N_18581,N_18835);
nor U19405 (N_19405,N_18903,N_18783);
or U19406 (N_19406,N_18987,N_18134);
or U19407 (N_19407,N_18702,N_18093);
xnor U19408 (N_19408,N_18005,N_18414);
xor U19409 (N_19409,N_18803,N_18939);
or U19410 (N_19410,N_18162,N_18268);
or U19411 (N_19411,N_18301,N_18337);
or U19412 (N_19412,N_18146,N_18408);
nand U19413 (N_19413,N_18800,N_18129);
xnor U19414 (N_19414,N_18433,N_18910);
or U19415 (N_19415,N_18263,N_18196);
and U19416 (N_19416,N_18743,N_18465);
nand U19417 (N_19417,N_18718,N_18900);
nand U19418 (N_19418,N_18289,N_18517);
or U19419 (N_19419,N_18472,N_18406);
or U19420 (N_19420,N_18923,N_18023);
and U19421 (N_19421,N_18020,N_18996);
nand U19422 (N_19422,N_18232,N_18754);
and U19423 (N_19423,N_18382,N_18145);
and U19424 (N_19424,N_18899,N_18340);
nor U19425 (N_19425,N_18753,N_18554);
and U19426 (N_19426,N_18842,N_18359);
nand U19427 (N_19427,N_18425,N_18829);
xnor U19428 (N_19428,N_18244,N_18275);
and U19429 (N_19429,N_18922,N_18386);
nor U19430 (N_19430,N_18888,N_18353);
nand U19431 (N_19431,N_18510,N_18751);
or U19432 (N_19432,N_18347,N_18439);
and U19433 (N_19433,N_18571,N_18319);
and U19434 (N_19434,N_18327,N_18022);
xor U19435 (N_19435,N_18462,N_18261);
and U19436 (N_19436,N_18499,N_18806);
nand U19437 (N_19437,N_18576,N_18358);
or U19438 (N_19438,N_18979,N_18767);
and U19439 (N_19439,N_18161,N_18640);
nand U19440 (N_19440,N_18667,N_18709);
xor U19441 (N_19441,N_18867,N_18153);
xor U19442 (N_19442,N_18539,N_18650);
or U19443 (N_19443,N_18627,N_18409);
xor U19444 (N_19444,N_18417,N_18973);
nor U19445 (N_19445,N_18613,N_18780);
nand U19446 (N_19446,N_18253,N_18637);
nor U19447 (N_19447,N_18731,N_18644);
xnor U19448 (N_19448,N_18254,N_18355);
nor U19449 (N_19449,N_18546,N_18175);
or U19450 (N_19450,N_18889,N_18547);
and U19451 (N_19451,N_18452,N_18225);
or U19452 (N_19452,N_18284,N_18342);
or U19453 (N_19453,N_18125,N_18403);
nand U19454 (N_19454,N_18295,N_18111);
and U19455 (N_19455,N_18732,N_18141);
and U19456 (N_19456,N_18449,N_18954);
or U19457 (N_19457,N_18684,N_18210);
or U19458 (N_19458,N_18148,N_18892);
and U19459 (N_19459,N_18865,N_18035);
and U19460 (N_19460,N_18201,N_18514);
nand U19461 (N_19461,N_18105,N_18737);
or U19462 (N_19462,N_18230,N_18935);
xor U19463 (N_19463,N_18728,N_18883);
nand U19464 (N_19464,N_18316,N_18239);
nand U19465 (N_19465,N_18972,N_18628);
or U19466 (N_19466,N_18722,N_18981);
or U19467 (N_19467,N_18527,N_18560);
and U19468 (N_19468,N_18810,N_18820);
or U19469 (N_19469,N_18940,N_18705);
or U19470 (N_19470,N_18366,N_18085);
nand U19471 (N_19471,N_18055,N_18902);
and U19472 (N_19472,N_18457,N_18805);
xnor U19473 (N_19473,N_18912,N_18194);
and U19474 (N_19474,N_18703,N_18561);
or U19475 (N_19475,N_18215,N_18072);
xnor U19476 (N_19476,N_18866,N_18834);
and U19477 (N_19477,N_18060,N_18943);
nand U19478 (N_19478,N_18159,N_18917);
nor U19479 (N_19479,N_18484,N_18609);
and U19480 (N_19480,N_18456,N_18029);
nand U19481 (N_19481,N_18558,N_18933);
nand U19482 (N_19482,N_18071,N_18955);
and U19483 (N_19483,N_18735,N_18179);
xor U19484 (N_19484,N_18802,N_18039);
nand U19485 (N_19485,N_18750,N_18998);
or U19486 (N_19486,N_18662,N_18211);
xnor U19487 (N_19487,N_18043,N_18507);
and U19488 (N_19488,N_18416,N_18518);
and U19489 (N_19489,N_18044,N_18377);
nor U19490 (N_19490,N_18712,N_18183);
nor U19491 (N_19491,N_18426,N_18719);
xnor U19492 (N_19492,N_18491,N_18498);
nand U19493 (N_19493,N_18271,N_18242);
nor U19494 (N_19494,N_18486,N_18583);
xnor U19495 (N_19495,N_18555,N_18807);
xnor U19496 (N_19496,N_18823,N_18602);
xor U19497 (N_19497,N_18081,N_18618);
nand U19498 (N_19498,N_18975,N_18140);
nor U19499 (N_19499,N_18151,N_18257);
nor U19500 (N_19500,N_18213,N_18841);
xor U19501 (N_19501,N_18965,N_18255);
xnor U19502 (N_19502,N_18352,N_18075);
nor U19503 (N_19503,N_18029,N_18636);
nand U19504 (N_19504,N_18541,N_18108);
nor U19505 (N_19505,N_18992,N_18494);
nand U19506 (N_19506,N_18564,N_18972);
or U19507 (N_19507,N_18424,N_18948);
and U19508 (N_19508,N_18512,N_18886);
nand U19509 (N_19509,N_18650,N_18161);
nand U19510 (N_19510,N_18162,N_18798);
xnor U19511 (N_19511,N_18931,N_18901);
or U19512 (N_19512,N_18372,N_18263);
or U19513 (N_19513,N_18932,N_18397);
and U19514 (N_19514,N_18281,N_18889);
nor U19515 (N_19515,N_18782,N_18799);
and U19516 (N_19516,N_18343,N_18458);
or U19517 (N_19517,N_18708,N_18439);
or U19518 (N_19518,N_18102,N_18041);
and U19519 (N_19519,N_18927,N_18850);
nor U19520 (N_19520,N_18329,N_18646);
xor U19521 (N_19521,N_18863,N_18425);
nor U19522 (N_19522,N_18363,N_18564);
xor U19523 (N_19523,N_18855,N_18979);
nand U19524 (N_19524,N_18426,N_18302);
or U19525 (N_19525,N_18031,N_18159);
and U19526 (N_19526,N_18375,N_18352);
nor U19527 (N_19527,N_18769,N_18522);
or U19528 (N_19528,N_18173,N_18251);
and U19529 (N_19529,N_18334,N_18693);
nand U19530 (N_19530,N_18767,N_18283);
nor U19531 (N_19531,N_18346,N_18752);
and U19532 (N_19532,N_18934,N_18014);
and U19533 (N_19533,N_18610,N_18690);
xnor U19534 (N_19534,N_18091,N_18123);
and U19535 (N_19535,N_18378,N_18711);
nor U19536 (N_19536,N_18454,N_18073);
xnor U19537 (N_19537,N_18233,N_18511);
xnor U19538 (N_19538,N_18198,N_18140);
and U19539 (N_19539,N_18574,N_18893);
xor U19540 (N_19540,N_18005,N_18409);
nand U19541 (N_19541,N_18471,N_18202);
and U19542 (N_19542,N_18229,N_18440);
xor U19543 (N_19543,N_18232,N_18535);
nand U19544 (N_19544,N_18273,N_18938);
and U19545 (N_19545,N_18854,N_18868);
and U19546 (N_19546,N_18042,N_18910);
nor U19547 (N_19547,N_18318,N_18498);
nand U19548 (N_19548,N_18027,N_18257);
and U19549 (N_19549,N_18408,N_18011);
xnor U19550 (N_19550,N_18969,N_18015);
xor U19551 (N_19551,N_18818,N_18675);
or U19552 (N_19552,N_18022,N_18379);
or U19553 (N_19553,N_18591,N_18628);
and U19554 (N_19554,N_18577,N_18011);
nor U19555 (N_19555,N_18136,N_18929);
and U19556 (N_19556,N_18604,N_18463);
or U19557 (N_19557,N_18826,N_18322);
or U19558 (N_19558,N_18410,N_18869);
or U19559 (N_19559,N_18098,N_18680);
nand U19560 (N_19560,N_18953,N_18297);
nand U19561 (N_19561,N_18872,N_18521);
nor U19562 (N_19562,N_18369,N_18039);
nand U19563 (N_19563,N_18246,N_18826);
or U19564 (N_19564,N_18230,N_18481);
xnor U19565 (N_19565,N_18795,N_18602);
xor U19566 (N_19566,N_18283,N_18231);
xor U19567 (N_19567,N_18075,N_18438);
and U19568 (N_19568,N_18984,N_18946);
and U19569 (N_19569,N_18363,N_18636);
and U19570 (N_19570,N_18069,N_18917);
or U19571 (N_19571,N_18312,N_18133);
and U19572 (N_19572,N_18936,N_18942);
xor U19573 (N_19573,N_18256,N_18979);
xnor U19574 (N_19574,N_18776,N_18875);
xnor U19575 (N_19575,N_18005,N_18691);
nor U19576 (N_19576,N_18125,N_18145);
nor U19577 (N_19577,N_18448,N_18823);
nor U19578 (N_19578,N_18536,N_18231);
nor U19579 (N_19579,N_18420,N_18193);
and U19580 (N_19580,N_18554,N_18542);
and U19581 (N_19581,N_18249,N_18101);
nand U19582 (N_19582,N_18159,N_18495);
nor U19583 (N_19583,N_18530,N_18374);
xnor U19584 (N_19584,N_18083,N_18619);
or U19585 (N_19585,N_18175,N_18035);
nor U19586 (N_19586,N_18479,N_18641);
xor U19587 (N_19587,N_18057,N_18436);
and U19588 (N_19588,N_18382,N_18690);
or U19589 (N_19589,N_18628,N_18558);
xnor U19590 (N_19590,N_18203,N_18643);
and U19591 (N_19591,N_18244,N_18477);
or U19592 (N_19592,N_18794,N_18416);
nor U19593 (N_19593,N_18855,N_18778);
xnor U19594 (N_19594,N_18541,N_18447);
and U19595 (N_19595,N_18489,N_18208);
nand U19596 (N_19596,N_18374,N_18174);
nor U19597 (N_19597,N_18660,N_18123);
or U19598 (N_19598,N_18478,N_18368);
and U19599 (N_19599,N_18757,N_18981);
nor U19600 (N_19600,N_18271,N_18658);
and U19601 (N_19601,N_18054,N_18404);
nor U19602 (N_19602,N_18856,N_18963);
xnor U19603 (N_19603,N_18898,N_18834);
nor U19604 (N_19604,N_18124,N_18235);
xnor U19605 (N_19605,N_18372,N_18032);
xor U19606 (N_19606,N_18468,N_18759);
nor U19607 (N_19607,N_18312,N_18241);
or U19608 (N_19608,N_18608,N_18924);
nand U19609 (N_19609,N_18201,N_18326);
nand U19610 (N_19610,N_18775,N_18179);
or U19611 (N_19611,N_18746,N_18729);
xnor U19612 (N_19612,N_18790,N_18843);
or U19613 (N_19613,N_18253,N_18186);
nor U19614 (N_19614,N_18838,N_18292);
nor U19615 (N_19615,N_18679,N_18434);
nand U19616 (N_19616,N_18838,N_18085);
nand U19617 (N_19617,N_18147,N_18749);
xor U19618 (N_19618,N_18013,N_18305);
and U19619 (N_19619,N_18182,N_18432);
nand U19620 (N_19620,N_18274,N_18998);
or U19621 (N_19621,N_18400,N_18978);
nand U19622 (N_19622,N_18943,N_18393);
nand U19623 (N_19623,N_18448,N_18484);
and U19624 (N_19624,N_18537,N_18084);
or U19625 (N_19625,N_18172,N_18862);
and U19626 (N_19626,N_18242,N_18895);
or U19627 (N_19627,N_18441,N_18042);
nand U19628 (N_19628,N_18519,N_18554);
nor U19629 (N_19629,N_18711,N_18412);
nor U19630 (N_19630,N_18049,N_18612);
and U19631 (N_19631,N_18688,N_18922);
or U19632 (N_19632,N_18421,N_18052);
nor U19633 (N_19633,N_18784,N_18486);
or U19634 (N_19634,N_18296,N_18563);
xor U19635 (N_19635,N_18104,N_18821);
and U19636 (N_19636,N_18371,N_18833);
or U19637 (N_19637,N_18192,N_18572);
xnor U19638 (N_19638,N_18158,N_18447);
or U19639 (N_19639,N_18179,N_18247);
or U19640 (N_19640,N_18991,N_18739);
or U19641 (N_19641,N_18263,N_18235);
nand U19642 (N_19642,N_18432,N_18260);
or U19643 (N_19643,N_18732,N_18598);
nor U19644 (N_19644,N_18072,N_18913);
xor U19645 (N_19645,N_18710,N_18316);
nor U19646 (N_19646,N_18418,N_18977);
nor U19647 (N_19647,N_18802,N_18568);
or U19648 (N_19648,N_18823,N_18933);
or U19649 (N_19649,N_18864,N_18220);
nand U19650 (N_19650,N_18581,N_18990);
or U19651 (N_19651,N_18213,N_18752);
xor U19652 (N_19652,N_18813,N_18396);
or U19653 (N_19653,N_18005,N_18900);
and U19654 (N_19654,N_18807,N_18620);
nor U19655 (N_19655,N_18384,N_18625);
nor U19656 (N_19656,N_18488,N_18830);
nand U19657 (N_19657,N_18100,N_18359);
nor U19658 (N_19658,N_18120,N_18555);
nand U19659 (N_19659,N_18123,N_18555);
nor U19660 (N_19660,N_18682,N_18493);
xor U19661 (N_19661,N_18574,N_18645);
and U19662 (N_19662,N_18726,N_18159);
nor U19663 (N_19663,N_18616,N_18991);
or U19664 (N_19664,N_18209,N_18666);
nand U19665 (N_19665,N_18669,N_18918);
nand U19666 (N_19666,N_18838,N_18228);
or U19667 (N_19667,N_18265,N_18488);
nand U19668 (N_19668,N_18679,N_18551);
xnor U19669 (N_19669,N_18343,N_18460);
nor U19670 (N_19670,N_18107,N_18480);
nand U19671 (N_19671,N_18856,N_18994);
nor U19672 (N_19672,N_18773,N_18379);
nand U19673 (N_19673,N_18124,N_18415);
nand U19674 (N_19674,N_18953,N_18124);
xnor U19675 (N_19675,N_18298,N_18149);
and U19676 (N_19676,N_18184,N_18666);
or U19677 (N_19677,N_18999,N_18972);
nor U19678 (N_19678,N_18668,N_18289);
nand U19679 (N_19679,N_18287,N_18206);
xnor U19680 (N_19680,N_18172,N_18023);
and U19681 (N_19681,N_18699,N_18459);
or U19682 (N_19682,N_18441,N_18587);
xor U19683 (N_19683,N_18123,N_18796);
nor U19684 (N_19684,N_18290,N_18458);
and U19685 (N_19685,N_18679,N_18348);
nor U19686 (N_19686,N_18835,N_18500);
or U19687 (N_19687,N_18048,N_18950);
nor U19688 (N_19688,N_18647,N_18359);
nor U19689 (N_19689,N_18867,N_18124);
or U19690 (N_19690,N_18691,N_18478);
or U19691 (N_19691,N_18353,N_18175);
xnor U19692 (N_19692,N_18804,N_18809);
xnor U19693 (N_19693,N_18633,N_18867);
and U19694 (N_19694,N_18367,N_18766);
or U19695 (N_19695,N_18172,N_18299);
nand U19696 (N_19696,N_18312,N_18753);
or U19697 (N_19697,N_18216,N_18974);
or U19698 (N_19698,N_18150,N_18430);
xor U19699 (N_19699,N_18559,N_18293);
nand U19700 (N_19700,N_18614,N_18972);
and U19701 (N_19701,N_18417,N_18457);
nor U19702 (N_19702,N_18646,N_18937);
or U19703 (N_19703,N_18572,N_18296);
or U19704 (N_19704,N_18252,N_18655);
xnor U19705 (N_19705,N_18574,N_18355);
nand U19706 (N_19706,N_18800,N_18691);
nor U19707 (N_19707,N_18695,N_18593);
xor U19708 (N_19708,N_18761,N_18810);
nand U19709 (N_19709,N_18019,N_18442);
nand U19710 (N_19710,N_18878,N_18543);
or U19711 (N_19711,N_18694,N_18003);
xor U19712 (N_19712,N_18589,N_18951);
nor U19713 (N_19713,N_18770,N_18476);
and U19714 (N_19714,N_18878,N_18830);
nor U19715 (N_19715,N_18115,N_18510);
nor U19716 (N_19716,N_18764,N_18437);
nor U19717 (N_19717,N_18958,N_18847);
nor U19718 (N_19718,N_18397,N_18227);
nand U19719 (N_19719,N_18681,N_18337);
and U19720 (N_19720,N_18770,N_18784);
or U19721 (N_19721,N_18306,N_18641);
or U19722 (N_19722,N_18989,N_18229);
nand U19723 (N_19723,N_18006,N_18525);
and U19724 (N_19724,N_18006,N_18731);
nor U19725 (N_19725,N_18171,N_18740);
nor U19726 (N_19726,N_18081,N_18358);
or U19727 (N_19727,N_18948,N_18915);
nor U19728 (N_19728,N_18836,N_18837);
nor U19729 (N_19729,N_18409,N_18541);
xnor U19730 (N_19730,N_18931,N_18993);
xnor U19731 (N_19731,N_18592,N_18451);
nor U19732 (N_19732,N_18002,N_18667);
and U19733 (N_19733,N_18874,N_18214);
xor U19734 (N_19734,N_18875,N_18258);
nand U19735 (N_19735,N_18833,N_18731);
or U19736 (N_19736,N_18840,N_18792);
and U19737 (N_19737,N_18012,N_18243);
nor U19738 (N_19738,N_18369,N_18246);
nor U19739 (N_19739,N_18817,N_18382);
nor U19740 (N_19740,N_18734,N_18480);
or U19741 (N_19741,N_18889,N_18348);
nand U19742 (N_19742,N_18598,N_18913);
nor U19743 (N_19743,N_18308,N_18971);
and U19744 (N_19744,N_18996,N_18165);
and U19745 (N_19745,N_18334,N_18626);
or U19746 (N_19746,N_18185,N_18328);
and U19747 (N_19747,N_18600,N_18372);
xnor U19748 (N_19748,N_18714,N_18500);
nor U19749 (N_19749,N_18260,N_18704);
or U19750 (N_19750,N_18199,N_18191);
or U19751 (N_19751,N_18766,N_18525);
nand U19752 (N_19752,N_18858,N_18927);
nor U19753 (N_19753,N_18935,N_18337);
xor U19754 (N_19754,N_18428,N_18412);
and U19755 (N_19755,N_18115,N_18782);
nor U19756 (N_19756,N_18050,N_18349);
nor U19757 (N_19757,N_18309,N_18639);
nand U19758 (N_19758,N_18565,N_18556);
nand U19759 (N_19759,N_18042,N_18823);
xor U19760 (N_19760,N_18135,N_18736);
xnor U19761 (N_19761,N_18357,N_18765);
xnor U19762 (N_19762,N_18808,N_18412);
xor U19763 (N_19763,N_18578,N_18132);
nand U19764 (N_19764,N_18774,N_18285);
and U19765 (N_19765,N_18079,N_18663);
and U19766 (N_19766,N_18168,N_18454);
nor U19767 (N_19767,N_18110,N_18289);
nand U19768 (N_19768,N_18382,N_18052);
and U19769 (N_19769,N_18380,N_18873);
nor U19770 (N_19770,N_18404,N_18196);
nand U19771 (N_19771,N_18920,N_18454);
xnor U19772 (N_19772,N_18883,N_18342);
nand U19773 (N_19773,N_18084,N_18890);
nand U19774 (N_19774,N_18692,N_18826);
xnor U19775 (N_19775,N_18184,N_18754);
nand U19776 (N_19776,N_18522,N_18946);
nand U19777 (N_19777,N_18365,N_18369);
or U19778 (N_19778,N_18807,N_18816);
xnor U19779 (N_19779,N_18862,N_18368);
nand U19780 (N_19780,N_18720,N_18573);
or U19781 (N_19781,N_18000,N_18235);
nand U19782 (N_19782,N_18850,N_18020);
nor U19783 (N_19783,N_18904,N_18360);
xnor U19784 (N_19784,N_18125,N_18270);
and U19785 (N_19785,N_18453,N_18669);
or U19786 (N_19786,N_18613,N_18809);
nand U19787 (N_19787,N_18005,N_18306);
nor U19788 (N_19788,N_18297,N_18734);
or U19789 (N_19789,N_18858,N_18387);
nor U19790 (N_19790,N_18359,N_18707);
nor U19791 (N_19791,N_18259,N_18797);
nand U19792 (N_19792,N_18871,N_18966);
and U19793 (N_19793,N_18206,N_18160);
nor U19794 (N_19794,N_18433,N_18703);
xnor U19795 (N_19795,N_18255,N_18361);
nand U19796 (N_19796,N_18671,N_18045);
nor U19797 (N_19797,N_18488,N_18460);
nand U19798 (N_19798,N_18932,N_18155);
xnor U19799 (N_19799,N_18013,N_18584);
and U19800 (N_19800,N_18794,N_18576);
nor U19801 (N_19801,N_18802,N_18557);
and U19802 (N_19802,N_18133,N_18733);
and U19803 (N_19803,N_18209,N_18898);
and U19804 (N_19804,N_18224,N_18548);
and U19805 (N_19805,N_18021,N_18551);
nand U19806 (N_19806,N_18178,N_18924);
xor U19807 (N_19807,N_18287,N_18516);
and U19808 (N_19808,N_18936,N_18273);
or U19809 (N_19809,N_18339,N_18516);
and U19810 (N_19810,N_18729,N_18668);
or U19811 (N_19811,N_18017,N_18439);
nand U19812 (N_19812,N_18482,N_18429);
and U19813 (N_19813,N_18976,N_18980);
nor U19814 (N_19814,N_18815,N_18694);
nor U19815 (N_19815,N_18322,N_18601);
or U19816 (N_19816,N_18033,N_18174);
xor U19817 (N_19817,N_18750,N_18566);
or U19818 (N_19818,N_18836,N_18121);
or U19819 (N_19819,N_18147,N_18928);
nand U19820 (N_19820,N_18184,N_18976);
or U19821 (N_19821,N_18942,N_18398);
or U19822 (N_19822,N_18640,N_18747);
and U19823 (N_19823,N_18140,N_18532);
xor U19824 (N_19824,N_18270,N_18441);
and U19825 (N_19825,N_18775,N_18500);
or U19826 (N_19826,N_18643,N_18360);
nand U19827 (N_19827,N_18030,N_18549);
or U19828 (N_19828,N_18293,N_18808);
or U19829 (N_19829,N_18663,N_18436);
xnor U19830 (N_19830,N_18788,N_18404);
and U19831 (N_19831,N_18998,N_18256);
nand U19832 (N_19832,N_18773,N_18279);
nor U19833 (N_19833,N_18502,N_18228);
nor U19834 (N_19834,N_18950,N_18150);
or U19835 (N_19835,N_18374,N_18432);
and U19836 (N_19836,N_18777,N_18471);
nor U19837 (N_19837,N_18734,N_18716);
nand U19838 (N_19838,N_18563,N_18674);
xor U19839 (N_19839,N_18115,N_18192);
nor U19840 (N_19840,N_18405,N_18452);
or U19841 (N_19841,N_18368,N_18224);
xor U19842 (N_19842,N_18631,N_18453);
nor U19843 (N_19843,N_18518,N_18984);
or U19844 (N_19844,N_18353,N_18459);
nand U19845 (N_19845,N_18167,N_18515);
xor U19846 (N_19846,N_18754,N_18712);
nand U19847 (N_19847,N_18530,N_18471);
xor U19848 (N_19848,N_18558,N_18083);
nor U19849 (N_19849,N_18529,N_18563);
nand U19850 (N_19850,N_18746,N_18900);
nor U19851 (N_19851,N_18342,N_18720);
nand U19852 (N_19852,N_18769,N_18317);
nand U19853 (N_19853,N_18377,N_18212);
or U19854 (N_19854,N_18998,N_18790);
nand U19855 (N_19855,N_18443,N_18220);
nor U19856 (N_19856,N_18589,N_18340);
nand U19857 (N_19857,N_18926,N_18978);
nand U19858 (N_19858,N_18118,N_18736);
nor U19859 (N_19859,N_18653,N_18198);
or U19860 (N_19860,N_18691,N_18628);
and U19861 (N_19861,N_18252,N_18325);
xnor U19862 (N_19862,N_18764,N_18752);
and U19863 (N_19863,N_18509,N_18087);
xnor U19864 (N_19864,N_18761,N_18220);
or U19865 (N_19865,N_18629,N_18483);
nand U19866 (N_19866,N_18701,N_18618);
nand U19867 (N_19867,N_18682,N_18945);
nor U19868 (N_19868,N_18151,N_18260);
nand U19869 (N_19869,N_18480,N_18442);
or U19870 (N_19870,N_18484,N_18074);
and U19871 (N_19871,N_18353,N_18305);
xnor U19872 (N_19872,N_18181,N_18625);
and U19873 (N_19873,N_18722,N_18507);
and U19874 (N_19874,N_18890,N_18196);
or U19875 (N_19875,N_18800,N_18505);
nand U19876 (N_19876,N_18935,N_18716);
nand U19877 (N_19877,N_18380,N_18980);
and U19878 (N_19878,N_18424,N_18741);
nor U19879 (N_19879,N_18275,N_18973);
xnor U19880 (N_19880,N_18078,N_18491);
xor U19881 (N_19881,N_18639,N_18056);
nor U19882 (N_19882,N_18490,N_18781);
nand U19883 (N_19883,N_18313,N_18197);
nor U19884 (N_19884,N_18631,N_18437);
nand U19885 (N_19885,N_18586,N_18891);
or U19886 (N_19886,N_18971,N_18583);
or U19887 (N_19887,N_18737,N_18194);
and U19888 (N_19888,N_18613,N_18412);
nor U19889 (N_19889,N_18906,N_18000);
and U19890 (N_19890,N_18447,N_18645);
and U19891 (N_19891,N_18227,N_18896);
or U19892 (N_19892,N_18132,N_18278);
nand U19893 (N_19893,N_18593,N_18682);
or U19894 (N_19894,N_18182,N_18814);
nand U19895 (N_19895,N_18312,N_18596);
or U19896 (N_19896,N_18664,N_18370);
xnor U19897 (N_19897,N_18495,N_18265);
nor U19898 (N_19898,N_18802,N_18603);
nor U19899 (N_19899,N_18626,N_18661);
or U19900 (N_19900,N_18703,N_18281);
or U19901 (N_19901,N_18973,N_18930);
and U19902 (N_19902,N_18658,N_18669);
xnor U19903 (N_19903,N_18233,N_18742);
and U19904 (N_19904,N_18192,N_18350);
nor U19905 (N_19905,N_18267,N_18841);
nor U19906 (N_19906,N_18339,N_18467);
and U19907 (N_19907,N_18893,N_18416);
nor U19908 (N_19908,N_18377,N_18568);
nand U19909 (N_19909,N_18507,N_18604);
and U19910 (N_19910,N_18073,N_18740);
or U19911 (N_19911,N_18783,N_18248);
xnor U19912 (N_19912,N_18568,N_18906);
nor U19913 (N_19913,N_18136,N_18371);
nor U19914 (N_19914,N_18324,N_18965);
nand U19915 (N_19915,N_18670,N_18168);
or U19916 (N_19916,N_18560,N_18491);
and U19917 (N_19917,N_18504,N_18625);
nand U19918 (N_19918,N_18331,N_18731);
nor U19919 (N_19919,N_18427,N_18998);
or U19920 (N_19920,N_18019,N_18992);
nor U19921 (N_19921,N_18077,N_18176);
nand U19922 (N_19922,N_18171,N_18808);
nand U19923 (N_19923,N_18540,N_18687);
xnor U19924 (N_19924,N_18900,N_18268);
xor U19925 (N_19925,N_18920,N_18179);
nand U19926 (N_19926,N_18346,N_18131);
xnor U19927 (N_19927,N_18813,N_18302);
nand U19928 (N_19928,N_18477,N_18126);
nor U19929 (N_19929,N_18793,N_18560);
and U19930 (N_19930,N_18764,N_18088);
or U19931 (N_19931,N_18539,N_18890);
nor U19932 (N_19932,N_18974,N_18189);
or U19933 (N_19933,N_18293,N_18064);
nor U19934 (N_19934,N_18588,N_18859);
nand U19935 (N_19935,N_18057,N_18051);
xnor U19936 (N_19936,N_18450,N_18713);
or U19937 (N_19937,N_18472,N_18355);
xor U19938 (N_19938,N_18881,N_18312);
nor U19939 (N_19939,N_18236,N_18406);
and U19940 (N_19940,N_18172,N_18204);
and U19941 (N_19941,N_18826,N_18577);
xor U19942 (N_19942,N_18747,N_18951);
xnor U19943 (N_19943,N_18431,N_18698);
nand U19944 (N_19944,N_18680,N_18795);
and U19945 (N_19945,N_18862,N_18389);
xnor U19946 (N_19946,N_18966,N_18059);
and U19947 (N_19947,N_18323,N_18802);
xnor U19948 (N_19948,N_18361,N_18043);
or U19949 (N_19949,N_18495,N_18183);
xnor U19950 (N_19950,N_18980,N_18453);
xor U19951 (N_19951,N_18531,N_18375);
nand U19952 (N_19952,N_18682,N_18069);
and U19953 (N_19953,N_18751,N_18701);
xnor U19954 (N_19954,N_18600,N_18093);
or U19955 (N_19955,N_18743,N_18432);
nor U19956 (N_19956,N_18886,N_18783);
or U19957 (N_19957,N_18261,N_18790);
xor U19958 (N_19958,N_18825,N_18729);
or U19959 (N_19959,N_18489,N_18007);
or U19960 (N_19960,N_18731,N_18895);
nand U19961 (N_19961,N_18550,N_18850);
or U19962 (N_19962,N_18225,N_18653);
xnor U19963 (N_19963,N_18761,N_18364);
nor U19964 (N_19964,N_18659,N_18485);
and U19965 (N_19965,N_18086,N_18633);
or U19966 (N_19966,N_18722,N_18321);
and U19967 (N_19967,N_18381,N_18302);
or U19968 (N_19968,N_18623,N_18612);
and U19969 (N_19969,N_18068,N_18605);
or U19970 (N_19970,N_18656,N_18648);
or U19971 (N_19971,N_18002,N_18271);
xor U19972 (N_19972,N_18008,N_18792);
nor U19973 (N_19973,N_18042,N_18943);
xnor U19974 (N_19974,N_18491,N_18945);
or U19975 (N_19975,N_18680,N_18131);
xnor U19976 (N_19976,N_18082,N_18039);
or U19977 (N_19977,N_18416,N_18263);
or U19978 (N_19978,N_18533,N_18641);
and U19979 (N_19979,N_18435,N_18065);
xor U19980 (N_19980,N_18250,N_18510);
and U19981 (N_19981,N_18992,N_18516);
nand U19982 (N_19982,N_18179,N_18441);
and U19983 (N_19983,N_18088,N_18625);
xnor U19984 (N_19984,N_18730,N_18942);
nor U19985 (N_19985,N_18169,N_18901);
xnor U19986 (N_19986,N_18569,N_18038);
nor U19987 (N_19987,N_18628,N_18998);
and U19988 (N_19988,N_18242,N_18554);
nor U19989 (N_19989,N_18252,N_18423);
or U19990 (N_19990,N_18847,N_18733);
or U19991 (N_19991,N_18402,N_18887);
xnor U19992 (N_19992,N_18828,N_18846);
xnor U19993 (N_19993,N_18607,N_18311);
and U19994 (N_19994,N_18410,N_18481);
and U19995 (N_19995,N_18207,N_18396);
and U19996 (N_19996,N_18780,N_18311);
and U19997 (N_19997,N_18696,N_18653);
and U19998 (N_19998,N_18531,N_18099);
nand U19999 (N_19999,N_18080,N_18137);
xor U20000 (N_20000,N_19739,N_19466);
or U20001 (N_20001,N_19259,N_19276);
nor U20002 (N_20002,N_19149,N_19371);
xnor U20003 (N_20003,N_19946,N_19881);
or U20004 (N_20004,N_19707,N_19724);
or U20005 (N_20005,N_19275,N_19550);
xor U20006 (N_20006,N_19215,N_19528);
xor U20007 (N_20007,N_19120,N_19570);
xnor U20008 (N_20008,N_19321,N_19091);
xnor U20009 (N_20009,N_19308,N_19362);
nand U20010 (N_20010,N_19110,N_19252);
xor U20011 (N_20011,N_19117,N_19541);
xnor U20012 (N_20012,N_19008,N_19061);
nand U20013 (N_20013,N_19535,N_19883);
or U20014 (N_20014,N_19831,N_19555);
and U20015 (N_20015,N_19886,N_19218);
or U20016 (N_20016,N_19426,N_19345);
or U20017 (N_20017,N_19048,N_19542);
nor U20018 (N_20018,N_19828,N_19403);
xnor U20019 (N_20019,N_19760,N_19441);
or U20020 (N_20020,N_19676,N_19728);
or U20021 (N_20021,N_19818,N_19517);
xor U20022 (N_20022,N_19579,N_19970);
or U20023 (N_20023,N_19556,N_19562);
or U20024 (N_20024,N_19755,N_19625);
nand U20025 (N_20025,N_19855,N_19102);
and U20026 (N_20026,N_19998,N_19282);
nor U20027 (N_20027,N_19750,N_19533);
or U20028 (N_20028,N_19880,N_19684);
nand U20029 (N_20029,N_19501,N_19040);
nor U20030 (N_20030,N_19078,N_19150);
or U20031 (N_20031,N_19730,N_19532);
nor U20032 (N_20032,N_19520,N_19599);
xnor U20033 (N_20033,N_19976,N_19774);
and U20034 (N_20034,N_19165,N_19159);
xnor U20035 (N_20035,N_19234,N_19978);
xnor U20036 (N_20036,N_19004,N_19446);
nand U20037 (N_20037,N_19757,N_19572);
nor U20038 (N_20038,N_19010,N_19055);
xor U20039 (N_20039,N_19648,N_19878);
xnor U20040 (N_20040,N_19833,N_19383);
nand U20041 (N_20041,N_19070,N_19433);
or U20042 (N_20042,N_19047,N_19458);
xor U20043 (N_20043,N_19289,N_19459);
nand U20044 (N_20044,N_19549,N_19935);
xnor U20045 (N_20045,N_19153,N_19546);
or U20046 (N_20046,N_19080,N_19134);
and U20047 (N_20047,N_19772,N_19361);
or U20048 (N_20048,N_19222,N_19493);
xnor U20049 (N_20049,N_19786,N_19644);
and U20050 (N_20050,N_19835,N_19598);
nand U20051 (N_20051,N_19398,N_19630);
and U20052 (N_20052,N_19847,N_19320);
nor U20053 (N_20053,N_19590,N_19177);
nor U20054 (N_20054,N_19233,N_19406);
xnor U20055 (N_20055,N_19206,N_19743);
or U20056 (N_20056,N_19767,N_19677);
xnor U20057 (N_20057,N_19701,N_19793);
or U20058 (N_20058,N_19489,N_19098);
xnor U20059 (N_20059,N_19999,N_19956);
and U20060 (N_20060,N_19508,N_19930);
nand U20061 (N_20061,N_19694,N_19203);
or U20062 (N_20062,N_19924,N_19964);
xnor U20063 (N_20063,N_19175,N_19666);
nand U20064 (N_20064,N_19604,N_19564);
nor U20065 (N_20065,N_19456,N_19805);
nor U20066 (N_20066,N_19011,N_19829);
and U20067 (N_20067,N_19210,N_19360);
nand U20068 (N_20068,N_19425,N_19619);
nor U20069 (N_20069,N_19997,N_19747);
and U20070 (N_20070,N_19926,N_19709);
and U20071 (N_20071,N_19936,N_19525);
nor U20072 (N_20072,N_19950,N_19776);
nor U20073 (N_20073,N_19436,N_19922);
or U20074 (N_20074,N_19605,N_19264);
and U20075 (N_20075,N_19453,N_19132);
xor U20076 (N_20076,N_19717,N_19814);
nand U20077 (N_20077,N_19434,N_19893);
or U20078 (N_20078,N_19601,N_19176);
nand U20079 (N_20079,N_19879,N_19748);
nand U20080 (N_20080,N_19813,N_19867);
and U20081 (N_20081,N_19028,N_19671);
nand U20082 (N_20082,N_19365,N_19791);
or U20083 (N_20083,N_19629,N_19650);
xor U20084 (N_20084,N_19292,N_19286);
xor U20085 (N_20085,N_19863,N_19511);
and U20086 (N_20086,N_19180,N_19049);
and U20087 (N_20087,N_19186,N_19278);
nor U20088 (N_20088,N_19913,N_19692);
and U20089 (N_20089,N_19636,N_19703);
nor U20090 (N_20090,N_19753,N_19375);
nand U20091 (N_20091,N_19868,N_19281);
or U20092 (N_20092,N_19530,N_19784);
nand U20093 (N_20093,N_19521,N_19557);
xnor U20094 (N_20094,N_19626,N_19460);
or U20095 (N_20095,N_19952,N_19302);
or U20096 (N_20096,N_19817,N_19735);
or U20097 (N_20097,N_19085,N_19563);
or U20098 (N_20098,N_19202,N_19343);
or U20099 (N_20099,N_19197,N_19096);
nor U20100 (N_20100,N_19690,N_19418);
and U20101 (N_20101,N_19971,N_19309);
nor U20102 (N_20102,N_19386,N_19337);
nand U20103 (N_20103,N_19440,N_19691);
xor U20104 (N_20104,N_19207,N_19079);
and U20105 (N_20105,N_19545,N_19819);
or U20106 (N_20106,N_19800,N_19189);
nor U20107 (N_20107,N_19733,N_19568);
and U20108 (N_20108,N_19063,N_19097);
nor U20109 (N_20109,N_19696,N_19140);
and U20110 (N_20110,N_19231,N_19645);
and U20111 (N_20111,N_19582,N_19888);
nor U20112 (N_20112,N_19909,N_19307);
nor U20113 (N_20113,N_19391,N_19088);
nor U20114 (N_20114,N_19243,N_19467);
and U20115 (N_20115,N_19890,N_19664);
nor U20116 (N_20116,N_19348,N_19811);
nand U20117 (N_20117,N_19616,N_19439);
nand U20118 (N_20118,N_19499,N_19194);
nand U20119 (N_20119,N_19699,N_19407);
and U20120 (N_20120,N_19591,N_19041);
xor U20121 (N_20121,N_19646,N_19781);
and U20122 (N_20122,N_19181,N_19548);
nand U20123 (N_20123,N_19849,N_19785);
or U20124 (N_20124,N_19109,N_19030);
xnor U20125 (N_20125,N_19857,N_19451);
nand U20126 (N_20126,N_19668,N_19914);
xnor U20127 (N_20127,N_19266,N_19712);
and U20128 (N_20128,N_19838,N_19751);
nor U20129 (N_20129,N_19538,N_19623);
nor U20130 (N_20130,N_19603,N_19864);
nand U20131 (N_20131,N_19704,N_19597);
xnor U20132 (N_20132,N_19363,N_19112);
nand U20133 (N_20133,N_19404,N_19992);
xor U20134 (N_20134,N_19973,N_19587);
nor U20135 (N_20135,N_19370,N_19339);
or U20136 (N_20136,N_19465,N_19066);
nand U20137 (N_20137,N_19839,N_19927);
and U20138 (N_20138,N_19351,N_19770);
nand U20139 (N_20139,N_19050,N_19795);
xor U20140 (N_20140,N_19798,N_19226);
nand U20141 (N_20141,N_19123,N_19042);
xor U20142 (N_20142,N_19141,N_19859);
nand U20143 (N_20143,N_19162,N_19421);
or U20144 (N_20144,N_19090,N_19799);
and U20145 (N_20145,N_19062,N_19283);
nand U20146 (N_20146,N_19214,N_19854);
xnor U20147 (N_20147,N_19801,N_19148);
and U20148 (N_20148,N_19900,N_19653);
nand U20149 (N_20149,N_19230,N_19665);
and U20150 (N_20150,N_19845,N_19155);
nor U20151 (N_20151,N_19114,N_19118);
or U20152 (N_20152,N_19933,N_19953);
or U20153 (N_20153,N_19934,N_19187);
xor U20154 (N_20154,N_19448,N_19746);
and U20155 (N_20155,N_19447,N_19480);
or U20156 (N_20156,N_19990,N_19792);
nor U20157 (N_20157,N_19212,N_19199);
nand U20158 (N_20158,N_19026,N_19469);
or U20159 (N_20159,N_19174,N_19350);
nor U20160 (N_20160,N_19737,N_19726);
nand U20161 (N_20161,N_19624,N_19144);
and U20162 (N_20162,N_19683,N_19216);
nand U20163 (N_20163,N_19412,N_19727);
xnor U20164 (N_20164,N_19399,N_19381);
nor U20165 (N_20165,N_19807,N_19510);
nor U20166 (N_20166,N_19674,N_19734);
nor U20167 (N_20167,N_19172,N_19262);
or U20168 (N_20168,N_19429,N_19325);
xor U20169 (N_20169,N_19200,N_19475);
and U20170 (N_20170,N_19569,N_19208);
nand U20171 (N_20171,N_19306,N_19595);
and U20172 (N_20172,N_19721,N_19167);
nand U20173 (N_20173,N_19269,N_19764);
xnor U20174 (N_20174,N_19505,N_19490);
nand U20175 (N_20175,N_19002,N_19225);
or U20176 (N_20176,N_19494,N_19183);
nor U20177 (N_20177,N_19482,N_19769);
or U20178 (N_20178,N_19198,N_19758);
and U20179 (N_20179,N_19850,N_19871);
or U20180 (N_20180,N_19393,N_19033);
nand U20181 (N_20181,N_19947,N_19506);
xor U20182 (N_20182,N_19100,N_19232);
and U20183 (N_20183,N_19672,N_19938);
or U20184 (N_20184,N_19217,N_19424);
xor U20185 (N_20185,N_19830,N_19223);
nor U20186 (N_20186,N_19586,N_19461);
or U20187 (N_20187,N_19290,N_19300);
nand U20188 (N_20188,N_19168,N_19113);
xor U20189 (N_20189,N_19745,N_19954);
nand U20190 (N_20190,N_19716,N_19824);
xnor U20191 (N_20191,N_19022,N_19497);
xor U20192 (N_20192,N_19977,N_19442);
or U20193 (N_20193,N_19614,N_19827);
and U20194 (N_20194,N_19382,N_19377);
nand U20195 (N_20195,N_19955,N_19897);
and U20196 (N_20196,N_19657,N_19870);
nor U20197 (N_20197,N_19736,N_19277);
or U20198 (N_20198,N_19413,N_19315);
and U20199 (N_20199,N_19613,N_19491);
and U20200 (N_20200,N_19647,N_19876);
nor U20201 (N_20201,N_19143,N_19023);
xnor U20202 (N_20202,N_19633,N_19777);
or U20203 (N_20203,N_19989,N_19488);
and U20204 (N_20204,N_19190,N_19058);
nand U20205 (N_20205,N_19072,N_19017);
and U20206 (N_20206,N_19069,N_19503);
and U20207 (N_20207,N_19108,N_19154);
xor U20208 (N_20208,N_19336,N_19711);
nor U20209 (N_20209,N_19334,N_19620);
or U20210 (N_20210,N_19037,N_19354);
nand U20211 (N_20211,N_19706,N_19679);
nor U20212 (N_20212,N_19009,N_19389);
xnor U20213 (N_20213,N_19156,N_19637);
xnor U20214 (N_20214,N_19732,N_19842);
or U20215 (N_20215,N_19323,N_19660);
or U20216 (N_20216,N_19584,N_19092);
and U20217 (N_20217,N_19941,N_19852);
or U20218 (N_20218,N_19152,N_19236);
nand U20219 (N_20219,N_19073,N_19869);
xor U20220 (N_20220,N_19255,N_19470);
or U20221 (N_20221,N_19116,N_19094);
nand U20222 (N_20222,N_19658,N_19963);
nand U20223 (N_20223,N_19693,N_19039);
or U20224 (N_20224,N_19554,N_19369);
nand U20225 (N_20225,N_19394,N_19103);
and U20226 (N_20226,N_19844,N_19607);
nand U20227 (N_20227,N_19642,N_19364);
nand U20228 (N_20228,N_19249,N_19659);
nor U20229 (N_20229,N_19596,N_19821);
and U20230 (N_20230,N_19722,N_19837);
nand U20231 (N_20231,N_19081,N_19543);
nand U20232 (N_20232,N_19654,N_19552);
and U20233 (N_20233,N_19279,N_19851);
nand U20234 (N_20234,N_19600,N_19430);
and U20235 (N_20235,N_19906,N_19287);
and U20236 (N_20236,N_19498,N_19133);
and U20237 (N_20237,N_19250,N_19898);
nor U20238 (N_20238,N_19787,N_19224);
or U20239 (N_20239,N_19184,N_19241);
or U20240 (N_20240,N_19916,N_19138);
xor U20241 (N_20241,N_19780,N_19661);
nor U20242 (N_20242,N_19247,N_19122);
nand U20243 (N_20243,N_19347,N_19872);
nor U20244 (N_20244,N_19071,N_19500);
xor U20245 (N_20245,N_19324,N_19875);
and U20246 (N_20246,N_19967,N_19944);
nand U20247 (N_20247,N_19067,N_19296);
or U20248 (N_20248,N_19937,N_19723);
nor U20249 (N_20249,N_19809,N_19298);
or U20250 (N_20250,N_19566,N_19411);
or U20251 (N_20251,N_19246,N_19128);
nor U20252 (N_20252,N_19432,N_19884);
xor U20253 (N_20253,N_19877,N_19702);
xnor U20254 (N_20254,N_19708,N_19788);
and U20255 (N_20255,N_19396,N_19720);
and U20256 (N_20256,N_19487,N_19068);
nand U20257 (N_20257,N_19054,N_19353);
and U20258 (N_20258,N_19248,N_19834);
nand U20259 (N_20259,N_19147,N_19327);
and U20260 (N_20260,N_19376,N_19910);
nor U20261 (N_20261,N_19681,N_19305);
and U20262 (N_20262,N_19822,N_19295);
xnor U20263 (N_20263,N_19211,N_19331);
and U20264 (N_20264,N_19558,N_19803);
nor U20265 (N_20265,N_19340,N_19126);
and U20266 (N_20266,N_19573,N_19332);
nand U20267 (N_20267,N_19422,N_19166);
xnor U20268 (N_20268,N_19046,N_19301);
or U20269 (N_20269,N_19127,N_19593);
or U20270 (N_20270,N_19949,N_19643);
xnor U20271 (N_20271,N_19485,N_19534);
nor U20272 (N_20272,N_19841,N_19794);
nor U20273 (N_20273,N_19729,N_19089);
and U20274 (N_20274,N_19789,N_19284);
and U20275 (N_20275,N_19136,N_19478);
and U20276 (N_20276,N_19994,N_19457);
xnor U20277 (N_20277,N_19205,N_19444);
nand U20278 (N_20278,N_19285,N_19638);
and U20279 (N_20279,N_19229,N_19529);
nor U20280 (N_20280,N_19602,N_19965);
nor U20281 (N_20281,N_19484,N_19895);
nor U20282 (N_20282,N_19220,N_19823);
nand U20283 (N_20283,N_19608,N_19227);
nor U20284 (N_20284,N_19239,N_19495);
nor U20285 (N_20285,N_19388,N_19536);
nand U20286 (N_20286,N_19891,N_19330);
nand U20287 (N_20287,N_19059,N_19816);
nor U20288 (N_20288,N_19065,N_19513);
nand U20289 (N_20289,N_19682,N_19966);
xnor U20290 (N_20290,N_19476,N_19471);
nand U20291 (N_20291,N_19316,N_19274);
xor U20292 (N_20292,N_19314,N_19640);
and U20293 (N_20293,N_19450,N_19961);
or U20294 (N_20294,N_19656,N_19996);
nor U20295 (N_20295,N_19044,N_19368);
nor U20296 (N_20296,N_19018,N_19843);
and U20297 (N_20297,N_19960,N_19609);
and U20298 (N_20298,N_19472,N_19991);
nand U20299 (N_20299,N_19718,N_19265);
xnor U20300 (N_20300,N_19449,N_19907);
nor U20301 (N_20301,N_19515,N_19559);
or U20302 (N_20302,N_19084,N_19585);
or U20303 (N_20303,N_19652,N_19235);
xnor U20304 (N_20304,N_19151,N_19341);
nor U20305 (N_20305,N_19826,N_19984);
xor U20306 (N_20306,N_19537,N_19512);
nand U20307 (N_20307,N_19796,N_19387);
nand U20308 (N_20308,N_19420,N_19680);
or U20309 (N_20309,N_19958,N_19052);
nand U20310 (N_20310,N_19612,N_19178);
nand U20311 (N_20311,N_19390,N_19075);
xor U20312 (N_20312,N_19483,N_19583);
and U20313 (N_20313,N_19161,N_19106);
nand U20314 (N_20314,N_19374,N_19917);
xor U20315 (N_20315,N_19105,N_19328);
nor U20316 (N_20316,N_19522,N_19775);
or U20317 (N_20317,N_19384,N_19565);
or U20318 (N_20318,N_19820,N_19409);
and U20319 (N_20319,N_19000,N_19477);
nor U20320 (N_20320,N_19064,N_19628);
or U20321 (N_20321,N_19815,N_19920);
nor U20322 (N_20322,N_19832,N_19021);
nand U20323 (N_20323,N_19311,N_19182);
and U20324 (N_20324,N_19929,N_19445);
xnor U20325 (N_20325,N_19519,N_19244);
and U20326 (N_20326,N_19940,N_19725);
nand U20327 (N_20327,N_19518,N_19082);
nor U20328 (N_20328,N_19812,N_19840);
and U20329 (N_20329,N_19468,N_19032);
nand U20330 (N_20330,N_19860,N_19678);
nor U20331 (N_20331,N_19710,N_19163);
nor U20332 (N_20332,N_19293,N_19051);
and U20333 (N_20333,N_19987,N_19257);
nand U20334 (N_20334,N_19754,N_19901);
nand U20335 (N_20335,N_19146,N_19346);
and U20336 (N_20336,N_19719,N_19288);
nor U20337 (N_20337,N_19270,N_19492);
xor U20338 (N_20338,N_19651,N_19020);
nand U20339 (N_20339,N_19188,N_19509);
nor U20340 (N_20340,N_19761,N_19975);
or U20341 (N_20341,N_19496,N_19372);
or U20342 (N_20342,N_19695,N_19349);
xor U20343 (N_20343,N_19771,N_19256);
or U20344 (N_20344,N_19782,N_19686);
and U20345 (N_20345,N_19083,N_19779);
nand U20346 (N_20346,N_19918,N_19763);
or U20347 (N_20347,N_19580,N_19762);
and U20348 (N_20348,N_19889,N_19939);
nor U20349 (N_20349,N_19303,N_19043);
or U20350 (N_20350,N_19539,N_19025);
nand U20351 (N_20351,N_19213,N_19111);
or U20352 (N_20352,N_19124,N_19036);
xnor U20353 (N_20353,N_19185,N_19254);
or U20354 (N_20354,N_19139,N_19145);
xnor U20355 (N_20355,N_19258,N_19925);
or U20356 (N_20356,N_19669,N_19291);
and U20357 (N_20357,N_19527,N_19479);
nand U20358 (N_20358,N_19627,N_19074);
nand U20359 (N_20359,N_19238,N_19342);
nand U20360 (N_20360,N_19423,N_19931);
xor U20361 (N_20361,N_19344,N_19806);
nand U20362 (N_20362,N_19988,N_19326);
or U20363 (N_20363,N_19474,N_19121);
nand U20364 (N_20364,N_19903,N_19209);
nand U20365 (N_20365,N_19095,N_19195);
nand U20366 (N_20366,N_19983,N_19738);
nor U20367 (N_20367,N_19299,N_19356);
or U20368 (N_20368,N_19621,N_19462);
nand U20369 (N_20369,N_19322,N_19027);
or U20370 (N_20370,N_19959,N_19639);
nand U20371 (N_20371,N_19908,N_19606);
nor U20372 (N_20372,N_19228,N_19401);
or U20373 (N_20373,N_19885,N_19874);
xor U20374 (N_20374,N_19358,N_19982);
nand U20375 (N_20375,N_19012,N_19915);
xnor U20376 (N_20376,N_19561,N_19400);
or U20377 (N_20377,N_19902,N_19431);
nand U20378 (N_20378,N_19853,N_19169);
nor U20379 (N_20379,N_19268,N_19240);
xnor U20380 (N_20380,N_19858,N_19504);
nand U20381 (N_20381,N_19414,N_19649);
and U20382 (N_20382,N_19366,N_19894);
nor U20383 (N_20383,N_19611,N_19700);
or U20384 (N_20384,N_19687,N_19848);
nor U20385 (N_20385,N_19921,N_19130);
or U20386 (N_20386,N_19003,N_19856);
or U20387 (N_20387,N_19663,N_19526);
nand U20388 (N_20388,N_19524,N_19576);
and U20389 (N_20389,N_19435,N_19865);
nor U20390 (N_20390,N_19179,N_19101);
nor U20391 (N_20391,N_19373,N_19896);
or U20392 (N_20392,N_19093,N_19191);
nor U20393 (N_20393,N_19313,N_19419);
and U20394 (N_20394,N_19981,N_19158);
nand U20395 (N_20395,N_19634,N_19945);
or U20396 (N_20396,N_19115,N_19379);
xor U20397 (N_20397,N_19980,N_19882);
or U20398 (N_20398,N_19547,N_19553);
xnor U20399 (N_20399,N_19567,N_19087);
or U20400 (N_20400,N_19797,N_19007);
nand U20401 (N_20401,N_19392,N_19312);
or U20402 (N_20402,N_19221,N_19029);
or U20403 (N_20403,N_19280,N_19006);
xor U20404 (N_20404,N_19273,N_19077);
nor U20405 (N_20405,N_19415,N_19986);
xnor U20406 (N_20406,N_19995,N_19455);
and U20407 (N_20407,N_19263,N_19355);
and U20408 (N_20408,N_19405,N_19675);
xnor U20409 (N_20409,N_19410,N_19662);
and U20410 (N_20410,N_19271,N_19086);
nor U20411 (N_20411,N_19667,N_19481);
and U20412 (N_20412,N_19802,N_19610);
nand U20413 (N_20413,N_19617,N_19862);
nor U20414 (N_20414,N_19454,N_19196);
or U20415 (N_20415,N_19107,N_19304);
xnor U20416 (N_20416,N_19076,N_19705);
nand U20417 (N_20417,N_19516,N_19622);
and U20418 (N_20418,N_19685,N_19928);
xnor U20419 (N_20419,N_19104,N_19804);
nor U20420 (N_20420,N_19057,N_19810);
nor U20421 (N_20421,N_19045,N_19766);
nor U20422 (N_20422,N_19592,N_19887);
nand U20423 (N_20423,N_19119,N_19790);
nand U20424 (N_20424,N_19486,N_19024);
nand U20425 (N_20425,N_19014,N_19272);
nand U20426 (N_20426,N_19594,N_19005);
or U20427 (N_20427,N_19756,N_19744);
nor U20428 (N_20428,N_19267,N_19261);
nand U20429 (N_20429,N_19416,N_19251);
nand U20430 (N_20430,N_19242,N_19053);
xor U20431 (N_20431,N_19329,N_19741);
nor U20432 (N_20432,N_19688,N_19408);
or U20433 (N_20433,N_19378,N_19531);
nor U20434 (N_20434,N_19164,N_19899);
nor U20435 (N_20435,N_19137,N_19581);
or U20436 (N_20436,N_19417,N_19673);
nor U20437 (N_20437,N_19979,N_19294);
xnor U20438 (N_20438,N_19773,N_19715);
nor U20439 (N_20439,N_19578,N_19099);
nand U20440 (N_20440,N_19001,N_19395);
nand U20441 (N_20441,N_19031,N_19574);
nand U20442 (N_20442,N_19507,N_19019);
xor U20443 (N_20443,N_19192,N_19338);
nor U20444 (N_20444,N_19540,N_19968);
nor U20445 (N_20445,N_19942,N_19428);
or U20446 (N_20446,N_19943,N_19740);
and U20447 (N_20447,N_19193,N_19905);
xnor U20448 (N_20448,N_19318,N_19615);
xnor U20449 (N_20449,N_19380,N_19951);
and U20450 (N_20450,N_19245,N_19904);
nor U20451 (N_20451,N_19427,N_19752);
xor U20452 (N_20452,N_19357,N_19333);
nand U20453 (N_20453,N_19237,N_19523);
nor U20454 (N_20454,N_19204,N_19016);
xnor U20455 (N_20455,N_19635,N_19135);
xnor U20456 (N_20456,N_19171,N_19731);
and U20457 (N_20457,N_19443,N_19577);
xor U20458 (N_20458,N_19142,N_19201);
or U20459 (N_20459,N_19575,N_19502);
nor U20460 (N_20460,N_19402,N_19985);
and U20461 (N_20461,N_19385,N_19873);
nor U20462 (N_20462,N_19034,N_19825);
and U20463 (N_20463,N_19125,N_19698);
nand U20464 (N_20464,N_19129,N_19713);
nand U20465 (N_20465,N_19352,N_19974);
nor U20466 (N_20466,N_19013,N_19560);
nand U20467 (N_20467,N_19655,N_19972);
nor U20468 (N_20468,N_19060,N_19514);
or U20469 (N_20469,N_19923,N_19367);
or U20470 (N_20470,N_19317,N_19714);
xor U20471 (N_20471,N_19697,N_19836);
xnor U20472 (N_20472,N_19589,N_19310);
nor U20473 (N_20473,N_19035,N_19015);
and U20474 (N_20474,N_19768,N_19962);
xor U20475 (N_20475,N_19463,N_19641);
nand U20476 (N_20476,N_19335,N_19260);
nand U20477 (N_20477,N_19588,N_19778);
or U20478 (N_20478,N_19464,N_19618);
or U20479 (N_20479,N_19319,N_19297);
and U20480 (N_20480,N_19993,N_19631);
xor U20481 (N_20481,N_19452,N_19544);
nor U20482 (N_20482,N_19253,N_19911);
nand U20483 (N_20483,N_19892,N_19783);
nand U20484 (N_20484,N_19551,N_19173);
xor U20485 (N_20485,N_19866,N_19749);
and U20486 (N_20486,N_19397,N_19670);
xnor U20487 (N_20487,N_19437,N_19932);
nor U20488 (N_20488,N_19157,N_19571);
nor U20489 (N_20489,N_19948,N_19957);
and U20490 (N_20490,N_19473,N_19742);
nand U20491 (N_20491,N_19170,N_19056);
xor U20492 (N_20492,N_19759,N_19632);
nand U20493 (N_20493,N_19438,N_19969);
nand U20494 (N_20494,N_19765,N_19359);
nor U20495 (N_20495,N_19689,N_19846);
nor U20496 (N_20496,N_19160,N_19131);
and U20497 (N_20497,N_19919,N_19861);
or U20498 (N_20498,N_19912,N_19219);
nand U20499 (N_20499,N_19038,N_19808);
or U20500 (N_20500,N_19058,N_19137);
xnor U20501 (N_20501,N_19471,N_19972);
xnor U20502 (N_20502,N_19289,N_19486);
nor U20503 (N_20503,N_19163,N_19730);
nor U20504 (N_20504,N_19885,N_19029);
nor U20505 (N_20505,N_19749,N_19058);
and U20506 (N_20506,N_19683,N_19259);
nand U20507 (N_20507,N_19551,N_19736);
or U20508 (N_20508,N_19506,N_19648);
xor U20509 (N_20509,N_19549,N_19987);
nand U20510 (N_20510,N_19524,N_19771);
xnor U20511 (N_20511,N_19714,N_19773);
and U20512 (N_20512,N_19869,N_19498);
or U20513 (N_20513,N_19833,N_19918);
or U20514 (N_20514,N_19512,N_19564);
and U20515 (N_20515,N_19033,N_19493);
or U20516 (N_20516,N_19674,N_19350);
nor U20517 (N_20517,N_19302,N_19898);
nand U20518 (N_20518,N_19534,N_19997);
xor U20519 (N_20519,N_19217,N_19150);
and U20520 (N_20520,N_19208,N_19110);
and U20521 (N_20521,N_19259,N_19171);
nor U20522 (N_20522,N_19631,N_19332);
xnor U20523 (N_20523,N_19969,N_19571);
nor U20524 (N_20524,N_19183,N_19695);
and U20525 (N_20525,N_19083,N_19097);
nand U20526 (N_20526,N_19636,N_19087);
xnor U20527 (N_20527,N_19099,N_19335);
or U20528 (N_20528,N_19085,N_19839);
nor U20529 (N_20529,N_19498,N_19201);
or U20530 (N_20530,N_19776,N_19418);
and U20531 (N_20531,N_19962,N_19463);
nor U20532 (N_20532,N_19391,N_19649);
and U20533 (N_20533,N_19226,N_19013);
xnor U20534 (N_20534,N_19760,N_19521);
nor U20535 (N_20535,N_19874,N_19602);
or U20536 (N_20536,N_19314,N_19355);
nor U20537 (N_20537,N_19794,N_19652);
or U20538 (N_20538,N_19935,N_19181);
or U20539 (N_20539,N_19557,N_19374);
nand U20540 (N_20540,N_19346,N_19688);
or U20541 (N_20541,N_19434,N_19921);
nand U20542 (N_20542,N_19923,N_19932);
nor U20543 (N_20543,N_19175,N_19936);
nand U20544 (N_20544,N_19021,N_19343);
nor U20545 (N_20545,N_19707,N_19556);
nand U20546 (N_20546,N_19184,N_19728);
and U20547 (N_20547,N_19966,N_19411);
xnor U20548 (N_20548,N_19731,N_19636);
and U20549 (N_20549,N_19236,N_19171);
and U20550 (N_20550,N_19137,N_19355);
xor U20551 (N_20551,N_19362,N_19414);
nor U20552 (N_20552,N_19471,N_19505);
nor U20553 (N_20553,N_19945,N_19661);
nor U20554 (N_20554,N_19428,N_19769);
and U20555 (N_20555,N_19977,N_19812);
and U20556 (N_20556,N_19582,N_19845);
xor U20557 (N_20557,N_19345,N_19393);
nor U20558 (N_20558,N_19026,N_19413);
xor U20559 (N_20559,N_19991,N_19879);
or U20560 (N_20560,N_19401,N_19483);
xnor U20561 (N_20561,N_19751,N_19551);
nor U20562 (N_20562,N_19644,N_19225);
nand U20563 (N_20563,N_19067,N_19119);
and U20564 (N_20564,N_19232,N_19722);
or U20565 (N_20565,N_19500,N_19755);
nand U20566 (N_20566,N_19362,N_19388);
and U20567 (N_20567,N_19145,N_19155);
xor U20568 (N_20568,N_19646,N_19653);
nor U20569 (N_20569,N_19966,N_19583);
or U20570 (N_20570,N_19856,N_19808);
xor U20571 (N_20571,N_19034,N_19757);
nor U20572 (N_20572,N_19677,N_19657);
nand U20573 (N_20573,N_19056,N_19611);
and U20574 (N_20574,N_19444,N_19950);
nor U20575 (N_20575,N_19077,N_19184);
nand U20576 (N_20576,N_19817,N_19259);
nor U20577 (N_20577,N_19817,N_19679);
or U20578 (N_20578,N_19488,N_19941);
or U20579 (N_20579,N_19068,N_19098);
or U20580 (N_20580,N_19349,N_19046);
nor U20581 (N_20581,N_19170,N_19828);
or U20582 (N_20582,N_19807,N_19716);
xnor U20583 (N_20583,N_19282,N_19658);
and U20584 (N_20584,N_19641,N_19605);
nor U20585 (N_20585,N_19660,N_19423);
xnor U20586 (N_20586,N_19999,N_19642);
nand U20587 (N_20587,N_19050,N_19190);
nand U20588 (N_20588,N_19241,N_19720);
xor U20589 (N_20589,N_19378,N_19567);
nand U20590 (N_20590,N_19166,N_19199);
nor U20591 (N_20591,N_19473,N_19874);
and U20592 (N_20592,N_19547,N_19911);
nor U20593 (N_20593,N_19953,N_19603);
and U20594 (N_20594,N_19918,N_19819);
nand U20595 (N_20595,N_19270,N_19680);
nand U20596 (N_20596,N_19594,N_19068);
nor U20597 (N_20597,N_19125,N_19975);
xnor U20598 (N_20598,N_19903,N_19858);
and U20599 (N_20599,N_19203,N_19876);
nand U20600 (N_20600,N_19109,N_19897);
xor U20601 (N_20601,N_19541,N_19516);
nor U20602 (N_20602,N_19410,N_19599);
xor U20603 (N_20603,N_19348,N_19085);
or U20604 (N_20604,N_19706,N_19962);
nor U20605 (N_20605,N_19117,N_19345);
and U20606 (N_20606,N_19803,N_19381);
nand U20607 (N_20607,N_19197,N_19239);
nand U20608 (N_20608,N_19338,N_19178);
nand U20609 (N_20609,N_19018,N_19608);
or U20610 (N_20610,N_19270,N_19152);
nor U20611 (N_20611,N_19034,N_19911);
and U20612 (N_20612,N_19125,N_19697);
and U20613 (N_20613,N_19367,N_19668);
nand U20614 (N_20614,N_19248,N_19868);
nor U20615 (N_20615,N_19703,N_19309);
or U20616 (N_20616,N_19203,N_19801);
nor U20617 (N_20617,N_19438,N_19626);
or U20618 (N_20618,N_19221,N_19060);
xor U20619 (N_20619,N_19013,N_19850);
nand U20620 (N_20620,N_19991,N_19029);
nand U20621 (N_20621,N_19672,N_19199);
nor U20622 (N_20622,N_19586,N_19852);
or U20623 (N_20623,N_19155,N_19313);
and U20624 (N_20624,N_19560,N_19223);
xnor U20625 (N_20625,N_19413,N_19586);
nand U20626 (N_20626,N_19903,N_19006);
nor U20627 (N_20627,N_19764,N_19388);
nor U20628 (N_20628,N_19860,N_19548);
xnor U20629 (N_20629,N_19515,N_19277);
nand U20630 (N_20630,N_19960,N_19545);
xor U20631 (N_20631,N_19328,N_19280);
nor U20632 (N_20632,N_19587,N_19292);
nand U20633 (N_20633,N_19450,N_19543);
nor U20634 (N_20634,N_19053,N_19850);
xnor U20635 (N_20635,N_19057,N_19511);
nand U20636 (N_20636,N_19807,N_19139);
and U20637 (N_20637,N_19897,N_19437);
xor U20638 (N_20638,N_19420,N_19565);
xor U20639 (N_20639,N_19622,N_19055);
nand U20640 (N_20640,N_19662,N_19043);
or U20641 (N_20641,N_19087,N_19277);
xnor U20642 (N_20642,N_19293,N_19795);
and U20643 (N_20643,N_19176,N_19155);
nand U20644 (N_20644,N_19370,N_19333);
nand U20645 (N_20645,N_19347,N_19308);
or U20646 (N_20646,N_19097,N_19667);
or U20647 (N_20647,N_19183,N_19856);
or U20648 (N_20648,N_19205,N_19001);
or U20649 (N_20649,N_19422,N_19879);
xor U20650 (N_20650,N_19308,N_19185);
nand U20651 (N_20651,N_19292,N_19591);
nor U20652 (N_20652,N_19050,N_19338);
or U20653 (N_20653,N_19887,N_19109);
nor U20654 (N_20654,N_19880,N_19193);
and U20655 (N_20655,N_19497,N_19292);
or U20656 (N_20656,N_19336,N_19233);
nand U20657 (N_20657,N_19838,N_19777);
or U20658 (N_20658,N_19525,N_19284);
nand U20659 (N_20659,N_19280,N_19854);
xor U20660 (N_20660,N_19340,N_19472);
xnor U20661 (N_20661,N_19365,N_19999);
nor U20662 (N_20662,N_19487,N_19163);
nand U20663 (N_20663,N_19781,N_19513);
xnor U20664 (N_20664,N_19684,N_19666);
nand U20665 (N_20665,N_19122,N_19840);
nor U20666 (N_20666,N_19752,N_19419);
nand U20667 (N_20667,N_19145,N_19304);
and U20668 (N_20668,N_19018,N_19752);
nand U20669 (N_20669,N_19781,N_19612);
and U20670 (N_20670,N_19076,N_19058);
nor U20671 (N_20671,N_19774,N_19903);
xor U20672 (N_20672,N_19704,N_19024);
xnor U20673 (N_20673,N_19613,N_19921);
nand U20674 (N_20674,N_19720,N_19021);
or U20675 (N_20675,N_19340,N_19213);
or U20676 (N_20676,N_19240,N_19172);
and U20677 (N_20677,N_19679,N_19448);
nand U20678 (N_20678,N_19275,N_19442);
xor U20679 (N_20679,N_19768,N_19639);
nand U20680 (N_20680,N_19661,N_19777);
and U20681 (N_20681,N_19995,N_19891);
and U20682 (N_20682,N_19623,N_19137);
nand U20683 (N_20683,N_19160,N_19999);
or U20684 (N_20684,N_19577,N_19851);
xor U20685 (N_20685,N_19614,N_19871);
and U20686 (N_20686,N_19997,N_19832);
and U20687 (N_20687,N_19841,N_19385);
xor U20688 (N_20688,N_19261,N_19860);
or U20689 (N_20689,N_19025,N_19628);
xnor U20690 (N_20690,N_19390,N_19488);
nand U20691 (N_20691,N_19096,N_19036);
xnor U20692 (N_20692,N_19554,N_19320);
xor U20693 (N_20693,N_19095,N_19776);
nand U20694 (N_20694,N_19978,N_19731);
nand U20695 (N_20695,N_19295,N_19316);
and U20696 (N_20696,N_19238,N_19947);
and U20697 (N_20697,N_19693,N_19914);
nand U20698 (N_20698,N_19534,N_19764);
and U20699 (N_20699,N_19049,N_19471);
and U20700 (N_20700,N_19303,N_19714);
nand U20701 (N_20701,N_19808,N_19869);
or U20702 (N_20702,N_19805,N_19766);
or U20703 (N_20703,N_19517,N_19194);
nand U20704 (N_20704,N_19465,N_19821);
xnor U20705 (N_20705,N_19809,N_19257);
and U20706 (N_20706,N_19538,N_19219);
xor U20707 (N_20707,N_19821,N_19678);
nor U20708 (N_20708,N_19697,N_19492);
or U20709 (N_20709,N_19540,N_19306);
or U20710 (N_20710,N_19311,N_19813);
nor U20711 (N_20711,N_19579,N_19265);
xor U20712 (N_20712,N_19479,N_19973);
nor U20713 (N_20713,N_19046,N_19681);
and U20714 (N_20714,N_19051,N_19977);
nand U20715 (N_20715,N_19173,N_19101);
nand U20716 (N_20716,N_19167,N_19285);
nand U20717 (N_20717,N_19487,N_19859);
and U20718 (N_20718,N_19612,N_19857);
nor U20719 (N_20719,N_19594,N_19868);
xnor U20720 (N_20720,N_19345,N_19161);
xnor U20721 (N_20721,N_19268,N_19758);
nor U20722 (N_20722,N_19788,N_19732);
xor U20723 (N_20723,N_19347,N_19511);
nor U20724 (N_20724,N_19325,N_19669);
or U20725 (N_20725,N_19983,N_19815);
or U20726 (N_20726,N_19014,N_19821);
xor U20727 (N_20727,N_19224,N_19189);
nand U20728 (N_20728,N_19025,N_19305);
nor U20729 (N_20729,N_19843,N_19393);
xor U20730 (N_20730,N_19985,N_19175);
nor U20731 (N_20731,N_19299,N_19870);
and U20732 (N_20732,N_19665,N_19446);
or U20733 (N_20733,N_19506,N_19908);
xnor U20734 (N_20734,N_19826,N_19496);
nor U20735 (N_20735,N_19023,N_19878);
xor U20736 (N_20736,N_19095,N_19257);
xnor U20737 (N_20737,N_19093,N_19745);
nor U20738 (N_20738,N_19861,N_19510);
nor U20739 (N_20739,N_19084,N_19644);
or U20740 (N_20740,N_19663,N_19114);
and U20741 (N_20741,N_19579,N_19596);
nor U20742 (N_20742,N_19640,N_19728);
and U20743 (N_20743,N_19265,N_19248);
xor U20744 (N_20744,N_19814,N_19971);
nor U20745 (N_20745,N_19136,N_19065);
or U20746 (N_20746,N_19640,N_19790);
or U20747 (N_20747,N_19793,N_19374);
nand U20748 (N_20748,N_19918,N_19647);
nand U20749 (N_20749,N_19295,N_19412);
nor U20750 (N_20750,N_19562,N_19700);
xnor U20751 (N_20751,N_19318,N_19516);
or U20752 (N_20752,N_19860,N_19845);
or U20753 (N_20753,N_19224,N_19353);
xor U20754 (N_20754,N_19927,N_19541);
and U20755 (N_20755,N_19597,N_19337);
xor U20756 (N_20756,N_19846,N_19177);
and U20757 (N_20757,N_19065,N_19635);
xor U20758 (N_20758,N_19777,N_19030);
xnor U20759 (N_20759,N_19023,N_19217);
xnor U20760 (N_20760,N_19373,N_19605);
xor U20761 (N_20761,N_19963,N_19946);
or U20762 (N_20762,N_19684,N_19015);
nand U20763 (N_20763,N_19996,N_19518);
xor U20764 (N_20764,N_19497,N_19569);
nor U20765 (N_20765,N_19152,N_19295);
nor U20766 (N_20766,N_19667,N_19850);
and U20767 (N_20767,N_19553,N_19343);
or U20768 (N_20768,N_19868,N_19123);
xor U20769 (N_20769,N_19895,N_19883);
xnor U20770 (N_20770,N_19120,N_19730);
nand U20771 (N_20771,N_19870,N_19814);
nand U20772 (N_20772,N_19275,N_19250);
xnor U20773 (N_20773,N_19878,N_19938);
nor U20774 (N_20774,N_19767,N_19621);
or U20775 (N_20775,N_19453,N_19820);
and U20776 (N_20776,N_19495,N_19695);
nor U20777 (N_20777,N_19075,N_19670);
or U20778 (N_20778,N_19084,N_19690);
xor U20779 (N_20779,N_19045,N_19421);
xor U20780 (N_20780,N_19546,N_19856);
nand U20781 (N_20781,N_19894,N_19554);
or U20782 (N_20782,N_19883,N_19410);
nor U20783 (N_20783,N_19419,N_19428);
and U20784 (N_20784,N_19527,N_19971);
nor U20785 (N_20785,N_19966,N_19581);
nor U20786 (N_20786,N_19377,N_19662);
xor U20787 (N_20787,N_19249,N_19234);
nor U20788 (N_20788,N_19714,N_19981);
nand U20789 (N_20789,N_19937,N_19737);
or U20790 (N_20790,N_19520,N_19080);
nand U20791 (N_20791,N_19548,N_19113);
nor U20792 (N_20792,N_19187,N_19902);
nand U20793 (N_20793,N_19760,N_19680);
xor U20794 (N_20794,N_19792,N_19623);
and U20795 (N_20795,N_19464,N_19815);
and U20796 (N_20796,N_19808,N_19042);
nor U20797 (N_20797,N_19861,N_19936);
xnor U20798 (N_20798,N_19233,N_19117);
xnor U20799 (N_20799,N_19116,N_19843);
or U20800 (N_20800,N_19095,N_19604);
and U20801 (N_20801,N_19465,N_19139);
xor U20802 (N_20802,N_19197,N_19257);
or U20803 (N_20803,N_19918,N_19636);
nand U20804 (N_20804,N_19751,N_19853);
nor U20805 (N_20805,N_19037,N_19745);
nor U20806 (N_20806,N_19316,N_19619);
xnor U20807 (N_20807,N_19993,N_19891);
and U20808 (N_20808,N_19264,N_19349);
xnor U20809 (N_20809,N_19350,N_19475);
nor U20810 (N_20810,N_19291,N_19136);
and U20811 (N_20811,N_19414,N_19019);
nand U20812 (N_20812,N_19141,N_19439);
nand U20813 (N_20813,N_19869,N_19853);
xor U20814 (N_20814,N_19896,N_19328);
or U20815 (N_20815,N_19959,N_19988);
nor U20816 (N_20816,N_19605,N_19011);
or U20817 (N_20817,N_19859,N_19536);
and U20818 (N_20818,N_19793,N_19954);
or U20819 (N_20819,N_19695,N_19769);
and U20820 (N_20820,N_19428,N_19681);
or U20821 (N_20821,N_19946,N_19479);
and U20822 (N_20822,N_19961,N_19831);
or U20823 (N_20823,N_19900,N_19155);
or U20824 (N_20824,N_19226,N_19966);
nor U20825 (N_20825,N_19597,N_19955);
nor U20826 (N_20826,N_19612,N_19333);
nor U20827 (N_20827,N_19072,N_19757);
and U20828 (N_20828,N_19819,N_19908);
nor U20829 (N_20829,N_19090,N_19752);
xor U20830 (N_20830,N_19061,N_19598);
nand U20831 (N_20831,N_19495,N_19287);
nor U20832 (N_20832,N_19269,N_19317);
and U20833 (N_20833,N_19697,N_19721);
nor U20834 (N_20834,N_19363,N_19762);
nor U20835 (N_20835,N_19201,N_19747);
or U20836 (N_20836,N_19977,N_19359);
nor U20837 (N_20837,N_19146,N_19976);
or U20838 (N_20838,N_19931,N_19421);
xnor U20839 (N_20839,N_19443,N_19745);
xnor U20840 (N_20840,N_19396,N_19147);
xor U20841 (N_20841,N_19186,N_19317);
and U20842 (N_20842,N_19387,N_19846);
and U20843 (N_20843,N_19352,N_19042);
or U20844 (N_20844,N_19303,N_19759);
nand U20845 (N_20845,N_19129,N_19634);
nand U20846 (N_20846,N_19918,N_19450);
nand U20847 (N_20847,N_19145,N_19296);
nand U20848 (N_20848,N_19921,N_19167);
nor U20849 (N_20849,N_19849,N_19265);
nand U20850 (N_20850,N_19854,N_19369);
and U20851 (N_20851,N_19200,N_19481);
or U20852 (N_20852,N_19887,N_19253);
xor U20853 (N_20853,N_19624,N_19481);
xnor U20854 (N_20854,N_19264,N_19396);
and U20855 (N_20855,N_19106,N_19818);
or U20856 (N_20856,N_19673,N_19239);
nor U20857 (N_20857,N_19467,N_19011);
and U20858 (N_20858,N_19011,N_19010);
nor U20859 (N_20859,N_19119,N_19116);
nor U20860 (N_20860,N_19626,N_19743);
or U20861 (N_20861,N_19393,N_19483);
xnor U20862 (N_20862,N_19606,N_19061);
xor U20863 (N_20863,N_19259,N_19664);
and U20864 (N_20864,N_19606,N_19558);
or U20865 (N_20865,N_19812,N_19425);
and U20866 (N_20866,N_19739,N_19132);
nand U20867 (N_20867,N_19353,N_19847);
or U20868 (N_20868,N_19853,N_19805);
xor U20869 (N_20869,N_19798,N_19772);
or U20870 (N_20870,N_19627,N_19095);
and U20871 (N_20871,N_19769,N_19017);
nand U20872 (N_20872,N_19206,N_19929);
xor U20873 (N_20873,N_19765,N_19242);
or U20874 (N_20874,N_19502,N_19413);
and U20875 (N_20875,N_19652,N_19644);
nor U20876 (N_20876,N_19070,N_19923);
nand U20877 (N_20877,N_19376,N_19568);
nand U20878 (N_20878,N_19161,N_19666);
or U20879 (N_20879,N_19041,N_19661);
and U20880 (N_20880,N_19624,N_19986);
and U20881 (N_20881,N_19422,N_19271);
xor U20882 (N_20882,N_19467,N_19411);
nor U20883 (N_20883,N_19155,N_19555);
nand U20884 (N_20884,N_19894,N_19165);
and U20885 (N_20885,N_19647,N_19031);
nor U20886 (N_20886,N_19025,N_19045);
and U20887 (N_20887,N_19148,N_19745);
xnor U20888 (N_20888,N_19852,N_19452);
nand U20889 (N_20889,N_19440,N_19235);
xor U20890 (N_20890,N_19650,N_19196);
nor U20891 (N_20891,N_19510,N_19921);
or U20892 (N_20892,N_19538,N_19349);
or U20893 (N_20893,N_19920,N_19650);
nor U20894 (N_20894,N_19172,N_19636);
xnor U20895 (N_20895,N_19369,N_19904);
nand U20896 (N_20896,N_19440,N_19523);
xor U20897 (N_20897,N_19192,N_19705);
nand U20898 (N_20898,N_19857,N_19746);
or U20899 (N_20899,N_19065,N_19903);
or U20900 (N_20900,N_19457,N_19954);
xnor U20901 (N_20901,N_19692,N_19415);
or U20902 (N_20902,N_19917,N_19930);
nor U20903 (N_20903,N_19212,N_19542);
and U20904 (N_20904,N_19682,N_19952);
and U20905 (N_20905,N_19201,N_19959);
nand U20906 (N_20906,N_19740,N_19199);
nor U20907 (N_20907,N_19213,N_19909);
and U20908 (N_20908,N_19472,N_19598);
or U20909 (N_20909,N_19870,N_19836);
and U20910 (N_20910,N_19321,N_19822);
nor U20911 (N_20911,N_19026,N_19799);
nand U20912 (N_20912,N_19586,N_19898);
nor U20913 (N_20913,N_19083,N_19039);
or U20914 (N_20914,N_19764,N_19585);
and U20915 (N_20915,N_19912,N_19854);
xor U20916 (N_20916,N_19911,N_19013);
and U20917 (N_20917,N_19052,N_19967);
or U20918 (N_20918,N_19170,N_19809);
and U20919 (N_20919,N_19419,N_19951);
nor U20920 (N_20920,N_19186,N_19563);
or U20921 (N_20921,N_19850,N_19419);
nor U20922 (N_20922,N_19860,N_19883);
and U20923 (N_20923,N_19258,N_19906);
xnor U20924 (N_20924,N_19127,N_19014);
or U20925 (N_20925,N_19826,N_19217);
xor U20926 (N_20926,N_19472,N_19028);
and U20927 (N_20927,N_19831,N_19232);
xor U20928 (N_20928,N_19134,N_19747);
xor U20929 (N_20929,N_19002,N_19992);
and U20930 (N_20930,N_19700,N_19971);
nor U20931 (N_20931,N_19049,N_19804);
nor U20932 (N_20932,N_19602,N_19196);
and U20933 (N_20933,N_19668,N_19937);
or U20934 (N_20934,N_19383,N_19256);
nand U20935 (N_20935,N_19973,N_19558);
nor U20936 (N_20936,N_19946,N_19884);
nor U20937 (N_20937,N_19820,N_19539);
and U20938 (N_20938,N_19605,N_19636);
nand U20939 (N_20939,N_19471,N_19874);
nor U20940 (N_20940,N_19864,N_19928);
nand U20941 (N_20941,N_19679,N_19513);
or U20942 (N_20942,N_19101,N_19620);
or U20943 (N_20943,N_19763,N_19803);
nor U20944 (N_20944,N_19419,N_19719);
nand U20945 (N_20945,N_19060,N_19084);
nand U20946 (N_20946,N_19692,N_19436);
or U20947 (N_20947,N_19917,N_19238);
and U20948 (N_20948,N_19028,N_19761);
and U20949 (N_20949,N_19279,N_19341);
nand U20950 (N_20950,N_19111,N_19732);
and U20951 (N_20951,N_19215,N_19401);
and U20952 (N_20952,N_19248,N_19129);
and U20953 (N_20953,N_19398,N_19532);
xnor U20954 (N_20954,N_19711,N_19318);
nor U20955 (N_20955,N_19845,N_19708);
or U20956 (N_20956,N_19900,N_19916);
xor U20957 (N_20957,N_19846,N_19005);
and U20958 (N_20958,N_19672,N_19760);
xor U20959 (N_20959,N_19193,N_19422);
and U20960 (N_20960,N_19650,N_19913);
and U20961 (N_20961,N_19847,N_19648);
xor U20962 (N_20962,N_19949,N_19084);
nand U20963 (N_20963,N_19203,N_19057);
and U20964 (N_20964,N_19670,N_19278);
nor U20965 (N_20965,N_19629,N_19172);
xor U20966 (N_20966,N_19150,N_19416);
nand U20967 (N_20967,N_19991,N_19368);
xnor U20968 (N_20968,N_19500,N_19290);
or U20969 (N_20969,N_19863,N_19498);
nor U20970 (N_20970,N_19624,N_19302);
nand U20971 (N_20971,N_19091,N_19134);
nor U20972 (N_20972,N_19209,N_19973);
nand U20973 (N_20973,N_19643,N_19727);
xor U20974 (N_20974,N_19809,N_19261);
and U20975 (N_20975,N_19076,N_19653);
and U20976 (N_20976,N_19030,N_19581);
nand U20977 (N_20977,N_19620,N_19526);
and U20978 (N_20978,N_19004,N_19195);
xor U20979 (N_20979,N_19956,N_19160);
nor U20980 (N_20980,N_19261,N_19426);
xnor U20981 (N_20981,N_19753,N_19783);
nand U20982 (N_20982,N_19546,N_19773);
nand U20983 (N_20983,N_19095,N_19735);
nand U20984 (N_20984,N_19718,N_19770);
or U20985 (N_20985,N_19732,N_19140);
nor U20986 (N_20986,N_19093,N_19168);
nand U20987 (N_20987,N_19205,N_19162);
nor U20988 (N_20988,N_19505,N_19110);
xnor U20989 (N_20989,N_19498,N_19455);
xor U20990 (N_20990,N_19685,N_19518);
and U20991 (N_20991,N_19985,N_19118);
xnor U20992 (N_20992,N_19902,N_19085);
nor U20993 (N_20993,N_19626,N_19270);
and U20994 (N_20994,N_19879,N_19082);
and U20995 (N_20995,N_19498,N_19846);
xnor U20996 (N_20996,N_19041,N_19141);
xor U20997 (N_20997,N_19319,N_19541);
xor U20998 (N_20998,N_19433,N_19502);
nand U20999 (N_20999,N_19644,N_19412);
nor U21000 (N_21000,N_20574,N_20468);
xor U21001 (N_21001,N_20753,N_20684);
and U21002 (N_21002,N_20436,N_20718);
nor U21003 (N_21003,N_20785,N_20817);
nor U21004 (N_21004,N_20671,N_20627);
or U21005 (N_21005,N_20114,N_20913);
nor U21006 (N_21006,N_20085,N_20779);
nor U21007 (N_21007,N_20935,N_20927);
and U21008 (N_21008,N_20771,N_20775);
nor U21009 (N_21009,N_20491,N_20189);
nor U21010 (N_21010,N_20645,N_20009);
nand U21011 (N_21011,N_20383,N_20682);
nand U21012 (N_21012,N_20283,N_20668);
nand U21013 (N_21013,N_20346,N_20267);
nand U21014 (N_21014,N_20939,N_20005);
or U21015 (N_21015,N_20665,N_20494);
xor U21016 (N_21016,N_20868,N_20632);
nand U21017 (N_21017,N_20359,N_20679);
or U21018 (N_21018,N_20381,N_20479);
xnor U21019 (N_21019,N_20783,N_20770);
nand U21020 (N_21020,N_20577,N_20920);
nand U21021 (N_21021,N_20037,N_20907);
nor U21022 (N_21022,N_20051,N_20995);
or U21023 (N_21023,N_20303,N_20235);
or U21024 (N_21024,N_20476,N_20286);
and U21025 (N_21025,N_20227,N_20421);
and U21026 (N_21026,N_20874,N_20678);
nor U21027 (N_21027,N_20312,N_20879);
or U21028 (N_21028,N_20640,N_20334);
and U21029 (N_21029,N_20357,N_20048);
and U21030 (N_21030,N_20274,N_20571);
or U21031 (N_21031,N_20113,N_20837);
nand U21032 (N_21032,N_20564,N_20495);
xnor U21033 (N_21033,N_20273,N_20938);
and U21034 (N_21034,N_20466,N_20960);
nand U21035 (N_21035,N_20097,N_20290);
nand U21036 (N_21036,N_20028,N_20991);
or U21037 (N_21037,N_20954,N_20689);
xor U21038 (N_21038,N_20726,N_20573);
nand U21039 (N_21039,N_20777,N_20500);
or U21040 (N_21040,N_20095,N_20597);
xnor U21041 (N_21041,N_20003,N_20801);
or U21042 (N_21042,N_20860,N_20845);
and U21043 (N_21043,N_20498,N_20743);
and U21044 (N_21044,N_20736,N_20833);
or U21045 (N_21045,N_20876,N_20630);
or U21046 (N_21046,N_20971,N_20952);
and U21047 (N_21047,N_20281,N_20546);
and U21048 (N_21048,N_20559,N_20297);
or U21049 (N_21049,N_20167,N_20490);
nor U21050 (N_21050,N_20258,N_20078);
and U21051 (N_21051,N_20412,N_20629);
and U21052 (N_21052,N_20467,N_20892);
xnor U21053 (N_21053,N_20165,N_20716);
xnor U21054 (N_21054,N_20996,N_20989);
nor U21055 (N_21055,N_20536,N_20272);
xnor U21056 (N_21056,N_20463,N_20317);
nand U21057 (N_21057,N_20262,N_20007);
nand U21058 (N_21058,N_20976,N_20061);
or U21059 (N_21059,N_20932,N_20634);
nor U21060 (N_21060,N_20812,N_20737);
or U21061 (N_21061,N_20740,N_20619);
nor U21062 (N_21062,N_20606,N_20620);
nor U21063 (N_21063,N_20150,N_20511);
and U21064 (N_21064,N_20374,N_20806);
and U21065 (N_21065,N_20683,N_20425);
nor U21066 (N_21066,N_20761,N_20756);
and U21067 (N_21067,N_20553,N_20196);
xnor U21068 (N_21068,N_20045,N_20228);
xor U21069 (N_21069,N_20291,N_20377);
nor U21070 (N_21070,N_20465,N_20276);
and U21071 (N_21071,N_20242,N_20790);
xnor U21072 (N_21072,N_20446,N_20527);
xor U21073 (N_21073,N_20888,N_20687);
nand U21074 (N_21074,N_20323,N_20504);
nor U21075 (N_21075,N_20526,N_20305);
nor U21076 (N_21076,N_20147,N_20613);
nand U21077 (N_21077,N_20881,N_20247);
or U21078 (N_21078,N_20271,N_20847);
xnor U21079 (N_21079,N_20125,N_20951);
xor U21080 (N_21080,N_20062,N_20379);
or U21081 (N_21081,N_20793,N_20131);
xnor U21082 (N_21082,N_20535,N_20561);
nor U21083 (N_21083,N_20731,N_20044);
nand U21084 (N_21084,N_20266,N_20730);
xnor U21085 (N_21085,N_20609,N_20117);
nor U21086 (N_21086,N_20575,N_20795);
or U21087 (N_21087,N_20369,N_20441);
nand U21088 (N_21088,N_20120,N_20586);
nand U21089 (N_21089,N_20341,N_20473);
xnor U21090 (N_21090,N_20414,N_20366);
and U21091 (N_21091,N_20254,N_20400);
xor U21092 (N_21092,N_20340,N_20893);
or U21093 (N_21093,N_20764,N_20091);
or U21094 (N_21094,N_20694,N_20532);
or U21095 (N_21095,N_20842,N_20349);
nand U21096 (N_21096,N_20862,N_20914);
nand U21097 (N_21097,N_20520,N_20175);
and U21098 (N_21098,N_20019,N_20799);
or U21099 (N_21099,N_20543,N_20864);
and U21100 (N_21100,N_20411,N_20533);
xnor U21101 (N_21101,N_20452,N_20127);
xnor U21102 (N_21102,N_20475,N_20481);
or U21103 (N_21103,N_20234,N_20884);
and U21104 (N_21104,N_20000,N_20675);
nor U21105 (N_21105,N_20655,N_20299);
nand U21106 (N_21106,N_20767,N_20482);
and U21107 (N_21107,N_20887,N_20439);
nand U21108 (N_21108,N_20081,N_20517);
or U21109 (N_21109,N_20278,N_20741);
xor U21110 (N_21110,N_20250,N_20398);
nand U21111 (N_21111,N_20318,N_20314);
or U21112 (N_21112,N_20157,N_20622);
nand U21113 (N_21113,N_20820,N_20941);
or U21114 (N_21114,N_20572,N_20408);
or U21115 (N_21115,N_20394,N_20814);
nand U21116 (N_21116,N_20100,N_20763);
and U21117 (N_21117,N_20469,N_20972);
or U21118 (N_21118,N_20263,N_20382);
xor U21119 (N_21119,N_20174,N_20852);
and U21120 (N_21120,N_20502,N_20364);
xor U21121 (N_21121,N_20988,N_20871);
nor U21122 (N_21122,N_20851,N_20449);
or U21123 (N_21123,N_20395,N_20990);
nor U21124 (N_21124,N_20738,N_20337);
xor U21125 (N_21125,N_20187,N_20946);
nor U21126 (N_21126,N_20919,N_20107);
or U21127 (N_21127,N_20173,N_20257);
or U21128 (N_21128,N_20092,N_20068);
or U21129 (N_21129,N_20245,N_20221);
or U21130 (N_21130,N_20739,N_20531);
or U21131 (N_21131,N_20385,N_20794);
xnor U21132 (N_21132,N_20184,N_20183);
xnor U21133 (N_21133,N_20405,N_20908);
nand U21134 (N_21134,N_20797,N_20215);
and U21135 (N_21135,N_20309,N_20455);
nor U21136 (N_21136,N_20616,N_20637);
xnor U21137 (N_21137,N_20453,N_20603);
xor U21138 (N_21138,N_20706,N_20894);
or U21139 (N_21139,N_20652,N_20590);
nand U21140 (N_21140,N_20975,N_20877);
or U21141 (N_21141,N_20474,N_20136);
nor U21142 (N_21142,N_20096,N_20524);
or U21143 (N_21143,N_20765,N_20461);
nand U21144 (N_21144,N_20389,N_20159);
nor U21145 (N_21145,N_20372,N_20327);
nand U21146 (N_21146,N_20470,N_20168);
xor U21147 (N_21147,N_20179,N_20973);
or U21148 (N_21148,N_20080,N_20534);
or U21149 (N_21149,N_20295,N_20004);
or U21150 (N_21150,N_20859,N_20966);
and U21151 (N_21151,N_20611,N_20647);
and U21152 (N_21152,N_20713,N_20734);
nand U21153 (N_21153,N_20224,N_20930);
or U21154 (N_21154,N_20945,N_20031);
nor U21155 (N_21155,N_20231,N_20241);
nor U21156 (N_21156,N_20915,N_20302);
nand U21157 (N_21157,N_20614,N_20135);
and U21158 (N_21158,N_20202,N_20899);
nand U21159 (N_21159,N_20707,N_20280);
xnor U21160 (N_21160,N_20448,N_20958);
and U21161 (N_21161,N_20831,N_20545);
nand U21162 (N_21162,N_20692,N_20288);
nor U21163 (N_21163,N_20926,N_20784);
nand U21164 (N_21164,N_20685,N_20270);
nor U21165 (N_21165,N_20501,N_20163);
and U21166 (N_21166,N_20145,N_20844);
nor U21167 (N_21167,N_20041,N_20677);
nand U21168 (N_21168,N_20156,N_20458);
nor U21169 (N_21169,N_20275,N_20013);
or U21170 (N_21170,N_20848,N_20496);
and U21171 (N_21171,N_20083,N_20001);
nand U21172 (N_21172,N_20759,N_20178);
nand U21173 (N_21173,N_20804,N_20699);
nor U21174 (N_21174,N_20982,N_20076);
nor U21175 (N_21175,N_20787,N_20418);
nor U21176 (N_21176,N_20898,N_20865);
nor U21177 (N_21177,N_20070,N_20343);
and U21178 (N_21178,N_20355,N_20508);
nor U21179 (N_21179,N_20977,N_20830);
xor U21180 (N_21180,N_20646,N_20727);
nand U21181 (N_21181,N_20615,N_20253);
xor U21182 (N_21182,N_20043,N_20774);
or U21183 (N_21183,N_20199,N_20803);
nand U21184 (N_21184,N_20955,N_20672);
xor U21185 (N_21185,N_20378,N_20654);
or U21186 (N_21186,N_20153,N_20399);
nand U21187 (N_21187,N_20503,N_20230);
nor U21188 (N_21188,N_20506,N_20049);
nor U21189 (N_21189,N_20151,N_20356);
nor U21190 (N_21190,N_20717,N_20375);
or U21191 (N_21191,N_20025,N_20653);
xor U21192 (N_21192,N_20827,N_20593);
nor U21193 (N_21193,N_20850,N_20633);
nor U21194 (N_21194,N_20657,N_20811);
nor U21195 (N_21195,N_20697,N_20431);
and U21196 (N_21196,N_20360,N_20021);
nand U21197 (N_21197,N_20891,N_20659);
nor U21198 (N_21198,N_20180,N_20370);
xnor U21199 (N_21199,N_20758,N_20434);
nor U21200 (N_21200,N_20711,N_20390);
nor U21201 (N_21201,N_20846,N_20686);
or U21202 (N_21202,N_20244,N_20749);
nand U21203 (N_21203,N_20587,N_20639);
nand U21204 (N_21204,N_20208,N_20248);
or U21205 (N_21205,N_20649,N_20006);
xor U21206 (N_21206,N_20552,N_20942);
or U21207 (N_21207,N_20791,N_20723);
and U21208 (N_21208,N_20433,N_20435);
nand U21209 (N_21209,N_20834,N_20485);
or U21210 (N_21210,N_20229,N_20195);
and U21211 (N_21211,N_20828,N_20002);
nand U21212 (N_21212,N_20052,N_20072);
nor U21213 (N_21213,N_20064,N_20424);
xnor U21214 (N_21214,N_20936,N_20030);
nor U21215 (N_21215,N_20073,N_20821);
xor U21216 (N_21216,N_20621,N_20916);
or U21217 (N_21217,N_20591,N_20556);
nand U21218 (N_21218,N_20917,N_20602);
nand U21219 (N_21219,N_20413,N_20011);
and U21220 (N_21220,N_20345,N_20330);
nor U21221 (N_21221,N_20328,N_20889);
nand U21222 (N_21222,N_20154,N_20038);
nand U21223 (N_21223,N_20443,N_20292);
and U21224 (N_21224,N_20137,N_20688);
or U21225 (N_21225,N_20704,N_20437);
nor U21226 (N_21226,N_20745,N_20093);
or U21227 (N_21227,N_20724,N_20998);
or U21228 (N_21228,N_20403,N_20957);
nand U21229 (N_21229,N_20315,N_20537);
xor U21230 (N_21230,N_20406,N_20896);
nand U21231 (N_21231,N_20836,N_20992);
nand U21232 (N_21232,N_20222,N_20947);
nor U21233 (N_21233,N_20800,N_20963);
or U21234 (N_21234,N_20223,N_20454);
nand U21235 (N_21235,N_20444,N_20752);
and U21236 (N_21236,N_20805,N_20900);
or U21237 (N_21237,N_20773,N_20829);
nand U21238 (N_21238,N_20319,N_20768);
and U21239 (N_21239,N_20909,N_20562);
or U21240 (N_21240,N_20046,N_20970);
and U21241 (N_21241,N_20595,N_20226);
xnor U21242 (N_21242,N_20933,N_20931);
and U21243 (N_21243,N_20256,N_20557);
xnor U21244 (N_21244,N_20259,N_20792);
nor U21245 (N_21245,N_20772,N_20509);
and U21246 (N_21246,N_20348,N_20339);
and U21247 (N_21247,N_20024,N_20538);
or U21248 (N_21248,N_20185,N_20442);
nor U21249 (N_21249,N_20279,N_20306);
or U21250 (N_21250,N_20522,N_20246);
or U21251 (N_21251,N_20880,N_20873);
nor U21252 (N_21252,N_20922,N_20505);
or U21253 (N_21253,N_20565,N_20566);
and U21254 (N_21254,N_20144,N_20911);
xor U21255 (N_21255,N_20802,N_20514);
xor U21256 (N_21256,N_20423,N_20525);
xnor U21257 (N_21257,N_20486,N_20077);
and U21258 (N_21258,N_20287,N_20832);
or U21259 (N_21259,N_20580,N_20440);
nor U21260 (N_21260,N_20929,N_20132);
or U21261 (N_21261,N_20895,N_20060);
nand U21262 (N_21262,N_20487,N_20255);
xnor U21263 (N_21263,N_20499,N_20693);
and U21264 (N_21264,N_20656,N_20109);
nor U21265 (N_21265,N_20182,N_20549);
nand U21266 (N_21266,N_20705,N_20404);
or U21267 (N_21267,N_20981,N_20944);
nor U21268 (N_21268,N_20643,N_20294);
and U21269 (N_21269,N_20581,N_20548);
xor U21270 (N_21270,N_20218,N_20325);
nor U21271 (N_21271,N_20519,N_20710);
nor U21272 (N_21272,N_20883,N_20747);
or U21273 (N_21273,N_20042,N_20979);
and U21274 (N_21274,N_20260,N_20497);
xor U21275 (N_21275,N_20225,N_20798);
xnor U21276 (N_21276,N_20123,N_20725);
nand U21277 (N_21277,N_20600,N_20240);
and U21278 (N_21278,N_20233,N_20329);
or U21279 (N_21279,N_20171,N_20540);
nor U21280 (N_21280,N_20464,N_20776);
xnor U21281 (N_21281,N_20358,N_20035);
and U21282 (N_21282,N_20569,N_20816);
and U21283 (N_21283,N_20069,N_20075);
xnor U21284 (N_21284,N_20650,N_20815);
or U21285 (N_21285,N_20192,N_20807);
and U21286 (N_21286,N_20601,N_20698);
xor U21287 (N_21287,N_20211,N_20017);
or U21288 (N_21288,N_20190,N_20863);
nor U21289 (N_21289,N_20612,N_20158);
nand U21290 (N_21290,N_20376,N_20387);
nand U21291 (N_21291,N_20198,N_20438);
nand U21292 (N_21292,N_20869,N_20786);
nand U21293 (N_21293,N_20948,N_20489);
or U21294 (N_21294,N_20719,N_20363);
nand U21295 (N_21295,N_20102,N_20885);
nand U21296 (N_21296,N_20338,N_20585);
xor U21297 (N_21297,N_20362,N_20188);
nand U21298 (N_21298,N_20265,N_20427);
or U21299 (N_21299,N_20149,N_20380);
nor U21300 (N_21300,N_20478,N_20809);
nor U21301 (N_21301,N_20721,N_20285);
nor U21302 (N_21302,N_20371,N_20928);
xor U21303 (N_21303,N_20401,N_20307);
or U21304 (N_21304,N_20744,N_20417);
xor U21305 (N_21305,N_20304,N_20121);
nor U21306 (N_21306,N_20084,N_20420);
or U21307 (N_21307,N_20690,N_20351);
or U21308 (N_21308,N_20116,N_20714);
and U21309 (N_21309,N_20943,N_20782);
nor U21310 (N_21310,N_20604,N_20742);
nor U21311 (N_21311,N_20623,N_20735);
and U21312 (N_21312,N_20071,N_20778);
or U21313 (N_21313,N_20617,N_20209);
nor U21314 (N_21314,N_20596,N_20762);
or U21315 (N_21315,N_20220,N_20967);
xnor U21316 (N_21316,N_20289,N_20959);
or U21317 (N_21317,N_20901,N_20961);
nor U21318 (N_21318,N_20513,N_20493);
and U21319 (N_21319,N_20923,N_20956);
xnor U21320 (N_21320,N_20708,N_20906);
nor U21321 (N_21321,N_20875,N_20904);
and U21322 (N_21322,N_20217,N_20176);
or U21323 (N_21323,N_20039,N_20119);
xor U21324 (N_21324,N_20104,N_20822);
xor U21325 (N_21325,N_20203,N_20086);
nand U21326 (N_21326,N_20133,N_20243);
nand U21327 (N_21327,N_20521,N_20890);
or U21328 (N_21328,N_20261,N_20870);
and U21329 (N_21329,N_20746,N_20997);
nand U21330 (N_21330,N_20018,N_20722);
nor U21331 (N_21331,N_20264,N_20141);
and U21332 (N_21332,N_20635,N_20676);
nand U21333 (N_21333,N_20662,N_20201);
or U21334 (N_21334,N_20016,N_20388);
and U21335 (N_21335,N_20701,N_20523);
and U21336 (N_21336,N_20249,N_20316);
nor U21337 (N_21337,N_20214,N_20098);
nor U21338 (N_21338,N_20397,N_20079);
or U21339 (N_21339,N_20516,N_20978);
nand U21340 (N_21340,N_20094,N_20840);
or U21341 (N_21341,N_20206,N_20130);
xor U21342 (N_21342,N_20352,N_20402);
and U21343 (N_21343,N_20667,N_20560);
xnor U21344 (N_21344,N_20968,N_20172);
nand U21345 (N_21345,N_20047,N_20036);
nor U21346 (N_21346,N_20232,N_20422);
nand U21347 (N_21347,N_20849,N_20651);
and U21348 (N_21348,N_20607,N_20570);
xor U21349 (N_21349,N_20530,N_20631);
xor U21350 (N_21350,N_20313,N_20056);
or U21351 (N_21351,N_20712,N_20866);
nor U21352 (N_21352,N_20155,N_20905);
xnor U21353 (N_21353,N_20128,N_20965);
or U21354 (N_21354,N_20057,N_20354);
xor U21355 (N_21355,N_20641,N_20451);
nor U21356 (N_21356,N_20709,N_20568);
and U21357 (N_21357,N_20660,N_20599);
and U21358 (N_21358,N_20949,N_20027);
or U21359 (N_21359,N_20324,N_20861);
xor U21360 (N_21360,N_20818,N_20367);
or U21361 (N_21361,N_20124,N_20022);
and U21362 (N_21362,N_20111,N_20148);
nand U21363 (N_21363,N_20554,N_20937);
xor U21364 (N_21364,N_20555,N_20810);
or U21365 (N_21365,N_20396,N_20194);
and U21366 (N_21366,N_20558,N_20789);
xnor U21367 (N_21367,N_20510,N_20483);
nor U21368 (N_21368,N_20980,N_20728);
nand U21369 (N_21369,N_20129,N_20541);
nor U21370 (N_21370,N_20472,N_20213);
or U21371 (N_21371,N_20122,N_20673);
nor U21372 (N_21372,N_20715,N_20032);
xor U21373 (N_21373,N_20074,N_20432);
or U21374 (N_21374,N_20426,N_20445);
and U21375 (N_21375,N_20336,N_20702);
nand U21376 (N_21376,N_20430,N_20142);
and U21377 (N_21377,N_20012,N_20428);
nor U21378 (N_21378,N_20311,N_20824);
nand U21379 (N_21379,N_20664,N_20015);
xor U21380 (N_21380,N_20087,N_20321);
and U21381 (N_21381,N_20029,N_20628);
nor U21382 (N_21382,N_20589,N_20384);
nor U21383 (N_21383,N_20732,N_20034);
or U21384 (N_21384,N_20191,N_20115);
xor U21385 (N_21385,N_20393,N_20924);
nor U21386 (N_21386,N_20769,N_20103);
nor U21387 (N_21387,N_20626,N_20813);
nor U21388 (N_21388,N_20386,N_20666);
nand U21389 (N_21389,N_20164,N_20331);
nand U21390 (N_21390,N_20088,N_20878);
or U21391 (N_21391,N_20670,N_20471);
or U21392 (N_21392,N_20644,N_20999);
and U21393 (N_21393,N_20964,N_20539);
nor U21394 (N_21394,N_20216,N_20910);
or U21395 (N_21395,N_20040,N_20326);
or U21396 (N_21396,N_20618,N_20583);
xnor U21397 (N_21397,N_20344,N_20720);
and U21398 (N_21398,N_20477,N_20450);
nor U21399 (N_21399,N_20166,N_20853);
nor U21400 (N_21400,N_20669,N_20757);
xnor U21401 (N_21401,N_20239,N_20320);
nand U21402 (N_21402,N_20480,N_20053);
or U21403 (N_21403,N_20542,N_20409);
or U21404 (N_21404,N_20985,N_20841);
nor U21405 (N_21405,N_20204,N_20161);
xor U21406 (N_21406,N_20118,N_20925);
xor U21407 (N_21407,N_20605,N_20680);
nor U21408 (N_21408,N_20026,N_20282);
nor U21409 (N_21409,N_20563,N_20050);
and U21410 (N_21410,N_20950,N_20912);
nand U21411 (N_21411,N_20181,N_20090);
nand U21412 (N_21412,N_20391,N_20236);
and U21413 (N_21413,N_20143,N_20365);
nand U21414 (N_21414,N_20856,N_20588);
nor U21415 (N_21415,N_20733,N_20993);
nand U21416 (N_21416,N_20700,N_20139);
and U21417 (N_21417,N_20082,N_20823);
nand U21418 (N_21418,N_20238,N_20826);
and U21419 (N_21419,N_20347,N_20636);
and U21420 (N_21420,N_20492,N_20008);
and U21421 (N_21421,N_20342,N_20547);
nor U21422 (N_21422,N_20984,N_20170);
xnor U21423 (N_21423,N_20152,N_20200);
nor U21424 (N_21424,N_20921,N_20300);
nor U21425 (N_21425,N_20101,N_20108);
or U21426 (N_21426,N_20033,N_20162);
nand U21427 (N_21427,N_20750,N_20838);
nor U21428 (N_21428,N_20277,N_20854);
xor U21429 (N_21429,N_20598,N_20186);
nor U21430 (N_21430,N_20788,N_20112);
xor U21431 (N_21431,N_20014,N_20332);
xnor U21432 (N_21432,N_20835,N_20781);
and U21433 (N_21433,N_20212,N_20407);
nand U21434 (N_21434,N_20140,N_20059);
nor U21435 (N_21435,N_20284,N_20579);
xnor U21436 (N_21436,N_20902,N_20592);
nor U21437 (N_21437,N_20886,N_20058);
and U21438 (N_21438,N_20020,N_20766);
nor U21439 (N_21439,N_20106,N_20368);
nand U21440 (N_21440,N_20843,N_20447);
nor U21441 (N_21441,N_20512,N_20416);
nor U21442 (N_21442,N_20624,N_20661);
or U21443 (N_21443,N_20333,N_20457);
xor U21444 (N_21444,N_20268,N_20550);
and U21445 (N_21445,N_20857,N_20610);
and U21446 (N_21446,N_20269,N_20658);
nand U21447 (N_21447,N_20703,N_20518);
and U21448 (N_21448,N_20310,N_20625);
nor U21449 (N_21449,N_20146,N_20974);
xnor U21450 (N_21450,N_20193,N_20023);
xnor U21451 (N_21451,N_20839,N_20748);
and U21452 (N_21452,N_20544,N_20529);
and U21453 (N_21453,N_20308,N_20808);
xor U21454 (N_21454,N_20134,N_20099);
nand U21455 (N_21455,N_20760,N_20484);
and U21456 (N_21456,N_20251,N_20460);
nor U21457 (N_21457,N_20065,N_20858);
nand U21458 (N_21458,N_20459,N_20576);
nor U21459 (N_21459,N_20934,N_20825);
nor U21460 (N_21460,N_20293,N_20754);
nand U21461 (N_21461,N_20169,N_20638);
xnor U21462 (N_21462,N_20160,N_20210);
nor U21463 (N_21463,N_20882,N_20903);
and U21464 (N_21464,N_20067,N_20674);
and U21465 (N_21465,N_20177,N_20582);
or U21466 (N_21466,N_20415,N_20353);
or U21467 (N_21467,N_20528,N_20696);
and U21468 (N_21468,N_20986,N_20419);
xnor U21469 (N_21469,N_20551,N_20301);
and U21470 (N_21470,N_20648,N_20962);
nor U21471 (N_21471,N_20855,N_20361);
or U21472 (N_21472,N_20105,N_20819);
xnor U21473 (N_21473,N_20110,N_20515);
and U21474 (N_21474,N_20207,N_20350);
nor U21475 (N_21475,N_20237,N_20322);
and U21476 (N_21476,N_20953,N_20867);
nand U21477 (N_21477,N_20063,N_20296);
and U21478 (N_21478,N_20642,N_20969);
nor U21479 (N_21479,N_20608,N_20796);
nand U21480 (N_21480,N_20994,N_20507);
nor U21481 (N_21481,N_20410,N_20054);
nand U21482 (N_21482,N_20695,N_20392);
nand U21483 (N_21483,N_20751,N_20066);
or U21484 (N_21484,N_20126,N_20488);
xnor U21485 (N_21485,N_20663,N_20197);
nand U21486 (N_21486,N_20755,N_20373);
nand U21487 (N_21487,N_20872,N_20983);
nor U21488 (N_21488,N_20578,N_20252);
or U21489 (N_21489,N_20567,N_20897);
nand U21490 (N_21490,N_20089,N_20462);
nand U21491 (N_21491,N_20298,N_20138);
xor U21492 (N_21492,N_20010,N_20055);
and U21493 (N_21493,N_20780,N_20918);
nand U21494 (N_21494,N_20987,N_20594);
and U21495 (N_21495,N_20729,N_20456);
xor U21496 (N_21496,N_20691,N_20681);
nor U21497 (N_21497,N_20335,N_20584);
or U21498 (N_21498,N_20429,N_20205);
nand U21499 (N_21499,N_20940,N_20219);
nand U21500 (N_21500,N_20984,N_20449);
nand U21501 (N_21501,N_20969,N_20070);
or U21502 (N_21502,N_20236,N_20609);
or U21503 (N_21503,N_20656,N_20271);
nor U21504 (N_21504,N_20386,N_20010);
or U21505 (N_21505,N_20170,N_20406);
or U21506 (N_21506,N_20415,N_20346);
nor U21507 (N_21507,N_20408,N_20920);
or U21508 (N_21508,N_20225,N_20128);
and U21509 (N_21509,N_20663,N_20416);
xnor U21510 (N_21510,N_20064,N_20222);
and U21511 (N_21511,N_20151,N_20892);
nand U21512 (N_21512,N_20730,N_20397);
xor U21513 (N_21513,N_20077,N_20614);
nand U21514 (N_21514,N_20689,N_20055);
xnor U21515 (N_21515,N_20982,N_20921);
nor U21516 (N_21516,N_20594,N_20470);
xor U21517 (N_21517,N_20241,N_20173);
or U21518 (N_21518,N_20190,N_20203);
xnor U21519 (N_21519,N_20717,N_20759);
xor U21520 (N_21520,N_20977,N_20919);
and U21521 (N_21521,N_20990,N_20151);
or U21522 (N_21522,N_20880,N_20495);
xor U21523 (N_21523,N_20273,N_20931);
and U21524 (N_21524,N_20834,N_20061);
nand U21525 (N_21525,N_20180,N_20770);
or U21526 (N_21526,N_20912,N_20048);
and U21527 (N_21527,N_20741,N_20456);
nor U21528 (N_21528,N_20031,N_20242);
nor U21529 (N_21529,N_20011,N_20385);
nand U21530 (N_21530,N_20180,N_20138);
or U21531 (N_21531,N_20967,N_20623);
or U21532 (N_21532,N_20406,N_20480);
nand U21533 (N_21533,N_20611,N_20844);
nand U21534 (N_21534,N_20363,N_20267);
xnor U21535 (N_21535,N_20822,N_20105);
nand U21536 (N_21536,N_20245,N_20080);
xor U21537 (N_21537,N_20116,N_20330);
xnor U21538 (N_21538,N_20219,N_20002);
and U21539 (N_21539,N_20459,N_20681);
xnor U21540 (N_21540,N_20187,N_20340);
nand U21541 (N_21541,N_20170,N_20241);
or U21542 (N_21542,N_20524,N_20414);
xor U21543 (N_21543,N_20460,N_20625);
or U21544 (N_21544,N_20588,N_20632);
xnor U21545 (N_21545,N_20303,N_20930);
nand U21546 (N_21546,N_20243,N_20347);
or U21547 (N_21547,N_20813,N_20991);
xnor U21548 (N_21548,N_20784,N_20081);
nor U21549 (N_21549,N_20620,N_20124);
nor U21550 (N_21550,N_20895,N_20693);
nor U21551 (N_21551,N_20265,N_20349);
nand U21552 (N_21552,N_20012,N_20805);
nor U21553 (N_21553,N_20663,N_20506);
or U21554 (N_21554,N_20562,N_20164);
nand U21555 (N_21555,N_20364,N_20270);
nor U21556 (N_21556,N_20198,N_20219);
and U21557 (N_21557,N_20050,N_20113);
or U21558 (N_21558,N_20700,N_20876);
and U21559 (N_21559,N_20128,N_20804);
nand U21560 (N_21560,N_20605,N_20421);
nor U21561 (N_21561,N_20072,N_20907);
nor U21562 (N_21562,N_20334,N_20922);
nor U21563 (N_21563,N_20173,N_20768);
nor U21564 (N_21564,N_20496,N_20212);
nor U21565 (N_21565,N_20291,N_20639);
and U21566 (N_21566,N_20523,N_20953);
xnor U21567 (N_21567,N_20797,N_20584);
nand U21568 (N_21568,N_20135,N_20109);
or U21569 (N_21569,N_20990,N_20722);
and U21570 (N_21570,N_20766,N_20590);
or U21571 (N_21571,N_20823,N_20446);
or U21572 (N_21572,N_20875,N_20751);
nor U21573 (N_21573,N_20212,N_20076);
or U21574 (N_21574,N_20085,N_20666);
or U21575 (N_21575,N_20657,N_20366);
and U21576 (N_21576,N_20194,N_20055);
and U21577 (N_21577,N_20074,N_20005);
xnor U21578 (N_21578,N_20298,N_20620);
and U21579 (N_21579,N_20403,N_20587);
and U21580 (N_21580,N_20600,N_20054);
nor U21581 (N_21581,N_20079,N_20959);
nand U21582 (N_21582,N_20247,N_20571);
nor U21583 (N_21583,N_20751,N_20084);
nor U21584 (N_21584,N_20729,N_20254);
or U21585 (N_21585,N_20037,N_20529);
and U21586 (N_21586,N_20068,N_20318);
and U21587 (N_21587,N_20200,N_20408);
or U21588 (N_21588,N_20056,N_20551);
nand U21589 (N_21589,N_20013,N_20948);
and U21590 (N_21590,N_20271,N_20273);
nor U21591 (N_21591,N_20508,N_20524);
or U21592 (N_21592,N_20897,N_20291);
nor U21593 (N_21593,N_20439,N_20311);
nand U21594 (N_21594,N_20706,N_20759);
nand U21595 (N_21595,N_20678,N_20937);
and U21596 (N_21596,N_20102,N_20891);
nand U21597 (N_21597,N_20229,N_20446);
and U21598 (N_21598,N_20813,N_20439);
and U21599 (N_21599,N_20398,N_20932);
and U21600 (N_21600,N_20247,N_20516);
and U21601 (N_21601,N_20596,N_20327);
and U21602 (N_21602,N_20108,N_20414);
nand U21603 (N_21603,N_20779,N_20334);
xor U21604 (N_21604,N_20323,N_20627);
or U21605 (N_21605,N_20832,N_20062);
nand U21606 (N_21606,N_20949,N_20018);
or U21607 (N_21607,N_20004,N_20877);
and U21608 (N_21608,N_20848,N_20569);
nor U21609 (N_21609,N_20634,N_20416);
and U21610 (N_21610,N_20245,N_20317);
nand U21611 (N_21611,N_20109,N_20379);
nor U21612 (N_21612,N_20337,N_20621);
or U21613 (N_21613,N_20785,N_20437);
and U21614 (N_21614,N_20585,N_20450);
or U21615 (N_21615,N_20937,N_20683);
or U21616 (N_21616,N_20073,N_20741);
and U21617 (N_21617,N_20096,N_20446);
or U21618 (N_21618,N_20502,N_20426);
nand U21619 (N_21619,N_20704,N_20110);
and U21620 (N_21620,N_20553,N_20732);
and U21621 (N_21621,N_20347,N_20887);
nand U21622 (N_21622,N_20680,N_20954);
or U21623 (N_21623,N_20032,N_20432);
and U21624 (N_21624,N_20627,N_20966);
nor U21625 (N_21625,N_20918,N_20040);
nor U21626 (N_21626,N_20996,N_20363);
nand U21627 (N_21627,N_20602,N_20199);
xor U21628 (N_21628,N_20906,N_20353);
nor U21629 (N_21629,N_20390,N_20852);
and U21630 (N_21630,N_20489,N_20284);
or U21631 (N_21631,N_20300,N_20977);
nor U21632 (N_21632,N_20775,N_20719);
nand U21633 (N_21633,N_20459,N_20144);
or U21634 (N_21634,N_20072,N_20337);
and U21635 (N_21635,N_20054,N_20268);
and U21636 (N_21636,N_20414,N_20789);
and U21637 (N_21637,N_20077,N_20305);
xnor U21638 (N_21638,N_20206,N_20768);
and U21639 (N_21639,N_20591,N_20008);
nand U21640 (N_21640,N_20191,N_20345);
xor U21641 (N_21641,N_20116,N_20397);
nor U21642 (N_21642,N_20819,N_20994);
nand U21643 (N_21643,N_20748,N_20708);
and U21644 (N_21644,N_20223,N_20519);
nand U21645 (N_21645,N_20644,N_20941);
nor U21646 (N_21646,N_20272,N_20969);
nand U21647 (N_21647,N_20439,N_20636);
and U21648 (N_21648,N_20203,N_20420);
or U21649 (N_21649,N_20953,N_20087);
and U21650 (N_21650,N_20520,N_20114);
and U21651 (N_21651,N_20426,N_20195);
or U21652 (N_21652,N_20251,N_20111);
xor U21653 (N_21653,N_20062,N_20570);
xor U21654 (N_21654,N_20759,N_20729);
nor U21655 (N_21655,N_20771,N_20952);
and U21656 (N_21656,N_20286,N_20183);
nor U21657 (N_21657,N_20728,N_20120);
nand U21658 (N_21658,N_20039,N_20191);
and U21659 (N_21659,N_20712,N_20640);
nor U21660 (N_21660,N_20744,N_20807);
or U21661 (N_21661,N_20316,N_20798);
or U21662 (N_21662,N_20966,N_20091);
or U21663 (N_21663,N_20704,N_20608);
nor U21664 (N_21664,N_20180,N_20500);
and U21665 (N_21665,N_20930,N_20611);
nand U21666 (N_21666,N_20092,N_20736);
xor U21667 (N_21667,N_20487,N_20167);
nor U21668 (N_21668,N_20362,N_20495);
xnor U21669 (N_21669,N_20958,N_20389);
xnor U21670 (N_21670,N_20113,N_20989);
and U21671 (N_21671,N_20894,N_20497);
and U21672 (N_21672,N_20734,N_20407);
and U21673 (N_21673,N_20559,N_20137);
and U21674 (N_21674,N_20036,N_20855);
xnor U21675 (N_21675,N_20621,N_20319);
nand U21676 (N_21676,N_20081,N_20765);
or U21677 (N_21677,N_20360,N_20875);
and U21678 (N_21678,N_20768,N_20663);
xor U21679 (N_21679,N_20475,N_20254);
or U21680 (N_21680,N_20607,N_20930);
or U21681 (N_21681,N_20949,N_20682);
and U21682 (N_21682,N_20518,N_20721);
nand U21683 (N_21683,N_20693,N_20864);
xor U21684 (N_21684,N_20690,N_20974);
nor U21685 (N_21685,N_20743,N_20036);
xnor U21686 (N_21686,N_20707,N_20537);
or U21687 (N_21687,N_20171,N_20389);
and U21688 (N_21688,N_20832,N_20392);
xor U21689 (N_21689,N_20585,N_20319);
nand U21690 (N_21690,N_20063,N_20682);
and U21691 (N_21691,N_20386,N_20260);
nand U21692 (N_21692,N_20046,N_20352);
nor U21693 (N_21693,N_20551,N_20957);
nand U21694 (N_21694,N_20990,N_20259);
and U21695 (N_21695,N_20317,N_20960);
nand U21696 (N_21696,N_20937,N_20443);
and U21697 (N_21697,N_20106,N_20606);
and U21698 (N_21698,N_20764,N_20892);
nor U21699 (N_21699,N_20714,N_20980);
and U21700 (N_21700,N_20786,N_20673);
xor U21701 (N_21701,N_20435,N_20350);
or U21702 (N_21702,N_20620,N_20120);
nor U21703 (N_21703,N_20518,N_20045);
or U21704 (N_21704,N_20712,N_20322);
xor U21705 (N_21705,N_20879,N_20394);
xnor U21706 (N_21706,N_20428,N_20536);
or U21707 (N_21707,N_20103,N_20446);
nand U21708 (N_21708,N_20564,N_20760);
or U21709 (N_21709,N_20363,N_20272);
and U21710 (N_21710,N_20554,N_20414);
and U21711 (N_21711,N_20562,N_20582);
or U21712 (N_21712,N_20559,N_20384);
nor U21713 (N_21713,N_20849,N_20063);
nor U21714 (N_21714,N_20773,N_20872);
or U21715 (N_21715,N_20675,N_20756);
nand U21716 (N_21716,N_20677,N_20535);
and U21717 (N_21717,N_20879,N_20289);
or U21718 (N_21718,N_20728,N_20946);
nor U21719 (N_21719,N_20489,N_20194);
xnor U21720 (N_21720,N_20309,N_20651);
xor U21721 (N_21721,N_20930,N_20654);
nand U21722 (N_21722,N_20406,N_20761);
or U21723 (N_21723,N_20088,N_20480);
nand U21724 (N_21724,N_20251,N_20850);
nand U21725 (N_21725,N_20753,N_20845);
xor U21726 (N_21726,N_20390,N_20065);
nor U21727 (N_21727,N_20907,N_20997);
or U21728 (N_21728,N_20403,N_20770);
nand U21729 (N_21729,N_20884,N_20466);
nor U21730 (N_21730,N_20641,N_20452);
nor U21731 (N_21731,N_20662,N_20183);
and U21732 (N_21732,N_20570,N_20677);
and U21733 (N_21733,N_20265,N_20783);
or U21734 (N_21734,N_20705,N_20837);
and U21735 (N_21735,N_20337,N_20273);
nand U21736 (N_21736,N_20798,N_20566);
xor U21737 (N_21737,N_20940,N_20810);
nand U21738 (N_21738,N_20193,N_20040);
and U21739 (N_21739,N_20136,N_20148);
or U21740 (N_21740,N_20833,N_20294);
nand U21741 (N_21741,N_20381,N_20080);
and U21742 (N_21742,N_20343,N_20864);
nand U21743 (N_21743,N_20671,N_20446);
nand U21744 (N_21744,N_20315,N_20610);
xor U21745 (N_21745,N_20349,N_20267);
xor U21746 (N_21746,N_20017,N_20705);
nor U21747 (N_21747,N_20262,N_20894);
and U21748 (N_21748,N_20451,N_20374);
and U21749 (N_21749,N_20985,N_20193);
or U21750 (N_21750,N_20207,N_20149);
xnor U21751 (N_21751,N_20267,N_20355);
nor U21752 (N_21752,N_20903,N_20414);
or U21753 (N_21753,N_20654,N_20763);
xnor U21754 (N_21754,N_20355,N_20531);
and U21755 (N_21755,N_20466,N_20305);
or U21756 (N_21756,N_20381,N_20901);
nand U21757 (N_21757,N_20959,N_20446);
and U21758 (N_21758,N_20053,N_20065);
and U21759 (N_21759,N_20497,N_20672);
nand U21760 (N_21760,N_20995,N_20956);
xor U21761 (N_21761,N_20251,N_20422);
xnor U21762 (N_21762,N_20865,N_20877);
and U21763 (N_21763,N_20093,N_20871);
nor U21764 (N_21764,N_20314,N_20557);
nand U21765 (N_21765,N_20194,N_20958);
and U21766 (N_21766,N_20272,N_20316);
and U21767 (N_21767,N_20037,N_20409);
and U21768 (N_21768,N_20237,N_20806);
xor U21769 (N_21769,N_20010,N_20807);
xor U21770 (N_21770,N_20651,N_20350);
and U21771 (N_21771,N_20591,N_20793);
and U21772 (N_21772,N_20000,N_20597);
nor U21773 (N_21773,N_20689,N_20780);
and U21774 (N_21774,N_20747,N_20919);
nand U21775 (N_21775,N_20372,N_20248);
nand U21776 (N_21776,N_20303,N_20206);
or U21777 (N_21777,N_20092,N_20299);
or U21778 (N_21778,N_20190,N_20084);
or U21779 (N_21779,N_20862,N_20028);
xnor U21780 (N_21780,N_20829,N_20191);
xor U21781 (N_21781,N_20569,N_20152);
xor U21782 (N_21782,N_20896,N_20397);
or U21783 (N_21783,N_20473,N_20109);
or U21784 (N_21784,N_20352,N_20035);
nor U21785 (N_21785,N_20614,N_20548);
nand U21786 (N_21786,N_20429,N_20251);
or U21787 (N_21787,N_20578,N_20984);
nor U21788 (N_21788,N_20464,N_20521);
or U21789 (N_21789,N_20015,N_20436);
nand U21790 (N_21790,N_20972,N_20833);
xor U21791 (N_21791,N_20201,N_20292);
nand U21792 (N_21792,N_20758,N_20691);
or U21793 (N_21793,N_20366,N_20800);
xnor U21794 (N_21794,N_20440,N_20029);
nor U21795 (N_21795,N_20184,N_20507);
and U21796 (N_21796,N_20278,N_20974);
or U21797 (N_21797,N_20207,N_20926);
and U21798 (N_21798,N_20035,N_20503);
or U21799 (N_21799,N_20620,N_20033);
nand U21800 (N_21800,N_20990,N_20842);
and U21801 (N_21801,N_20095,N_20195);
or U21802 (N_21802,N_20443,N_20782);
xnor U21803 (N_21803,N_20539,N_20785);
or U21804 (N_21804,N_20479,N_20147);
xor U21805 (N_21805,N_20106,N_20558);
nand U21806 (N_21806,N_20809,N_20177);
nor U21807 (N_21807,N_20752,N_20379);
xor U21808 (N_21808,N_20664,N_20642);
nor U21809 (N_21809,N_20592,N_20735);
nand U21810 (N_21810,N_20347,N_20333);
and U21811 (N_21811,N_20418,N_20284);
and U21812 (N_21812,N_20586,N_20919);
xnor U21813 (N_21813,N_20513,N_20966);
nor U21814 (N_21814,N_20013,N_20219);
xor U21815 (N_21815,N_20760,N_20434);
and U21816 (N_21816,N_20013,N_20621);
nand U21817 (N_21817,N_20198,N_20002);
or U21818 (N_21818,N_20559,N_20268);
nand U21819 (N_21819,N_20365,N_20243);
nand U21820 (N_21820,N_20339,N_20676);
and U21821 (N_21821,N_20202,N_20857);
or U21822 (N_21822,N_20466,N_20880);
xnor U21823 (N_21823,N_20502,N_20645);
nand U21824 (N_21824,N_20872,N_20867);
or U21825 (N_21825,N_20382,N_20601);
or U21826 (N_21826,N_20984,N_20673);
and U21827 (N_21827,N_20699,N_20232);
nor U21828 (N_21828,N_20412,N_20152);
nor U21829 (N_21829,N_20324,N_20335);
and U21830 (N_21830,N_20655,N_20828);
nor U21831 (N_21831,N_20337,N_20465);
or U21832 (N_21832,N_20378,N_20082);
xor U21833 (N_21833,N_20542,N_20450);
or U21834 (N_21834,N_20951,N_20784);
and U21835 (N_21835,N_20159,N_20169);
or U21836 (N_21836,N_20626,N_20227);
nor U21837 (N_21837,N_20248,N_20635);
nor U21838 (N_21838,N_20055,N_20401);
nand U21839 (N_21839,N_20678,N_20326);
or U21840 (N_21840,N_20758,N_20780);
nor U21841 (N_21841,N_20882,N_20612);
xnor U21842 (N_21842,N_20672,N_20902);
xnor U21843 (N_21843,N_20688,N_20868);
or U21844 (N_21844,N_20653,N_20554);
nor U21845 (N_21845,N_20702,N_20858);
nor U21846 (N_21846,N_20544,N_20283);
nor U21847 (N_21847,N_20649,N_20924);
xor U21848 (N_21848,N_20372,N_20780);
nand U21849 (N_21849,N_20151,N_20793);
or U21850 (N_21850,N_20165,N_20217);
nor U21851 (N_21851,N_20305,N_20440);
xnor U21852 (N_21852,N_20573,N_20940);
nor U21853 (N_21853,N_20754,N_20438);
or U21854 (N_21854,N_20363,N_20522);
and U21855 (N_21855,N_20693,N_20760);
xor U21856 (N_21856,N_20020,N_20018);
nor U21857 (N_21857,N_20039,N_20856);
nor U21858 (N_21858,N_20790,N_20254);
xor U21859 (N_21859,N_20120,N_20813);
nand U21860 (N_21860,N_20524,N_20297);
or U21861 (N_21861,N_20539,N_20696);
nand U21862 (N_21862,N_20092,N_20156);
nand U21863 (N_21863,N_20213,N_20313);
or U21864 (N_21864,N_20906,N_20270);
nand U21865 (N_21865,N_20623,N_20419);
nor U21866 (N_21866,N_20773,N_20572);
nor U21867 (N_21867,N_20251,N_20494);
nor U21868 (N_21868,N_20725,N_20639);
nand U21869 (N_21869,N_20884,N_20376);
nor U21870 (N_21870,N_20764,N_20742);
or U21871 (N_21871,N_20525,N_20327);
nor U21872 (N_21872,N_20528,N_20562);
or U21873 (N_21873,N_20218,N_20423);
nand U21874 (N_21874,N_20897,N_20832);
and U21875 (N_21875,N_20289,N_20908);
nor U21876 (N_21876,N_20326,N_20023);
nand U21877 (N_21877,N_20677,N_20596);
or U21878 (N_21878,N_20516,N_20535);
nand U21879 (N_21879,N_20075,N_20828);
or U21880 (N_21880,N_20102,N_20518);
xor U21881 (N_21881,N_20756,N_20578);
nor U21882 (N_21882,N_20433,N_20784);
nor U21883 (N_21883,N_20598,N_20481);
xnor U21884 (N_21884,N_20084,N_20040);
and U21885 (N_21885,N_20053,N_20974);
nand U21886 (N_21886,N_20834,N_20583);
nand U21887 (N_21887,N_20843,N_20429);
nor U21888 (N_21888,N_20893,N_20294);
nor U21889 (N_21889,N_20935,N_20123);
xnor U21890 (N_21890,N_20992,N_20994);
nor U21891 (N_21891,N_20661,N_20891);
or U21892 (N_21892,N_20677,N_20297);
xnor U21893 (N_21893,N_20622,N_20896);
nand U21894 (N_21894,N_20065,N_20863);
nor U21895 (N_21895,N_20388,N_20855);
and U21896 (N_21896,N_20633,N_20737);
or U21897 (N_21897,N_20795,N_20004);
xor U21898 (N_21898,N_20049,N_20056);
and U21899 (N_21899,N_20163,N_20220);
xor U21900 (N_21900,N_20941,N_20582);
or U21901 (N_21901,N_20657,N_20137);
nor U21902 (N_21902,N_20192,N_20647);
xnor U21903 (N_21903,N_20905,N_20697);
xor U21904 (N_21904,N_20240,N_20222);
nand U21905 (N_21905,N_20469,N_20778);
nor U21906 (N_21906,N_20447,N_20891);
or U21907 (N_21907,N_20873,N_20032);
nand U21908 (N_21908,N_20887,N_20565);
nor U21909 (N_21909,N_20375,N_20960);
xnor U21910 (N_21910,N_20453,N_20142);
nand U21911 (N_21911,N_20146,N_20631);
or U21912 (N_21912,N_20447,N_20607);
nand U21913 (N_21913,N_20610,N_20876);
or U21914 (N_21914,N_20800,N_20100);
xor U21915 (N_21915,N_20957,N_20741);
xor U21916 (N_21916,N_20157,N_20185);
or U21917 (N_21917,N_20206,N_20457);
and U21918 (N_21918,N_20487,N_20697);
and U21919 (N_21919,N_20813,N_20622);
or U21920 (N_21920,N_20277,N_20183);
xnor U21921 (N_21921,N_20104,N_20269);
and U21922 (N_21922,N_20006,N_20724);
nand U21923 (N_21923,N_20834,N_20692);
and U21924 (N_21924,N_20309,N_20654);
and U21925 (N_21925,N_20085,N_20262);
xor U21926 (N_21926,N_20177,N_20455);
and U21927 (N_21927,N_20048,N_20077);
nor U21928 (N_21928,N_20362,N_20805);
xor U21929 (N_21929,N_20928,N_20433);
xnor U21930 (N_21930,N_20056,N_20944);
xnor U21931 (N_21931,N_20902,N_20101);
nand U21932 (N_21932,N_20888,N_20169);
and U21933 (N_21933,N_20968,N_20093);
nand U21934 (N_21934,N_20427,N_20343);
nor U21935 (N_21935,N_20123,N_20312);
or U21936 (N_21936,N_20464,N_20182);
nor U21937 (N_21937,N_20926,N_20673);
nor U21938 (N_21938,N_20732,N_20507);
and U21939 (N_21939,N_20531,N_20215);
or U21940 (N_21940,N_20181,N_20450);
or U21941 (N_21941,N_20375,N_20885);
xnor U21942 (N_21942,N_20018,N_20061);
and U21943 (N_21943,N_20108,N_20052);
or U21944 (N_21944,N_20709,N_20725);
or U21945 (N_21945,N_20875,N_20145);
xnor U21946 (N_21946,N_20745,N_20120);
xor U21947 (N_21947,N_20201,N_20242);
nor U21948 (N_21948,N_20242,N_20235);
or U21949 (N_21949,N_20385,N_20991);
nand U21950 (N_21950,N_20860,N_20384);
xnor U21951 (N_21951,N_20553,N_20762);
nor U21952 (N_21952,N_20902,N_20950);
xor U21953 (N_21953,N_20265,N_20490);
or U21954 (N_21954,N_20950,N_20338);
xor U21955 (N_21955,N_20508,N_20992);
nand U21956 (N_21956,N_20708,N_20136);
and U21957 (N_21957,N_20878,N_20646);
xnor U21958 (N_21958,N_20884,N_20882);
or U21959 (N_21959,N_20425,N_20230);
and U21960 (N_21960,N_20880,N_20489);
and U21961 (N_21961,N_20436,N_20921);
and U21962 (N_21962,N_20656,N_20191);
nand U21963 (N_21963,N_20644,N_20314);
and U21964 (N_21964,N_20075,N_20658);
xnor U21965 (N_21965,N_20161,N_20943);
nand U21966 (N_21966,N_20403,N_20794);
nor U21967 (N_21967,N_20637,N_20159);
and U21968 (N_21968,N_20596,N_20475);
and U21969 (N_21969,N_20398,N_20374);
or U21970 (N_21970,N_20108,N_20614);
and U21971 (N_21971,N_20184,N_20101);
nand U21972 (N_21972,N_20886,N_20266);
and U21973 (N_21973,N_20679,N_20696);
and U21974 (N_21974,N_20829,N_20496);
xor U21975 (N_21975,N_20391,N_20149);
nor U21976 (N_21976,N_20336,N_20856);
or U21977 (N_21977,N_20816,N_20793);
nor U21978 (N_21978,N_20109,N_20090);
nor U21979 (N_21979,N_20438,N_20983);
nor U21980 (N_21980,N_20730,N_20595);
or U21981 (N_21981,N_20936,N_20572);
nand U21982 (N_21982,N_20707,N_20427);
or U21983 (N_21983,N_20213,N_20342);
nor U21984 (N_21984,N_20488,N_20352);
nor U21985 (N_21985,N_20773,N_20351);
and U21986 (N_21986,N_20242,N_20134);
xnor U21987 (N_21987,N_20701,N_20422);
nor U21988 (N_21988,N_20346,N_20572);
nand U21989 (N_21989,N_20145,N_20907);
or U21990 (N_21990,N_20596,N_20114);
or U21991 (N_21991,N_20559,N_20472);
nand U21992 (N_21992,N_20087,N_20516);
xor U21993 (N_21993,N_20919,N_20952);
or U21994 (N_21994,N_20093,N_20996);
or U21995 (N_21995,N_20017,N_20388);
and U21996 (N_21996,N_20913,N_20872);
and U21997 (N_21997,N_20253,N_20754);
nand U21998 (N_21998,N_20862,N_20757);
and U21999 (N_21999,N_20391,N_20011);
nand U22000 (N_22000,N_21915,N_21939);
nand U22001 (N_22001,N_21794,N_21152);
or U22002 (N_22002,N_21027,N_21405);
nand U22003 (N_22003,N_21746,N_21907);
or U22004 (N_22004,N_21838,N_21795);
nor U22005 (N_22005,N_21367,N_21873);
nand U22006 (N_22006,N_21100,N_21351);
nor U22007 (N_22007,N_21228,N_21604);
or U22008 (N_22008,N_21964,N_21408);
and U22009 (N_22009,N_21602,N_21893);
nand U22010 (N_22010,N_21242,N_21350);
nor U22011 (N_22011,N_21155,N_21861);
or U22012 (N_22012,N_21081,N_21678);
or U22013 (N_22013,N_21841,N_21262);
and U22014 (N_22014,N_21600,N_21785);
xnor U22015 (N_22015,N_21721,N_21134);
nand U22016 (N_22016,N_21680,N_21454);
and U22017 (N_22017,N_21388,N_21821);
xor U22018 (N_22018,N_21653,N_21187);
nor U22019 (N_22019,N_21220,N_21806);
xor U22020 (N_22020,N_21807,N_21896);
or U22021 (N_22021,N_21269,N_21993);
nor U22022 (N_22022,N_21518,N_21591);
nor U22023 (N_22023,N_21411,N_21022);
nor U22024 (N_22024,N_21484,N_21120);
nor U22025 (N_22025,N_21357,N_21267);
xnor U22026 (N_22026,N_21249,N_21998);
nor U22027 (N_22027,N_21528,N_21648);
and U22028 (N_22028,N_21299,N_21483);
xor U22029 (N_22029,N_21019,N_21361);
and U22030 (N_22030,N_21194,N_21193);
nand U22031 (N_22031,N_21307,N_21223);
nor U22032 (N_22032,N_21979,N_21898);
or U22033 (N_22033,N_21103,N_21966);
xor U22034 (N_22034,N_21215,N_21564);
nand U22035 (N_22035,N_21595,N_21895);
and U22036 (N_22036,N_21497,N_21149);
and U22037 (N_22037,N_21627,N_21329);
nor U22038 (N_22038,N_21649,N_21894);
xor U22039 (N_22039,N_21396,N_21079);
or U22040 (N_22040,N_21264,N_21859);
or U22041 (N_22041,N_21168,N_21551);
nor U22042 (N_22042,N_21769,N_21363);
xnor U22043 (N_22043,N_21513,N_21020);
nand U22044 (N_22044,N_21401,N_21008);
nand U22045 (N_22045,N_21904,N_21224);
xor U22046 (N_22046,N_21382,N_21071);
nand U22047 (N_22047,N_21478,N_21852);
xor U22048 (N_22048,N_21125,N_21694);
or U22049 (N_22049,N_21707,N_21280);
nor U22050 (N_22050,N_21856,N_21384);
nor U22051 (N_22051,N_21586,N_21308);
or U22052 (N_22052,N_21098,N_21573);
nand U22053 (N_22053,N_21538,N_21677);
nand U22054 (N_22054,N_21963,N_21397);
nor U22055 (N_22055,N_21569,N_21559);
nor U22056 (N_22056,N_21212,N_21706);
and U22057 (N_22057,N_21863,N_21309);
and U22058 (N_22058,N_21684,N_21037);
nor U22059 (N_22059,N_21668,N_21550);
nor U22060 (N_22060,N_21912,N_21923);
nand U22061 (N_22061,N_21186,N_21687);
xnor U22062 (N_22062,N_21990,N_21034);
nor U22063 (N_22063,N_21655,N_21878);
nor U22064 (N_22064,N_21747,N_21886);
nand U22065 (N_22065,N_21272,N_21960);
xor U22066 (N_22066,N_21069,N_21651);
and U22067 (N_22067,N_21466,N_21461);
or U22068 (N_22068,N_21410,N_21250);
and U22069 (N_22069,N_21734,N_21084);
or U22070 (N_22070,N_21750,N_21984);
or U22071 (N_22071,N_21953,N_21201);
nand U22072 (N_22072,N_21509,N_21144);
and U22073 (N_22073,N_21441,N_21185);
nor U22074 (N_22074,N_21537,N_21415);
nand U22075 (N_22075,N_21216,N_21502);
and U22076 (N_22076,N_21047,N_21266);
or U22077 (N_22077,N_21700,N_21645);
nand U22078 (N_22078,N_21636,N_21942);
nor U22079 (N_22079,N_21183,N_21395);
nor U22080 (N_22080,N_21713,N_21536);
and U22081 (N_22081,N_21468,N_21161);
and U22082 (N_22082,N_21697,N_21469);
or U22083 (N_22083,N_21652,N_21446);
xor U22084 (N_22084,N_21891,N_21634);
nand U22085 (N_22085,N_21630,N_21941);
xor U22086 (N_22086,N_21780,N_21801);
xnor U22087 (N_22087,N_21174,N_21567);
and U22088 (N_22088,N_21312,N_21608);
xnor U22089 (N_22089,N_21799,N_21371);
and U22090 (N_22090,N_21742,N_21880);
nor U22091 (N_22091,N_21903,N_21711);
xor U22092 (N_22092,N_21989,N_21414);
xor U22093 (N_22093,N_21305,N_21531);
nand U22094 (N_22094,N_21784,N_21864);
or U22095 (N_22095,N_21115,N_21511);
nand U22096 (N_22096,N_21260,N_21050);
or U22097 (N_22097,N_21210,N_21119);
nor U22098 (N_22098,N_21804,N_21259);
and U22099 (N_22099,N_21944,N_21337);
nand U22100 (N_22100,N_21127,N_21251);
or U22101 (N_22101,N_21849,N_21080);
and U22102 (N_22102,N_21688,N_21965);
and U22103 (N_22103,N_21736,N_21368);
nor U22104 (N_22104,N_21096,N_21741);
and U22105 (N_22105,N_21973,N_21541);
xor U22106 (N_22106,N_21535,N_21610);
or U22107 (N_22107,N_21580,N_21418);
nand U22108 (N_22108,N_21777,N_21114);
nor U22109 (N_22109,N_21974,N_21045);
nor U22110 (N_22110,N_21885,N_21876);
and U22111 (N_22111,N_21376,N_21954);
nand U22112 (N_22112,N_21934,N_21837);
nor U22113 (N_22113,N_21874,N_21135);
xor U22114 (N_22114,N_21563,N_21407);
xor U22115 (N_22115,N_21715,N_21254);
nand U22116 (N_22116,N_21670,N_21510);
or U22117 (N_22117,N_21360,N_21031);
or U22118 (N_22118,N_21703,N_21546);
xnor U22119 (N_22119,N_21151,N_21459);
xnor U22120 (N_22120,N_21802,N_21381);
nand U22121 (N_22121,N_21994,N_21179);
nand U22122 (N_22122,N_21204,N_21409);
nand U22123 (N_22123,N_21579,N_21091);
nand U22124 (N_22124,N_21393,N_21596);
or U22125 (N_22125,N_21659,N_21727);
nand U22126 (N_22126,N_21805,N_21158);
or U22127 (N_22127,N_21024,N_21004);
and U22128 (N_22128,N_21951,N_21032);
xnor U22129 (N_22129,N_21798,N_21871);
or U22130 (N_22130,N_21137,N_21203);
or U22131 (N_22131,N_21975,N_21237);
nor U22132 (N_22132,N_21824,N_21631);
nand U22133 (N_22133,N_21673,N_21489);
and U22134 (N_22134,N_21702,N_21000);
or U22135 (N_22135,N_21916,N_21773);
or U22136 (N_22136,N_21054,N_21012);
nand U22137 (N_22137,N_21021,N_21553);
or U22138 (N_22138,N_21171,N_21017);
and U22139 (N_22139,N_21705,N_21763);
nor U22140 (N_22140,N_21301,N_21815);
xnor U22141 (N_22141,N_21331,N_21180);
nand U22142 (N_22142,N_21731,N_21279);
nand U22143 (N_22143,N_21496,N_21315);
nand U22144 (N_22144,N_21474,N_21218);
nand U22145 (N_22145,N_21060,N_21162);
nor U22146 (N_22146,N_21525,N_21028);
nor U22147 (N_22147,N_21901,N_21853);
nor U22148 (N_22148,N_21882,N_21790);
and U22149 (N_22149,N_21978,N_21530);
and U22150 (N_22150,N_21503,N_21689);
xnor U22151 (N_22151,N_21199,N_21486);
and U22152 (N_22152,N_21517,N_21850);
nand U22153 (N_22153,N_21759,N_21992);
and U22154 (N_22154,N_21356,N_21416);
or U22155 (N_22155,N_21319,N_21172);
nand U22156 (N_22156,N_21438,N_21547);
nand U22157 (N_22157,N_21555,N_21450);
and U22158 (N_22158,N_21048,N_21198);
xnor U22159 (N_22159,N_21839,N_21313);
or U22160 (N_22160,N_21226,N_21002);
xnor U22161 (N_22161,N_21825,N_21040);
or U22162 (N_22162,N_21906,N_21059);
or U22163 (N_22163,N_21585,N_21255);
nand U22164 (N_22164,N_21442,N_21811);
nor U22165 (N_22165,N_21933,N_21888);
xnor U22166 (N_22166,N_21189,N_21845);
nand U22167 (N_22167,N_21128,N_21744);
or U22168 (N_22168,N_21093,N_21112);
nor U22169 (N_22169,N_21222,N_21813);
xnor U22170 (N_22170,N_21075,N_21529);
nor U22171 (N_22171,N_21866,N_21641);
and U22172 (N_22172,N_21905,N_21877);
nor U22173 (N_22173,N_21003,N_21061);
nand U22174 (N_22174,N_21730,N_21138);
or U22175 (N_22175,N_21111,N_21423);
xor U22176 (N_22176,N_21462,N_21330);
nor U22177 (N_22177,N_21320,N_21967);
nor U22178 (N_22178,N_21449,N_21872);
xnor U22179 (N_22179,N_21437,N_21899);
nand U22180 (N_22180,N_21487,N_21221);
nand U22181 (N_22181,N_21686,N_21936);
nand U22182 (N_22182,N_21326,N_21751);
nor U22183 (N_22183,N_21661,N_21412);
or U22184 (N_22184,N_21584,N_21427);
nand U22185 (N_22185,N_21399,N_21614);
xnor U22186 (N_22186,N_21922,N_21665);
or U22187 (N_22187,N_21052,N_21136);
and U22188 (N_22188,N_21667,N_21160);
xor U22189 (N_22189,N_21229,N_21778);
xor U22190 (N_22190,N_21341,N_21398);
and U22191 (N_22191,N_21304,N_21757);
nor U22192 (N_22192,N_21295,N_21285);
and U22193 (N_22193,N_21981,N_21006);
or U22194 (N_22194,N_21745,N_21911);
nand U22195 (N_22195,N_21113,N_21930);
or U22196 (N_22196,N_21150,N_21797);
and U22197 (N_22197,N_21810,N_21090);
or U22198 (N_22198,N_21372,N_21302);
nor U22199 (N_22199,N_21521,N_21338);
or U22200 (N_22200,N_21347,N_21765);
nor U22201 (N_22201,N_21833,N_21758);
or U22202 (N_22202,N_21991,N_21129);
or U22203 (N_22203,N_21656,N_21683);
xor U22204 (N_22204,N_21364,N_21914);
or U22205 (N_22205,N_21325,N_21523);
and U22206 (N_22206,N_21380,N_21840);
or U22207 (N_22207,N_21495,N_21465);
or U22208 (N_22208,N_21755,N_21719);
nor U22209 (N_22209,N_21800,N_21265);
or U22210 (N_22210,N_21718,N_21246);
nor U22211 (N_22211,N_21464,N_21327);
xnor U22212 (N_22212,N_21597,N_21879);
nand U22213 (N_22213,N_21188,N_21995);
nor U22214 (N_22214,N_21419,N_21714);
xnor U22215 (N_22215,N_21952,N_21732);
or U22216 (N_22216,N_21147,N_21165);
and U22217 (N_22217,N_21029,N_21725);
or U22218 (N_22218,N_21917,N_21178);
and U22219 (N_22219,N_21753,N_21383);
or U22220 (N_22220,N_21067,N_21533);
and U22221 (N_22221,N_21622,N_21344);
nand U22222 (N_22222,N_21077,N_21240);
nand U22223 (N_22223,N_21348,N_21016);
or U22224 (N_22224,N_21268,N_21576);
nand U22225 (N_22225,N_21572,N_21516);
nand U22226 (N_22226,N_21480,N_21154);
nand U22227 (N_22227,N_21182,N_21925);
xnor U22228 (N_22228,N_21498,N_21776);
or U22229 (N_22229,N_21787,N_21403);
xnor U22230 (N_22230,N_21654,N_21094);
nand U22231 (N_22231,N_21752,N_21558);
nand U22232 (N_22232,N_21682,N_21760);
nand U22233 (N_22233,N_21349,N_21213);
xnor U22234 (N_22234,N_21292,N_21104);
and U22235 (N_22235,N_21664,N_21791);
nor U22236 (N_22236,N_21574,N_21190);
nand U22237 (N_22237,N_21286,N_21789);
xor U22238 (N_22238,N_21107,N_21290);
nand U22239 (N_22239,N_21297,N_21812);
nor U22240 (N_22240,N_21662,N_21253);
or U22241 (N_22241,N_21733,N_21606);
nand U22242 (N_22242,N_21832,N_21184);
and U22243 (N_22243,N_21458,N_21448);
xor U22244 (N_22244,N_21287,N_21157);
xor U22245 (N_22245,N_21962,N_21261);
nand U22246 (N_22246,N_21053,N_21532);
and U22247 (N_22247,N_21311,N_21858);
or U22248 (N_22248,N_21406,N_21010);
and U22249 (N_22249,N_21615,N_21926);
or U22250 (N_22250,N_21566,N_21601);
nand U22251 (N_22251,N_21013,N_21842);
and U22252 (N_22252,N_21626,N_21018);
nand U22253 (N_22253,N_21823,N_21972);
xnor U22254 (N_22254,N_21712,N_21870);
or U22255 (N_22255,N_21507,N_21083);
or U22256 (N_22256,N_21835,N_21007);
or U22257 (N_22257,N_21435,N_21314);
nand U22258 (N_22258,N_21803,N_21938);
or U22259 (N_22259,N_21549,N_21628);
xor U22260 (N_22260,N_21303,N_21639);
and U22261 (N_22261,N_21704,N_21488);
nand U22262 (N_22262,N_21116,N_21969);
xnor U22263 (N_22263,N_21754,N_21353);
nand U22264 (N_22264,N_21726,N_21339);
xnor U22265 (N_22265,N_21560,N_21781);
nor U22266 (N_22266,N_21200,N_21657);
nand U22267 (N_22267,N_21793,N_21514);
nand U22268 (N_22268,N_21310,N_21623);
or U22269 (N_22269,N_21208,N_21177);
xnor U22270 (N_22270,N_21666,N_21475);
nand U22271 (N_22271,N_21556,N_21082);
xnor U22272 (N_22272,N_21695,N_21336);
and U22273 (N_22273,N_21211,N_21543);
or U22274 (N_22274,N_21425,N_21582);
or U22275 (N_22275,N_21515,N_21782);
nand U22276 (N_22276,N_21851,N_21997);
nor U22277 (N_22277,N_21023,N_21940);
nand U22278 (N_22278,N_21971,N_21625);
xor U22279 (N_22279,N_21479,N_21571);
nand U22280 (N_22280,N_21918,N_21501);
nand U22281 (N_22281,N_21039,N_21477);
nand U22282 (N_22282,N_21690,N_21430);
and U22283 (N_22283,N_21044,N_21142);
and U22284 (N_22284,N_21494,N_21463);
or U22285 (N_22285,N_21522,N_21389);
xnor U22286 (N_22286,N_21500,N_21354);
and U22287 (N_22287,N_21176,N_21252);
xor U22288 (N_22288,N_21982,N_21232);
xor U22289 (N_22289,N_21089,N_21692);
xnor U22290 (N_22290,N_21121,N_21554);
and U22291 (N_22291,N_21701,N_21927);
nand U22292 (N_22292,N_21593,N_21238);
and U22293 (N_22293,N_21598,N_21605);
xnor U22294 (N_22294,N_21035,N_21544);
and U22295 (N_22295,N_21629,N_21524);
or U22296 (N_22296,N_21470,N_21085);
nand U22297 (N_22297,N_21064,N_21101);
nand U22298 (N_22298,N_21961,N_21456);
and U22299 (N_22299,N_21424,N_21439);
nor U22300 (N_22300,N_21033,N_21374);
and U22301 (N_22301,N_21729,N_21072);
nand U22302 (N_22302,N_21959,N_21207);
nor U22303 (N_22303,N_21696,N_21378);
or U22304 (N_22304,N_21088,N_21637);
xor U22305 (N_22305,N_21740,N_21830);
or U22306 (N_22306,N_21445,N_21175);
xnor U22307 (N_22307,N_21482,N_21011);
nor U22308 (N_22308,N_21428,N_21334);
nand U22309 (N_22309,N_21041,N_21996);
nor U22310 (N_22310,N_21433,N_21256);
or U22311 (N_22311,N_21170,N_21455);
or U22312 (N_22312,N_21476,N_21950);
and U22313 (N_22313,N_21577,N_21913);
xor U22314 (N_22314,N_21291,N_21693);
xnor U22315 (N_22315,N_21947,N_21362);
nor U22316 (N_22316,N_21685,N_21117);
nor U22317 (N_22317,N_21768,N_21771);
xor U22318 (N_22318,N_21248,N_21046);
or U22319 (N_22319,N_21457,N_21214);
nor U22320 (N_22320,N_21390,N_21365);
or U22321 (N_22321,N_21087,N_21352);
xor U22322 (N_22322,N_21908,N_21073);
xnor U22323 (N_22323,N_21831,N_21328);
or U22324 (N_22324,N_21646,N_21788);
and U22325 (N_22325,N_21369,N_21066);
or U22326 (N_22326,N_21391,N_21206);
xnor U22327 (N_22327,N_21743,N_21400);
xnor U22328 (N_22328,N_21471,N_21335);
nand U22329 (N_22329,N_21650,N_21043);
and U22330 (N_22330,N_21321,N_21735);
xnor U22331 (N_22331,N_21025,N_21057);
and U22332 (N_22332,N_21583,N_21422);
or U22333 (N_22333,N_21030,N_21698);
and U22334 (N_22334,N_21300,N_21599);
and U22335 (N_22335,N_21834,N_21062);
and U22336 (N_22336,N_21676,N_21619);
xor U22337 (N_22337,N_21792,N_21594);
and U22338 (N_22338,N_21884,N_21526);
nor U22339 (N_22339,N_21846,N_21404);
or U22340 (N_22340,N_21542,N_21239);
nand U22341 (N_22341,N_21283,N_21889);
nand U22342 (N_22342,N_21985,N_21843);
and U22343 (N_22343,N_21281,N_21263);
nor U22344 (N_22344,N_21491,N_21472);
and U22345 (N_22345,N_21658,N_21289);
xor U22346 (N_22346,N_21058,N_21426);
or U22347 (N_22347,N_21820,N_21274);
or U22348 (N_22348,N_21921,N_21231);
xor U22349 (N_22349,N_21722,N_21828);
xnor U22350 (N_22350,N_21724,N_21796);
and U22351 (N_22351,N_21153,N_21716);
and U22352 (N_22352,N_21481,N_21429);
and U22353 (N_22353,N_21130,N_21562);
or U22354 (N_22354,N_21230,N_21588);
nor U22355 (N_22355,N_21099,N_21737);
and U22356 (N_22356,N_21143,N_21946);
and U22357 (N_22357,N_21860,N_21146);
nand U22358 (N_22358,N_21490,N_21275);
nor U22359 (N_22359,N_21026,N_21163);
xor U22360 (N_22360,N_21009,N_21244);
nor U22361 (N_22361,N_21192,N_21643);
or U22362 (N_22362,N_21774,N_21862);
xnor U22363 (N_22363,N_21123,N_21294);
nand U22364 (N_22364,N_21519,N_21633);
nand U22365 (N_22365,N_21106,N_21855);
and U22366 (N_22366,N_21575,N_21865);
nor U22367 (N_22367,N_21346,N_21931);
nor U22368 (N_22368,N_21370,N_21443);
nor U22369 (N_22369,N_21209,N_21306);
nor U22370 (N_22370,N_21282,N_21097);
xnor U22371 (N_22371,N_21417,N_21674);
or U22372 (N_22372,N_21108,N_21890);
nand U22373 (N_22373,N_21051,N_21068);
nor U22374 (N_22374,N_21557,N_21568);
xor U22375 (N_22375,N_21392,N_21976);
or U22376 (N_22376,N_21005,N_21723);
nand U22377 (N_22377,N_21166,N_21247);
nand U22378 (N_22378,N_21647,N_21420);
nor U22379 (N_22379,N_21609,N_21520);
xor U22380 (N_22380,N_21988,N_21968);
and U22381 (N_22381,N_21355,N_21775);
and U22382 (N_22382,N_21540,N_21063);
xor U22383 (N_22383,N_21095,N_21958);
nand U22384 (N_22384,N_21049,N_21679);
nand U22385 (N_22385,N_21822,N_21772);
nor U22386 (N_22386,N_21561,N_21202);
and U22387 (N_22387,N_21955,N_21273);
xnor U22388 (N_22388,N_21590,N_21373);
nor U22389 (N_22389,N_21139,N_21332);
nand U22390 (N_22390,N_21739,N_21014);
xor U22391 (N_22391,N_21225,N_21159);
nor U22392 (N_22392,N_21900,N_21074);
nand U22393 (N_22393,N_21783,N_21296);
xnor U22394 (N_22394,N_21548,N_21945);
and U22395 (N_22395,N_21245,N_21847);
nand U22396 (N_22396,N_21042,N_21432);
and U22397 (N_22397,N_21819,N_21038);
xor U22398 (N_22398,N_21434,N_21808);
nor U22399 (N_22399,N_21581,N_21887);
nor U22400 (N_22400,N_21883,N_21640);
or U22401 (N_22401,N_21875,N_21708);
or U22402 (N_22402,N_21243,N_21829);
nand U22403 (N_22403,N_21169,N_21452);
nand U22404 (N_22404,N_21132,N_21316);
xnor U22405 (N_22405,N_21762,N_21492);
xor U22406 (N_22406,N_21140,N_21848);
and U22407 (N_22407,N_21191,N_21620);
and U22408 (N_22408,N_21956,N_21317);
and U22409 (N_22409,N_21618,N_21977);
xor U22410 (N_22410,N_21366,N_21818);
xnor U22411 (N_22411,N_21671,N_21324);
nor U22412 (N_22412,N_21709,N_21728);
or U22413 (N_22413,N_21611,N_21276);
nand U22414 (N_22414,N_21816,N_21133);
nor U22415 (N_22415,N_21681,N_21892);
and U22416 (N_22416,N_21980,N_21506);
or U22417 (N_22417,N_21578,N_21748);
and U22418 (N_22418,N_21375,N_21638);
or U22419 (N_22419,N_21570,N_21126);
nand U22420 (N_22420,N_21131,N_21485);
or U22421 (N_22421,N_21691,N_21493);
and U22422 (N_22422,N_21987,N_21141);
nand U22423 (N_22423,N_21910,N_21761);
nand U22424 (N_22424,N_21957,N_21219);
or U22425 (N_22425,N_21413,N_21451);
xnor U22426 (N_22426,N_21612,N_21015);
xnor U22427 (N_22427,N_21539,N_21056);
xnor U22428 (N_22428,N_21181,N_21340);
nor U22429 (N_22429,N_21675,N_21227);
nor U22430 (N_22430,N_21814,N_21277);
nand U22431 (N_22431,N_21999,N_21738);
and U22432 (N_22432,N_21779,N_21756);
xor U22433 (N_22433,N_21065,N_21786);
nor U22434 (N_22434,N_21644,N_21770);
and U22435 (N_22435,N_21453,N_21358);
nand U22436 (N_22436,N_21270,N_21616);
and U22437 (N_22437,N_21909,N_21512);
and U22438 (N_22438,N_21983,N_21589);
nor U22439 (N_22439,N_21937,N_21402);
xnor U22440 (N_22440,N_21672,N_21233);
xor U22441 (N_22441,N_21817,N_21467);
nor U22442 (N_22442,N_21387,N_21343);
xor U22443 (N_22443,N_21421,N_21499);
or U22444 (N_22444,N_21924,N_21284);
nand U22445 (N_22445,N_21444,N_21298);
xnor U22446 (N_22446,N_21164,N_21935);
and U22447 (N_22447,N_21613,N_21236);
nand U22448 (N_22448,N_21001,N_21070);
xnor U22449 (N_22449,N_21844,N_21271);
nor U22450 (N_22450,N_21447,N_21436);
and U22451 (N_22451,N_21948,N_21460);
xnor U22452 (N_22452,N_21869,N_21929);
or U22453 (N_22453,N_21986,N_21318);
and U22454 (N_22454,N_21867,N_21086);
and U22455 (N_22455,N_21110,N_21505);
nand U22456 (N_22456,N_21767,N_21145);
or U22457 (N_22457,N_21076,N_21809);
nor U22458 (N_22458,N_21624,N_21109);
nand U22459 (N_22459,N_21122,N_21868);
xnor U22460 (N_22460,N_21196,N_21217);
xor U22461 (N_22461,N_21766,N_21920);
and U22462 (N_22462,N_21385,N_21592);
nand U22463 (N_22463,N_21173,N_21603);
and U22464 (N_22464,N_21635,N_21970);
xor U22465 (N_22465,N_21102,N_21826);
or U22466 (N_22466,N_21545,N_21534);
nand U22467 (N_22467,N_21377,N_21431);
and U22468 (N_22468,N_21587,N_21148);
nor U22469 (N_22469,N_21386,N_21293);
nor U22470 (N_22470,N_21167,N_21234);
nand U22471 (N_22471,N_21928,N_21607);
and U22472 (N_22472,N_21124,N_21565);
nand U22473 (N_22473,N_21394,N_21943);
nand U22474 (N_22474,N_21197,N_21717);
nand U22475 (N_22475,N_21258,N_21379);
and U22476 (N_22476,N_21235,N_21323);
nand U22477 (N_22477,N_21949,N_21919);
xnor U22478 (N_22478,N_21359,N_21617);
and U22479 (N_22479,N_21345,N_21078);
or U22480 (N_22480,N_21710,N_21932);
nor U22481 (N_22481,N_21241,N_21827);
xor U22482 (N_22482,N_21504,N_21552);
or U22483 (N_22483,N_21257,N_21902);
xor U22484 (N_22484,N_21473,N_21836);
or U22485 (N_22485,N_21092,N_21632);
nand U22486 (N_22486,N_21105,N_21195);
nor U22487 (N_22487,N_21897,N_21621);
or U22488 (N_22488,N_21333,N_21508);
nand U22489 (N_22489,N_21118,N_21854);
nand U22490 (N_22490,N_21663,N_21036);
xnor U22491 (N_22491,N_21660,N_21322);
nor U22492 (N_22492,N_21699,N_21288);
nand U22493 (N_22493,N_21527,N_21440);
nor U22494 (N_22494,N_21055,N_21205);
xor U22495 (N_22495,N_21278,N_21720);
and U22496 (N_22496,N_21342,N_21881);
or U22497 (N_22497,N_21857,N_21156);
and U22498 (N_22498,N_21764,N_21669);
and U22499 (N_22499,N_21642,N_21749);
nand U22500 (N_22500,N_21585,N_21021);
nand U22501 (N_22501,N_21443,N_21582);
or U22502 (N_22502,N_21122,N_21126);
nor U22503 (N_22503,N_21429,N_21960);
nor U22504 (N_22504,N_21624,N_21882);
and U22505 (N_22505,N_21113,N_21240);
xor U22506 (N_22506,N_21843,N_21871);
nand U22507 (N_22507,N_21010,N_21699);
nor U22508 (N_22508,N_21986,N_21818);
nand U22509 (N_22509,N_21015,N_21661);
nand U22510 (N_22510,N_21505,N_21132);
nor U22511 (N_22511,N_21034,N_21012);
and U22512 (N_22512,N_21864,N_21635);
and U22513 (N_22513,N_21281,N_21202);
xnor U22514 (N_22514,N_21556,N_21559);
nand U22515 (N_22515,N_21569,N_21534);
and U22516 (N_22516,N_21083,N_21364);
or U22517 (N_22517,N_21506,N_21562);
nor U22518 (N_22518,N_21647,N_21268);
or U22519 (N_22519,N_21489,N_21363);
or U22520 (N_22520,N_21218,N_21935);
nor U22521 (N_22521,N_21118,N_21506);
or U22522 (N_22522,N_21367,N_21727);
nor U22523 (N_22523,N_21170,N_21747);
nand U22524 (N_22524,N_21902,N_21284);
xnor U22525 (N_22525,N_21918,N_21403);
and U22526 (N_22526,N_21591,N_21851);
nor U22527 (N_22527,N_21426,N_21325);
and U22528 (N_22528,N_21789,N_21867);
or U22529 (N_22529,N_21276,N_21863);
xor U22530 (N_22530,N_21004,N_21702);
or U22531 (N_22531,N_21152,N_21496);
xor U22532 (N_22532,N_21562,N_21362);
nand U22533 (N_22533,N_21502,N_21084);
or U22534 (N_22534,N_21352,N_21060);
or U22535 (N_22535,N_21038,N_21829);
xor U22536 (N_22536,N_21845,N_21870);
or U22537 (N_22537,N_21428,N_21738);
xor U22538 (N_22538,N_21699,N_21898);
or U22539 (N_22539,N_21320,N_21310);
nor U22540 (N_22540,N_21197,N_21128);
and U22541 (N_22541,N_21871,N_21979);
and U22542 (N_22542,N_21575,N_21185);
nor U22543 (N_22543,N_21740,N_21766);
and U22544 (N_22544,N_21803,N_21337);
nand U22545 (N_22545,N_21762,N_21768);
nand U22546 (N_22546,N_21635,N_21213);
nand U22547 (N_22547,N_21487,N_21962);
xnor U22548 (N_22548,N_21152,N_21827);
xor U22549 (N_22549,N_21583,N_21952);
nand U22550 (N_22550,N_21890,N_21171);
and U22551 (N_22551,N_21409,N_21339);
or U22552 (N_22552,N_21523,N_21121);
and U22553 (N_22553,N_21488,N_21277);
nor U22554 (N_22554,N_21472,N_21006);
and U22555 (N_22555,N_21514,N_21715);
xor U22556 (N_22556,N_21330,N_21766);
and U22557 (N_22557,N_21705,N_21562);
xor U22558 (N_22558,N_21301,N_21390);
nand U22559 (N_22559,N_21658,N_21681);
xnor U22560 (N_22560,N_21824,N_21559);
or U22561 (N_22561,N_21589,N_21809);
or U22562 (N_22562,N_21201,N_21370);
and U22563 (N_22563,N_21697,N_21459);
nand U22564 (N_22564,N_21043,N_21443);
nand U22565 (N_22565,N_21974,N_21293);
and U22566 (N_22566,N_21030,N_21340);
or U22567 (N_22567,N_21001,N_21806);
nand U22568 (N_22568,N_21255,N_21987);
or U22569 (N_22569,N_21168,N_21621);
nand U22570 (N_22570,N_21261,N_21326);
nor U22571 (N_22571,N_21837,N_21509);
nand U22572 (N_22572,N_21376,N_21090);
xnor U22573 (N_22573,N_21722,N_21732);
and U22574 (N_22574,N_21965,N_21812);
xor U22575 (N_22575,N_21694,N_21530);
xor U22576 (N_22576,N_21200,N_21976);
xnor U22577 (N_22577,N_21977,N_21299);
nand U22578 (N_22578,N_21273,N_21435);
or U22579 (N_22579,N_21431,N_21333);
xnor U22580 (N_22580,N_21996,N_21741);
xor U22581 (N_22581,N_21832,N_21825);
nor U22582 (N_22582,N_21120,N_21481);
nor U22583 (N_22583,N_21699,N_21537);
nor U22584 (N_22584,N_21543,N_21328);
and U22585 (N_22585,N_21113,N_21879);
xnor U22586 (N_22586,N_21612,N_21683);
xor U22587 (N_22587,N_21310,N_21082);
xor U22588 (N_22588,N_21472,N_21221);
nor U22589 (N_22589,N_21927,N_21386);
and U22590 (N_22590,N_21337,N_21731);
or U22591 (N_22591,N_21385,N_21402);
or U22592 (N_22592,N_21676,N_21869);
or U22593 (N_22593,N_21038,N_21924);
xnor U22594 (N_22594,N_21062,N_21387);
nand U22595 (N_22595,N_21565,N_21097);
xnor U22596 (N_22596,N_21603,N_21908);
or U22597 (N_22597,N_21535,N_21998);
and U22598 (N_22598,N_21253,N_21622);
nand U22599 (N_22599,N_21430,N_21740);
nor U22600 (N_22600,N_21562,N_21779);
nand U22601 (N_22601,N_21987,N_21079);
nor U22602 (N_22602,N_21121,N_21272);
and U22603 (N_22603,N_21782,N_21232);
and U22604 (N_22604,N_21842,N_21068);
xor U22605 (N_22605,N_21835,N_21858);
or U22606 (N_22606,N_21658,N_21962);
nand U22607 (N_22607,N_21203,N_21779);
and U22608 (N_22608,N_21637,N_21700);
or U22609 (N_22609,N_21142,N_21156);
xor U22610 (N_22610,N_21935,N_21415);
nor U22611 (N_22611,N_21294,N_21980);
xnor U22612 (N_22612,N_21124,N_21708);
xor U22613 (N_22613,N_21079,N_21820);
or U22614 (N_22614,N_21109,N_21321);
xnor U22615 (N_22615,N_21741,N_21924);
or U22616 (N_22616,N_21389,N_21723);
nand U22617 (N_22617,N_21288,N_21006);
and U22618 (N_22618,N_21133,N_21339);
and U22619 (N_22619,N_21919,N_21182);
and U22620 (N_22620,N_21144,N_21949);
or U22621 (N_22621,N_21997,N_21200);
nor U22622 (N_22622,N_21135,N_21414);
xnor U22623 (N_22623,N_21587,N_21483);
xor U22624 (N_22624,N_21530,N_21516);
nand U22625 (N_22625,N_21165,N_21924);
xor U22626 (N_22626,N_21434,N_21022);
or U22627 (N_22627,N_21686,N_21444);
xnor U22628 (N_22628,N_21163,N_21779);
nand U22629 (N_22629,N_21289,N_21742);
or U22630 (N_22630,N_21262,N_21774);
nor U22631 (N_22631,N_21165,N_21620);
nand U22632 (N_22632,N_21795,N_21140);
xor U22633 (N_22633,N_21379,N_21030);
and U22634 (N_22634,N_21952,N_21741);
nor U22635 (N_22635,N_21134,N_21254);
or U22636 (N_22636,N_21471,N_21716);
and U22637 (N_22637,N_21955,N_21541);
and U22638 (N_22638,N_21387,N_21781);
nand U22639 (N_22639,N_21152,N_21647);
nand U22640 (N_22640,N_21093,N_21912);
or U22641 (N_22641,N_21207,N_21316);
nor U22642 (N_22642,N_21131,N_21950);
nand U22643 (N_22643,N_21304,N_21031);
nand U22644 (N_22644,N_21655,N_21074);
and U22645 (N_22645,N_21176,N_21571);
nand U22646 (N_22646,N_21874,N_21217);
xor U22647 (N_22647,N_21642,N_21620);
xor U22648 (N_22648,N_21156,N_21638);
xor U22649 (N_22649,N_21279,N_21064);
nor U22650 (N_22650,N_21749,N_21268);
xnor U22651 (N_22651,N_21357,N_21367);
and U22652 (N_22652,N_21982,N_21777);
and U22653 (N_22653,N_21880,N_21791);
nand U22654 (N_22654,N_21302,N_21853);
or U22655 (N_22655,N_21692,N_21449);
nand U22656 (N_22656,N_21876,N_21971);
and U22657 (N_22657,N_21206,N_21356);
and U22658 (N_22658,N_21622,N_21063);
nand U22659 (N_22659,N_21330,N_21554);
or U22660 (N_22660,N_21457,N_21369);
xor U22661 (N_22661,N_21114,N_21343);
nand U22662 (N_22662,N_21202,N_21452);
or U22663 (N_22663,N_21398,N_21796);
nor U22664 (N_22664,N_21064,N_21937);
nand U22665 (N_22665,N_21193,N_21522);
nor U22666 (N_22666,N_21210,N_21851);
or U22667 (N_22667,N_21525,N_21098);
nor U22668 (N_22668,N_21904,N_21767);
xor U22669 (N_22669,N_21888,N_21214);
or U22670 (N_22670,N_21558,N_21665);
or U22671 (N_22671,N_21016,N_21139);
nor U22672 (N_22672,N_21738,N_21945);
nand U22673 (N_22673,N_21479,N_21573);
or U22674 (N_22674,N_21850,N_21240);
nand U22675 (N_22675,N_21275,N_21207);
or U22676 (N_22676,N_21905,N_21890);
and U22677 (N_22677,N_21239,N_21297);
nand U22678 (N_22678,N_21521,N_21395);
xnor U22679 (N_22679,N_21460,N_21924);
or U22680 (N_22680,N_21570,N_21388);
xnor U22681 (N_22681,N_21748,N_21092);
xnor U22682 (N_22682,N_21477,N_21729);
xnor U22683 (N_22683,N_21912,N_21664);
nor U22684 (N_22684,N_21863,N_21767);
or U22685 (N_22685,N_21309,N_21509);
or U22686 (N_22686,N_21855,N_21320);
xor U22687 (N_22687,N_21300,N_21322);
and U22688 (N_22688,N_21160,N_21785);
and U22689 (N_22689,N_21158,N_21080);
xor U22690 (N_22690,N_21033,N_21417);
nor U22691 (N_22691,N_21597,N_21881);
nand U22692 (N_22692,N_21925,N_21347);
nor U22693 (N_22693,N_21349,N_21610);
nor U22694 (N_22694,N_21400,N_21755);
and U22695 (N_22695,N_21428,N_21809);
nor U22696 (N_22696,N_21369,N_21588);
nand U22697 (N_22697,N_21714,N_21942);
and U22698 (N_22698,N_21647,N_21881);
xor U22699 (N_22699,N_21914,N_21396);
or U22700 (N_22700,N_21546,N_21937);
nor U22701 (N_22701,N_21823,N_21678);
nand U22702 (N_22702,N_21387,N_21678);
nor U22703 (N_22703,N_21845,N_21139);
or U22704 (N_22704,N_21336,N_21284);
nor U22705 (N_22705,N_21618,N_21939);
nor U22706 (N_22706,N_21197,N_21941);
or U22707 (N_22707,N_21474,N_21335);
nand U22708 (N_22708,N_21942,N_21718);
xor U22709 (N_22709,N_21531,N_21083);
nand U22710 (N_22710,N_21422,N_21108);
xor U22711 (N_22711,N_21964,N_21417);
nand U22712 (N_22712,N_21667,N_21223);
nor U22713 (N_22713,N_21711,N_21444);
and U22714 (N_22714,N_21717,N_21049);
or U22715 (N_22715,N_21037,N_21214);
and U22716 (N_22716,N_21594,N_21645);
xor U22717 (N_22717,N_21971,N_21246);
nor U22718 (N_22718,N_21137,N_21278);
nand U22719 (N_22719,N_21429,N_21229);
and U22720 (N_22720,N_21866,N_21542);
nor U22721 (N_22721,N_21983,N_21183);
nand U22722 (N_22722,N_21273,N_21105);
nand U22723 (N_22723,N_21944,N_21949);
and U22724 (N_22724,N_21774,N_21822);
xnor U22725 (N_22725,N_21150,N_21964);
and U22726 (N_22726,N_21861,N_21436);
xor U22727 (N_22727,N_21974,N_21141);
nand U22728 (N_22728,N_21427,N_21123);
and U22729 (N_22729,N_21917,N_21274);
nand U22730 (N_22730,N_21259,N_21654);
or U22731 (N_22731,N_21341,N_21335);
nand U22732 (N_22732,N_21393,N_21080);
xnor U22733 (N_22733,N_21749,N_21403);
nand U22734 (N_22734,N_21735,N_21881);
nor U22735 (N_22735,N_21542,N_21839);
nand U22736 (N_22736,N_21839,N_21575);
nor U22737 (N_22737,N_21337,N_21892);
nor U22738 (N_22738,N_21531,N_21184);
xnor U22739 (N_22739,N_21496,N_21614);
nor U22740 (N_22740,N_21185,N_21414);
nor U22741 (N_22741,N_21423,N_21561);
or U22742 (N_22742,N_21576,N_21874);
xor U22743 (N_22743,N_21161,N_21774);
xnor U22744 (N_22744,N_21110,N_21349);
nor U22745 (N_22745,N_21115,N_21277);
nor U22746 (N_22746,N_21677,N_21706);
and U22747 (N_22747,N_21294,N_21514);
nor U22748 (N_22748,N_21720,N_21362);
nand U22749 (N_22749,N_21326,N_21972);
or U22750 (N_22750,N_21028,N_21337);
nor U22751 (N_22751,N_21284,N_21271);
nor U22752 (N_22752,N_21965,N_21391);
nor U22753 (N_22753,N_21338,N_21692);
xnor U22754 (N_22754,N_21540,N_21246);
nor U22755 (N_22755,N_21709,N_21832);
and U22756 (N_22756,N_21341,N_21507);
nor U22757 (N_22757,N_21990,N_21321);
or U22758 (N_22758,N_21092,N_21386);
nand U22759 (N_22759,N_21609,N_21197);
nand U22760 (N_22760,N_21974,N_21815);
nand U22761 (N_22761,N_21050,N_21180);
or U22762 (N_22762,N_21619,N_21227);
xor U22763 (N_22763,N_21764,N_21115);
nand U22764 (N_22764,N_21887,N_21616);
xnor U22765 (N_22765,N_21164,N_21485);
or U22766 (N_22766,N_21125,N_21746);
xnor U22767 (N_22767,N_21869,N_21867);
and U22768 (N_22768,N_21660,N_21154);
xnor U22769 (N_22769,N_21332,N_21646);
nor U22770 (N_22770,N_21391,N_21705);
and U22771 (N_22771,N_21710,N_21365);
nor U22772 (N_22772,N_21772,N_21714);
nand U22773 (N_22773,N_21005,N_21514);
or U22774 (N_22774,N_21841,N_21386);
and U22775 (N_22775,N_21174,N_21232);
or U22776 (N_22776,N_21830,N_21605);
nand U22777 (N_22777,N_21732,N_21356);
xnor U22778 (N_22778,N_21633,N_21637);
or U22779 (N_22779,N_21911,N_21449);
or U22780 (N_22780,N_21828,N_21380);
nand U22781 (N_22781,N_21793,N_21199);
nand U22782 (N_22782,N_21045,N_21655);
nand U22783 (N_22783,N_21966,N_21285);
nor U22784 (N_22784,N_21770,N_21075);
nand U22785 (N_22785,N_21836,N_21548);
or U22786 (N_22786,N_21196,N_21608);
nand U22787 (N_22787,N_21182,N_21729);
nor U22788 (N_22788,N_21669,N_21577);
nand U22789 (N_22789,N_21157,N_21996);
nor U22790 (N_22790,N_21188,N_21644);
nand U22791 (N_22791,N_21632,N_21211);
nand U22792 (N_22792,N_21046,N_21802);
xnor U22793 (N_22793,N_21074,N_21717);
nor U22794 (N_22794,N_21013,N_21925);
nand U22795 (N_22795,N_21501,N_21640);
or U22796 (N_22796,N_21076,N_21738);
nand U22797 (N_22797,N_21481,N_21421);
nor U22798 (N_22798,N_21917,N_21241);
and U22799 (N_22799,N_21308,N_21204);
xnor U22800 (N_22800,N_21900,N_21750);
nor U22801 (N_22801,N_21138,N_21051);
xnor U22802 (N_22802,N_21338,N_21667);
or U22803 (N_22803,N_21521,N_21316);
and U22804 (N_22804,N_21605,N_21562);
nand U22805 (N_22805,N_21991,N_21085);
nand U22806 (N_22806,N_21727,N_21582);
xor U22807 (N_22807,N_21010,N_21355);
or U22808 (N_22808,N_21051,N_21287);
and U22809 (N_22809,N_21954,N_21753);
nand U22810 (N_22810,N_21699,N_21070);
and U22811 (N_22811,N_21093,N_21256);
nor U22812 (N_22812,N_21926,N_21453);
xnor U22813 (N_22813,N_21108,N_21657);
or U22814 (N_22814,N_21136,N_21099);
or U22815 (N_22815,N_21637,N_21264);
nor U22816 (N_22816,N_21490,N_21702);
nor U22817 (N_22817,N_21610,N_21312);
nand U22818 (N_22818,N_21980,N_21329);
or U22819 (N_22819,N_21839,N_21303);
nor U22820 (N_22820,N_21987,N_21478);
nand U22821 (N_22821,N_21454,N_21103);
xnor U22822 (N_22822,N_21316,N_21949);
nand U22823 (N_22823,N_21969,N_21158);
nor U22824 (N_22824,N_21897,N_21301);
xor U22825 (N_22825,N_21581,N_21327);
nand U22826 (N_22826,N_21838,N_21921);
xor U22827 (N_22827,N_21579,N_21038);
xor U22828 (N_22828,N_21317,N_21659);
nand U22829 (N_22829,N_21166,N_21924);
or U22830 (N_22830,N_21860,N_21449);
nor U22831 (N_22831,N_21875,N_21071);
and U22832 (N_22832,N_21850,N_21465);
and U22833 (N_22833,N_21039,N_21277);
nand U22834 (N_22834,N_21393,N_21710);
and U22835 (N_22835,N_21252,N_21489);
nand U22836 (N_22836,N_21195,N_21945);
xor U22837 (N_22837,N_21237,N_21664);
xnor U22838 (N_22838,N_21818,N_21645);
xnor U22839 (N_22839,N_21237,N_21308);
and U22840 (N_22840,N_21387,N_21487);
and U22841 (N_22841,N_21746,N_21496);
and U22842 (N_22842,N_21371,N_21145);
or U22843 (N_22843,N_21800,N_21013);
xnor U22844 (N_22844,N_21968,N_21549);
and U22845 (N_22845,N_21298,N_21805);
xnor U22846 (N_22846,N_21741,N_21440);
nand U22847 (N_22847,N_21406,N_21850);
nand U22848 (N_22848,N_21860,N_21206);
nand U22849 (N_22849,N_21219,N_21315);
xor U22850 (N_22850,N_21329,N_21725);
nor U22851 (N_22851,N_21962,N_21363);
xnor U22852 (N_22852,N_21128,N_21176);
and U22853 (N_22853,N_21557,N_21162);
nor U22854 (N_22854,N_21250,N_21523);
nand U22855 (N_22855,N_21654,N_21683);
nand U22856 (N_22856,N_21405,N_21173);
and U22857 (N_22857,N_21684,N_21424);
xor U22858 (N_22858,N_21280,N_21428);
xor U22859 (N_22859,N_21726,N_21233);
nor U22860 (N_22860,N_21536,N_21042);
nor U22861 (N_22861,N_21916,N_21986);
nor U22862 (N_22862,N_21461,N_21710);
and U22863 (N_22863,N_21003,N_21692);
nand U22864 (N_22864,N_21722,N_21436);
nor U22865 (N_22865,N_21330,N_21703);
xnor U22866 (N_22866,N_21228,N_21870);
or U22867 (N_22867,N_21300,N_21436);
nand U22868 (N_22868,N_21166,N_21509);
and U22869 (N_22869,N_21092,N_21871);
or U22870 (N_22870,N_21720,N_21022);
xor U22871 (N_22871,N_21323,N_21084);
or U22872 (N_22872,N_21597,N_21579);
nor U22873 (N_22873,N_21905,N_21210);
nor U22874 (N_22874,N_21602,N_21218);
xor U22875 (N_22875,N_21046,N_21827);
xor U22876 (N_22876,N_21311,N_21355);
nor U22877 (N_22877,N_21091,N_21199);
nor U22878 (N_22878,N_21475,N_21026);
and U22879 (N_22879,N_21367,N_21086);
or U22880 (N_22880,N_21985,N_21710);
xnor U22881 (N_22881,N_21010,N_21425);
nand U22882 (N_22882,N_21410,N_21462);
and U22883 (N_22883,N_21419,N_21370);
and U22884 (N_22884,N_21984,N_21418);
and U22885 (N_22885,N_21509,N_21113);
or U22886 (N_22886,N_21852,N_21450);
nor U22887 (N_22887,N_21479,N_21320);
or U22888 (N_22888,N_21405,N_21204);
xnor U22889 (N_22889,N_21530,N_21687);
nor U22890 (N_22890,N_21556,N_21992);
nand U22891 (N_22891,N_21767,N_21759);
or U22892 (N_22892,N_21207,N_21441);
or U22893 (N_22893,N_21077,N_21616);
nor U22894 (N_22894,N_21205,N_21317);
nor U22895 (N_22895,N_21432,N_21409);
nand U22896 (N_22896,N_21489,N_21976);
nor U22897 (N_22897,N_21602,N_21636);
xor U22898 (N_22898,N_21041,N_21229);
nand U22899 (N_22899,N_21693,N_21667);
and U22900 (N_22900,N_21201,N_21088);
and U22901 (N_22901,N_21276,N_21934);
nor U22902 (N_22902,N_21823,N_21014);
nand U22903 (N_22903,N_21668,N_21979);
and U22904 (N_22904,N_21120,N_21526);
nand U22905 (N_22905,N_21370,N_21123);
or U22906 (N_22906,N_21428,N_21822);
or U22907 (N_22907,N_21764,N_21464);
nor U22908 (N_22908,N_21186,N_21792);
and U22909 (N_22909,N_21323,N_21245);
and U22910 (N_22910,N_21281,N_21779);
nand U22911 (N_22911,N_21370,N_21237);
or U22912 (N_22912,N_21068,N_21891);
and U22913 (N_22913,N_21768,N_21080);
nand U22914 (N_22914,N_21847,N_21366);
or U22915 (N_22915,N_21663,N_21138);
xor U22916 (N_22916,N_21932,N_21985);
or U22917 (N_22917,N_21651,N_21313);
and U22918 (N_22918,N_21212,N_21915);
or U22919 (N_22919,N_21683,N_21071);
and U22920 (N_22920,N_21312,N_21662);
nor U22921 (N_22921,N_21434,N_21170);
nand U22922 (N_22922,N_21275,N_21416);
nand U22923 (N_22923,N_21951,N_21359);
and U22924 (N_22924,N_21322,N_21144);
nand U22925 (N_22925,N_21217,N_21087);
xnor U22926 (N_22926,N_21500,N_21865);
or U22927 (N_22927,N_21704,N_21403);
nor U22928 (N_22928,N_21012,N_21278);
nand U22929 (N_22929,N_21160,N_21987);
or U22930 (N_22930,N_21038,N_21092);
xnor U22931 (N_22931,N_21735,N_21958);
or U22932 (N_22932,N_21955,N_21742);
nor U22933 (N_22933,N_21557,N_21934);
or U22934 (N_22934,N_21865,N_21032);
nand U22935 (N_22935,N_21677,N_21200);
nor U22936 (N_22936,N_21076,N_21523);
xor U22937 (N_22937,N_21743,N_21961);
xor U22938 (N_22938,N_21974,N_21956);
nand U22939 (N_22939,N_21747,N_21045);
nand U22940 (N_22940,N_21545,N_21066);
xnor U22941 (N_22941,N_21643,N_21739);
xor U22942 (N_22942,N_21352,N_21491);
nand U22943 (N_22943,N_21948,N_21491);
nor U22944 (N_22944,N_21619,N_21205);
nand U22945 (N_22945,N_21640,N_21172);
and U22946 (N_22946,N_21335,N_21087);
nand U22947 (N_22947,N_21309,N_21921);
and U22948 (N_22948,N_21536,N_21916);
xnor U22949 (N_22949,N_21702,N_21654);
or U22950 (N_22950,N_21980,N_21798);
nand U22951 (N_22951,N_21162,N_21048);
nand U22952 (N_22952,N_21422,N_21051);
nand U22953 (N_22953,N_21732,N_21429);
or U22954 (N_22954,N_21791,N_21360);
or U22955 (N_22955,N_21156,N_21778);
xor U22956 (N_22956,N_21769,N_21466);
xnor U22957 (N_22957,N_21375,N_21218);
or U22958 (N_22958,N_21723,N_21103);
or U22959 (N_22959,N_21735,N_21926);
or U22960 (N_22960,N_21514,N_21859);
or U22961 (N_22961,N_21047,N_21804);
xor U22962 (N_22962,N_21106,N_21605);
xor U22963 (N_22963,N_21460,N_21849);
nor U22964 (N_22964,N_21504,N_21175);
nor U22965 (N_22965,N_21082,N_21481);
nor U22966 (N_22966,N_21122,N_21934);
nand U22967 (N_22967,N_21583,N_21541);
xor U22968 (N_22968,N_21025,N_21004);
and U22969 (N_22969,N_21257,N_21088);
and U22970 (N_22970,N_21304,N_21148);
and U22971 (N_22971,N_21856,N_21659);
nand U22972 (N_22972,N_21899,N_21845);
or U22973 (N_22973,N_21812,N_21622);
nand U22974 (N_22974,N_21265,N_21396);
nor U22975 (N_22975,N_21927,N_21731);
xor U22976 (N_22976,N_21041,N_21040);
nand U22977 (N_22977,N_21066,N_21945);
and U22978 (N_22978,N_21775,N_21978);
or U22979 (N_22979,N_21749,N_21173);
or U22980 (N_22980,N_21649,N_21963);
and U22981 (N_22981,N_21018,N_21905);
nor U22982 (N_22982,N_21936,N_21721);
and U22983 (N_22983,N_21216,N_21069);
nor U22984 (N_22984,N_21455,N_21993);
xnor U22985 (N_22985,N_21509,N_21905);
and U22986 (N_22986,N_21939,N_21383);
xnor U22987 (N_22987,N_21024,N_21992);
and U22988 (N_22988,N_21656,N_21545);
xor U22989 (N_22989,N_21565,N_21449);
nor U22990 (N_22990,N_21066,N_21891);
or U22991 (N_22991,N_21732,N_21807);
nor U22992 (N_22992,N_21150,N_21326);
or U22993 (N_22993,N_21632,N_21747);
nand U22994 (N_22994,N_21519,N_21880);
and U22995 (N_22995,N_21427,N_21862);
xor U22996 (N_22996,N_21896,N_21770);
or U22997 (N_22997,N_21175,N_21118);
nand U22998 (N_22998,N_21942,N_21723);
or U22999 (N_22999,N_21752,N_21223);
or U23000 (N_23000,N_22599,N_22969);
or U23001 (N_23001,N_22267,N_22815);
nand U23002 (N_23002,N_22806,N_22503);
nand U23003 (N_23003,N_22122,N_22347);
or U23004 (N_23004,N_22209,N_22318);
nor U23005 (N_23005,N_22457,N_22178);
nor U23006 (N_23006,N_22295,N_22970);
or U23007 (N_23007,N_22140,N_22587);
nand U23008 (N_23008,N_22926,N_22066);
and U23009 (N_23009,N_22842,N_22498);
xor U23010 (N_23010,N_22586,N_22026);
or U23011 (N_23011,N_22488,N_22365);
xor U23012 (N_23012,N_22594,N_22652);
nor U23013 (N_23013,N_22024,N_22975);
nand U23014 (N_23014,N_22808,N_22007);
xor U23015 (N_23015,N_22037,N_22568);
and U23016 (N_23016,N_22034,N_22962);
nand U23017 (N_23017,N_22788,N_22293);
or U23018 (N_23018,N_22598,N_22524);
nand U23019 (N_23019,N_22288,N_22383);
and U23020 (N_23020,N_22338,N_22069);
nand U23021 (N_23021,N_22637,N_22520);
xnor U23022 (N_23022,N_22054,N_22106);
xor U23023 (N_23023,N_22933,N_22690);
nor U23024 (N_23024,N_22636,N_22857);
nand U23025 (N_23025,N_22978,N_22455);
or U23026 (N_23026,N_22574,N_22584);
or U23027 (N_23027,N_22811,N_22805);
nand U23028 (N_23028,N_22150,N_22307);
nor U23029 (N_23029,N_22084,N_22005);
nor U23030 (N_23030,N_22166,N_22740);
or U23031 (N_23031,N_22316,N_22127);
and U23032 (N_23032,N_22987,N_22360);
and U23033 (N_23033,N_22146,N_22532);
nand U23034 (N_23034,N_22905,N_22554);
and U23035 (N_23035,N_22137,N_22816);
xor U23036 (N_23036,N_22050,N_22278);
nand U23037 (N_23037,N_22612,N_22351);
nand U23038 (N_23038,N_22979,N_22733);
nand U23039 (N_23039,N_22666,N_22681);
nor U23040 (N_23040,N_22180,N_22063);
or U23041 (N_23041,N_22653,N_22971);
or U23042 (N_23042,N_22371,N_22775);
or U23043 (N_23043,N_22530,N_22849);
nor U23044 (N_23044,N_22792,N_22261);
nand U23045 (N_23045,N_22560,N_22623);
nand U23046 (N_23046,N_22280,N_22044);
or U23047 (N_23047,N_22443,N_22853);
xor U23048 (N_23048,N_22947,N_22534);
nand U23049 (N_23049,N_22829,N_22107);
nor U23050 (N_23050,N_22302,N_22262);
xnor U23051 (N_23051,N_22898,N_22450);
nor U23052 (N_23052,N_22670,N_22985);
nor U23053 (N_23053,N_22296,N_22257);
nand U23054 (N_23054,N_22441,N_22750);
nor U23055 (N_23055,N_22776,N_22650);
nand U23056 (N_23056,N_22566,N_22613);
and U23057 (N_23057,N_22895,N_22770);
or U23058 (N_23058,N_22115,N_22845);
and U23059 (N_23059,N_22203,N_22921);
nand U23060 (N_23060,N_22188,N_22284);
or U23061 (N_23061,N_22513,N_22606);
nor U23062 (N_23062,N_22839,N_22361);
nor U23063 (N_23063,N_22630,N_22263);
and U23064 (N_23064,N_22832,N_22247);
or U23065 (N_23065,N_22350,N_22795);
or U23066 (N_23066,N_22927,N_22105);
or U23067 (N_23067,N_22710,N_22780);
and U23068 (N_23068,N_22675,N_22592);
xnor U23069 (N_23069,N_22642,N_22936);
nand U23070 (N_23070,N_22499,N_22241);
and U23071 (N_23071,N_22693,N_22285);
and U23072 (N_23072,N_22470,N_22382);
and U23073 (N_23073,N_22010,N_22569);
or U23074 (N_23074,N_22860,N_22194);
nand U23075 (N_23075,N_22438,N_22425);
and U23076 (N_23076,N_22237,N_22268);
nor U23077 (N_23077,N_22583,N_22892);
xnor U23078 (N_23078,N_22659,N_22414);
nor U23079 (N_23079,N_22939,N_22030);
or U23080 (N_23080,N_22781,N_22689);
nor U23081 (N_23081,N_22992,N_22250);
xor U23082 (N_23082,N_22923,N_22447);
and U23083 (N_23083,N_22144,N_22461);
nand U23084 (N_23084,N_22607,N_22121);
or U23085 (N_23085,N_22761,N_22528);
or U23086 (N_23086,N_22784,N_22516);
xnor U23087 (N_23087,N_22326,N_22621);
nor U23088 (N_23088,N_22960,N_22311);
xnor U23089 (N_23089,N_22673,N_22315);
xor U23090 (N_23090,N_22549,N_22877);
or U23091 (N_23091,N_22133,N_22785);
and U23092 (N_23092,N_22373,N_22899);
and U23093 (N_23093,N_22334,N_22935);
or U23094 (N_23094,N_22094,N_22605);
nand U23095 (N_23095,N_22906,N_22109);
or U23096 (N_23096,N_22230,N_22712);
and U23097 (N_23097,N_22938,N_22075);
nor U23098 (N_23098,N_22492,N_22511);
nand U23099 (N_23099,N_22497,N_22369);
xnor U23100 (N_23100,N_22682,N_22798);
and U23101 (N_23101,N_22844,N_22787);
nand U23102 (N_23102,N_22852,N_22240);
and U23103 (N_23103,N_22897,N_22793);
and U23104 (N_23104,N_22234,N_22125);
nor U23105 (N_23105,N_22378,N_22778);
or U23106 (N_23106,N_22223,N_22872);
and U23107 (N_23107,N_22381,N_22277);
xor U23108 (N_23108,N_22996,N_22032);
xnor U23109 (N_23109,N_22177,N_22449);
or U23110 (N_23110,N_22191,N_22977);
xnor U23111 (N_23111,N_22972,N_22081);
nand U23112 (N_23112,N_22635,N_22523);
and U23113 (N_23113,N_22655,N_22271);
nand U23114 (N_23114,N_22796,N_22922);
or U23115 (N_23115,N_22840,N_22973);
xor U23116 (N_23116,N_22102,N_22462);
nor U23117 (N_23117,N_22739,N_22819);
nor U23118 (N_23118,N_22423,N_22402);
or U23119 (N_23119,N_22256,N_22998);
nand U23120 (N_23120,N_22370,N_22465);
and U23121 (N_23121,N_22981,N_22494);
xnor U23122 (N_23122,N_22814,N_22559);
xnor U23123 (N_23123,N_22611,N_22843);
nand U23124 (N_23124,N_22184,N_22907);
and U23125 (N_23125,N_22061,N_22476);
nor U23126 (N_23126,N_22343,N_22570);
xnor U23127 (N_23127,N_22940,N_22397);
xor U23128 (N_23128,N_22664,N_22353);
nand U23129 (N_23129,N_22047,N_22158);
or U23130 (N_23130,N_22841,N_22167);
and U23131 (N_23131,N_22432,N_22509);
or U23132 (N_23132,N_22722,N_22442);
and U23133 (N_23133,N_22189,N_22434);
and U23134 (N_23134,N_22640,N_22580);
nor U23135 (N_23135,N_22747,N_22968);
or U23136 (N_23136,N_22110,N_22751);
nand U23137 (N_23137,N_22415,N_22638);
xor U23138 (N_23138,N_22164,N_22916);
nand U23139 (N_23139,N_22573,N_22013);
nand U23140 (N_23140,N_22298,N_22401);
nand U23141 (N_23141,N_22526,N_22108);
nor U23142 (N_23142,N_22802,N_22555);
xor U23143 (N_23143,N_22471,N_22038);
and U23144 (N_23144,N_22252,N_22826);
nand U23145 (N_23145,N_22505,N_22345);
and U23146 (N_23146,N_22019,N_22474);
and U23147 (N_23147,N_22201,N_22965);
xnor U23148 (N_23148,N_22327,N_22136);
xnor U23149 (N_23149,N_22961,N_22305);
and U23150 (N_23150,N_22764,N_22768);
nor U23151 (N_23151,N_22290,N_22422);
nand U23152 (N_23152,N_22325,N_22260);
or U23153 (N_23153,N_22012,N_22887);
or U23154 (N_23154,N_22858,N_22909);
nand U23155 (N_23155,N_22138,N_22394);
or U23156 (N_23156,N_22301,N_22046);
nand U23157 (N_23157,N_22027,N_22088);
xor U23158 (N_23158,N_22654,N_22595);
nand U23159 (N_23159,N_22691,N_22582);
xor U23160 (N_23160,N_22219,N_22779);
nand U23161 (N_23161,N_22911,N_22855);
xnor U23162 (N_23162,N_22539,N_22868);
and U23163 (N_23163,N_22067,N_22479);
xor U23164 (N_23164,N_22195,N_22745);
xnor U23165 (N_23165,N_22702,N_22453);
nand U23166 (N_23166,N_22258,N_22604);
nand U23167 (N_23167,N_22649,N_22152);
nand U23168 (N_23168,N_22056,N_22091);
or U23169 (N_23169,N_22428,N_22215);
nand U23170 (N_23170,N_22255,N_22648);
or U23171 (N_23171,N_22339,N_22163);
and U23172 (N_23172,N_22071,N_22807);
nand U23173 (N_23173,N_22454,N_22708);
nand U23174 (N_23174,N_22797,N_22873);
and U23175 (N_23175,N_22221,N_22727);
and U23176 (N_23176,N_22342,N_22487);
or U23177 (N_23177,N_22048,N_22344);
and U23178 (N_23178,N_22082,N_22542);
xor U23179 (N_23179,N_22641,N_22329);
xnor U23180 (N_23180,N_22856,N_22292);
nand U23181 (N_23181,N_22002,N_22510);
nor U23182 (N_23182,N_22726,N_22874);
nand U23183 (N_23183,N_22896,N_22132);
nor U23184 (N_23184,N_22435,N_22309);
and U23185 (N_23185,N_22571,N_22009);
xnor U23186 (N_23186,N_22974,N_22810);
and U23187 (N_23187,N_22244,N_22190);
nand U23188 (N_23188,N_22155,N_22676);
xnor U23189 (N_23189,N_22362,N_22943);
or U23190 (N_23190,N_22060,N_22229);
and U23191 (N_23191,N_22495,N_22116);
nor U23192 (N_23192,N_22424,N_22303);
and U23193 (N_23193,N_22162,N_22882);
nand U23194 (N_23194,N_22375,N_22953);
nand U23195 (N_23195,N_22838,N_22399);
xnor U23196 (N_23196,N_22986,N_22589);
or U23197 (N_23197,N_22512,N_22291);
xnor U23198 (N_23198,N_22161,N_22608);
nand U23199 (N_23199,N_22719,N_22870);
nor U23200 (N_23200,N_22165,N_22556);
or U23201 (N_23201,N_22021,N_22614);
and U23202 (N_23202,N_22945,N_22593);
xnor U23203 (N_23203,N_22813,N_22072);
xor U23204 (N_23204,N_22772,N_22439);
nor U23205 (N_23205,N_22557,N_22426);
nand U23206 (N_23206,N_22590,N_22491);
or U23207 (N_23207,N_22039,N_22828);
xnor U23208 (N_23208,N_22192,N_22801);
nor U23209 (N_23209,N_22738,N_22119);
and U23210 (N_23210,N_22395,N_22224);
and U23211 (N_23211,N_22774,N_22579);
and U23212 (N_23212,N_22893,N_22323);
nor U23213 (N_23213,N_22762,N_22728);
and U23214 (N_23214,N_22396,N_22276);
nand U23215 (N_23215,N_22736,N_22118);
or U23216 (N_23216,N_22660,N_22226);
nor U23217 (N_23217,N_22760,N_22620);
and U23218 (N_23218,N_22235,N_22550);
nand U23219 (N_23219,N_22332,N_22651);
xor U23220 (N_23220,N_22238,N_22865);
and U23221 (N_23221,N_22924,N_22742);
nand U23222 (N_23222,N_22861,N_22427);
xor U23223 (N_23223,N_22357,N_22767);
and U23224 (N_23224,N_22942,N_22758);
and U23225 (N_23225,N_22891,N_22051);
nor U23226 (N_23226,N_22634,N_22212);
and U23227 (N_23227,N_22954,N_22233);
nor U23228 (N_23228,N_22912,N_22662);
xnor U23229 (N_23229,N_22576,N_22251);
nor U23230 (N_23230,N_22880,N_22701);
and U23231 (N_23231,N_22830,N_22359);
or U23232 (N_23232,N_22320,N_22446);
or U23233 (N_23233,N_22486,N_22884);
nand U23234 (N_23234,N_22416,N_22929);
xor U23235 (N_23235,N_22430,N_22076);
nor U23236 (N_23236,N_22404,N_22444);
nor U23237 (N_23237,N_22078,N_22473);
or U23238 (N_23238,N_22312,N_22777);
xnor U23239 (N_23239,N_22931,N_22406);
and U23240 (N_23240,N_22354,N_22259);
nor U23241 (N_23241,N_22506,N_22817);
xnor U23242 (N_23242,N_22988,N_22367);
nand U23243 (N_23243,N_22757,N_22065);
nor U23244 (N_23244,N_22948,N_22324);
nor U23245 (N_23245,N_22544,N_22688);
nand U23246 (N_23246,N_22862,N_22368);
nand U23247 (N_23247,N_22588,N_22677);
or U23248 (N_23248,N_22680,N_22147);
or U23249 (N_23249,N_22716,N_22964);
nand U23250 (N_23250,N_22322,N_22099);
nand U23251 (N_23251,N_22086,N_22419);
nand U23252 (N_23252,N_22304,N_22403);
nor U23253 (N_23253,N_22848,N_22040);
or U23254 (N_23254,N_22448,N_22095);
xnor U23255 (N_23255,N_22308,N_22143);
nand U23256 (N_23256,N_22098,N_22431);
and U23257 (N_23257,N_22643,N_22794);
xor U23258 (N_23258,N_22199,N_22822);
xnor U23259 (N_23259,N_22313,N_22626);
xor U23260 (N_23260,N_22142,N_22522);
xor U23261 (N_23261,N_22881,N_22270);
xor U23262 (N_23262,N_22265,N_22213);
or U23263 (N_23263,N_22668,N_22068);
and U23264 (N_23264,N_22658,N_22545);
nand U23265 (N_23265,N_22889,N_22390);
nor U23266 (N_23266,N_22467,N_22043);
and U23267 (N_23267,N_22991,N_22591);
and U23268 (N_23268,N_22341,N_22692);
and U23269 (N_23269,N_22031,N_22173);
xor U23270 (N_23270,N_22851,N_22011);
nor U23271 (N_23271,N_22440,N_22731);
xor U23272 (N_23272,N_22997,N_22236);
nor U23273 (N_23273,N_22124,N_22741);
nand U23274 (N_23274,N_22617,N_22782);
xor U23275 (N_23275,N_22346,N_22602);
or U23276 (N_23276,N_22123,N_22686);
and U23277 (N_23277,N_22279,N_22956);
or U23278 (N_23278,N_22976,N_22243);
nor U23279 (N_23279,N_22249,N_22466);
or U23280 (N_23280,N_22958,N_22624);
xnor U23281 (N_23281,N_22765,N_22160);
and U23282 (N_23282,N_22533,N_22321);
xnor U23283 (N_23283,N_22200,N_22697);
xor U23284 (N_23284,N_22477,N_22663);
nor U23285 (N_23285,N_22661,N_22734);
nand U23286 (N_23286,N_22883,N_22041);
and U23287 (N_23287,N_22600,N_22913);
nor U23288 (N_23288,N_22218,N_22149);
and U23289 (N_23289,N_22274,N_22714);
nor U23290 (N_23290,N_22696,N_22101);
xnor U23291 (N_23291,N_22205,N_22482);
nor U23292 (N_23292,N_22633,N_22168);
or U23293 (N_23293,N_22748,N_22536);
nand U23294 (N_23294,N_22951,N_22789);
or U23295 (N_23295,N_22493,N_22578);
nor U23296 (N_23296,N_22452,N_22863);
nor U23297 (N_23297,N_22331,N_22306);
and U23298 (N_23298,N_22089,N_22480);
xnor U23299 (N_23299,N_22104,N_22299);
nor U23300 (N_23300,N_22871,N_22206);
nand U23301 (N_23301,N_22057,N_22103);
or U23302 (N_23302,N_22483,N_22337);
xor U23303 (N_23303,N_22721,N_22087);
xor U23304 (N_23304,N_22363,N_22210);
xnor U23305 (N_23305,N_22092,N_22340);
nand U23306 (N_23306,N_22159,N_22097);
nand U23307 (N_23307,N_22847,N_22821);
nor U23308 (N_23308,N_22335,N_22366);
and U23309 (N_23309,N_22902,N_22080);
nand U23310 (N_23310,N_22558,N_22372);
and U23311 (N_23311,N_22894,N_22131);
xnor U23312 (N_23312,N_22625,N_22699);
xnor U23313 (N_23313,N_22328,N_22272);
nand U23314 (N_23314,N_22193,N_22410);
nand U23315 (N_23315,N_22672,N_22198);
nor U23316 (N_23316,N_22242,N_22083);
or U23317 (N_23317,N_22752,N_22478);
nand U23318 (N_23318,N_22197,N_22695);
xnor U23319 (N_23319,N_22629,N_22148);
or U23320 (N_23320,N_22903,N_22684);
or U23321 (N_23321,N_22910,N_22900);
nor U23322 (N_23322,N_22538,N_22531);
and U23323 (N_23323,N_22786,N_22245);
and U23324 (N_23324,N_22398,N_22561);
and U23325 (N_23325,N_22800,N_22100);
or U23326 (N_23326,N_22489,N_22836);
and U23327 (N_23327,N_22529,N_22824);
nor U23328 (N_23328,N_22519,N_22317);
and U23329 (N_23329,N_22518,N_22207);
nor U23330 (N_23330,N_22723,N_22639);
or U23331 (N_23331,N_22172,N_22707);
nor U23332 (N_23332,N_22886,N_22827);
and U23333 (N_23333,N_22451,N_22385);
nand U23334 (N_23334,N_22955,N_22820);
xor U23335 (N_23335,N_22790,N_22475);
nand U23336 (N_23336,N_22227,N_22185);
nand U23337 (N_23337,N_22049,N_22963);
and U23338 (N_23338,N_22349,N_22387);
or U23339 (N_23339,N_22959,N_22901);
and U23340 (N_23340,N_22281,N_22720);
xnor U23341 (N_23341,N_22551,N_22208);
xor U23342 (N_23342,N_22273,N_22804);
nand U23343 (N_23343,N_22564,N_22458);
nand U23344 (N_23344,N_22269,N_22437);
and U23345 (N_23345,N_22704,N_22181);
and U23346 (N_23346,N_22756,N_22846);
nand U23347 (N_23347,N_22202,N_22391);
and U23348 (N_23348,N_22709,N_22074);
and U23349 (N_23349,N_22597,N_22217);
or U23350 (N_23350,N_22114,N_22490);
nand U23351 (N_23351,N_22003,N_22145);
xor U23352 (N_23352,N_22888,N_22264);
xnor U23353 (N_23353,N_22156,N_22525);
and U23354 (N_23354,N_22412,N_22380);
xnor U23355 (N_23355,N_22941,N_22755);
or U23356 (N_23356,N_22552,N_22139);
nand U23357 (N_23357,N_22171,N_22678);
xnor U23358 (N_23358,N_22055,N_22175);
nor U23359 (N_23359,N_22388,N_22799);
nand U23360 (N_23360,N_22484,N_22500);
xnor U23361 (N_23361,N_22096,N_22336);
or U23362 (N_23362,N_22685,N_22456);
nor U23363 (N_23363,N_22854,N_22508);
nor U23364 (N_23364,N_22015,N_22045);
xnor U23365 (N_23365,N_22129,N_22222);
nor U23366 (N_23366,N_22646,N_22698);
nor U23367 (N_23367,N_22502,N_22632);
and U23368 (N_23368,N_22562,N_22433);
xnor U23369 (N_23369,N_22254,N_22718);
and U23370 (N_23370,N_22875,N_22117);
and U23371 (N_23371,N_22950,N_22683);
or U23372 (N_23372,N_22581,N_22090);
nand U23373 (N_23373,N_22348,N_22966);
nand U23374 (N_23374,N_22364,N_22610);
nor U23375 (N_23375,N_22429,N_22377);
xnor U23376 (N_23376,N_22501,N_22812);
and U23377 (N_23377,N_22724,N_22017);
xnor U23378 (N_23378,N_22737,N_22266);
nor U23379 (N_23379,N_22409,N_22535);
and U23380 (N_23380,N_22521,N_22990);
nand U23381 (N_23381,N_22379,N_22547);
or U23382 (N_23382,N_22994,N_22713);
xor U23383 (N_23383,N_22211,N_22983);
nand U23384 (N_23384,N_22711,N_22537);
nor U23385 (N_23385,N_22232,N_22619);
xor U23386 (N_23386,N_22062,N_22374);
nand U23387 (N_23387,N_22384,N_22674);
and U23388 (N_23388,N_22400,N_22603);
nand U23389 (N_23389,N_22036,N_22743);
xor U23390 (N_23390,N_22485,N_22999);
or U23391 (N_23391,N_22514,N_22572);
nand U23392 (N_23392,N_22920,N_22179);
nor U23393 (N_23393,N_22980,N_22628);
nor U23394 (N_23394,N_22546,N_22809);
nand U23395 (N_23395,N_22176,N_22783);
nand U23396 (N_23396,N_22064,N_22667);
nor U23397 (N_23397,N_22818,N_22463);
or U23398 (N_23398,N_22831,N_22216);
xor U23399 (N_23399,N_22744,N_22878);
nor U23400 (N_23400,N_22700,N_22004);
xnor U23401 (N_23401,N_22042,N_22228);
and U23402 (N_23402,N_22481,N_22869);
nor U23403 (N_23403,N_22282,N_22957);
nor U23404 (N_23404,N_22715,N_22093);
nor U23405 (N_23405,N_22355,N_22058);
xnor U23406 (N_23406,N_22705,N_22914);
or U23407 (N_23407,N_22527,N_22294);
or U23408 (N_23408,N_22771,N_22053);
or U23409 (N_23409,N_22928,N_22890);
nor U23410 (N_23410,N_22248,N_22763);
nand U23411 (N_23411,N_22864,N_22615);
nor U23412 (N_23412,N_22085,N_22746);
or U23413 (N_23413,N_22436,N_22930);
nor U23414 (N_23414,N_22174,N_22006);
and U23415 (N_23415,N_22669,N_22286);
nor U23416 (N_23416,N_22445,N_22472);
and U23417 (N_23417,N_22001,N_22879);
nor U23418 (N_23418,N_22949,N_22706);
and U23419 (N_23419,N_22885,N_22128);
nor U23420 (N_23420,N_22239,N_22644);
and U23421 (N_23421,N_22833,N_22022);
nand U23422 (N_23422,N_22314,N_22952);
xnor U23423 (N_23423,N_22297,N_22029);
and U23424 (N_23424,N_22919,N_22850);
xor U23425 (N_23425,N_22386,N_22729);
or U23426 (N_23426,N_22154,N_22289);
xnor U23427 (N_23427,N_22946,N_22565);
nor U23428 (N_23428,N_22577,N_22008);
or U23429 (N_23429,N_22464,N_22754);
nand U23430 (N_23430,N_22609,N_22627);
xnor U23431 (N_23431,N_22420,N_22287);
and U23432 (N_23432,N_22730,N_22915);
or U23433 (N_23433,N_22204,N_22111);
or U23434 (N_23434,N_22225,N_22393);
nor U23435 (N_23435,N_22407,N_22866);
nor U23436 (N_23436,N_22246,N_22169);
or U23437 (N_23437,N_22967,N_22504);
and U23438 (N_23438,N_22214,N_22126);
xor U23439 (N_23439,N_22141,N_22120);
xor U23440 (N_23440,N_22025,N_22310);
nor U23441 (N_23441,N_22059,N_22413);
or U23442 (N_23442,N_22182,N_22052);
or U23443 (N_23443,N_22196,N_22469);
and U23444 (N_23444,N_22585,N_22671);
nor U23445 (N_23445,N_22934,N_22113);
and U23446 (N_23446,N_22725,N_22077);
xor U23447 (N_23447,N_22616,N_22319);
nand U23448 (N_23448,N_22540,N_22112);
or U23449 (N_23449,N_22622,N_22596);
nor U23450 (N_23450,N_22618,N_22837);
nor U23451 (N_23451,N_22543,N_22468);
nor U23452 (N_23452,N_22016,N_22773);
and U23453 (N_23453,N_22908,N_22356);
nor U23454 (N_23454,N_22300,N_22679);
nor U23455 (N_23455,N_22984,N_22876);
nand U23456 (N_23456,N_22352,N_22657);
nand U23457 (N_23457,N_22358,N_22079);
nand U23458 (N_23458,N_22803,N_22418);
nor U23459 (N_23459,N_22575,N_22753);
nor U23460 (N_23460,N_22135,N_22023);
nand U23461 (N_23461,N_22130,N_22417);
nand U23462 (N_23462,N_22231,N_22834);
nor U23463 (N_23463,N_22993,N_22070);
nand U23464 (N_23464,N_22791,N_22917);
nand U23465 (N_23465,N_22567,N_22631);
nand U23466 (N_23466,N_22157,N_22035);
xnor U23467 (N_23467,N_22937,N_22151);
nand U23468 (N_23468,N_22018,N_22014);
and U23469 (N_23469,N_22220,N_22859);
xnor U23470 (N_23470,N_22073,N_22496);
nor U23471 (N_23471,N_22283,N_22153);
nor U23472 (N_23472,N_22507,N_22333);
xnor U23473 (N_23473,N_22925,N_22769);
nand U23474 (N_23474,N_22376,N_22918);
xor U23475 (N_23475,N_22687,N_22694);
or U23476 (N_23476,N_22183,N_22459);
or U23477 (N_23477,N_22932,N_22253);
and U23478 (N_23478,N_22170,N_22823);
or U23479 (N_23479,N_22553,N_22411);
and U23480 (N_23480,N_22904,N_22515);
nand U23481 (N_23481,N_22460,N_22187);
and U23482 (N_23482,N_22665,N_22647);
and U23483 (N_23483,N_22000,N_22548);
or U23484 (N_23484,N_22517,N_22703);
and U23485 (N_23485,N_22134,N_22645);
xor U23486 (N_23486,N_22717,N_22835);
nand U23487 (N_23487,N_22541,N_22186);
xnor U23488 (N_23488,N_22330,N_22995);
nor U23489 (N_23489,N_22656,N_22421);
nor U23490 (N_23490,N_22982,N_22563);
nor U23491 (N_23491,N_22028,N_22389);
xor U23492 (N_23492,N_22735,N_22020);
xnor U23493 (N_23493,N_22825,N_22601);
and U23494 (N_23494,N_22867,N_22749);
or U23495 (N_23495,N_22275,N_22405);
nand U23496 (N_23496,N_22408,N_22759);
nor U23497 (N_23497,N_22944,N_22392);
nand U23498 (N_23498,N_22033,N_22766);
xnor U23499 (N_23499,N_22732,N_22989);
and U23500 (N_23500,N_22254,N_22217);
or U23501 (N_23501,N_22137,N_22500);
nor U23502 (N_23502,N_22732,N_22482);
and U23503 (N_23503,N_22133,N_22016);
xor U23504 (N_23504,N_22001,N_22140);
and U23505 (N_23505,N_22289,N_22546);
xor U23506 (N_23506,N_22448,N_22294);
nand U23507 (N_23507,N_22052,N_22332);
and U23508 (N_23508,N_22478,N_22110);
and U23509 (N_23509,N_22641,N_22802);
nor U23510 (N_23510,N_22880,N_22950);
xnor U23511 (N_23511,N_22551,N_22090);
nand U23512 (N_23512,N_22407,N_22642);
xnor U23513 (N_23513,N_22704,N_22260);
or U23514 (N_23514,N_22624,N_22048);
xnor U23515 (N_23515,N_22798,N_22429);
or U23516 (N_23516,N_22567,N_22720);
nand U23517 (N_23517,N_22241,N_22719);
and U23518 (N_23518,N_22601,N_22375);
nor U23519 (N_23519,N_22068,N_22614);
and U23520 (N_23520,N_22767,N_22101);
xnor U23521 (N_23521,N_22297,N_22896);
xor U23522 (N_23522,N_22693,N_22135);
and U23523 (N_23523,N_22646,N_22759);
xnor U23524 (N_23524,N_22854,N_22510);
nand U23525 (N_23525,N_22454,N_22705);
xor U23526 (N_23526,N_22940,N_22055);
or U23527 (N_23527,N_22821,N_22265);
or U23528 (N_23528,N_22735,N_22551);
or U23529 (N_23529,N_22005,N_22234);
nand U23530 (N_23530,N_22918,N_22131);
nand U23531 (N_23531,N_22730,N_22077);
nand U23532 (N_23532,N_22440,N_22454);
or U23533 (N_23533,N_22285,N_22027);
nand U23534 (N_23534,N_22290,N_22084);
nand U23535 (N_23535,N_22086,N_22639);
and U23536 (N_23536,N_22395,N_22874);
or U23537 (N_23537,N_22005,N_22746);
nor U23538 (N_23538,N_22155,N_22777);
nor U23539 (N_23539,N_22492,N_22005);
nor U23540 (N_23540,N_22225,N_22307);
nor U23541 (N_23541,N_22977,N_22104);
xnor U23542 (N_23542,N_22663,N_22494);
and U23543 (N_23543,N_22710,N_22589);
and U23544 (N_23544,N_22252,N_22709);
nand U23545 (N_23545,N_22365,N_22790);
or U23546 (N_23546,N_22339,N_22586);
nor U23547 (N_23547,N_22196,N_22908);
nand U23548 (N_23548,N_22570,N_22140);
nor U23549 (N_23549,N_22274,N_22843);
nor U23550 (N_23550,N_22976,N_22405);
and U23551 (N_23551,N_22943,N_22478);
xor U23552 (N_23552,N_22906,N_22812);
nor U23553 (N_23553,N_22190,N_22002);
nand U23554 (N_23554,N_22139,N_22174);
nand U23555 (N_23555,N_22387,N_22020);
and U23556 (N_23556,N_22369,N_22139);
and U23557 (N_23557,N_22162,N_22328);
or U23558 (N_23558,N_22111,N_22963);
nor U23559 (N_23559,N_22429,N_22009);
nand U23560 (N_23560,N_22585,N_22777);
nand U23561 (N_23561,N_22750,N_22731);
or U23562 (N_23562,N_22308,N_22360);
and U23563 (N_23563,N_22923,N_22638);
nor U23564 (N_23564,N_22105,N_22080);
or U23565 (N_23565,N_22054,N_22192);
xor U23566 (N_23566,N_22823,N_22941);
and U23567 (N_23567,N_22861,N_22321);
xnor U23568 (N_23568,N_22495,N_22709);
nand U23569 (N_23569,N_22727,N_22780);
or U23570 (N_23570,N_22613,N_22071);
nand U23571 (N_23571,N_22985,N_22139);
or U23572 (N_23572,N_22539,N_22509);
or U23573 (N_23573,N_22895,N_22091);
and U23574 (N_23574,N_22546,N_22792);
xnor U23575 (N_23575,N_22385,N_22125);
nor U23576 (N_23576,N_22788,N_22216);
or U23577 (N_23577,N_22552,N_22556);
and U23578 (N_23578,N_22790,N_22937);
xnor U23579 (N_23579,N_22046,N_22282);
nand U23580 (N_23580,N_22434,N_22107);
nor U23581 (N_23581,N_22454,N_22873);
xor U23582 (N_23582,N_22437,N_22256);
nor U23583 (N_23583,N_22675,N_22518);
or U23584 (N_23584,N_22996,N_22371);
nor U23585 (N_23585,N_22976,N_22798);
and U23586 (N_23586,N_22954,N_22246);
nand U23587 (N_23587,N_22139,N_22828);
or U23588 (N_23588,N_22448,N_22638);
xor U23589 (N_23589,N_22743,N_22019);
xor U23590 (N_23590,N_22239,N_22047);
and U23591 (N_23591,N_22699,N_22351);
nor U23592 (N_23592,N_22203,N_22270);
or U23593 (N_23593,N_22665,N_22267);
or U23594 (N_23594,N_22178,N_22307);
xor U23595 (N_23595,N_22346,N_22262);
and U23596 (N_23596,N_22501,N_22612);
and U23597 (N_23597,N_22161,N_22235);
nor U23598 (N_23598,N_22086,N_22298);
xnor U23599 (N_23599,N_22257,N_22122);
xnor U23600 (N_23600,N_22127,N_22941);
and U23601 (N_23601,N_22509,N_22686);
or U23602 (N_23602,N_22380,N_22523);
nor U23603 (N_23603,N_22004,N_22239);
xnor U23604 (N_23604,N_22797,N_22144);
or U23605 (N_23605,N_22649,N_22161);
and U23606 (N_23606,N_22160,N_22383);
and U23607 (N_23607,N_22515,N_22522);
xor U23608 (N_23608,N_22254,N_22338);
or U23609 (N_23609,N_22806,N_22589);
and U23610 (N_23610,N_22846,N_22131);
or U23611 (N_23611,N_22883,N_22008);
nor U23612 (N_23612,N_22300,N_22785);
xnor U23613 (N_23613,N_22795,N_22835);
and U23614 (N_23614,N_22222,N_22325);
nor U23615 (N_23615,N_22357,N_22220);
and U23616 (N_23616,N_22076,N_22754);
nor U23617 (N_23617,N_22274,N_22831);
nor U23618 (N_23618,N_22035,N_22818);
nand U23619 (N_23619,N_22593,N_22631);
or U23620 (N_23620,N_22648,N_22001);
nand U23621 (N_23621,N_22380,N_22478);
xor U23622 (N_23622,N_22594,N_22792);
xnor U23623 (N_23623,N_22725,N_22113);
nand U23624 (N_23624,N_22953,N_22078);
or U23625 (N_23625,N_22582,N_22006);
xor U23626 (N_23626,N_22809,N_22864);
xnor U23627 (N_23627,N_22328,N_22468);
nand U23628 (N_23628,N_22605,N_22085);
and U23629 (N_23629,N_22464,N_22034);
or U23630 (N_23630,N_22341,N_22079);
nor U23631 (N_23631,N_22963,N_22730);
xnor U23632 (N_23632,N_22744,N_22999);
xnor U23633 (N_23633,N_22901,N_22716);
or U23634 (N_23634,N_22406,N_22530);
or U23635 (N_23635,N_22712,N_22587);
xnor U23636 (N_23636,N_22224,N_22049);
or U23637 (N_23637,N_22214,N_22053);
nor U23638 (N_23638,N_22129,N_22969);
or U23639 (N_23639,N_22908,N_22335);
nand U23640 (N_23640,N_22580,N_22806);
and U23641 (N_23641,N_22866,N_22295);
nand U23642 (N_23642,N_22024,N_22138);
xor U23643 (N_23643,N_22821,N_22073);
or U23644 (N_23644,N_22618,N_22976);
xnor U23645 (N_23645,N_22168,N_22827);
nor U23646 (N_23646,N_22773,N_22163);
and U23647 (N_23647,N_22381,N_22347);
or U23648 (N_23648,N_22113,N_22810);
nor U23649 (N_23649,N_22836,N_22632);
nand U23650 (N_23650,N_22955,N_22440);
and U23651 (N_23651,N_22021,N_22809);
nand U23652 (N_23652,N_22622,N_22656);
or U23653 (N_23653,N_22878,N_22563);
nor U23654 (N_23654,N_22504,N_22295);
or U23655 (N_23655,N_22294,N_22284);
and U23656 (N_23656,N_22877,N_22115);
nor U23657 (N_23657,N_22298,N_22801);
and U23658 (N_23658,N_22545,N_22778);
nand U23659 (N_23659,N_22909,N_22517);
and U23660 (N_23660,N_22469,N_22599);
and U23661 (N_23661,N_22820,N_22866);
nor U23662 (N_23662,N_22231,N_22303);
nor U23663 (N_23663,N_22943,N_22468);
nand U23664 (N_23664,N_22723,N_22547);
or U23665 (N_23665,N_22916,N_22546);
or U23666 (N_23666,N_22699,N_22431);
and U23667 (N_23667,N_22453,N_22802);
nand U23668 (N_23668,N_22881,N_22229);
xnor U23669 (N_23669,N_22195,N_22400);
or U23670 (N_23670,N_22583,N_22198);
nand U23671 (N_23671,N_22000,N_22430);
or U23672 (N_23672,N_22774,N_22796);
and U23673 (N_23673,N_22647,N_22332);
and U23674 (N_23674,N_22846,N_22993);
and U23675 (N_23675,N_22712,N_22884);
nor U23676 (N_23676,N_22621,N_22180);
and U23677 (N_23677,N_22630,N_22853);
xor U23678 (N_23678,N_22666,N_22949);
and U23679 (N_23679,N_22207,N_22489);
and U23680 (N_23680,N_22206,N_22816);
or U23681 (N_23681,N_22500,N_22893);
and U23682 (N_23682,N_22399,N_22865);
and U23683 (N_23683,N_22820,N_22197);
or U23684 (N_23684,N_22975,N_22611);
or U23685 (N_23685,N_22256,N_22609);
and U23686 (N_23686,N_22128,N_22667);
nor U23687 (N_23687,N_22915,N_22698);
and U23688 (N_23688,N_22999,N_22629);
nor U23689 (N_23689,N_22276,N_22612);
xnor U23690 (N_23690,N_22529,N_22432);
and U23691 (N_23691,N_22865,N_22441);
nand U23692 (N_23692,N_22910,N_22545);
nand U23693 (N_23693,N_22733,N_22982);
and U23694 (N_23694,N_22759,N_22856);
xor U23695 (N_23695,N_22973,N_22497);
nand U23696 (N_23696,N_22966,N_22622);
nor U23697 (N_23697,N_22161,N_22797);
nand U23698 (N_23698,N_22291,N_22126);
nor U23699 (N_23699,N_22365,N_22170);
xnor U23700 (N_23700,N_22771,N_22825);
or U23701 (N_23701,N_22466,N_22032);
nand U23702 (N_23702,N_22744,N_22592);
nand U23703 (N_23703,N_22309,N_22493);
nand U23704 (N_23704,N_22917,N_22304);
xor U23705 (N_23705,N_22671,N_22589);
nand U23706 (N_23706,N_22748,N_22124);
or U23707 (N_23707,N_22780,N_22966);
nor U23708 (N_23708,N_22788,N_22962);
or U23709 (N_23709,N_22124,N_22021);
and U23710 (N_23710,N_22599,N_22786);
or U23711 (N_23711,N_22593,N_22592);
nand U23712 (N_23712,N_22961,N_22725);
or U23713 (N_23713,N_22426,N_22113);
nand U23714 (N_23714,N_22157,N_22152);
xor U23715 (N_23715,N_22391,N_22750);
nor U23716 (N_23716,N_22397,N_22650);
and U23717 (N_23717,N_22566,N_22961);
or U23718 (N_23718,N_22417,N_22412);
nand U23719 (N_23719,N_22973,N_22576);
nand U23720 (N_23720,N_22158,N_22319);
and U23721 (N_23721,N_22293,N_22445);
xnor U23722 (N_23722,N_22964,N_22730);
xor U23723 (N_23723,N_22492,N_22718);
nand U23724 (N_23724,N_22072,N_22100);
nor U23725 (N_23725,N_22468,N_22963);
xnor U23726 (N_23726,N_22888,N_22119);
and U23727 (N_23727,N_22509,N_22774);
and U23728 (N_23728,N_22216,N_22138);
xnor U23729 (N_23729,N_22555,N_22452);
nand U23730 (N_23730,N_22432,N_22831);
nand U23731 (N_23731,N_22713,N_22796);
and U23732 (N_23732,N_22827,N_22078);
or U23733 (N_23733,N_22748,N_22591);
or U23734 (N_23734,N_22370,N_22377);
and U23735 (N_23735,N_22977,N_22647);
xor U23736 (N_23736,N_22509,N_22840);
nand U23737 (N_23737,N_22891,N_22006);
nand U23738 (N_23738,N_22601,N_22004);
nand U23739 (N_23739,N_22993,N_22686);
nor U23740 (N_23740,N_22486,N_22133);
nand U23741 (N_23741,N_22768,N_22486);
nand U23742 (N_23742,N_22920,N_22580);
nor U23743 (N_23743,N_22928,N_22426);
or U23744 (N_23744,N_22372,N_22003);
xnor U23745 (N_23745,N_22074,N_22664);
nor U23746 (N_23746,N_22948,N_22058);
nor U23747 (N_23747,N_22346,N_22202);
nand U23748 (N_23748,N_22329,N_22219);
and U23749 (N_23749,N_22290,N_22356);
xnor U23750 (N_23750,N_22804,N_22314);
and U23751 (N_23751,N_22917,N_22628);
and U23752 (N_23752,N_22179,N_22251);
nor U23753 (N_23753,N_22072,N_22622);
nand U23754 (N_23754,N_22177,N_22586);
or U23755 (N_23755,N_22904,N_22865);
xor U23756 (N_23756,N_22725,N_22201);
nand U23757 (N_23757,N_22957,N_22675);
xnor U23758 (N_23758,N_22323,N_22738);
and U23759 (N_23759,N_22356,N_22071);
nand U23760 (N_23760,N_22030,N_22865);
and U23761 (N_23761,N_22945,N_22012);
or U23762 (N_23762,N_22584,N_22991);
nor U23763 (N_23763,N_22863,N_22195);
nor U23764 (N_23764,N_22741,N_22491);
xnor U23765 (N_23765,N_22234,N_22298);
and U23766 (N_23766,N_22467,N_22070);
nand U23767 (N_23767,N_22460,N_22579);
or U23768 (N_23768,N_22079,N_22401);
xor U23769 (N_23769,N_22757,N_22019);
xor U23770 (N_23770,N_22378,N_22193);
and U23771 (N_23771,N_22404,N_22891);
or U23772 (N_23772,N_22206,N_22229);
or U23773 (N_23773,N_22578,N_22194);
and U23774 (N_23774,N_22967,N_22297);
or U23775 (N_23775,N_22876,N_22868);
and U23776 (N_23776,N_22051,N_22358);
nand U23777 (N_23777,N_22749,N_22850);
nor U23778 (N_23778,N_22866,N_22125);
or U23779 (N_23779,N_22822,N_22371);
nand U23780 (N_23780,N_22378,N_22492);
and U23781 (N_23781,N_22759,N_22983);
and U23782 (N_23782,N_22607,N_22690);
nor U23783 (N_23783,N_22365,N_22798);
or U23784 (N_23784,N_22648,N_22549);
or U23785 (N_23785,N_22275,N_22746);
and U23786 (N_23786,N_22477,N_22489);
xor U23787 (N_23787,N_22524,N_22881);
or U23788 (N_23788,N_22367,N_22262);
nand U23789 (N_23789,N_22345,N_22835);
nor U23790 (N_23790,N_22401,N_22427);
xor U23791 (N_23791,N_22668,N_22042);
nand U23792 (N_23792,N_22164,N_22972);
xnor U23793 (N_23793,N_22618,N_22023);
and U23794 (N_23794,N_22581,N_22609);
xor U23795 (N_23795,N_22943,N_22787);
xnor U23796 (N_23796,N_22766,N_22473);
nor U23797 (N_23797,N_22137,N_22414);
xnor U23798 (N_23798,N_22508,N_22817);
nor U23799 (N_23799,N_22230,N_22265);
xnor U23800 (N_23800,N_22757,N_22634);
or U23801 (N_23801,N_22874,N_22074);
nand U23802 (N_23802,N_22206,N_22639);
nand U23803 (N_23803,N_22499,N_22815);
xor U23804 (N_23804,N_22689,N_22867);
or U23805 (N_23805,N_22311,N_22895);
xnor U23806 (N_23806,N_22088,N_22899);
xor U23807 (N_23807,N_22329,N_22264);
xnor U23808 (N_23808,N_22470,N_22706);
or U23809 (N_23809,N_22217,N_22198);
nor U23810 (N_23810,N_22521,N_22577);
xnor U23811 (N_23811,N_22677,N_22695);
or U23812 (N_23812,N_22591,N_22472);
nor U23813 (N_23813,N_22502,N_22082);
xnor U23814 (N_23814,N_22727,N_22811);
or U23815 (N_23815,N_22442,N_22653);
and U23816 (N_23816,N_22133,N_22626);
nand U23817 (N_23817,N_22301,N_22241);
nor U23818 (N_23818,N_22444,N_22615);
or U23819 (N_23819,N_22979,N_22157);
nand U23820 (N_23820,N_22141,N_22855);
nand U23821 (N_23821,N_22892,N_22597);
nand U23822 (N_23822,N_22045,N_22305);
nand U23823 (N_23823,N_22657,N_22010);
and U23824 (N_23824,N_22065,N_22303);
and U23825 (N_23825,N_22230,N_22890);
nor U23826 (N_23826,N_22022,N_22095);
and U23827 (N_23827,N_22200,N_22505);
and U23828 (N_23828,N_22334,N_22620);
nor U23829 (N_23829,N_22677,N_22462);
nor U23830 (N_23830,N_22381,N_22149);
or U23831 (N_23831,N_22975,N_22920);
xor U23832 (N_23832,N_22156,N_22667);
or U23833 (N_23833,N_22212,N_22948);
xor U23834 (N_23834,N_22605,N_22621);
xor U23835 (N_23835,N_22005,N_22152);
and U23836 (N_23836,N_22478,N_22055);
nor U23837 (N_23837,N_22104,N_22644);
nor U23838 (N_23838,N_22316,N_22372);
nor U23839 (N_23839,N_22260,N_22994);
or U23840 (N_23840,N_22479,N_22013);
nor U23841 (N_23841,N_22444,N_22423);
and U23842 (N_23842,N_22102,N_22180);
and U23843 (N_23843,N_22459,N_22179);
nand U23844 (N_23844,N_22089,N_22647);
nand U23845 (N_23845,N_22503,N_22139);
or U23846 (N_23846,N_22406,N_22602);
nand U23847 (N_23847,N_22904,N_22204);
nand U23848 (N_23848,N_22497,N_22883);
nor U23849 (N_23849,N_22368,N_22064);
nand U23850 (N_23850,N_22265,N_22099);
or U23851 (N_23851,N_22186,N_22181);
nor U23852 (N_23852,N_22310,N_22627);
or U23853 (N_23853,N_22760,N_22895);
nand U23854 (N_23854,N_22746,N_22097);
xor U23855 (N_23855,N_22037,N_22462);
nand U23856 (N_23856,N_22600,N_22209);
xor U23857 (N_23857,N_22714,N_22552);
xor U23858 (N_23858,N_22505,N_22510);
nor U23859 (N_23859,N_22198,N_22605);
or U23860 (N_23860,N_22215,N_22040);
nand U23861 (N_23861,N_22596,N_22972);
nand U23862 (N_23862,N_22813,N_22808);
and U23863 (N_23863,N_22806,N_22137);
xor U23864 (N_23864,N_22282,N_22231);
nand U23865 (N_23865,N_22037,N_22100);
nor U23866 (N_23866,N_22889,N_22901);
and U23867 (N_23867,N_22760,N_22143);
and U23868 (N_23868,N_22880,N_22035);
or U23869 (N_23869,N_22314,N_22407);
xnor U23870 (N_23870,N_22392,N_22415);
xor U23871 (N_23871,N_22470,N_22642);
or U23872 (N_23872,N_22232,N_22141);
nor U23873 (N_23873,N_22935,N_22961);
nand U23874 (N_23874,N_22947,N_22603);
xnor U23875 (N_23875,N_22153,N_22699);
xnor U23876 (N_23876,N_22829,N_22397);
xnor U23877 (N_23877,N_22682,N_22549);
nor U23878 (N_23878,N_22322,N_22767);
nand U23879 (N_23879,N_22959,N_22417);
nor U23880 (N_23880,N_22484,N_22864);
or U23881 (N_23881,N_22260,N_22137);
xnor U23882 (N_23882,N_22066,N_22071);
or U23883 (N_23883,N_22320,N_22195);
xnor U23884 (N_23884,N_22542,N_22482);
nand U23885 (N_23885,N_22710,N_22343);
nand U23886 (N_23886,N_22951,N_22880);
nor U23887 (N_23887,N_22879,N_22937);
and U23888 (N_23888,N_22534,N_22046);
nand U23889 (N_23889,N_22735,N_22842);
nor U23890 (N_23890,N_22396,N_22624);
and U23891 (N_23891,N_22334,N_22849);
nand U23892 (N_23892,N_22076,N_22384);
nand U23893 (N_23893,N_22056,N_22429);
nand U23894 (N_23894,N_22838,N_22438);
or U23895 (N_23895,N_22303,N_22131);
and U23896 (N_23896,N_22776,N_22682);
xor U23897 (N_23897,N_22972,N_22525);
nor U23898 (N_23898,N_22286,N_22976);
nand U23899 (N_23899,N_22365,N_22434);
nand U23900 (N_23900,N_22088,N_22369);
nand U23901 (N_23901,N_22780,N_22565);
nand U23902 (N_23902,N_22652,N_22456);
nand U23903 (N_23903,N_22436,N_22354);
nor U23904 (N_23904,N_22549,N_22566);
and U23905 (N_23905,N_22071,N_22664);
and U23906 (N_23906,N_22886,N_22385);
xnor U23907 (N_23907,N_22939,N_22766);
nand U23908 (N_23908,N_22724,N_22712);
and U23909 (N_23909,N_22970,N_22187);
nand U23910 (N_23910,N_22909,N_22893);
nand U23911 (N_23911,N_22021,N_22376);
xnor U23912 (N_23912,N_22017,N_22426);
nand U23913 (N_23913,N_22698,N_22199);
nand U23914 (N_23914,N_22631,N_22184);
or U23915 (N_23915,N_22999,N_22457);
nor U23916 (N_23916,N_22980,N_22117);
nor U23917 (N_23917,N_22323,N_22191);
xor U23918 (N_23918,N_22212,N_22983);
or U23919 (N_23919,N_22308,N_22747);
and U23920 (N_23920,N_22382,N_22093);
nor U23921 (N_23921,N_22234,N_22815);
or U23922 (N_23922,N_22586,N_22641);
nor U23923 (N_23923,N_22620,N_22610);
and U23924 (N_23924,N_22243,N_22622);
nor U23925 (N_23925,N_22027,N_22037);
and U23926 (N_23926,N_22143,N_22051);
xnor U23927 (N_23927,N_22231,N_22586);
xnor U23928 (N_23928,N_22390,N_22009);
nand U23929 (N_23929,N_22728,N_22975);
xnor U23930 (N_23930,N_22690,N_22770);
and U23931 (N_23931,N_22075,N_22937);
nand U23932 (N_23932,N_22350,N_22525);
and U23933 (N_23933,N_22506,N_22609);
and U23934 (N_23934,N_22096,N_22103);
and U23935 (N_23935,N_22105,N_22971);
nor U23936 (N_23936,N_22316,N_22986);
or U23937 (N_23937,N_22472,N_22698);
xor U23938 (N_23938,N_22433,N_22578);
nand U23939 (N_23939,N_22729,N_22019);
nor U23940 (N_23940,N_22260,N_22739);
nor U23941 (N_23941,N_22033,N_22647);
or U23942 (N_23942,N_22507,N_22668);
or U23943 (N_23943,N_22716,N_22520);
nand U23944 (N_23944,N_22072,N_22500);
and U23945 (N_23945,N_22416,N_22014);
or U23946 (N_23946,N_22084,N_22888);
nor U23947 (N_23947,N_22383,N_22423);
nor U23948 (N_23948,N_22681,N_22409);
xnor U23949 (N_23949,N_22525,N_22196);
xor U23950 (N_23950,N_22353,N_22601);
or U23951 (N_23951,N_22557,N_22356);
xnor U23952 (N_23952,N_22292,N_22590);
and U23953 (N_23953,N_22979,N_22328);
nor U23954 (N_23954,N_22087,N_22985);
xnor U23955 (N_23955,N_22146,N_22977);
nand U23956 (N_23956,N_22012,N_22254);
nor U23957 (N_23957,N_22271,N_22909);
nand U23958 (N_23958,N_22717,N_22701);
nor U23959 (N_23959,N_22056,N_22325);
nand U23960 (N_23960,N_22043,N_22327);
or U23961 (N_23961,N_22017,N_22383);
or U23962 (N_23962,N_22006,N_22879);
and U23963 (N_23963,N_22230,N_22646);
nor U23964 (N_23964,N_22570,N_22764);
nor U23965 (N_23965,N_22155,N_22055);
or U23966 (N_23966,N_22926,N_22038);
nor U23967 (N_23967,N_22995,N_22657);
and U23968 (N_23968,N_22272,N_22261);
nor U23969 (N_23969,N_22741,N_22108);
nand U23970 (N_23970,N_22561,N_22269);
nor U23971 (N_23971,N_22611,N_22579);
nor U23972 (N_23972,N_22754,N_22168);
xor U23973 (N_23973,N_22069,N_22086);
and U23974 (N_23974,N_22840,N_22921);
nand U23975 (N_23975,N_22950,N_22048);
xor U23976 (N_23976,N_22635,N_22196);
nor U23977 (N_23977,N_22928,N_22728);
nor U23978 (N_23978,N_22870,N_22040);
and U23979 (N_23979,N_22689,N_22776);
nor U23980 (N_23980,N_22623,N_22795);
nor U23981 (N_23981,N_22406,N_22898);
or U23982 (N_23982,N_22064,N_22926);
xnor U23983 (N_23983,N_22873,N_22100);
nand U23984 (N_23984,N_22864,N_22222);
or U23985 (N_23985,N_22036,N_22922);
or U23986 (N_23986,N_22917,N_22796);
or U23987 (N_23987,N_22124,N_22422);
or U23988 (N_23988,N_22403,N_22581);
or U23989 (N_23989,N_22548,N_22325);
xnor U23990 (N_23990,N_22670,N_22206);
xnor U23991 (N_23991,N_22384,N_22354);
nor U23992 (N_23992,N_22830,N_22666);
xnor U23993 (N_23993,N_22252,N_22119);
or U23994 (N_23994,N_22882,N_22271);
or U23995 (N_23995,N_22140,N_22435);
or U23996 (N_23996,N_22533,N_22552);
xnor U23997 (N_23997,N_22143,N_22693);
xor U23998 (N_23998,N_22854,N_22821);
or U23999 (N_23999,N_22328,N_22821);
nand U24000 (N_24000,N_23484,N_23018);
xor U24001 (N_24001,N_23246,N_23764);
xor U24002 (N_24002,N_23918,N_23297);
xnor U24003 (N_24003,N_23170,N_23848);
or U24004 (N_24004,N_23895,N_23458);
nor U24005 (N_24005,N_23131,N_23964);
nand U24006 (N_24006,N_23881,N_23664);
nor U24007 (N_24007,N_23326,N_23619);
nand U24008 (N_24008,N_23858,N_23691);
nand U24009 (N_24009,N_23553,N_23041);
and U24010 (N_24010,N_23751,N_23332);
and U24011 (N_24011,N_23993,N_23483);
nor U24012 (N_24012,N_23634,N_23707);
nand U24013 (N_24013,N_23862,N_23894);
nand U24014 (N_24014,N_23050,N_23731);
nand U24015 (N_24015,N_23824,N_23815);
or U24016 (N_24016,N_23058,N_23254);
xnor U24017 (N_24017,N_23531,N_23430);
xnor U24018 (N_24018,N_23437,N_23885);
nor U24019 (N_24019,N_23009,N_23435);
nand U24020 (N_24020,N_23126,N_23793);
or U24021 (N_24021,N_23721,N_23842);
or U24022 (N_24022,N_23156,N_23564);
and U24023 (N_24023,N_23275,N_23620);
nor U24024 (N_24024,N_23747,N_23537);
xnor U24025 (N_24025,N_23729,N_23528);
nand U24026 (N_24026,N_23549,N_23414);
or U24027 (N_24027,N_23578,N_23561);
xor U24028 (N_24028,N_23724,N_23580);
and U24029 (N_24029,N_23251,N_23078);
or U24030 (N_24030,N_23904,N_23569);
and U24031 (N_24031,N_23119,N_23139);
xnor U24032 (N_24032,N_23014,N_23514);
nor U24033 (N_24033,N_23916,N_23114);
nor U24034 (N_24034,N_23714,N_23345);
nand U24035 (N_24035,N_23287,N_23750);
nor U24036 (N_24036,N_23442,N_23380);
nor U24037 (N_24037,N_23028,N_23941);
xnor U24038 (N_24038,N_23718,N_23221);
or U24039 (N_24039,N_23302,N_23261);
and U24040 (N_24040,N_23543,N_23796);
nand U24041 (N_24041,N_23276,N_23850);
nand U24042 (N_24042,N_23010,N_23915);
or U24043 (N_24043,N_23797,N_23185);
nor U24044 (N_24044,N_23847,N_23165);
nand U24045 (N_24045,N_23845,N_23097);
xnor U24046 (N_24046,N_23044,N_23337);
nor U24047 (N_24047,N_23982,N_23662);
nor U24048 (N_24048,N_23944,N_23667);
xor U24049 (N_24049,N_23213,N_23831);
nand U24050 (N_24050,N_23612,N_23004);
or U24051 (N_24051,N_23048,N_23826);
nand U24052 (N_24052,N_23777,N_23113);
or U24053 (N_24053,N_23681,N_23379);
nand U24054 (N_24054,N_23683,N_23348);
and U24055 (N_24055,N_23931,N_23364);
or U24056 (N_24056,N_23960,N_23997);
nor U24057 (N_24057,N_23638,N_23659);
or U24058 (N_24058,N_23601,N_23935);
or U24059 (N_24059,N_23525,N_23937);
xor U24060 (N_24060,N_23618,N_23095);
nand U24061 (N_24061,N_23782,N_23273);
xor U24062 (N_24062,N_23534,N_23889);
nand U24063 (N_24063,N_23307,N_23128);
nor U24064 (N_24064,N_23057,N_23675);
xor U24065 (N_24065,N_23849,N_23837);
nor U24066 (N_24066,N_23748,N_23653);
xor U24067 (N_24067,N_23648,N_23296);
xor U24068 (N_24068,N_23791,N_23350);
and U24069 (N_24069,N_23053,N_23392);
nor U24070 (N_24070,N_23539,N_23868);
nand U24071 (N_24071,N_23157,N_23737);
nor U24072 (N_24072,N_23652,N_23116);
or U24073 (N_24073,N_23344,N_23519);
and U24074 (N_24074,N_23477,N_23354);
nand U24075 (N_24075,N_23112,N_23196);
and U24076 (N_24076,N_23533,N_23907);
nor U24077 (N_24077,N_23329,N_23952);
nand U24078 (N_24078,N_23927,N_23186);
and U24079 (N_24079,N_23175,N_23237);
nand U24080 (N_24080,N_23702,N_23220);
nand U24081 (N_24081,N_23841,N_23579);
or U24082 (N_24082,N_23144,N_23371);
nor U24083 (N_24083,N_23900,N_23860);
and U24084 (N_24084,N_23037,N_23926);
nand U24085 (N_24085,N_23390,N_23523);
or U24086 (N_24086,N_23809,N_23076);
nor U24087 (N_24087,N_23779,N_23411);
nand U24088 (N_24088,N_23000,N_23930);
nor U24089 (N_24089,N_23038,N_23256);
nor U24090 (N_24090,N_23384,N_23631);
nor U24091 (N_24091,N_23577,N_23395);
and U24092 (N_24092,N_23173,N_23229);
xor U24093 (N_24093,N_23783,N_23558);
xor U24094 (N_24094,N_23509,N_23190);
xor U24095 (N_24095,N_23184,N_23066);
and U24096 (N_24096,N_23554,N_23011);
and U24097 (N_24097,N_23020,N_23285);
xor U24098 (N_24098,N_23607,N_23636);
or U24099 (N_24099,N_23559,N_23034);
and U24100 (N_24100,N_23954,N_23298);
xor U24101 (N_24101,N_23291,N_23265);
nand U24102 (N_24102,N_23166,N_23966);
and U24103 (N_24103,N_23505,N_23466);
and U24104 (N_24104,N_23283,N_23030);
or U24105 (N_24105,N_23310,N_23616);
nor U24106 (N_24106,N_23465,N_23370);
or U24107 (N_24107,N_23753,N_23773);
nand U24108 (N_24108,N_23940,N_23710);
nor U24109 (N_24109,N_23589,N_23270);
xnor U24110 (N_24110,N_23162,N_23544);
and U24111 (N_24111,N_23150,N_23624);
and U24112 (N_24112,N_23836,N_23540);
nor U24113 (N_24113,N_23467,N_23594);
nor U24114 (N_24114,N_23650,N_23046);
or U24115 (N_24115,N_23804,N_23225);
or U24116 (N_24116,N_23381,N_23194);
or U24117 (N_24117,N_23602,N_23176);
nand U24118 (N_24118,N_23851,N_23970);
nand U24119 (N_24119,N_23304,N_23195);
nor U24120 (N_24120,N_23167,N_23476);
nand U24121 (N_24121,N_23906,N_23378);
and U24122 (N_24122,N_23955,N_23921);
nand U24123 (N_24123,N_23356,N_23665);
xor U24124 (N_24124,N_23306,N_23154);
and U24125 (N_24125,N_23591,N_23385);
xnor U24126 (N_24126,N_23948,N_23410);
or U24127 (N_24127,N_23049,N_23932);
nand U24128 (N_24128,N_23663,N_23064);
and U24129 (N_24129,N_23887,N_23153);
nor U24130 (N_24130,N_23141,N_23716);
and U24131 (N_24131,N_23174,N_23677);
xor U24132 (N_24132,N_23867,N_23210);
nor U24133 (N_24133,N_23468,N_23262);
xor U24134 (N_24134,N_23013,N_23812);
nor U24135 (N_24135,N_23775,N_23497);
xnor U24136 (N_24136,N_23208,N_23857);
nand U24137 (N_24137,N_23408,N_23433);
and U24138 (N_24138,N_23883,N_23216);
and U24139 (N_24139,N_23277,N_23143);
or U24140 (N_24140,N_23403,N_23440);
and U24141 (N_24141,N_23682,N_23822);
and U24142 (N_24142,N_23086,N_23043);
and U24143 (N_24143,N_23349,N_23968);
or U24144 (N_24144,N_23054,N_23890);
nor U24145 (N_24145,N_23321,N_23572);
xor U24146 (N_24146,N_23230,N_23219);
xor U24147 (N_24147,N_23375,N_23398);
and U24148 (N_24148,N_23448,N_23980);
nand U24149 (N_24149,N_23622,N_23888);
nor U24150 (N_24150,N_23203,N_23127);
and U24151 (N_24151,N_23872,N_23072);
nand U24152 (N_24152,N_23546,N_23260);
or U24153 (N_24153,N_23766,N_23995);
and U24154 (N_24154,N_23294,N_23590);
nand U24155 (N_24155,N_23778,N_23137);
nor U24156 (N_24156,N_23409,N_23991);
nand U24157 (N_24157,N_23617,N_23300);
or U24158 (N_24158,N_23402,N_23340);
xnor U24159 (N_24159,N_23293,N_23145);
xor U24160 (N_24160,N_23263,N_23025);
or U24161 (N_24161,N_23122,N_23094);
nor U24162 (N_24162,N_23532,N_23084);
nand U24163 (N_24163,N_23103,N_23420);
or U24164 (N_24164,N_23319,N_23801);
nand U24165 (N_24165,N_23279,N_23994);
nor U24166 (N_24166,N_23161,N_23258);
nor U24167 (N_24167,N_23024,N_23715);
nand U24168 (N_24168,N_23576,N_23623);
and U24169 (N_24169,N_23003,N_23556);
and U24170 (N_24170,N_23882,N_23934);
or U24171 (N_24171,N_23939,N_23852);
nor U24172 (N_24172,N_23647,N_23768);
nor U24173 (N_24173,N_23875,N_23956);
and U24174 (N_24174,N_23450,N_23343);
and U24175 (N_24175,N_23586,N_23908);
xor U24176 (N_24176,N_23198,N_23642);
xnor U24177 (N_24177,N_23295,N_23099);
nand U24178 (N_24178,N_23938,N_23239);
or U24179 (N_24179,N_23690,N_23517);
nor U24180 (N_24180,N_23820,N_23012);
or U24181 (N_24181,N_23516,N_23227);
xor U24182 (N_24182,N_23530,N_23827);
nor U24183 (N_24183,N_23447,N_23091);
or U24184 (N_24184,N_23118,N_23763);
xor U24185 (N_24185,N_23723,N_23774);
nor U24186 (N_24186,N_23999,N_23432);
nor U24187 (N_24187,N_23093,N_23898);
nor U24188 (N_24188,N_23325,N_23282);
xor U24189 (N_24189,N_23016,N_23686);
nor U24190 (N_24190,N_23100,N_23794);
or U24191 (N_24191,N_23761,N_23660);
nand U24192 (N_24192,N_23083,N_23903);
xnor U24193 (N_24193,N_23788,N_23641);
nor U24194 (N_24194,N_23206,N_23606);
xnor U24195 (N_24195,N_23864,N_23023);
nor U24196 (N_24196,N_23799,N_23207);
and U24197 (N_24197,N_23893,N_23351);
nor U24198 (N_24198,N_23637,N_23767);
and U24199 (N_24199,N_23059,N_23096);
nor U24200 (N_24200,N_23322,N_23922);
nor U24201 (N_24201,N_23699,N_23280);
or U24202 (N_24202,N_23446,N_23396);
and U24203 (N_24203,N_23651,N_23147);
nand U24204 (N_24204,N_23473,N_23518);
or U24205 (N_24205,N_23241,N_23626);
nor U24206 (N_24206,N_23758,N_23386);
or U24207 (N_24207,N_23462,N_23292);
nand U24208 (N_24208,N_23436,N_23897);
and U24209 (N_24209,N_23305,N_23338);
and U24210 (N_24210,N_23694,N_23136);
nor U24211 (N_24211,N_23829,N_23355);
or U24212 (N_24212,N_23661,N_23204);
nand U24213 (N_24213,N_23744,N_23189);
nor U24214 (N_24214,N_23742,N_23950);
or U24215 (N_24215,N_23785,N_23979);
and U24216 (N_24216,N_23062,N_23457);
or U24217 (N_24217,N_23479,N_23856);
nand U24218 (N_24218,N_23192,N_23089);
or U24219 (N_24219,N_23913,N_23047);
or U24220 (N_24220,N_23202,N_23792);
nand U24221 (N_24221,N_23706,N_23268);
nand U24222 (N_24222,N_23649,N_23490);
or U24223 (N_24223,N_23722,N_23474);
or U24224 (N_24224,N_23599,N_23526);
nor U24225 (N_24225,N_23115,N_23346);
nor U24226 (N_24226,N_23101,N_23222);
and U24227 (N_24227,N_23936,N_23557);
and U24228 (N_24228,N_23963,N_23823);
and U24229 (N_24229,N_23772,N_23353);
or U24230 (N_24230,N_23133,N_23584);
and U24231 (N_24231,N_23444,N_23308);
and U24232 (N_24232,N_23901,N_23816);
or U24233 (N_24233,N_23121,N_23975);
nor U24234 (N_24234,N_23749,N_23179);
and U24235 (N_24235,N_23709,N_23209);
or U24236 (N_24236,N_23211,N_23629);
xnor U24237 (N_24237,N_23461,N_23504);
or U24238 (N_24238,N_23290,N_23672);
xor U24239 (N_24239,N_23281,N_23668);
and U24240 (N_24240,N_23565,N_23008);
or U24241 (N_24241,N_23567,N_23803);
and U24242 (N_24242,N_23055,N_23676);
nor U24243 (N_24243,N_23102,N_23324);
and U24244 (N_24244,N_23428,N_23107);
nor U24245 (N_24245,N_23090,N_23452);
or U24246 (N_24246,N_23377,N_23309);
or U24247 (N_24247,N_23670,N_23389);
nand U24248 (N_24248,N_23771,N_23743);
or U24249 (N_24249,N_23223,N_23861);
xor U24250 (N_24250,N_23738,N_23806);
nand U24251 (N_24251,N_23445,N_23639);
nor U24252 (N_24252,N_23967,N_23988);
nor U24253 (N_24253,N_23976,N_23713);
and U24254 (N_24254,N_23026,N_23032);
nand U24255 (N_24255,N_23695,N_23286);
nor U24256 (N_24256,N_23854,N_23303);
or U24257 (N_24257,N_23658,N_23592);
or U24258 (N_24258,N_23005,N_23512);
nor U24259 (N_24259,N_23407,N_23568);
or U24260 (N_24260,N_23896,N_23455);
and U24261 (N_24261,N_23920,N_23105);
and U24262 (N_24262,N_23615,N_23910);
and U24263 (N_24263,N_23600,N_23814);
nand U24264 (N_24264,N_23808,N_23705);
or U24265 (N_24265,N_23248,N_23805);
xnor U24266 (N_24266,N_23387,N_23951);
nor U24267 (N_24267,N_23825,N_23063);
xnor U24268 (N_24268,N_23065,N_23529);
or U24269 (N_24269,N_23314,N_23911);
nand U24270 (N_24270,N_23051,N_23765);
or U24271 (N_24271,N_23376,N_23374);
nand U24272 (N_24272,N_23736,N_23886);
or U24273 (N_24273,N_23798,N_23391);
xnor U24274 (N_24274,N_23819,N_23593);
xor U24275 (N_24275,N_23511,N_23891);
xor U24276 (N_24276,N_23077,N_23109);
nand U24277 (N_24277,N_23342,N_23168);
nand U24278 (N_24278,N_23522,N_23720);
nor U24279 (N_24279,N_23366,N_23717);
nor U24280 (N_24280,N_23178,N_23146);
xor U24281 (N_24281,N_23266,N_23595);
or U24282 (N_24282,N_23187,N_23575);
nor U24283 (N_24283,N_23274,N_23740);
or U24284 (N_24284,N_23313,N_23844);
and U24285 (N_24285,N_23135,N_23817);
nand U24286 (N_24286,N_23719,N_23871);
xor U24287 (N_24287,N_23703,N_23243);
nor U24288 (N_24288,N_23070,N_23789);
and U24289 (N_24289,N_23978,N_23401);
nor U24290 (N_24290,N_23605,N_23899);
xor U24291 (N_24291,N_23909,N_23085);
xor U24292 (N_24292,N_23547,N_23563);
nor U24293 (N_24293,N_23417,N_23134);
xor U24294 (N_24294,N_23962,N_23315);
xor U24295 (N_24295,N_23002,N_23657);
or U24296 (N_24296,N_23360,N_23985);
nand U24297 (N_24297,N_23245,N_23708);
nor U24298 (N_24298,N_23874,N_23188);
and U24299 (N_24299,N_23859,N_23481);
and U24300 (N_24300,N_23124,N_23671);
nand U24301 (N_24301,N_23503,N_23625);
nor U24302 (N_24302,N_23361,N_23320);
nand U24303 (N_24303,N_23813,N_23006);
or U24304 (N_24304,N_23171,N_23866);
nor U24305 (N_24305,N_23191,N_23098);
and U24306 (N_24306,N_23802,N_23397);
nand U24307 (N_24307,N_23197,N_23684);
or U24308 (N_24308,N_23946,N_23233);
nand U24309 (N_24309,N_23746,N_23855);
nor U24310 (N_24310,N_23033,N_23902);
and U24311 (N_24311,N_23499,N_23164);
nand U24312 (N_24312,N_23235,N_23482);
xnor U24313 (N_24313,N_23865,N_23787);
nand U24314 (N_24314,N_23502,N_23040);
nor U24315 (N_24315,N_23451,N_23132);
nor U24316 (N_24316,N_23613,N_23339);
nor U24317 (N_24317,N_23604,N_23507);
xor U24318 (N_24318,N_23971,N_23218);
and U24319 (N_24319,N_23770,N_23693);
and U24320 (N_24320,N_23680,N_23182);
nor U24321 (N_24321,N_23369,N_23289);
xnor U24322 (N_24322,N_23491,N_23608);
nand U24323 (N_24323,N_23784,N_23635);
or U24324 (N_24324,N_23566,N_23125);
xnor U24325 (N_24325,N_23487,N_23597);
nor U24326 (N_24326,N_23596,N_23075);
nor U24327 (N_24327,N_23943,N_23045);
and U24328 (N_24328,N_23762,N_23312);
xor U24329 (N_24329,N_23501,N_23019);
nor U24330 (N_24330,N_23654,N_23830);
or U24331 (N_24331,N_23924,N_23400);
xor U24332 (N_24332,N_23585,N_23253);
or U24333 (N_24333,N_23264,N_23341);
nor U24334 (N_24334,N_23998,N_23431);
or U24335 (N_24335,N_23311,N_23080);
or U24336 (N_24336,N_23470,N_23416);
nor U24337 (N_24337,N_23551,N_23987);
and U24338 (N_24338,N_23795,N_23177);
nor U24339 (N_24339,N_23728,N_23495);
xor U24340 (N_24340,N_23628,N_23800);
or U24341 (N_24341,N_23212,N_23163);
or U24342 (N_24342,N_23358,N_23029);
or U24343 (N_24343,N_23733,N_23160);
or U24344 (N_24344,N_23535,N_23524);
nand U24345 (N_24345,N_23087,N_23228);
xnor U24346 (N_24346,N_23469,N_23232);
and U24347 (N_24347,N_23073,N_23581);
nor U24348 (N_24348,N_23552,N_23240);
nand U24349 (N_24349,N_23538,N_23735);
and U24350 (N_24350,N_23427,N_23510);
xor U24351 (N_24351,N_23953,N_23106);
and U24352 (N_24352,N_23082,N_23609);
or U24353 (N_24353,N_23074,N_23007);
and U24354 (N_24354,N_23574,N_23560);
xnor U24355 (N_24355,N_23301,N_23317);
and U24356 (N_24356,N_23520,N_23630);
or U24357 (N_24357,N_23422,N_23821);
nor U24358 (N_24358,N_23679,N_23739);
or U24359 (N_24359,N_23284,N_23081);
and U24360 (N_24360,N_23238,N_23692);
nand U24361 (N_24361,N_23061,N_23666);
xnor U24362 (N_24362,N_23541,N_23035);
or U24363 (N_24363,N_23015,N_23947);
xnor U24364 (N_24364,N_23627,N_23712);
nor U24365 (N_24365,N_23786,N_23917);
and U24366 (N_24366,N_23244,N_23498);
and U24367 (N_24367,N_23323,N_23949);
and U24368 (N_24368,N_23426,N_23697);
nand U24369 (N_24369,N_23878,N_23129);
and U24370 (N_24370,N_23357,N_23996);
nor U24371 (N_24371,N_23372,N_23990);
xor U24372 (N_24372,N_23500,N_23536);
nand U24373 (N_24373,N_23421,N_23621);
or U24374 (N_24374,N_23542,N_23732);
nor U24375 (N_24375,N_23234,N_23299);
or U24376 (N_24376,N_23673,N_23199);
xor U24377 (N_24377,N_23912,N_23646);
nor U24378 (N_24378,N_23255,N_23333);
or U24379 (N_24379,N_23352,N_23404);
xor U24380 (N_24380,N_23570,N_23036);
and U24381 (N_24381,N_23471,N_23942);
nand U24382 (N_24382,N_23459,N_23496);
xor U24383 (N_24383,N_23478,N_23678);
xor U24384 (N_24384,N_23067,N_23250);
nor U24385 (N_24385,N_23905,N_23027);
nor U24386 (N_24386,N_23017,N_23869);
xnor U24387 (N_24387,N_23200,N_23527);
or U24388 (N_24388,N_23521,N_23181);
xnor U24389 (N_24389,N_23870,N_23151);
xnor U24390 (N_24390,N_23328,N_23700);
nor U24391 (N_24391,N_23486,N_23992);
and U24392 (N_24392,N_23021,N_23363);
or U24393 (N_24393,N_23393,N_23923);
and U24394 (N_24394,N_23969,N_23278);
and U24395 (N_24395,N_23696,N_23614);
and U24396 (N_24396,N_23880,N_23863);
or U24397 (N_24397,N_23644,N_23506);
nor U24398 (N_24398,N_23973,N_23236);
nand U24399 (N_24399,N_23042,N_23494);
or U24400 (N_24400,N_23945,N_23224);
nor U24401 (N_24401,N_23643,N_23656);
or U24402 (N_24402,N_23368,N_23688);
and U24403 (N_24403,N_23079,N_23790);
or U24404 (N_24404,N_23711,N_23704);
or U24405 (N_24405,N_23441,N_23148);
nand U24406 (N_24406,N_23423,N_23674);
or U24407 (N_24407,N_23645,N_23362);
nor U24408 (N_24408,N_23914,N_23548);
nor U24409 (N_24409,N_23434,N_23810);
nand U24410 (N_24410,N_23060,N_23347);
nor U24411 (N_24411,N_23475,N_23449);
nand U24412 (N_24412,N_23562,N_23180);
xnor U24413 (N_24413,N_23725,N_23961);
or U24414 (N_24414,N_23149,N_23843);
xnor U24415 (N_24415,N_23545,N_23439);
nor U24416 (N_24416,N_23231,N_23846);
or U24417 (N_24417,N_23587,N_23588);
or U24418 (N_24418,N_23472,N_23365);
or U24419 (N_24419,N_23205,N_23933);
and U24420 (N_24420,N_23925,N_23069);
or U24421 (N_24421,N_23685,N_23140);
nor U24422 (N_24422,N_23052,N_23776);
xor U24423 (N_24423,N_23730,N_23142);
nor U24424 (N_24424,N_23359,N_23201);
or U24425 (N_24425,N_23734,N_23123);
nor U24426 (N_24426,N_23111,N_23807);
nand U24427 (N_24427,N_23818,N_23130);
or U24428 (N_24428,N_23633,N_23873);
and U24429 (N_24429,N_23756,N_23769);
xnor U24430 (N_24430,N_23488,N_23088);
nand U24431 (N_24431,N_23981,N_23415);
nor U24432 (N_24432,N_23193,N_23687);
xor U24433 (N_24433,N_23839,N_23781);
and U24434 (N_24434,N_23876,N_23443);
nand U24435 (N_24435,N_23834,N_23959);
or U24436 (N_24436,N_23336,N_23159);
and U24437 (N_24437,N_23919,N_23071);
nand U24438 (N_24438,N_23485,N_23571);
nor U24439 (N_24439,N_23252,N_23438);
and U24440 (N_24440,N_23555,N_23453);
nor U24441 (N_24441,N_23513,N_23877);
and U24442 (N_24442,N_23760,N_23335);
xor U24443 (N_24443,N_23752,N_23669);
and U24444 (N_24444,N_23388,N_23318);
or U24445 (N_24445,N_23271,N_23972);
or U24446 (N_24446,N_23104,N_23155);
and U24447 (N_24447,N_23492,N_23316);
and U24448 (N_24448,N_23424,N_23984);
nor U24449 (N_24449,N_23331,N_23832);
nor U24450 (N_24450,N_23288,N_23986);
nand U24451 (N_24451,N_23989,N_23169);
xor U24452 (N_24452,N_23022,N_23958);
nand U24453 (N_24453,N_23217,N_23429);
nor U24454 (N_24454,N_23413,N_23373);
nor U24455 (N_24455,N_23828,N_23757);
nor U24456 (N_24456,N_23454,N_23573);
xnor U24457 (N_24457,N_23726,N_23327);
nand U24458 (N_24458,N_23267,N_23929);
or U24459 (N_24459,N_23835,N_23158);
nand U24460 (N_24460,N_23259,N_23412);
nor U24461 (N_24461,N_23249,N_23983);
nor U24462 (N_24462,N_23853,N_23463);
or U24463 (N_24463,N_23183,N_23745);
nor U24464 (N_24464,N_23269,N_23698);
nand U24465 (N_24465,N_23598,N_23056);
and U24466 (N_24466,N_23092,N_23138);
nor U24467 (N_24467,N_23039,N_23515);
xor U24468 (N_24468,N_23480,N_23840);
or U24469 (N_24469,N_23456,N_23214);
nand U24470 (N_24470,N_23068,N_23689);
and U24471 (N_24471,N_23418,N_23811);
or U24472 (N_24472,N_23977,N_23965);
nand U24473 (N_24473,N_23382,N_23215);
nand U24474 (N_24474,N_23383,N_23741);
nor U24475 (N_24475,N_23405,N_23508);
xor U24476 (N_24476,N_23974,N_23242);
and U24477 (N_24477,N_23001,N_23582);
nor U24478 (N_24478,N_23701,N_23226);
or U24479 (N_24479,N_23603,N_23838);
xnor U24480 (N_24480,N_23425,N_23394);
and U24481 (N_24481,N_23780,N_23110);
or U24482 (N_24482,N_23172,N_23399);
xnor U24483 (N_24483,N_23754,N_23247);
or U24484 (N_24484,N_23330,N_23892);
nor U24485 (N_24485,N_23632,N_23406);
or U24486 (N_24486,N_23884,N_23334);
xnor U24487 (N_24487,N_23928,N_23727);
nand U24488 (N_24488,N_23460,N_23655);
nand U24489 (N_24489,N_23489,N_23272);
or U24490 (N_24490,N_23755,N_23257);
nor U24491 (N_24491,N_23031,N_23957);
nand U24492 (N_24492,N_23550,N_23152);
nor U24493 (N_24493,N_23610,N_23640);
nand U24494 (N_24494,N_23833,N_23419);
or U24495 (N_24495,N_23759,N_23108);
xor U24496 (N_24496,N_23120,N_23583);
and U24497 (N_24497,N_23879,N_23611);
xor U24498 (N_24498,N_23464,N_23117);
and U24499 (N_24499,N_23493,N_23367);
and U24500 (N_24500,N_23401,N_23157);
or U24501 (N_24501,N_23095,N_23208);
or U24502 (N_24502,N_23127,N_23548);
xnor U24503 (N_24503,N_23811,N_23497);
and U24504 (N_24504,N_23901,N_23297);
nand U24505 (N_24505,N_23705,N_23654);
nor U24506 (N_24506,N_23670,N_23319);
nor U24507 (N_24507,N_23027,N_23742);
nand U24508 (N_24508,N_23728,N_23140);
nand U24509 (N_24509,N_23636,N_23555);
nand U24510 (N_24510,N_23556,N_23360);
nor U24511 (N_24511,N_23444,N_23974);
nor U24512 (N_24512,N_23307,N_23482);
xnor U24513 (N_24513,N_23855,N_23229);
nand U24514 (N_24514,N_23000,N_23405);
or U24515 (N_24515,N_23106,N_23742);
and U24516 (N_24516,N_23700,N_23261);
nand U24517 (N_24517,N_23541,N_23078);
nand U24518 (N_24518,N_23962,N_23984);
nand U24519 (N_24519,N_23441,N_23704);
xnor U24520 (N_24520,N_23525,N_23121);
nor U24521 (N_24521,N_23300,N_23319);
xnor U24522 (N_24522,N_23799,N_23017);
xor U24523 (N_24523,N_23526,N_23431);
xor U24524 (N_24524,N_23451,N_23110);
nand U24525 (N_24525,N_23235,N_23787);
xnor U24526 (N_24526,N_23428,N_23833);
xnor U24527 (N_24527,N_23797,N_23212);
xnor U24528 (N_24528,N_23491,N_23567);
or U24529 (N_24529,N_23876,N_23929);
nand U24530 (N_24530,N_23297,N_23593);
and U24531 (N_24531,N_23958,N_23162);
or U24532 (N_24532,N_23017,N_23977);
nor U24533 (N_24533,N_23908,N_23180);
and U24534 (N_24534,N_23052,N_23431);
or U24535 (N_24535,N_23069,N_23672);
or U24536 (N_24536,N_23553,N_23202);
xor U24537 (N_24537,N_23026,N_23223);
nand U24538 (N_24538,N_23105,N_23881);
nand U24539 (N_24539,N_23050,N_23110);
or U24540 (N_24540,N_23354,N_23679);
nand U24541 (N_24541,N_23163,N_23583);
or U24542 (N_24542,N_23977,N_23866);
nand U24543 (N_24543,N_23342,N_23729);
or U24544 (N_24544,N_23620,N_23415);
nor U24545 (N_24545,N_23651,N_23252);
and U24546 (N_24546,N_23856,N_23185);
and U24547 (N_24547,N_23151,N_23440);
and U24548 (N_24548,N_23253,N_23011);
nor U24549 (N_24549,N_23030,N_23411);
and U24550 (N_24550,N_23445,N_23952);
or U24551 (N_24551,N_23036,N_23644);
or U24552 (N_24552,N_23124,N_23612);
and U24553 (N_24553,N_23027,N_23311);
and U24554 (N_24554,N_23487,N_23951);
xnor U24555 (N_24555,N_23214,N_23762);
xnor U24556 (N_24556,N_23895,N_23473);
nor U24557 (N_24557,N_23666,N_23633);
and U24558 (N_24558,N_23352,N_23108);
xor U24559 (N_24559,N_23871,N_23614);
nand U24560 (N_24560,N_23921,N_23471);
nand U24561 (N_24561,N_23405,N_23837);
or U24562 (N_24562,N_23624,N_23734);
or U24563 (N_24563,N_23866,N_23308);
and U24564 (N_24564,N_23922,N_23248);
nand U24565 (N_24565,N_23309,N_23391);
or U24566 (N_24566,N_23463,N_23651);
nor U24567 (N_24567,N_23113,N_23261);
nand U24568 (N_24568,N_23625,N_23022);
nor U24569 (N_24569,N_23774,N_23056);
xnor U24570 (N_24570,N_23768,N_23401);
nor U24571 (N_24571,N_23728,N_23255);
xor U24572 (N_24572,N_23087,N_23627);
xnor U24573 (N_24573,N_23818,N_23637);
and U24574 (N_24574,N_23540,N_23053);
and U24575 (N_24575,N_23336,N_23946);
nor U24576 (N_24576,N_23144,N_23431);
xor U24577 (N_24577,N_23411,N_23899);
nand U24578 (N_24578,N_23609,N_23176);
nand U24579 (N_24579,N_23207,N_23543);
nor U24580 (N_24580,N_23258,N_23938);
and U24581 (N_24581,N_23996,N_23035);
xor U24582 (N_24582,N_23583,N_23119);
xnor U24583 (N_24583,N_23930,N_23521);
nor U24584 (N_24584,N_23671,N_23968);
nor U24585 (N_24585,N_23907,N_23433);
nor U24586 (N_24586,N_23866,N_23383);
or U24587 (N_24587,N_23073,N_23325);
and U24588 (N_24588,N_23108,N_23150);
nor U24589 (N_24589,N_23607,N_23838);
or U24590 (N_24590,N_23240,N_23229);
nand U24591 (N_24591,N_23220,N_23006);
or U24592 (N_24592,N_23277,N_23202);
or U24593 (N_24593,N_23534,N_23790);
xor U24594 (N_24594,N_23134,N_23372);
nor U24595 (N_24595,N_23763,N_23733);
nand U24596 (N_24596,N_23583,N_23151);
or U24597 (N_24597,N_23920,N_23972);
nor U24598 (N_24598,N_23130,N_23086);
nor U24599 (N_24599,N_23183,N_23849);
xnor U24600 (N_24600,N_23282,N_23487);
nand U24601 (N_24601,N_23978,N_23845);
and U24602 (N_24602,N_23319,N_23583);
nand U24603 (N_24603,N_23126,N_23048);
and U24604 (N_24604,N_23070,N_23767);
or U24605 (N_24605,N_23127,N_23011);
nor U24606 (N_24606,N_23754,N_23362);
or U24607 (N_24607,N_23190,N_23283);
nor U24608 (N_24608,N_23094,N_23373);
nor U24609 (N_24609,N_23746,N_23720);
or U24610 (N_24610,N_23695,N_23020);
nor U24611 (N_24611,N_23012,N_23649);
nor U24612 (N_24612,N_23751,N_23798);
nand U24613 (N_24613,N_23392,N_23414);
xor U24614 (N_24614,N_23515,N_23695);
nand U24615 (N_24615,N_23195,N_23267);
nand U24616 (N_24616,N_23772,N_23594);
nand U24617 (N_24617,N_23975,N_23162);
nand U24618 (N_24618,N_23965,N_23886);
and U24619 (N_24619,N_23674,N_23380);
nor U24620 (N_24620,N_23495,N_23217);
and U24621 (N_24621,N_23362,N_23884);
nor U24622 (N_24622,N_23013,N_23890);
xor U24623 (N_24623,N_23252,N_23312);
and U24624 (N_24624,N_23428,N_23218);
nand U24625 (N_24625,N_23500,N_23022);
xnor U24626 (N_24626,N_23393,N_23971);
nand U24627 (N_24627,N_23159,N_23655);
xnor U24628 (N_24628,N_23778,N_23226);
nor U24629 (N_24629,N_23076,N_23993);
or U24630 (N_24630,N_23883,N_23179);
xnor U24631 (N_24631,N_23003,N_23795);
nor U24632 (N_24632,N_23112,N_23717);
nand U24633 (N_24633,N_23710,N_23461);
nand U24634 (N_24634,N_23533,N_23502);
or U24635 (N_24635,N_23512,N_23801);
xor U24636 (N_24636,N_23380,N_23939);
xnor U24637 (N_24637,N_23927,N_23798);
nand U24638 (N_24638,N_23958,N_23357);
nand U24639 (N_24639,N_23567,N_23769);
nand U24640 (N_24640,N_23852,N_23018);
or U24641 (N_24641,N_23529,N_23310);
or U24642 (N_24642,N_23410,N_23108);
xor U24643 (N_24643,N_23198,N_23258);
nor U24644 (N_24644,N_23097,N_23022);
nand U24645 (N_24645,N_23598,N_23521);
and U24646 (N_24646,N_23105,N_23967);
and U24647 (N_24647,N_23075,N_23507);
and U24648 (N_24648,N_23703,N_23254);
nor U24649 (N_24649,N_23272,N_23734);
nor U24650 (N_24650,N_23029,N_23167);
nand U24651 (N_24651,N_23441,N_23472);
and U24652 (N_24652,N_23313,N_23117);
or U24653 (N_24653,N_23360,N_23688);
xnor U24654 (N_24654,N_23871,N_23799);
and U24655 (N_24655,N_23748,N_23931);
nand U24656 (N_24656,N_23123,N_23239);
nand U24657 (N_24657,N_23451,N_23440);
nor U24658 (N_24658,N_23197,N_23972);
or U24659 (N_24659,N_23200,N_23182);
nor U24660 (N_24660,N_23047,N_23186);
xnor U24661 (N_24661,N_23579,N_23295);
xor U24662 (N_24662,N_23264,N_23623);
nand U24663 (N_24663,N_23621,N_23060);
xor U24664 (N_24664,N_23622,N_23076);
and U24665 (N_24665,N_23443,N_23731);
nand U24666 (N_24666,N_23093,N_23718);
nor U24667 (N_24667,N_23886,N_23039);
and U24668 (N_24668,N_23029,N_23354);
nor U24669 (N_24669,N_23597,N_23156);
and U24670 (N_24670,N_23540,N_23311);
nor U24671 (N_24671,N_23589,N_23116);
and U24672 (N_24672,N_23576,N_23036);
nand U24673 (N_24673,N_23553,N_23887);
nand U24674 (N_24674,N_23534,N_23302);
nand U24675 (N_24675,N_23651,N_23601);
nand U24676 (N_24676,N_23972,N_23901);
xnor U24677 (N_24677,N_23505,N_23383);
or U24678 (N_24678,N_23897,N_23773);
nand U24679 (N_24679,N_23691,N_23307);
xnor U24680 (N_24680,N_23453,N_23689);
and U24681 (N_24681,N_23346,N_23167);
nand U24682 (N_24682,N_23529,N_23819);
or U24683 (N_24683,N_23827,N_23497);
xnor U24684 (N_24684,N_23850,N_23727);
nand U24685 (N_24685,N_23625,N_23151);
xnor U24686 (N_24686,N_23974,N_23303);
xor U24687 (N_24687,N_23033,N_23717);
nor U24688 (N_24688,N_23152,N_23164);
and U24689 (N_24689,N_23827,N_23750);
xnor U24690 (N_24690,N_23902,N_23071);
nor U24691 (N_24691,N_23820,N_23752);
nor U24692 (N_24692,N_23780,N_23564);
xor U24693 (N_24693,N_23430,N_23937);
and U24694 (N_24694,N_23096,N_23905);
or U24695 (N_24695,N_23139,N_23984);
and U24696 (N_24696,N_23162,N_23913);
and U24697 (N_24697,N_23499,N_23562);
nand U24698 (N_24698,N_23573,N_23410);
or U24699 (N_24699,N_23914,N_23663);
or U24700 (N_24700,N_23962,N_23085);
or U24701 (N_24701,N_23333,N_23033);
nor U24702 (N_24702,N_23780,N_23900);
nand U24703 (N_24703,N_23976,N_23909);
nor U24704 (N_24704,N_23348,N_23983);
or U24705 (N_24705,N_23176,N_23810);
xor U24706 (N_24706,N_23185,N_23531);
nand U24707 (N_24707,N_23865,N_23688);
and U24708 (N_24708,N_23065,N_23791);
nand U24709 (N_24709,N_23673,N_23164);
and U24710 (N_24710,N_23998,N_23143);
and U24711 (N_24711,N_23974,N_23637);
xnor U24712 (N_24712,N_23670,N_23809);
or U24713 (N_24713,N_23338,N_23972);
nand U24714 (N_24714,N_23722,N_23701);
nand U24715 (N_24715,N_23621,N_23340);
xnor U24716 (N_24716,N_23866,N_23846);
nand U24717 (N_24717,N_23610,N_23617);
or U24718 (N_24718,N_23165,N_23648);
and U24719 (N_24719,N_23511,N_23564);
or U24720 (N_24720,N_23500,N_23044);
and U24721 (N_24721,N_23191,N_23755);
and U24722 (N_24722,N_23341,N_23976);
nor U24723 (N_24723,N_23434,N_23296);
nor U24724 (N_24724,N_23356,N_23277);
or U24725 (N_24725,N_23663,N_23256);
or U24726 (N_24726,N_23378,N_23606);
nor U24727 (N_24727,N_23281,N_23420);
and U24728 (N_24728,N_23630,N_23654);
or U24729 (N_24729,N_23475,N_23561);
nand U24730 (N_24730,N_23424,N_23039);
nor U24731 (N_24731,N_23562,N_23779);
and U24732 (N_24732,N_23165,N_23544);
xnor U24733 (N_24733,N_23675,N_23910);
and U24734 (N_24734,N_23087,N_23223);
nor U24735 (N_24735,N_23290,N_23215);
xnor U24736 (N_24736,N_23254,N_23647);
or U24737 (N_24737,N_23751,N_23169);
or U24738 (N_24738,N_23867,N_23467);
nor U24739 (N_24739,N_23917,N_23603);
nor U24740 (N_24740,N_23915,N_23986);
nand U24741 (N_24741,N_23681,N_23079);
or U24742 (N_24742,N_23648,N_23914);
xnor U24743 (N_24743,N_23834,N_23839);
and U24744 (N_24744,N_23258,N_23535);
or U24745 (N_24745,N_23294,N_23160);
or U24746 (N_24746,N_23001,N_23657);
nand U24747 (N_24747,N_23350,N_23005);
nand U24748 (N_24748,N_23178,N_23157);
and U24749 (N_24749,N_23742,N_23575);
nor U24750 (N_24750,N_23429,N_23135);
or U24751 (N_24751,N_23898,N_23609);
xor U24752 (N_24752,N_23471,N_23984);
nand U24753 (N_24753,N_23829,N_23549);
or U24754 (N_24754,N_23649,N_23946);
nand U24755 (N_24755,N_23181,N_23026);
nor U24756 (N_24756,N_23441,N_23768);
nor U24757 (N_24757,N_23694,N_23189);
or U24758 (N_24758,N_23439,N_23151);
xor U24759 (N_24759,N_23991,N_23535);
or U24760 (N_24760,N_23314,N_23015);
nor U24761 (N_24761,N_23735,N_23606);
or U24762 (N_24762,N_23929,N_23061);
or U24763 (N_24763,N_23908,N_23259);
or U24764 (N_24764,N_23465,N_23845);
xor U24765 (N_24765,N_23371,N_23560);
and U24766 (N_24766,N_23393,N_23367);
nand U24767 (N_24767,N_23889,N_23443);
or U24768 (N_24768,N_23598,N_23789);
nand U24769 (N_24769,N_23408,N_23996);
or U24770 (N_24770,N_23077,N_23434);
and U24771 (N_24771,N_23649,N_23742);
or U24772 (N_24772,N_23375,N_23184);
nand U24773 (N_24773,N_23087,N_23433);
nand U24774 (N_24774,N_23732,N_23175);
or U24775 (N_24775,N_23285,N_23845);
xor U24776 (N_24776,N_23787,N_23137);
nand U24777 (N_24777,N_23353,N_23867);
nor U24778 (N_24778,N_23096,N_23709);
nor U24779 (N_24779,N_23135,N_23885);
xnor U24780 (N_24780,N_23941,N_23067);
and U24781 (N_24781,N_23876,N_23111);
or U24782 (N_24782,N_23403,N_23162);
and U24783 (N_24783,N_23308,N_23811);
and U24784 (N_24784,N_23784,N_23857);
nor U24785 (N_24785,N_23094,N_23286);
and U24786 (N_24786,N_23542,N_23963);
and U24787 (N_24787,N_23821,N_23542);
xor U24788 (N_24788,N_23363,N_23999);
nor U24789 (N_24789,N_23705,N_23460);
and U24790 (N_24790,N_23756,N_23369);
xor U24791 (N_24791,N_23091,N_23394);
nand U24792 (N_24792,N_23392,N_23989);
or U24793 (N_24793,N_23039,N_23390);
and U24794 (N_24794,N_23220,N_23959);
xor U24795 (N_24795,N_23631,N_23005);
nand U24796 (N_24796,N_23309,N_23335);
xor U24797 (N_24797,N_23736,N_23467);
nand U24798 (N_24798,N_23517,N_23848);
xor U24799 (N_24799,N_23287,N_23571);
nand U24800 (N_24800,N_23620,N_23946);
xnor U24801 (N_24801,N_23833,N_23775);
or U24802 (N_24802,N_23383,N_23075);
xor U24803 (N_24803,N_23361,N_23352);
nand U24804 (N_24804,N_23469,N_23015);
and U24805 (N_24805,N_23176,N_23689);
xor U24806 (N_24806,N_23903,N_23370);
or U24807 (N_24807,N_23234,N_23879);
xor U24808 (N_24808,N_23593,N_23843);
xor U24809 (N_24809,N_23778,N_23958);
xnor U24810 (N_24810,N_23225,N_23087);
or U24811 (N_24811,N_23072,N_23118);
or U24812 (N_24812,N_23474,N_23970);
and U24813 (N_24813,N_23482,N_23552);
or U24814 (N_24814,N_23936,N_23533);
or U24815 (N_24815,N_23188,N_23719);
xor U24816 (N_24816,N_23510,N_23835);
or U24817 (N_24817,N_23359,N_23845);
and U24818 (N_24818,N_23078,N_23306);
nor U24819 (N_24819,N_23680,N_23428);
nand U24820 (N_24820,N_23779,N_23555);
and U24821 (N_24821,N_23131,N_23762);
nor U24822 (N_24822,N_23609,N_23515);
nand U24823 (N_24823,N_23350,N_23388);
nor U24824 (N_24824,N_23528,N_23315);
xnor U24825 (N_24825,N_23954,N_23544);
nor U24826 (N_24826,N_23231,N_23034);
and U24827 (N_24827,N_23062,N_23984);
xnor U24828 (N_24828,N_23102,N_23263);
nor U24829 (N_24829,N_23857,N_23193);
nand U24830 (N_24830,N_23955,N_23017);
nand U24831 (N_24831,N_23386,N_23811);
nor U24832 (N_24832,N_23619,N_23057);
nand U24833 (N_24833,N_23967,N_23400);
or U24834 (N_24834,N_23825,N_23633);
xnor U24835 (N_24835,N_23719,N_23046);
xnor U24836 (N_24836,N_23769,N_23456);
nand U24837 (N_24837,N_23334,N_23865);
nand U24838 (N_24838,N_23415,N_23126);
xor U24839 (N_24839,N_23804,N_23384);
and U24840 (N_24840,N_23513,N_23371);
nand U24841 (N_24841,N_23125,N_23094);
nand U24842 (N_24842,N_23750,N_23596);
nand U24843 (N_24843,N_23536,N_23514);
and U24844 (N_24844,N_23717,N_23885);
xnor U24845 (N_24845,N_23829,N_23898);
nor U24846 (N_24846,N_23611,N_23425);
nand U24847 (N_24847,N_23482,N_23312);
xnor U24848 (N_24848,N_23504,N_23065);
nand U24849 (N_24849,N_23438,N_23253);
nand U24850 (N_24850,N_23056,N_23388);
nor U24851 (N_24851,N_23477,N_23239);
and U24852 (N_24852,N_23225,N_23987);
nand U24853 (N_24853,N_23285,N_23053);
nand U24854 (N_24854,N_23856,N_23241);
nor U24855 (N_24855,N_23695,N_23519);
nor U24856 (N_24856,N_23966,N_23818);
and U24857 (N_24857,N_23341,N_23443);
or U24858 (N_24858,N_23721,N_23402);
nor U24859 (N_24859,N_23473,N_23630);
and U24860 (N_24860,N_23110,N_23058);
or U24861 (N_24861,N_23572,N_23698);
xor U24862 (N_24862,N_23470,N_23160);
or U24863 (N_24863,N_23458,N_23010);
nand U24864 (N_24864,N_23557,N_23157);
xor U24865 (N_24865,N_23057,N_23719);
or U24866 (N_24866,N_23752,N_23222);
xor U24867 (N_24867,N_23344,N_23602);
nor U24868 (N_24868,N_23163,N_23277);
nor U24869 (N_24869,N_23821,N_23625);
or U24870 (N_24870,N_23096,N_23989);
and U24871 (N_24871,N_23950,N_23792);
and U24872 (N_24872,N_23421,N_23099);
and U24873 (N_24873,N_23613,N_23577);
and U24874 (N_24874,N_23983,N_23797);
nor U24875 (N_24875,N_23923,N_23022);
nand U24876 (N_24876,N_23063,N_23655);
xnor U24877 (N_24877,N_23270,N_23000);
nand U24878 (N_24878,N_23282,N_23756);
or U24879 (N_24879,N_23950,N_23504);
nor U24880 (N_24880,N_23163,N_23795);
xnor U24881 (N_24881,N_23269,N_23566);
or U24882 (N_24882,N_23194,N_23092);
and U24883 (N_24883,N_23683,N_23569);
and U24884 (N_24884,N_23505,N_23587);
xnor U24885 (N_24885,N_23434,N_23975);
xnor U24886 (N_24886,N_23683,N_23546);
nand U24887 (N_24887,N_23611,N_23055);
xor U24888 (N_24888,N_23961,N_23760);
and U24889 (N_24889,N_23168,N_23884);
nand U24890 (N_24890,N_23069,N_23313);
or U24891 (N_24891,N_23676,N_23156);
and U24892 (N_24892,N_23653,N_23849);
nand U24893 (N_24893,N_23712,N_23351);
and U24894 (N_24894,N_23776,N_23961);
nand U24895 (N_24895,N_23219,N_23580);
or U24896 (N_24896,N_23077,N_23113);
or U24897 (N_24897,N_23798,N_23756);
xor U24898 (N_24898,N_23897,N_23466);
and U24899 (N_24899,N_23482,N_23274);
xor U24900 (N_24900,N_23435,N_23979);
nand U24901 (N_24901,N_23181,N_23479);
xor U24902 (N_24902,N_23679,N_23757);
xnor U24903 (N_24903,N_23518,N_23970);
nor U24904 (N_24904,N_23956,N_23966);
nand U24905 (N_24905,N_23046,N_23440);
or U24906 (N_24906,N_23097,N_23205);
xor U24907 (N_24907,N_23255,N_23689);
nand U24908 (N_24908,N_23916,N_23389);
or U24909 (N_24909,N_23917,N_23901);
or U24910 (N_24910,N_23670,N_23631);
nor U24911 (N_24911,N_23181,N_23059);
and U24912 (N_24912,N_23386,N_23759);
nor U24913 (N_24913,N_23100,N_23361);
xor U24914 (N_24914,N_23570,N_23614);
nor U24915 (N_24915,N_23304,N_23192);
or U24916 (N_24916,N_23708,N_23917);
nor U24917 (N_24917,N_23128,N_23258);
or U24918 (N_24918,N_23015,N_23937);
nand U24919 (N_24919,N_23391,N_23797);
xnor U24920 (N_24920,N_23149,N_23971);
nand U24921 (N_24921,N_23131,N_23686);
nand U24922 (N_24922,N_23397,N_23981);
or U24923 (N_24923,N_23288,N_23095);
nand U24924 (N_24924,N_23221,N_23409);
and U24925 (N_24925,N_23894,N_23166);
xnor U24926 (N_24926,N_23705,N_23926);
nand U24927 (N_24927,N_23642,N_23033);
and U24928 (N_24928,N_23012,N_23568);
nor U24929 (N_24929,N_23085,N_23517);
xor U24930 (N_24930,N_23685,N_23384);
and U24931 (N_24931,N_23205,N_23087);
nand U24932 (N_24932,N_23683,N_23973);
nand U24933 (N_24933,N_23794,N_23009);
and U24934 (N_24934,N_23487,N_23432);
xnor U24935 (N_24935,N_23595,N_23980);
nand U24936 (N_24936,N_23291,N_23654);
and U24937 (N_24937,N_23570,N_23966);
nor U24938 (N_24938,N_23192,N_23488);
xor U24939 (N_24939,N_23687,N_23943);
and U24940 (N_24940,N_23481,N_23291);
nor U24941 (N_24941,N_23863,N_23576);
nand U24942 (N_24942,N_23569,N_23503);
and U24943 (N_24943,N_23439,N_23218);
and U24944 (N_24944,N_23556,N_23052);
nor U24945 (N_24945,N_23728,N_23303);
xnor U24946 (N_24946,N_23587,N_23966);
or U24947 (N_24947,N_23040,N_23417);
xor U24948 (N_24948,N_23744,N_23961);
nor U24949 (N_24949,N_23253,N_23890);
nor U24950 (N_24950,N_23815,N_23408);
nor U24951 (N_24951,N_23880,N_23369);
xor U24952 (N_24952,N_23141,N_23645);
nor U24953 (N_24953,N_23689,N_23534);
or U24954 (N_24954,N_23528,N_23961);
xor U24955 (N_24955,N_23171,N_23412);
and U24956 (N_24956,N_23047,N_23410);
and U24957 (N_24957,N_23430,N_23542);
and U24958 (N_24958,N_23453,N_23916);
xor U24959 (N_24959,N_23828,N_23912);
and U24960 (N_24960,N_23453,N_23408);
nand U24961 (N_24961,N_23069,N_23622);
and U24962 (N_24962,N_23135,N_23899);
or U24963 (N_24963,N_23596,N_23031);
and U24964 (N_24964,N_23252,N_23381);
xor U24965 (N_24965,N_23914,N_23670);
or U24966 (N_24966,N_23885,N_23819);
and U24967 (N_24967,N_23812,N_23097);
or U24968 (N_24968,N_23320,N_23467);
or U24969 (N_24969,N_23337,N_23777);
xor U24970 (N_24970,N_23224,N_23070);
xnor U24971 (N_24971,N_23151,N_23606);
and U24972 (N_24972,N_23651,N_23849);
and U24973 (N_24973,N_23618,N_23232);
nor U24974 (N_24974,N_23486,N_23402);
and U24975 (N_24975,N_23991,N_23172);
and U24976 (N_24976,N_23379,N_23778);
and U24977 (N_24977,N_23982,N_23055);
nor U24978 (N_24978,N_23186,N_23359);
and U24979 (N_24979,N_23682,N_23149);
xor U24980 (N_24980,N_23403,N_23166);
or U24981 (N_24981,N_23493,N_23783);
xnor U24982 (N_24982,N_23486,N_23435);
or U24983 (N_24983,N_23443,N_23276);
or U24984 (N_24984,N_23660,N_23972);
nor U24985 (N_24985,N_23116,N_23547);
nand U24986 (N_24986,N_23532,N_23944);
and U24987 (N_24987,N_23853,N_23764);
and U24988 (N_24988,N_23431,N_23620);
and U24989 (N_24989,N_23743,N_23429);
nand U24990 (N_24990,N_23342,N_23657);
or U24991 (N_24991,N_23960,N_23071);
and U24992 (N_24992,N_23249,N_23845);
or U24993 (N_24993,N_23773,N_23230);
and U24994 (N_24994,N_23387,N_23307);
xnor U24995 (N_24995,N_23131,N_23418);
nand U24996 (N_24996,N_23537,N_23037);
nand U24997 (N_24997,N_23813,N_23517);
and U24998 (N_24998,N_23983,N_23022);
xor U24999 (N_24999,N_23222,N_23475);
or UO_0 (O_0,N_24371,N_24273);
and UO_1 (O_1,N_24598,N_24465);
xnor UO_2 (O_2,N_24986,N_24332);
nor UO_3 (O_3,N_24917,N_24216);
nand UO_4 (O_4,N_24961,N_24594);
nand UO_5 (O_5,N_24888,N_24788);
nor UO_6 (O_6,N_24786,N_24797);
nor UO_7 (O_7,N_24923,N_24787);
xor UO_8 (O_8,N_24068,N_24637);
and UO_9 (O_9,N_24079,N_24102);
nor UO_10 (O_10,N_24973,N_24744);
or UO_11 (O_11,N_24354,N_24632);
xor UO_12 (O_12,N_24702,N_24568);
nand UO_13 (O_13,N_24667,N_24946);
xnor UO_14 (O_14,N_24051,N_24010);
and UO_15 (O_15,N_24883,N_24101);
nand UO_16 (O_16,N_24860,N_24827);
nor UO_17 (O_17,N_24967,N_24815);
nand UO_18 (O_18,N_24331,N_24731);
or UO_19 (O_19,N_24446,N_24935);
nor UO_20 (O_20,N_24028,N_24413);
and UO_21 (O_21,N_24498,N_24355);
or UO_22 (O_22,N_24211,N_24109);
and UO_23 (O_23,N_24557,N_24049);
xnor UO_24 (O_24,N_24151,N_24514);
nand UO_25 (O_25,N_24839,N_24877);
nand UO_26 (O_26,N_24255,N_24714);
xnor UO_27 (O_27,N_24018,N_24526);
nor UO_28 (O_28,N_24031,N_24662);
xor UO_29 (O_29,N_24328,N_24751);
and UO_30 (O_30,N_24416,N_24892);
xor UO_31 (O_31,N_24444,N_24604);
and UO_32 (O_32,N_24197,N_24295);
xor UO_33 (O_33,N_24811,N_24750);
and UO_34 (O_34,N_24174,N_24466);
xnor UO_35 (O_35,N_24482,N_24324);
xnor UO_36 (O_36,N_24554,N_24025);
nand UO_37 (O_37,N_24265,N_24032);
nand UO_38 (O_38,N_24403,N_24696);
xor UO_39 (O_39,N_24183,N_24645);
nor UO_40 (O_40,N_24358,N_24312);
nor UO_41 (O_41,N_24374,N_24362);
or UO_42 (O_42,N_24175,N_24301);
or UO_43 (O_43,N_24424,N_24882);
or UO_44 (O_44,N_24959,N_24274);
or UO_45 (O_45,N_24707,N_24552);
or UO_46 (O_46,N_24014,N_24932);
or UO_47 (O_47,N_24812,N_24726);
or UO_48 (O_48,N_24740,N_24529);
nand UO_49 (O_49,N_24123,N_24914);
nand UO_50 (O_50,N_24422,N_24437);
xnor UO_51 (O_51,N_24075,N_24414);
xor UO_52 (O_52,N_24614,N_24131);
or UO_53 (O_53,N_24067,N_24962);
nand UO_54 (O_54,N_24640,N_24804);
or UO_55 (O_55,N_24938,N_24314);
nor UO_56 (O_56,N_24921,N_24375);
nor UO_57 (O_57,N_24347,N_24343);
xor UO_58 (O_58,N_24583,N_24166);
nand UO_59 (O_59,N_24236,N_24539);
nor UO_60 (O_60,N_24542,N_24323);
and UO_61 (O_61,N_24623,N_24538);
xor UO_62 (O_62,N_24289,N_24567);
and UO_63 (O_63,N_24344,N_24098);
and UO_64 (O_64,N_24257,N_24810);
or UO_65 (O_65,N_24243,N_24758);
or UO_66 (O_66,N_24103,N_24125);
nand UO_67 (O_67,N_24580,N_24991);
nand UO_68 (O_68,N_24821,N_24115);
nand UO_69 (O_69,N_24525,N_24412);
or UO_70 (O_70,N_24199,N_24763);
or UO_71 (O_71,N_24579,N_24220);
nand UO_72 (O_72,N_24884,N_24681);
nand UO_73 (O_73,N_24384,N_24288);
xor UO_74 (O_74,N_24572,N_24137);
or UO_75 (O_75,N_24253,N_24974);
and UO_76 (O_76,N_24352,N_24616);
nor UO_77 (O_77,N_24448,N_24447);
and UO_78 (O_78,N_24369,N_24474);
nand UO_79 (O_79,N_24957,N_24370);
and UO_80 (O_80,N_24613,N_24864);
nand UO_81 (O_81,N_24802,N_24041);
and UO_82 (O_82,N_24820,N_24644);
and UO_83 (O_83,N_24895,N_24890);
and UO_84 (O_84,N_24182,N_24309);
nor UO_85 (O_85,N_24718,N_24672);
nor UO_86 (O_86,N_24022,N_24953);
nor UO_87 (O_87,N_24776,N_24187);
or UO_88 (O_88,N_24795,N_24478);
xnor UO_89 (O_89,N_24642,N_24249);
or UO_90 (O_90,N_24473,N_24631);
nand UO_91 (O_91,N_24655,N_24300);
and UO_92 (O_92,N_24509,N_24879);
and UO_93 (O_93,N_24052,N_24082);
nand UO_94 (O_94,N_24303,N_24336);
and UO_95 (O_95,N_24210,N_24649);
nor UO_96 (O_96,N_24924,N_24907);
xor UO_97 (O_97,N_24784,N_24972);
and UO_98 (O_98,N_24545,N_24831);
nand UO_99 (O_99,N_24927,N_24195);
nor UO_100 (O_100,N_24268,N_24334);
and UO_101 (O_101,N_24673,N_24984);
xnor UO_102 (O_102,N_24368,N_24517);
and UO_103 (O_103,N_24327,N_24144);
nand UO_104 (O_104,N_24227,N_24700);
nor UO_105 (O_105,N_24979,N_24765);
xor UO_106 (O_106,N_24126,N_24593);
or UO_107 (O_107,N_24335,N_24162);
nand UO_108 (O_108,N_24149,N_24925);
nor UO_109 (O_109,N_24852,N_24348);
nand UO_110 (O_110,N_24383,N_24597);
nor UO_111 (O_111,N_24987,N_24377);
and UO_112 (O_112,N_24099,N_24430);
nand UO_113 (O_113,N_24004,N_24484);
and UO_114 (O_114,N_24639,N_24290);
nand UO_115 (O_115,N_24070,N_24163);
nand UO_116 (O_116,N_24218,N_24767);
nor UO_117 (O_117,N_24558,N_24318);
and UO_118 (O_118,N_24942,N_24706);
and UO_119 (O_119,N_24676,N_24873);
and UO_120 (O_120,N_24561,N_24061);
nand UO_121 (O_121,N_24592,N_24179);
xor UO_122 (O_122,N_24747,N_24503);
and UO_123 (O_123,N_24191,N_24445);
or UO_124 (O_124,N_24398,N_24760);
xor UO_125 (O_125,N_24746,N_24741);
and UO_126 (O_126,N_24634,N_24536);
and UO_127 (O_127,N_24922,N_24993);
or UO_128 (O_128,N_24994,N_24002);
or UO_129 (O_129,N_24172,N_24429);
and UO_130 (O_130,N_24160,N_24408);
nand UO_131 (O_131,N_24678,N_24133);
nor UO_132 (O_132,N_24563,N_24512);
xnor UO_133 (O_133,N_24724,N_24748);
xnor UO_134 (O_134,N_24511,N_24493);
or UO_135 (O_135,N_24845,N_24073);
xor UO_136 (O_136,N_24038,N_24796);
nor UO_137 (O_137,N_24366,N_24725);
xnor UO_138 (O_138,N_24194,N_24854);
nand UO_139 (O_139,N_24752,N_24341);
or UO_140 (O_140,N_24995,N_24527);
nor UO_141 (O_141,N_24338,N_24768);
nand UO_142 (O_142,N_24564,N_24190);
and UO_143 (O_143,N_24277,N_24252);
xor UO_144 (O_144,N_24982,N_24515);
and UO_145 (O_145,N_24584,N_24628);
or UO_146 (O_146,N_24799,N_24200);
nor UO_147 (O_147,N_24705,N_24127);
nor UO_148 (O_148,N_24985,N_24933);
and UO_149 (O_149,N_24822,N_24129);
and UO_150 (O_150,N_24944,N_24235);
or UO_151 (O_151,N_24035,N_24048);
or UO_152 (O_152,N_24231,N_24260);
nor UO_153 (O_153,N_24086,N_24629);
and UO_154 (O_154,N_24855,N_24307);
xor UO_155 (O_155,N_24222,N_24588);
nor UO_156 (O_156,N_24105,N_24550);
nor UO_157 (O_157,N_24551,N_24945);
or UO_158 (O_158,N_24510,N_24116);
xor UO_159 (O_159,N_24999,N_24606);
or UO_160 (O_160,N_24089,N_24248);
nor UO_161 (O_161,N_24697,N_24192);
nand UO_162 (O_162,N_24169,N_24060);
nor UO_163 (O_163,N_24980,N_24113);
xor UO_164 (O_164,N_24595,N_24427);
or UO_165 (O_165,N_24139,N_24459);
xnor UO_166 (O_166,N_24836,N_24963);
and UO_167 (O_167,N_24045,N_24057);
nand UO_168 (O_168,N_24023,N_24516);
or UO_169 (O_169,N_24769,N_24150);
nand UO_170 (O_170,N_24544,N_24078);
and UO_171 (O_171,N_24585,N_24528);
and UO_172 (O_172,N_24540,N_24017);
nor UO_173 (O_173,N_24997,N_24012);
xnor UO_174 (O_174,N_24739,N_24112);
or UO_175 (O_175,N_24766,N_24793);
and UO_176 (O_176,N_24059,N_24443);
or UO_177 (O_177,N_24117,N_24615);
or UO_178 (O_178,N_24165,N_24330);
or UO_179 (O_179,N_24633,N_24256);
and UO_180 (O_180,N_24781,N_24915);
or UO_181 (O_181,N_24505,N_24055);
and UO_182 (O_182,N_24770,N_24759);
nor UO_183 (O_183,N_24656,N_24651);
or UO_184 (O_184,N_24727,N_24612);
nand UO_185 (O_185,N_24212,N_24148);
or UO_186 (O_186,N_24111,N_24899);
or UO_187 (O_187,N_24990,N_24833);
xnor UO_188 (O_188,N_24738,N_24381);
nor UO_189 (O_189,N_24054,N_24847);
nor UO_190 (O_190,N_24620,N_24617);
xor UO_191 (O_191,N_24684,N_24680);
and UO_192 (O_192,N_24607,N_24134);
or UO_193 (O_193,N_24161,N_24842);
and UO_194 (O_194,N_24121,N_24704);
nor UO_195 (O_195,N_24521,N_24805);
and UO_196 (O_196,N_24732,N_24547);
xor UO_197 (O_197,N_24896,N_24610);
or UO_198 (O_198,N_24287,N_24889);
nand UO_199 (O_199,N_24088,N_24155);
xnor UO_200 (O_200,N_24723,N_24185);
nor UO_201 (O_201,N_24382,N_24909);
nand UO_202 (O_202,N_24954,N_24494);
or UO_203 (O_203,N_24306,N_24351);
or UO_204 (O_204,N_24659,N_24830);
or UO_205 (O_205,N_24092,N_24988);
or UO_206 (O_206,N_24270,N_24170);
nor UO_207 (O_207,N_24001,N_24221);
or UO_208 (O_208,N_24091,N_24874);
nor UO_209 (O_209,N_24489,N_24589);
and UO_210 (O_210,N_24152,N_24006);
xnor UO_211 (O_211,N_24504,N_24138);
xor UO_212 (O_212,N_24215,N_24244);
xor UO_213 (O_213,N_24910,N_24817);
or UO_214 (O_214,N_24020,N_24457);
or UO_215 (O_215,N_24276,N_24154);
and UO_216 (O_216,N_24479,N_24213);
nand UO_217 (O_217,N_24428,N_24124);
xor UO_218 (O_218,N_24357,N_24066);
nor UO_219 (O_219,N_24771,N_24208);
nand UO_220 (O_220,N_24407,N_24657);
and UO_221 (O_221,N_24838,N_24562);
or UO_222 (O_222,N_24904,N_24928);
and UO_223 (O_223,N_24167,N_24500);
nor UO_224 (O_224,N_24887,N_24581);
nor UO_225 (O_225,N_24491,N_24431);
and UO_226 (O_226,N_24916,N_24626);
nand UO_227 (O_227,N_24173,N_24027);
nor UO_228 (O_228,N_24559,N_24966);
and UO_229 (O_229,N_24378,N_24016);
nand UO_230 (O_230,N_24843,N_24577);
and UO_231 (O_231,N_24549,N_24029);
nor UO_232 (O_232,N_24764,N_24685);
xnor UO_233 (O_233,N_24201,N_24261);
nor UO_234 (O_234,N_24266,N_24326);
xnor UO_235 (O_235,N_24828,N_24141);
nand UO_236 (O_236,N_24095,N_24541);
and UO_237 (O_237,N_24578,N_24044);
nor UO_238 (O_238,N_24114,N_24247);
xor UO_239 (O_239,N_24647,N_24468);
and UO_240 (O_240,N_24275,N_24271);
xor UO_241 (O_241,N_24453,N_24926);
xor UO_242 (O_242,N_24147,N_24069);
or UO_243 (O_243,N_24209,N_24686);
nand UO_244 (O_244,N_24469,N_24872);
xor UO_245 (O_245,N_24841,N_24813);
and UO_246 (O_246,N_24906,N_24886);
and UO_247 (O_247,N_24450,N_24780);
nand UO_248 (O_248,N_24792,N_24036);
nor UO_249 (O_249,N_24600,N_24322);
nand UO_250 (O_250,N_24865,N_24533);
nor UO_251 (O_251,N_24046,N_24423);
nor UO_252 (O_252,N_24761,N_24483);
or UO_253 (O_253,N_24436,N_24487);
and UO_254 (O_254,N_24868,N_24292);
xnor UO_255 (O_255,N_24043,N_24867);
or UO_256 (O_256,N_24958,N_24778);
nor UO_257 (O_257,N_24388,N_24693);
nor UO_258 (O_258,N_24376,N_24464);
xnor UO_259 (O_259,N_24880,N_24385);
nor UO_260 (O_260,N_24230,N_24263);
xnor UO_261 (O_261,N_24107,N_24128);
nand UO_262 (O_262,N_24785,N_24941);
nand UO_263 (O_263,N_24602,N_24421);
nor UO_264 (O_264,N_24582,N_24294);
nand UO_265 (O_265,N_24721,N_24219);
or UO_266 (O_266,N_24586,N_24232);
nand UO_267 (O_267,N_24308,N_24319);
xor UO_268 (O_268,N_24217,N_24021);
or UO_269 (O_269,N_24814,N_24406);
and UO_270 (O_270,N_24948,N_24519);
nand UO_271 (O_271,N_24096,N_24456);
nand UO_272 (O_272,N_24432,N_24142);
or UO_273 (O_273,N_24524,N_24901);
nor UO_274 (O_274,N_24665,N_24492);
xnor UO_275 (O_275,N_24898,N_24729);
nand UO_276 (O_276,N_24861,N_24463);
and UO_277 (O_277,N_24159,N_24790);
and UO_278 (O_278,N_24692,N_24798);
nor UO_279 (O_279,N_24844,N_24866);
nand UO_280 (O_280,N_24284,N_24690);
xnor UO_281 (O_281,N_24005,N_24264);
or UO_282 (O_282,N_24819,N_24522);
or UO_283 (O_283,N_24574,N_24543);
and UO_284 (O_284,N_24238,N_24507);
nor UO_285 (O_285,N_24053,N_24703);
nor UO_286 (O_286,N_24998,N_24699);
xor UO_287 (O_287,N_24401,N_24283);
and UO_288 (O_288,N_24698,N_24900);
nor UO_289 (O_289,N_24392,N_24387);
xor UO_290 (O_290,N_24304,N_24791);
nand UO_291 (O_291,N_24203,N_24919);
or UO_292 (O_292,N_24342,N_24080);
and UO_293 (O_293,N_24871,N_24609);
xor UO_294 (O_294,N_24461,N_24772);
xor UO_295 (O_295,N_24119,N_24030);
nor UO_296 (O_296,N_24939,N_24940);
nor UO_297 (O_297,N_24426,N_24736);
and UO_298 (O_298,N_24269,N_24710);
and UO_299 (O_299,N_24278,N_24638);
or UO_300 (O_300,N_24019,N_24011);
and UO_301 (O_301,N_24625,N_24390);
nor UO_302 (O_302,N_24094,N_24876);
nand UO_303 (O_303,N_24809,N_24630);
nand UO_304 (O_304,N_24960,N_24816);
and UO_305 (O_305,N_24618,N_24186);
or UO_306 (O_306,N_24688,N_24789);
and UO_307 (O_307,N_24571,N_24653);
xnor UO_308 (O_308,N_24202,N_24346);
and UO_309 (O_309,N_24291,N_24952);
nand UO_310 (O_310,N_24003,N_24272);
nor UO_311 (O_311,N_24237,N_24196);
nand UO_312 (O_312,N_24970,N_24885);
nor UO_313 (O_313,N_24850,N_24929);
and UO_314 (O_314,N_24118,N_24405);
or UO_315 (O_315,N_24320,N_24989);
nand UO_316 (O_316,N_24480,N_24008);
nand UO_317 (O_317,N_24379,N_24333);
and UO_318 (O_318,N_24259,N_24176);
xor UO_319 (O_319,N_24394,N_24675);
nand UO_320 (O_320,N_24282,N_24846);
or UO_321 (O_321,N_24762,N_24189);
nor UO_322 (O_322,N_24496,N_24104);
xnor UO_323 (O_323,N_24683,N_24591);
nand UO_324 (O_324,N_24267,N_24110);
nand UO_325 (O_325,N_24757,N_24532);
nand UO_326 (O_326,N_24576,N_24039);
and UO_327 (O_327,N_24878,N_24977);
xnor UO_328 (O_328,N_24475,N_24404);
or UO_329 (O_329,N_24367,N_24730);
xnor UO_330 (O_330,N_24783,N_24353);
nor UO_331 (O_331,N_24090,N_24438);
or UO_332 (O_332,N_24801,N_24951);
nor UO_333 (O_333,N_24596,N_24477);
and UO_334 (O_334,N_24298,N_24490);
or UO_335 (O_335,N_24937,N_24229);
and UO_336 (O_336,N_24184,N_24902);
nand UO_337 (O_337,N_24824,N_24402);
nor UO_338 (O_338,N_24250,N_24207);
nand UO_339 (O_339,N_24181,N_24934);
or UO_340 (O_340,N_24233,N_24978);
xor UO_341 (O_341,N_24755,N_24299);
nor UO_342 (O_342,N_24848,N_24835);
or UO_343 (O_343,N_24666,N_24223);
nor UO_344 (O_344,N_24992,N_24800);
xnor UO_345 (O_345,N_24063,N_24132);
nor UO_346 (O_346,N_24495,N_24565);
and UO_347 (O_347,N_24968,N_24599);
nand UO_348 (O_348,N_24034,N_24246);
or UO_349 (O_349,N_24439,N_24071);
nand UO_350 (O_350,N_24621,N_24360);
nand UO_351 (O_351,N_24100,N_24520);
and UO_352 (O_352,N_24782,N_24745);
xnor UO_353 (O_353,N_24773,N_24411);
and UO_354 (O_354,N_24140,N_24711);
or UO_355 (O_355,N_24654,N_24000);
xor UO_356 (O_356,N_24234,N_24316);
nor UO_357 (O_357,N_24349,N_24420);
or UO_358 (O_358,N_24911,N_24258);
nor UO_359 (O_359,N_24410,N_24310);
nor UO_360 (O_360,N_24241,N_24826);
and UO_361 (O_361,N_24168,N_24534);
nand UO_362 (O_362,N_24779,N_24449);
xnor UO_363 (O_363,N_24513,N_24863);
xor UO_364 (O_364,N_24661,N_24930);
or UO_365 (O_365,N_24084,N_24396);
xor UO_366 (O_366,N_24971,N_24329);
xor UO_367 (O_367,N_24658,N_24712);
nand UO_368 (O_368,N_24587,N_24857);
or UO_369 (O_369,N_24689,N_24364);
and UO_370 (O_370,N_24254,N_24156);
or UO_371 (O_371,N_24013,N_24774);
xnor UO_372 (O_372,N_24452,N_24840);
nand UO_373 (O_373,N_24476,N_24546);
xor UO_374 (O_374,N_24918,N_24501);
nor UO_375 (O_375,N_24389,N_24239);
xor UO_376 (O_376,N_24713,N_24359);
xor UO_377 (O_377,N_24337,N_24743);
nand UO_378 (O_378,N_24636,N_24064);
or UO_379 (O_379,N_24499,N_24646);
xnor UO_380 (O_380,N_24419,N_24893);
nor UO_381 (O_381,N_24749,N_24380);
and UO_382 (O_382,N_24891,N_24641);
nor UO_383 (O_383,N_24093,N_24603);
or UO_384 (O_384,N_24471,N_24807);
or UO_385 (O_385,N_24853,N_24262);
nor UO_386 (O_386,N_24363,N_24734);
nor UO_387 (O_387,N_24399,N_24671);
nand UO_388 (O_388,N_24733,N_24936);
nor UO_389 (O_389,N_24317,N_24856);
xor UO_390 (O_390,N_24417,N_24293);
nand UO_391 (O_391,N_24719,N_24566);
or UO_392 (O_392,N_24350,N_24981);
and UO_393 (O_393,N_24903,N_24386);
nor UO_394 (O_394,N_24440,N_24074);
xnor UO_395 (O_395,N_24722,N_24135);
or UO_396 (O_396,N_24481,N_24775);
and UO_397 (O_397,N_24570,N_24643);
and UO_398 (O_398,N_24302,N_24920);
and UO_399 (O_399,N_24130,N_24619);
nand UO_400 (O_400,N_24556,N_24040);
nor UO_401 (O_401,N_24434,N_24305);
nor UO_402 (O_402,N_24047,N_24224);
and UO_403 (O_403,N_24669,N_24897);
nand UO_404 (O_404,N_24315,N_24026);
nor UO_405 (O_405,N_24087,N_24829);
nor UO_406 (O_406,N_24859,N_24969);
nand UO_407 (O_407,N_24530,N_24372);
xor UO_408 (O_408,N_24356,N_24171);
or UO_409 (O_409,N_24297,N_24339);
or UO_410 (O_410,N_24754,N_24691);
nor UO_411 (O_411,N_24393,N_24679);
and UO_412 (O_412,N_24214,N_24056);
nand UO_413 (O_413,N_24949,N_24321);
or UO_414 (O_414,N_24996,N_24177);
and UO_415 (O_415,N_24240,N_24225);
or UO_416 (O_416,N_24205,N_24875);
xnor UO_417 (O_417,N_24687,N_24286);
or UO_418 (O_418,N_24818,N_24956);
nor UO_419 (O_419,N_24143,N_24664);
nor UO_420 (O_420,N_24083,N_24905);
or UO_421 (O_421,N_24106,N_24881);
or UO_422 (O_422,N_24590,N_24180);
and UO_423 (O_423,N_24279,N_24024);
and UO_424 (O_424,N_24467,N_24870);
xnor UO_425 (O_425,N_24825,N_24497);
xor UO_426 (O_426,N_24553,N_24442);
or UO_427 (O_427,N_24136,N_24280);
and UO_428 (O_428,N_24325,N_24108);
xor UO_429 (O_429,N_24085,N_24837);
nand UO_430 (O_430,N_24983,N_24573);
nor UO_431 (O_431,N_24146,N_24508);
or UO_432 (O_432,N_24397,N_24622);
nand UO_433 (O_433,N_24624,N_24009);
nor UO_434 (O_434,N_24178,N_24803);
nor UO_435 (O_435,N_24608,N_24976);
or UO_436 (O_436,N_24373,N_24455);
nand UO_437 (O_437,N_24834,N_24122);
or UO_438 (O_438,N_24648,N_24943);
nand UO_439 (O_439,N_24451,N_24204);
and UO_440 (O_440,N_24652,N_24157);
and UO_441 (O_441,N_24361,N_24605);
xor UO_442 (O_442,N_24964,N_24296);
xor UO_443 (O_443,N_24717,N_24228);
nand UO_444 (O_444,N_24913,N_24145);
and UO_445 (O_445,N_24502,N_24715);
or UO_446 (O_446,N_24081,N_24735);
xnor UO_447 (O_447,N_24164,N_24832);
xor UO_448 (O_448,N_24947,N_24472);
and UO_449 (O_449,N_24756,N_24097);
or UO_450 (O_450,N_24415,N_24535);
or UO_451 (O_451,N_24950,N_24486);
and UO_452 (O_452,N_24340,N_24242);
nor UO_453 (O_453,N_24742,N_24050);
xor UO_454 (O_454,N_24708,N_24460);
xnor UO_455 (O_455,N_24753,N_24650);
nor UO_456 (O_456,N_24458,N_24077);
nand UO_457 (O_457,N_24120,N_24462);
nand UO_458 (O_458,N_24226,N_24931);
nand UO_459 (O_459,N_24193,N_24033);
xnor UO_460 (O_460,N_24670,N_24965);
or UO_461 (O_461,N_24015,N_24668);
nand UO_462 (O_462,N_24058,N_24794);
or UO_463 (O_463,N_24548,N_24485);
nor UO_464 (O_464,N_24007,N_24285);
and UO_465 (O_465,N_24065,N_24400);
nand UO_466 (O_466,N_24206,N_24869);
or UO_467 (O_467,N_24635,N_24601);
nor UO_468 (O_468,N_24042,N_24806);
nand UO_469 (O_469,N_24158,N_24955);
or UO_470 (O_470,N_24720,N_24409);
or UO_471 (O_471,N_24076,N_24858);
or UO_472 (O_472,N_24518,N_24808);
and UO_473 (O_473,N_24488,N_24777);
nor UO_474 (O_474,N_24365,N_24345);
and UO_475 (O_475,N_24245,N_24062);
xor UO_476 (O_476,N_24523,N_24531);
or UO_477 (O_477,N_24709,N_24894);
xnor UO_478 (O_478,N_24441,N_24454);
or UO_479 (O_479,N_24701,N_24037);
or UO_480 (O_480,N_24569,N_24418);
nor UO_481 (O_481,N_24072,N_24823);
nor UO_482 (O_482,N_24575,N_24311);
and UO_483 (O_483,N_24682,N_24313);
nand UO_484 (O_484,N_24660,N_24851);
nor UO_485 (O_485,N_24716,N_24849);
nand UO_486 (O_486,N_24627,N_24611);
nand UO_487 (O_487,N_24728,N_24663);
xor UO_488 (O_488,N_24391,N_24435);
xnor UO_489 (O_489,N_24737,N_24694);
and UO_490 (O_490,N_24395,N_24198);
xor UO_491 (O_491,N_24251,N_24506);
xor UO_492 (O_492,N_24433,N_24555);
or UO_493 (O_493,N_24537,N_24470);
xnor UO_494 (O_494,N_24677,N_24560);
and UO_495 (O_495,N_24912,N_24153);
xnor UO_496 (O_496,N_24674,N_24188);
or UO_497 (O_497,N_24281,N_24862);
xor UO_498 (O_498,N_24908,N_24425);
nand UO_499 (O_499,N_24975,N_24695);
nand UO_500 (O_500,N_24004,N_24771);
xor UO_501 (O_501,N_24330,N_24206);
nor UO_502 (O_502,N_24676,N_24779);
nor UO_503 (O_503,N_24802,N_24988);
xnor UO_504 (O_504,N_24855,N_24402);
or UO_505 (O_505,N_24615,N_24761);
nand UO_506 (O_506,N_24699,N_24460);
and UO_507 (O_507,N_24019,N_24176);
or UO_508 (O_508,N_24672,N_24046);
xor UO_509 (O_509,N_24079,N_24893);
nand UO_510 (O_510,N_24666,N_24997);
nor UO_511 (O_511,N_24216,N_24370);
or UO_512 (O_512,N_24659,N_24375);
xor UO_513 (O_513,N_24267,N_24873);
xnor UO_514 (O_514,N_24021,N_24278);
or UO_515 (O_515,N_24139,N_24185);
or UO_516 (O_516,N_24764,N_24224);
or UO_517 (O_517,N_24375,N_24875);
nand UO_518 (O_518,N_24507,N_24642);
and UO_519 (O_519,N_24406,N_24531);
or UO_520 (O_520,N_24306,N_24590);
and UO_521 (O_521,N_24875,N_24539);
nor UO_522 (O_522,N_24540,N_24532);
and UO_523 (O_523,N_24038,N_24175);
or UO_524 (O_524,N_24895,N_24309);
nor UO_525 (O_525,N_24233,N_24306);
and UO_526 (O_526,N_24519,N_24779);
and UO_527 (O_527,N_24996,N_24980);
nand UO_528 (O_528,N_24906,N_24468);
xor UO_529 (O_529,N_24100,N_24990);
nand UO_530 (O_530,N_24408,N_24414);
and UO_531 (O_531,N_24011,N_24643);
nor UO_532 (O_532,N_24702,N_24660);
nor UO_533 (O_533,N_24489,N_24334);
nor UO_534 (O_534,N_24575,N_24018);
or UO_535 (O_535,N_24615,N_24574);
xnor UO_536 (O_536,N_24885,N_24076);
and UO_537 (O_537,N_24172,N_24971);
nor UO_538 (O_538,N_24622,N_24968);
nand UO_539 (O_539,N_24939,N_24783);
nor UO_540 (O_540,N_24656,N_24392);
or UO_541 (O_541,N_24790,N_24123);
and UO_542 (O_542,N_24170,N_24051);
nor UO_543 (O_543,N_24457,N_24889);
nor UO_544 (O_544,N_24764,N_24781);
nand UO_545 (O_545,N_24742,N_24775);
or UO_546 (O_546,N_24747,N_24319);
or UO_547 (O_547,N_24813,N_24432);
xor UO_548 (O_548,N_24018,N_24413);
nand UO_549 (O_549,N_24767,N_24314);
nor UO_550 (O_550,N_24078,N_24581);
or UO_551 (O_551,N_24917,N_24063);
and UO_552 (O_552,N_24291,N_24299);
or UO_553 (O_553,N_24781,N_24863);
and UO_554 (O_554,N_24864,N_24319);
and UO_555 (O_555,N_24160,N_24666);
nor UO_556 (O_556,N_24050,N_24856);
and UO_557 (O_557,N_24224,N_24253);
xnor UO_558 (O_558,N_24359,N_24417);
nor UO_559 (O_559,N_24474,N_24135);
or UO_560 (O_560,N_24372,N_24763);
nor UO_561 (O_561,N_24157,N_24999);
and UO_562 (O_562,N_24012,N_24522);
xor UO_563 (O_563,N_24152,N_24825);
and UO_564 (O_564,N_24156,N_24841);
xor UO_565 (O_565,N_24831,N_24254);
nand UO_566 (O_566,N_24279,N_24188);
nor UO_567 (O_567,N_24333,N_24071);
nor UO_568 (O_568,N_24700,N_24107);
or UO_569 (O_569,N_24192,N_24631);
xnor UO_570 (O_570,N_24363,N_24213);
xor UO_571 (O_571,N_24244,N_24384);
xor UO_572 (O_572,N_24571,N_24481);
xor UO_573 (O_573,N_24558,N_24572);
xor UO_574 (O_574,N_24692,N_24116);
or UO_575 (O_575,N_24781,N_24689);
and UO_576 (O_576,N_24206,N_24953);
or UO_577 (O_577,N_24354,N_24218);
xor UO_578 (O_578,N_24286,N_24521);
or UO_579 (O_579,N_24664,N_24071);
nand UO_580 (O_580,N_24076,N_24542);
and UO_581 (O_581,N_24551,N_24439);
or UO_582 (O_582,N_24759,N_24612);
or UO_583 (O_583,N_24913,N_24574);
or UO_584 (O_584,N_24244,N_24914);
nand UO_585 (O_585,N_24187,N_24661);
xor UO_586 (O_586,N_24207,N_24553);
or UO_587 (O_587,N_24709,N_24324);
nor UO_588 (O_588,N_24239,N_24196);
xnor UO_589 (O_589,N_24591,N_24219);
xor UO_590 (O_590,N_24019,N_24098);
xor UO_591 (O_591,N_24252,N_24098);
nor UO_592 (O_592,N_24943,N_24426);
xnor UO_593 (O_593,N_24557,N_24834);
or UO_594 (O_594,N_24736,N_24879);
or UO_595 (O_595,N_24268,N_24828);
nand UO_596 (O_596,N_24323,N_24163);
and UO_597 (O_597,N_24543,N_24678);
nor UO_598 (O_598,N_24669,N_24132);
xor UO_599 (O_599,N_24866,N_24155);
xnor UO_600 (O_600,N_24247,N_24487);
or UO_601 (O_601,N_24513,N_24368);
or UO_602 (O_602,N_24656,N_24814);
nor UO_603 (O_603,N_24063,N_24657);
nor UO_604 (O_604,N_24849,N_24616);
or UO_605 (O_605,N_24098,N_24164);
or UO_606 (O_606,N_24063,N_24311);
nor UO_607 (O_607,N_24313,N_24008);
nor UO_608 (O_608,N_24118,N_24613);
and UO_609 (O_609,N_24481,N_24356);
nand UO_610 (O_610,N_24710,N_24292);
or UO_611 (O_611,N_24326,N_24709);
xor UO_612 (O_612,N_24436,N_24454);
or UO_613 (O_613,N_24897,N_24812);
xnor UO_614 (O_614,N_24942,N_24083);
and UO_615 (O_615,N_24225,N_24992);
or UO_616 (O_616,N_24099,N_24703);
nor UO_617 (O_617,N_24540,N_24007);
nor UO_618 (O_618,N_24500,N_24710);
or UO_619 (O_619,N_24518,N_24762);
nor UO_620 (O_620,N_24104,N_24135);
xor UO_621 (O_621,N_24929,N_24390);
and UO_622 (O_622,N_24207,N_24029);
and UO_623 (O_623,N_24196,N_24370);
nor UO_624 (O_624,N_24331,N_24018);
nand UO_625 (O_625,N_24893,N_24958);
xnor UO_626 (O_626,N_24821,N_24587);
nand UO_627 (O_627,N_24379,N_24803);
or UO_628 (O_628,N_24709,N_24958);
and UO_629 (O_629,N_24493,N_24681);
nor UO_630 (O_630,N_24062,N_24704);
xor UO_631 (O_631,N_24717,N_24518);
nand UO_632 (O_632,N_24995,N_24805);
and UO_633 (O_633,N_24335,N_24811);
and UO_634 (O_634,N_24583,N_24289);
xor UO_635 (O_635,N_24012,N_24941);
nand UO_636 (O_636,N_24483,N_24955);
nor UO_637 (O_637,N_24492,N_24613);
and UO_638 (O_638,N_24938,N_24055);
or UO_639 (O_639,N_24704,N_24815);
nand UO_640 (O_640,N_24472,N_24439);
and UO_641 (O_641,N_24415,N_24948);
nand UO_642 (O_642,N_24613,N_24354);
and UO_643 (O_643,N_24520,N_24651);
or UO_644 (O_644,N_24997,N_24950);
nor UO_645 (O_645,N_24670,N_24415);
nor UO_646 (O_646,N_24335,N_24248);
or UO_647 (O_647,N_24254,N_24700);
or UO_648 (O_648,N_24206,N_24483);
nor UO_649 (O_649,N_24024,N_24668);
nor UO_650 (O_650,N_24658,N_24650);
xnor UO_651 (O_651,N_24291,N_24548);
nor UO_652 (O_652,N_24049,N_24646);
xnor UO_653 (O_653,N_24077,N_24444);
and UO_654 (O_654,N_24353,N_24523);
or UO_655 (O_655,N_24815,N_24596);
nand UO_656 (O_656,N_24826,N_24618);
or UO_657 (O_657,N_24858,N_24176);
or UO_658 (O_658,N_24929,N_24894);
and UO_659 (O_659,N_24307,N_24981);
nand UO_660 (O_660,N_24291,N_24073);
nor UO_661 (O_661,N_24394,N_24782);
nor UO_662 (O_662,N_24791,N_24650);
nand UO_663 (O_663,N_24417,N_24757);
xor UO_664 (O_664,N_24546,N_24211);
nand UO_665 (O_665,N_24769,N_24028);
nor UO_666 (O_666,N_24756,N_24623);
or UO_667 (O_667,N_24580,N_24931);
xor UO_668 (O_668,N_24986,N_24365);
and UO_669 (O_669,N_24877,N_24433);
nor UO_670 (O_670,N_24613,N_24415);
nand UO_671 (O_671,N_24616,N_24838);
nand UO_672 (O_672,N_24105,N_24130);
nor UO_673 (O_673,N_24936,N_24739);
or UO_674 (O_674,N_24077,N_24603);
nor UO_675 (O_675,N_24565,N_24364);
xnor UO_676 (O_676,N_24177,N_24218);
nor UO_677 (O_677,N_24982,N_24031);
and UO_678 (O_678,N_24052,N_24978);
nor UO_679 (O_679,N_24404,N_24306);
xnor UO_680 (O_680,N_24260,N_24216);
xnor UO_681 (O_681,N_24999,N_24906);
or UO_682 (O_682,N_24106,N_24841);
nor UO_683 (O_683,N_24460,N_24005);
xnor UO_684 (O_684,N_24139,N_24835);
and UO_685 (O_685,N_24757,N_24879);
nand UO_686 (O_686,N_24032,N_24241);
nand UO_687 (O_687,N_24260,N_24752);
nor UO_688 (O_688,N_24442,N_24091);
nor UO_689 (O_689,N_24479,N_24849);
nor UO_690 (O_690,N_24946,N_24194);
nor UO_691 (O_691,N_24456,N_24386);
xor UO_692 (O_692,N_24102,N_24852);
and UO_693 (O_693,N_24847,N_24125);
nand UO_694 (O_694,N_24282,N_24959);
or UO_695 (O_695,N_24706,N_24053);
or UO_696 (O_696,N_24034,N_24867);
or UO_697 (O_697,N_24159,N_24698);
and UO_698 (O_698,N_24095,N_24005);
xor UO_699 (O_699,N_24708,N_24161);
nor UO_700 (O_700,N_24202,N_24033);
or UO_701 (O_701,N_24677,N_24092);
nor UO_702 (O_702,N_24780,N_24557);
or UO_703 (O_703,N_24975,N_24894);
xnor UO_704 (O_704,N_24398,N_24316);
nand UO_705 (O_705,N_24964,N_24925);
nor UO_706 (O_706,N_24280,N_24861);
and UO_707 (O_707,N_24063,N_24827);
and UO_708 (O_708,N_24575,N_24739);
and UO_709 (O_709,N_24299,N_24210);
and UO_710 (O_710,N_24131,N_24104);
nand UO_711 (O_711,N_24225,N_24101);
and UO_712 (O_712,N_24577,N_24960);
or UO_713 (O_713,N_24980,N_24875);
and UO_714 (O_714,N_24734,N_24199);
or UO_715 (O_715,N_24110,N_24276);
xor UO_716 (O_716,N_24714,N_24967);
nand UO_717 (O_717,N_24475,N_24768);
xnor UO_718 (O_718,N_24506,N_24170);
nor UO_719 (O_719,N_24858,N_24692);
xnor UO_720 (O_720,N_24696,N_24265);
and UO_721 (O_721,N_24362,N_24849);
nand UO_722 (O_722,N_24195,N_24679);
nor UO_723 (O_723,N_24709,N_24357);
or UO_724 (O_724,N_24436,N_24888);
and UO_725 (O_725,N_24673,N_24708);
and UO_726 (O_726,N_24427,N_24022);
nand UO_727 (O_727,N_24787,N_24038);
nor UO_728 (O_728,N_24727,N_24941);
xor UO_729 (O_729,N_24432,N_24830);
and UO_730 (O_730,N_24743,N_24440);
nand UO_731 (O_731,N_24851,N_24018);
and UO_732 (O_732,N_24166,N_24147);
nor UO_733 (O_733,N_24180,N_24227);
or UO_734 (O_734,N_24714,N_24378);
nor UO_735 (O_735,N_24203,N_24272);
nor UO_736 (O_736,N_24645,N_24377);
nor UO_737 (O_737,N_24091,N_24331);
nand UO_738 (O_738,N_24226,N_24724);
nand UO_739 (O_739,N_24020,N_24916);
nor UO_740 (O_740,N_24810,N_24332);
nor UO_741 (O_741,N_24264,N_24944);
xor UO_742 (O_742,N_24446,N_24821);
nor UO_743 (O_743,N_24935,N_24723);
nand UO_744 (O_744,N_24015,N_24301);
nor UO_745 (O_745,N_24799,N_24782);
xor UO_746 (O_746,N_24761,N_24275);
nor UO_747 (O_747,N_24039,N_24199);
nor UO_748 (O_748,N_24599,N_24754);
or UO_749 (O_749,N_24036,N_24173);
and UO_750 (O_750,N_24372,N_24315);
nand UO_751 (O_751,N_24143,N_24259);
nand UO_752 (O_752,N_24997,N_24024);
xor UO_753 (O_753,N_24914,N_24921);
nand UO_754 (O_754,N_24882,N_24112);
nand UO_755 (O_755,N_24973,N_24934);
nor UO_756 (O_756,N_24865,N_24470);
and UO_757 (O_757,N_24522,N_24120);
xor UO_758 (O_758,N_24900,N_24014);
nor UO_759 (O_759,N_24901,N_24604);
nor UO_760 (O_760,N_24844,N_24155);
nand UO_761 (O_761,N_24568,N_24912);
nor UO_762 (O_762,N_24045,N_24660);
and UO_763 (O_763,N_24970,N_24366);
nor UO_764 (O_764,N_24397,N_24334);
nand UO_765 (O_765,N_24740,N_24618);
or UO_766 (O_766,N_24798,N_24282);
nand UO_767 (O_767,N_24881,N_24777);
or UO_768 (O_768,N_24156,N_24453);
xor UO_769 (O_769,N_24569,N_24096);
nand UO_770 (O_770,N_24608,N_24724);
nand UO_771 (O_771,N_24728,N_24682);
or UO_772 (O_772,N_24927,N_24538);
nand UO_773 (O_773,N_24656,N_24826);
nand UO_774 (O_774,N_24517,N_24246);
nand UO_775 (O_775,N_24908,N_24656);
nand UO_776 (O_776,N_24725,N_24184);
or UO_777 (O_777,N_24605,N_24333);
xnor UO_778 (O_778,N_24410,N_24432);
nor UO_779 (O_779,N_24745,N_24873);
or UO_780 (O_780,N_24708,N_24398);
xnor UO_781 (O_781,N_24740,N_24310);
or UO_782 (O_782,N_24689,N_24861);
nor UO_783 (O_783,N_24212,N_24922);
nand UO_784 (O_784,N_24141,N_24243);
xor UO_785 (O_785,N_24627,N_24888);
xnor UO_786 (O_786,N_24879,N_24839);
nand UO_787 (O_787,N_24804,N_24429);
or UO_788 (O_788,N_24536,N_24537);
xnor UO_789 (O_789,N_24553,N_24668);
nor UO_790 (O_790,N_24372,N_24494);
nand UO_791 (O_791,N_24858,N_24960);
and UO_792 (O_792,N_24697,N_24666);
or UO_793 (O_793,N_24828,N_24253);
or UO_794 (O_794,N_24048,N_24818);
xnor UO_795 (O_795,N_24481,N_24787);
nor UO_796 (O_796,N_24436,N_24240);
or UO_797 (O_797,N_24142,N_24138);
nor UO_798 (O_798,N_24742,N_24503);
xor UO_799 (O_799,N_24262,N_24338);
xnor UO_800 (O_800,N_24749,N_24049);
xor UO_801 (O_801,N_24195,N_24801);
nand UO_802 (O_802,N_24949,N_24752);
or UO_803 (O_803,N_24969,N_24334);
nand UO_804 (O_804,N_24421,N_24671);
xor UO_805 (O_805,N_24950,N_24829);
and UO_806 (O_806,N_24597,N_24681);
or UO_807 (O_807,N_24515,N_24606);
or UO_808 (O_808,N_24865,N_24967);
nor UO_809 (O_809,N_24464,N_24107);
nand UO_810 (O_810,N_24500,N_24542);
nor UO_811 (O_811,N_24353,N_24681);
nor UO_812 (O_812,N_24136,N_24452);
or UO_813 (O_813,N_24456,N_24656);
nor UO_814 (O_814,N_24515,N_24888);
nand UO_815 (O_815,N_24205,N_24677);
and UO_816 (O_816,N_24375,N_24454);
and UO_817 (O_817,N_24682,N_24787);
nand UO_818 (O_818,N_24426,N_24036);
xnor UO_819 (O_819,N_24321,N_24601);
nor UO_820 (O_820,N_24980,N_24546);
nand UO_821 (O_821,N_24490,N_24418);
nor UO_822 (O_822,N_24360,N_24261);
and UO_823 (O_823,N_24115,N_24682);
and UO_824 (O_824,N_24721,N_24580);
xor UO_825 (O_825,N_24138,N_24086);
nor UO_826 (O_826,N_24528,N_24618);
nand UO_827 (O_827,N_24756,N_24926);
nand UO_828 (O_828,N_24376,N_24969);
nor UO_829 (O_829,N_24038,N_24955);
nand UO_830 (O_830,N_24357,N_24409);
xnor UO_831 (O_831,N_24510,N_24136);
or UO_832 (O_832,N_24402,N_24730);
and UO_833 (O_833,N_24923,N_24093);
and UO_834 (O_834,N_24787,N_24788);
nand UO_835 (O_835,N_24076,N_24769);
or UO_836 (O_836,N_24981,N_24598);
nand UO_837 (O_837,N_24285,N_24580);
and UO_838 (O_838,N_24958,N_24373);
nand UO_839 (O_839,N_24056,N_24479);
nand UO_840 (O_840,N_24407,N_24709);
nand UO_841 (O_841,N_24753,N_24384);
nand UO_842 (O_842,N_24588,N_24477);
xor UO_843 (O_843,N_24619,N_24774);
and UO_844 (O_844,N_24323,N_24633);
xnor UO_845 (O_845,N_24360,N_24584);
or UO_846 (O_846,N_24223,N_24070);
or UO_847 (O_847,N_24236,N_24921);
or UO_848 (O_848,N_24251,N_24289);
nor UO_849 (O_849,N_24821,N_24768);
and UO_850 (O_850,N_24418,N_24389);
nor UO_851 (O_851,N_24583,N_24688);
xor UO_852 (O_852,N_24354,N_24679);
nand UO_853 (O_853,N_24287,N_24786);
or UO_854 (O_854,N_24622,N_24842);
or UO_855 (O_855,N_24754,N_24823);
and UO_856 (O_856,N_24027,N_24375);
and UO_857 (O_857,N_24241,N_24187);
or UO_858 (O_858,N_24201,N_24637);
and UO_859 (O_859,N_24886,N_24230);
or UO_860 (O_860,N_24347,N_24931);
xor UO_861 (O_861,N_24789,N_24335);
xor UO_862 (O_862,N_24998,N_24574);
xnor UO_863 (O_863,N_24596,N_24138);
and UO_864 (O_864,N_24647,N_24617);
or UO_865 (O_865,N_24886,N_24152);
and UO_866 (O_866,N_24740,N_24435);
or UO_867 (O_867,N_24862,N_24156);
nor UO_868 (O_868,N_24534,N_24225);
and UO_869 (O_869,N_24399,N_24087);
nor UO_870 (O_870,N_24933,N_24514);
nor UO_871 (O_871,N_24264,N_24536);
or UO_872 (O_872,N_24148,N_24348);
and UO_873 (O_873,N_24243,N_24161);
nor UO_874 (O_874,N_24566,N_24727);
nand UO_875 (O_875,N_24829,N_24044);
or UO_876 (O_876,N_24185,N_24427);
nand UO_877 (O_877,N_24747,N_24339);
nand UO_878 (O_878,N_24943,N_24378);
and UO_879 (O_879,N_24507,N_24849);
and UO_880 (O_880,N_24165,N_24754);
or UO_881 (O_881,N_24574,N_24426);
nor UO_882 (O_882,N_24703,N_24190);
xnor UO_883 (O_883,N_24797,N_24540);
xor UO_884 (O_884,N_24319,N_24023);
xnor UO_885 (O_885,N_24643,N_24887);
and UO_886 (O_886,N_24117,N_24710);
and UO_887 (O_887,N_24711,N_24378);
nand UO_888 (O_888,N_24473,N_24112);
and UO_889 (O_889,N_24507,N_24580);
nand UO_890 (O_890,N_24551,N_24393);
or UO_891 (O_891,N_24349,N_24900);
xnor UO_892 (O_892,N_24342,N_24984);
or UO_893 (O_893,N_24078,N_24077);
xor UO_894 (O_894,N_24065,N_24004);
or UO_895 (O_895,N_24726,N_24839);
or UO_896 (O_896,N_24599,N_24752);
and UO_897 (O_897,N_24815,N_24299);
or UO_898 (O_898,N_24429,N_24514);
or UO_899 (O_899,N_24552,N_24566);
nand UO_900 (O_900,N_24982,N_24532);
nand UO_901 (O_901,N_24403,N_24163);
nand UO_902 (O_902,N_24496,N_24623);
nor UO_903 (O_903,N_24984,N_24193);
and UO_904 (O_904,N_24539,N_24587);
or UO_905 (O_905,N_24193,N_24735);
xor UO_906 (O_906,N_24908,N_24550);
nand UO_907 (O_907,N_24742,N_24733);
nand UO_908 (O_908,N_24515,N_24304);
and UO_909 (O_909,N_24831,N_24671);
nand UO_910 (O_910,N_24583,N_24027);
and UO_911 (O_911,N_24400,N_24144);
and UO_912 (O_912,N_24448,N_24171);
nor UO_913 (O_913,N_24659,N_24008);
and UO_914 (O_914,N_24299,N_24931);
or UO_915 (O_915,N_24170,N_24543);
or UO_916 (O_916,N_24114,N_24036);
xnor UO_917 (O_917,N_24965,N_24752);
xor UO_918 (O_918,N_24649,N_24300);
or UO_919 (O_919,N_24658,N_24186);
or UO_920 (O_920,N_24419,N_24727);
or UO_921 (O_921,N_24317,N_24415);
xor UO_922 (O_922,N_24252,N_24511);
xor UO_923 (O_923,N_24793,N_24113);
or UO_924 (O_924,N_24933,N_24753);
and UO_925 (O_925,N_24696,N_24594);
or UO_926 (O_926,N_24423,N_24706);
nand UO_927 (O_927,N_24594,N_24634);
xor UO_928 (O_928,N_24430,N_24460);
nand UO_929 (O_929,N_24726,N_24546);
nor UO_930 (O_930,N_24187,N_24111);
xnor UO_931 (O_931,N_24863,N_24288);
and UO_932 (O_932,N_24560,N_24465);
or UO_933 (O_933,N_24746,N_24050);
nand UO_934 (O_934,N_24597,N_24764);
nand UO_935 (O_935,N_24335,N_24064);
or UO_936 (O_936,N_24743,N_24351);
xnor UO_937 (O_937,N_24731,N_24481);
nor UO_938 (O_938,N_24610,N_24775);
xnor UO_939 (O_939,N_24979,N_24836);
nand UO_940 (O_940,N_24590,N_24799);
or UO_941 (O_941,N_24926,N_24829);
nand UO_942 (O_942,N_24077,N_24312);
and UO_943 (O_943,N_24366,N_24830);
and UO_944 (O_944,N_24130,N_24691);
xor UO_945 (O_945,N_24972,N_24805);
nor UO_946 (O_946,N_24392,N_24648);
or UO_947 (O_947,N_24907,N_24585);
and UO_948 (O_948,N_24166,N_24313);
or UO_949 (O_949,N_24079,N_24522);
or UO_950 (O_950,N_24137,N_24805);
or UO_951 (O_951,N_24784,N_24262);
or UO_952 (O_952,N_24940,N_24331);
nor UO_953 (O_953,N_24646,N_24226);
nand UO_954 (O_954,N_24740,N_24482);
nand UO_955 (O_955,N_24131,N_24971);
nor UO_956 (O_956,N_24997,N_24225);
nor UO_957 (O_957,N_24020,N_24076);
and UO_958 (O_958,N_24502,N_24705);
xor UO_959 (O_959,N_24190,N_24405);
nor UO_960 (O_960,N_24871,N_24210);
nor UO_961 (O_961,N_24904,N_24689);
and UO_962 (O_962,N_24234,N_24950);
and UO_963 (O_963,N_24454,N_24057);
and UO_964 (O_964,N_24413,N_24381);
and UO_965 (O_965,N_24258,N_24275);
or UO_966 (O_966,N_24245,N_24244);
and UO_967 (O_967,N_24305,N_24587);
xor UO_968 (O_968,N_24655,N_24526);
xor UO_969 (O_969,N_24832,N_24195);
and UO_970 (O_970,N_24642,N_24983);
and UO_971 (O_971,N_24351,N_24037);
nor UO_972 (O_972,N_24575,N_24411);
xnor UO_973 (O_973,N_24015,N_24702);
or UO_974 (O_974,N_24333,N_24896);
xor UO_975 (O_975,N_24400,N_24138);
and UO_976 (O_976,N_24699,N_24764);
nand UO_977 (O_977,N_24829,N_24115);
nor UO_978 (O_978,N_24364,N_24555);
or UO_979 (O_979,N_24579,N_24042);
xor UO_980 (O_980,N_24625,N_24669);
nand UO_981 (O_981,N_24909,N_24977);
nand UO_982 (O_982,N_24162,N_24777);
nand UO_983 (O_983,N_24145,N_24071);
and UO_984 (O_984,N_24133,N_24474);
nand UO_985 (O_985,N_24410,N_24892);
or UO_986 (O_986,N_24876,N_24531);
xor UO_987 (O_987,N_24772,N_24882);
or UO_988 (O_988,N_24829,N_24937);
nand UO_989 (O_989,N_24829,N_24000);
and UO_990 (O_990,N_24591,N_24824);
and UO_991 (O_991,N_24571,N_24295);
nor UO_992 (O_992,N_24605,N_24634);
and UO_993 (O_993,N_24104,N_24290);
and UO_994 (O_994,N_24146,N_24939);
nand UO_995 (O_995,N_24808,N_24466);
nand UO_996 (O_996,N_24252,N_24109);
nor UO_997 (O_997,N_24691,N_24210);
nor UO_998 (O_998,N_24438,N_24113);
xnor UO_999 (O_999,N_24943,N_24205);
nor UO_1000 (O_1000,N_24447,N_24729);
nand UO_1001 (O_1001,N_24079,N_24917);
nand UO_1002 (O_1002,N_24577,N_24076);
nand UO_1003 (O_1003,N_24825,N_24331);
xor UO_1004 (O_1004,N_24388,N_24749);
xor UO_1005 (O_1005,N_24027,N_24566);
and UO_1006 (O_1006,N_24339,N_24692);
or UO_1007 (O_1007,N_24893,N_24796);
and UO_1008 (O_1008,N_24745,N_24999);
nand UO_1009 (O_1009,N_24958,N_24126);
nand UO_1010 (O_1010,N_24061,N_24553);
nand UO_1011 (O_1011,N_24009,N_24704);
or UO_1012 (O_1012,N_24140,N_24330);
xnor UO_1013 (O_1013,N_24229,N_24521);
or UO_1014 (O_1014,N_24647,N_24248);
or UO_1015 (O_1015,N_24545,N_24120);
nor UO_1016 (O_1016,N_24775,N_24398);
nor UO_1017 (O_1017,N_24026,N_24555);
or UO_1018 (O_1018,N_24468,N_24167);
and UO_1019 (O_1019,N_24695,N_24039);
xnor UO_1020 (O_1020,N_24806,N_24599);
and UO_1021 (O_1021,N_24840,N_24229);
xor UO_1022 (O_1022,N_24732,N_24978);
and UO_1023 (O_1023,N_24211,N_24087);
or UO_1024 (O_1024,N_24615,N_24903);
nand UO_1025 (O_1025,N_24546,N_24513);
or UO_1026 (O_1026,N_24459,N_24693);
nand UO_1027 (O_1027,N_24576,N_24241);
nor UO_1028 (O_1028,N_24141,N_24260);
nand UO_1029 (O_1029,N_24941,N_24186);
nand UO_1030 (O_1030,N_24912,N_24060);
nor UO_1031 (O_1031,N_24517,N_24102);
nor UO_1032 (O_1032,N_24204,N_24724);
xor UO_1033 (O_1033,N_24028,N_24998);
nand UO_1034 (O_1034,N_24887,N_24213);
nand UO_1035 (O_1035,N_24564,N_24840);
nor UO_1036 (O_1036,N_24773,N_24378);
or UO_1037 (O_1037,N_24594,N_24686);
nor UO_1038 (O_1038,N_24211,N_24206);
and UO_1039 (O_1039,N_24755,N_24109);
and UO_1040 (O_1040,N_24440,N_24526);
xnor UO_1041 (O_1041,N_24056,N_24173);
and UO_1042 (O_1042,N_24505,N_24369);
and UO_1043 (O_1043,N_24597,N_24881);
nand UO_1044 (O_1044,N_24285,N_24420);
nor UO_1045 (O_1045,N_24677,N_24111);
xnor UO_1046 (O_1046,N_24010,N_24442);
nor UO_1047 (O_1047,N_24385,N_24853);
and UO_1048 (O_1048,N_24720,N_24231);
nor UO_1049 (O_1049,N_24227,N_24868);
xor UO_1050 (O_1050,N_24687,N_24713);
nand UO_1051 (O_1051,N_24749,N_24485);
nand UO_1052 (O_1052,N_24416,N_24147);
nor UO_1053 (O_1053,N_24535,N_24784);
xor UO_1054 (O_1054,N_24189,N_24885);
nand UO_1055 (O_1055,N_24223,N_24942);
nor UO_1056 (O_1056,N_24929,N_24893);
and UO_1057 (O_1057,N_24421,N_24408);
and UO_1058 (O_1058,N_24522,N_24064);
or UO_1059 (O_1059,N_24184,N_24819);
nor UO_1060 (O_1060,N_24839,N_24632);
or UO_1061 (O_1061,N_24091,N_24639);
nand UO_1062 (O_1062,N_24987,N_24367);
nand UO_1063 (O_1063,N_24409,N_24918);
and UO_1064 (O_1064,N_24359,N_24682);
nor UO_1065 (O_1065,N_24530,N_24469);
nand UO_1066 (O_1066,N_24028,N_24546);
nor UO_1067 (O_1067,N_24163,N_24555);
and UO_1068 (O_1068,N_24630,N_24776);
xnor UO_1069 (O_1069,N_24418,N_24960);
xnor UO_1070 (O_1070,N_24361,N_24805);
and UO_1071 (O_1071,N_24935,N_24337);
xor UO_1072 (O_1072,N_24544,N_24838);
or UO_1073 (O_1073,N_24902,N_24621);
xnor UO_1074 (O_1074,N_24111,N_24166);
and UO_1075 (O_1075,N_24049,N_24949);
nand UO_1076 (O_1076,N_24818,N_24114);
nor UO_1077 (O_1077,N_24577,N_24442);
nand UO_1078 (O_1078,N_24978,N_24297);
xnor UO_1079 (O_1079,N_24604,N_24332);
or UO_1080 (O_1080,N_24623,N_24718);
xnor UO_1081 (O_1081,N_24734,N_24807);
or UO_1082 (O_1082,N_24008,N_24066);
and UO_1083 (O_1083,N_24534,N_24118);
or UO_1084 (O_1084,N_24438,N_24983);
xor UO_1085 (O_1085,N_24594,N_24653);
or UO_1086 (O_1086,N_24156,N_24102);
and UO_1087 (O_1087,N_24253,N_24871);
and UO_1088 (O_1088,N_24783,N_24038);
nand UO_1089 (O_1089,N_24175,N_24728);
xnor UO_1090 (O_1090,N_24132,N_24350);
nor UO_1091 (O_1091,N_24587,N_24197);
nor UO_1092 (O_1092,N_24587,N_24286);
xor UO_1093 (O_1093,N_24013,N_24343);
or UO_1094 (O_1094,N_24622,N_24934);
or UO_1095 (O_1095,N_24948,N_24202);
or UO_1096 (O_1096,N_24004,N_24469);
xor UO_1097 (O_1097,N_24945,N_24756);
or UO_1098 (O_1098,N_24165,N_24323);
nand UO_1099 (O_1099,N_24974,N_24195);
nor UO_1100 (O_1100,N_24235,N_24774);
or UO_1101 (O_1101,N_24051,N_24201);
xor UO_1102 (O_1102,N_24352,N_24423);
or UO_1103 (O_1103,N_24383,N_24584);
or UO_1104 (O_1104,N_24434,N_24872);
nand UO_1105 (O_1105,N_24863,N_24965);
and UO_1106 (O_1106,N_24053,N_24764);
nor UO_1107 (O_1107,N_24768,N_24732);
and UO_1108 (O_1108,N_24010,N_24657);
nor UO_1109 (O_1109,N_24439,N_24881);
or UO_1110 (O_1110,N_24883,N_24485);
xor UO_1111 (O_1111,N_24396,N_24922);
or UO_1112 (O_1112,N_24695,N_24673);
nor UO_1113 (O_1113,N_24259,N_24991);
nand UO_1114 (O_1114,N_24884,N_24629);
or UO_1115 (O_1115,N_24720,N_24200);
xnor UO_1116 (O_1116,N_24344,N_24464);
and UO_1117 (O_1117,N_24680,N_24787);
xnor UO_1118 (O_1118,N_24273,N_24382);
xnor UO_1119 (O_1119,N_24007,N_24027);
xnor UO_1120 (O_1120,N_24876,N_24720);
xor UO_1121 (O_1121,N_24951,N_24673);
and UO_1122 (O_1122,N_24361,N_24607);
and UO_1123 (O_1123,N_24518,N_24259);
nand UO_1124 (O_1124,N_24830,N_24676);
or UO_1125 (O_1125,N_24320,N_24735);
nor UO_1126 (O_1126,N_24066,N_24248);
or UO_1127 (O_1127,N_24381,N_24169);
xor UO_1128 (O_1128,N_24442,N_24205);
or UO_1129 (O_1129,N_24381,N_24290);
nand UO_1130 (O_1130,N_24186,N_24728);
or UO_1131 (O_1131,N_24352,N_24139);
and UO_1132 (O_1132,N_24716,N_24803);
nand UO_1133 (O_1133,N_24890,N_24755);
xor UO_1134 (O_1134,N_24296,N_24240);
nand UO_1135 (O_1135,N_24610,N_24321);
nand UO_1136 (O_1136,N_24354,N_24943);
and UO_1137 (O_1137,N_24961,N_24765);
and UO_1138 (O_1138,N_24775,N_24299);
or UO_1139 (O_1139,N_24348,N_24335);
nor UO_1140 (O_1140,N_24284,N_24831);
nor UO_1141 (O_1141,N_24766,N_24564);
or UO_1142 (O_1142,N_24332,N_24487);
xnor UO_1143 (O_1143,N_24790,N_24495);
xnor UO_1144 (O_1144,N_24346,N_24052);
nor UO_1145 (O_1145,N_24655,N_24793);
nor UO_1146 (O_1146,N_24952,N_24534);
and UO_1147 (O_1147,N_24119,N_24331);
and UO_1148 (O_1148,N_24726,N_24428);
or UO_1149 (O_1149,N_24501,N_24437);
nand UO_1150 (O_1150,N_24943,N_24012);
nor UO_1151 (O_1151,N_24732,N_24238);
nand UO_1152 (O_1152,N_24082,N_24454);
or UO_1153 (O_1153,N_24124,N_24020);
xnor UO_1154 (O_1154,N_24356,N_24277);
nand UO_1155 (O_1155,N_24961,N_24837);
nor UO_1156 (O_1156,N_24729,N_24189);
nand UO_1157 (O_1157,N_24185,N_24070);
nand UO_1158 (O_1158,N_24380,N_24417);
and UO_1159 (O_1159,N_24840,N_24885);
nand UO_1160 (O_1160,N_24379,N_24347);
nor UO_1161 (O_1161,N_24493,N_24571);
nand UO_1162 (O_1162,N_24932,N_24953);
nor UO_1163 (O_1163,N_24109,N_24810);
nand UO_1164 (O_1164,N_24345,N_24610);
xor UO_1165 (O_1165,N_24535,N_24207);
nor UO_1166 (O_1166,N_24009,N_24538);
nor UO_1167 (O_1167,N_24195,N_24165);
and UO_1168 (O_1168,N_24175,N_24503);
and UO_1169 (O_1169,N_24727,N_24711);
nand UO_1170 (O_1170,N_24511,N_24000);
and UO_1171 (O_1171,N_24344,N_24107);
and UO_1172 (O_1172,N_24624,N_24046);
or UO_1173 (O_1173,N_24451,N_24301);
or UO_1174 (O_1174,N_24675,N_24525);
nand UO_1175 (O_1175,N_24833,N_24135);
and UO_1176 (O_1176,N_24475,N_24566);
or UO_1177 (O_1177,N_24322,N_24252);
nand UO_1178 (O_1178,N_24661,N_24035);
xnor UO_1179 (O_1179,N_24658,N_24619);
nor UO_1180 (O_1180,N_24431,N_24920);
or UO_1181 (O_1181,N_24179,N_24304);
nor UO_1182 (O_1182,N_24272,N_24977);
xnor UO_1183 (O_1183,N_24630,N_24555);
and UO_1184 (O_1184,N_24247,N_24565);
xor UO_1185 (O_1185,N_24980,N_24743);
nor UO_1186 (O_1186,N_24048,N_24057);
nand UO_1187 (O_1187,N_24395,N_24113);
or UO_1188 (O_1188,N_24838,N_24658);
and UO_1189 (O_1189,N_24745,N_24466);
or UO_1190 (O_1190,N_24202,N_24074);
nor UO_1191 (O_1191,N_24610,N_24505);
xnor UO_1192 (O_1192,N_24652,N_24770);
nand UO_1193 (O_1193,N_24483,N_24019);
nand UO_1194 (O_1194,N_24021,N_24335);
or UO_1195 (O_1195,N_24464,N_24319);
nand UO_1196 (O_1196,N_24889,N_24884);
and UO_1197 (O_1197,N_24461,N_24659);
xnor UO_1198 (O_1198,N_24078,N_24386);
xnor UO_1199 (O_1199,N_24877,N_24369);
nor UO_1200 (O_1200,N_24797,N_24274);
and UO_1201 (O_1201,N_24293,N_24001);
or UO_1202 (O_1202,N_24270,N_24222);
nand UO_1203 (O_1203,N_24525,N_24733);
nand UO_1204 (O_1204,N_24022,N_24010);
nand UO_1205 (O_1205,N_24429,N_24832);
and UO_1206 (O_1206,N_24808,N_24832);
or UO_1207 (O_1207,N_24587,N_24125);
and UO_1208 (O_1208,N_24585,N_24349);
or UO_1209 (O_1209,N_24233,N_24365);
nor UO_1210 (O_1210,N_24621,N_24741);
or UO_1211 (O_1211,N_24752,N_24530);
nand UO_1212 (O_1212,N_24180,N_24231);
and UO_1213 (O_1213,N_24867,N_24614);
or UO_1214 (O_1214,N_24537,N_24452);
nand UO_1215 (O_1215,N_24451,N_24103);
or UO_1216 (O_1216,N_24363,N_24881);
xnor UO_1217 (O_1217,N_24838,N_24830);
nand UO_1218 (O_1218,N_24797,N_24947);
nand UO_1219 (O_1219,N_24426,N_24053);
xnor UO_1220 (O_1220,N_24774,N_24385);
and UO_1221 (O_1221,N_24974,N_24125);
and UO_1222 (O_1222,N_24615,N_24270);
nor UO_1223 (O_1223,N_24768,N_24577);
and UO_1224 (O_1224,N_24244,N_24292);
and UO_1225 (O_1225,N_24982,N_24307);
nand UO_1226 (O_1226,N_24555,N_24421);
or UO_1227 (O_1227,N_24778,N_24027);
xor UO_1228 (O_1228,N_24008,N_24998);
nor UO_1229 (O_1229,N_24069,N_24824);
nand UO_1230 (O_1230,N_24771,N_24560);
nand UO_1231 (O_1231,N_24114,N_24358);
nor UO_1232 (O_1232,N_24654,N_24727);
or UO_1233 (O_1233,N_24176,N_24930);
and UO_1234 (O_1234,N_24634,N_24371);
nand UO_1235 (O_1235,N_24581,N_24575);
nand UO_1236 (O_1236,N_24906,N_24151);
nor UO_1237 (O_1237,N_24637,N_24802);
nor UO_1238 (O_1238,N_24000,N_24811);
or UO_1239 (O_1239,N_24782,N_24415);
nand UO_1240 (O_1240,N_24196,N_24542);
nand UO_1241 (O_1241,N_24523,N_24904);
nor UO_1242 (O_1242,N_24787,N_24744);
xor UO_1243 (O_1243,N_24398,N_24908);
and UO_1244 (O_1244,N_24879,N_24861);
nor UO_1245 (O_1245,N_24935,N_24467);
or UO_1246 (O_1246,N_24521,N_24116);
and UO_1247 (O_1247,N_24790,N_24129);
and UO_1248 (O_1248,N_24383,N_24433);
xnor UO_1249 (O_1249,N_24806,N_24152);
nor UO_1250 (O_1250,N_24832,N_24522);
and UO_1251 (O_1251,N_24349,N_24084);
or UO_1252 (O_1252,N_24918,N_24012);
or UO_1253 (O_1253,N_24443,N_24055);
and UO_1254 (O_1254,N_24833,N_24440);
xnor UO_1255 (O_1255,N_24243,N_24700);
nand UO_1256 (O_1256,N_24830,N_24411);
nand UO_1257 (O_1257,N_24009,N_24857);
nor UO_1258 (O_1258,N_24952,N_24134);
nand UO_1259 (O_1259,N_24350,N_24865);
nor UO_1260 (O_1260,N_24398,N_24357);
and UO_1261 (O_1261,N_24834,N_24947);
nor UO_1262 (O_1262,N_24698,N_24980);
and UO_1263 (O_1263,N_24968,N_24366);
and UO_1264 (O_1264,N_24276,N_24376);
or UO_1265 (O_1265,N_24979,N_24964);
and UO_1266 (O_1266,N_24900,N_24957);
or UO_1267 (O_1267,N_24157,N_24256);
nor UO_1268 (O_1268,N_24308,N_24920);
nor UO_1269 (O_1269,N_24136,N_24982);
xor UO_1270 (O_1270,N_24093,N_24352);
and UO_1271 (O_1271,N_24154,N_24475);
nand UO_1272 (O_1272,N_24513,N_24820);
xnor UO_1273 (O_1273,N_24080,N_24722);
and UO_1274 (O_1274,N_24721,N_24780);
or UO_1275 (O_1275,N_24089,N_24558);
xor UO_1276 (O_1276,N_24281,N_24181);
or UO_1277 (O_1277,N_24873,N_24912);
xnor UO_1278 (O_1278,N_24881,N_24833);
xor UO_1279 (O_1279,N_24330,N_24369);
nor UO_1280 (O_1280,N_24479,N_24063);
xnor UO_1281 (O_1281,N_24404,N_24459);
and UO_1282 (O_1282,N_24287,N_24438);
xor UO_1283 (O_1283,N_24558,N_24865);
xnor UO_1284 (O_1284,N_24418,N_24647);
and UO_1285 (O_1285,N_24377,N_24538);
nand UO_1286 (O_1286,N_24488,N_24916);
xnor UO_1287 (O_1287,N_24379,N_24099);
nor UO_1288 (O_1288,N_24552,N_24778);
nor UO_1289 (O_1289,N_24934,N_24195);
nand UO_1290 (O_1290,N_24085,N_24548);
or UO_1291 (O_1291,N_24741,N_24623);
or UO_1292 (O_1292,N_24490,N_24272);
or UO_1293 (O_1293,N_24094,N_24666);
or UO_1294 (O_1294,N_24395,N_24055);
or UO_1295 (O_1295,N_24452,N_24051);
or UO_1296 (O_1296,N_24074,N_24085);
nand UO_1297 (O_1297,N_24161,N_24023);
nor UO_1298 (O_1298,N_24502,N_24216);
or UO_1299 (O_1299,N_24322,N_24130);
xor UO_1300 (O_1300,N_24504,N_24911);
and UO_1301 (O_1301,N_24281,N_24006);
nor UO_1302 (O_1302,N_24797,N_24046);
nor UO_1303 (O_1303,N_24235,N_24763);
nor UO_1304 (O_1304,N_24715,N_24985);
or UO_1305 (O_1305,N_24153,N_24157);
nor UO_1306 (O_1306,N_24293,N_24300);
xnor UO_1307 (O_1307,N_24085,N_24228);
or UO_1308 (O_1308,N_24468,N_24266);
nor UO_1309 (O_1309,N_24587,N_24033);
nor UO_1310 (O_1310,N_24820,N_24664);
nand UO_1311 (O_1311,N_24232,N_24333);
nor UO_1312 (O_1312,N_24304,N_24280);
xnor UO_1313 (O_1313,N_24393,N_24965);
or UO_1314 (O_1314,N_24038,N_24551);
nor UO_1315 (O_1315,N_24571,N_24059);
nor UO_1316 (O_1316,N_24932,N_24716);
nand UO_1317 (O_1317,N_24041,N_24434);
nor UO_1318 (O_1318,N_24718,N_24543);
and UO_1319 (O_1319,N_24734,N_24107);
nand UO_1320 (O_1320,N_24228,N_24852);
and UO_1321 (O_1321,N_24935,N_24013);
and UO_1322 (O_1322,N_24675,N_24518);
xnor UO_1323 (O_1323,N_24683,N_24029);
xor UO_1324 (O_1324,N_24083,N_24036);
xor UO_1325 (O_1325,N_24146,N_24892);
xor UO_1326 (O_1326,N_24864,N_24342);
or UO_1327 (O_1327,N_24875,N_24857);
nand UO_1328 (O_1328,N_24730,N_24324);
or UO_1329 (O_1329,N_24428,N_24021);
and UO_1330 (O_1330,N_24011,N_24091);
xnor UO_1331 (O_1331,N_24566,N_24947);
and UO_1332 (O_1332,N_24274,N_24775);
nor UO_1333 (O_1333,N_24329,N_24743);
or UO_1334 (O_1334,N_24256,N_24099);
nor UO_1335 (O_1335,N_24737,N_24458);
xor UO_1336 (O_1336,N_24268,N_24976);
and UO_1337 (O_1337,N_24677,N_24963);
and UO_1338 (O_1338,N_24882,N_24867);
nor UO_1339 (O_1339,N_24548,N_24591);
or UO_1340 (O_1340,N_24526,N_24894);
nand UO_1341 (O_1341,N_24584,N_24983);
nand UO_1342 (O_1342,N_24074,N_24061);
and UO_1343 (O_1343,N_24774,N_24969);
nand UO_1344 (O_1344,N_24431,N_24448);
or UO_1345 (O_1345,N_24835,N_24346);
and UO_1346 (O_1346,N_24415,N_24236);
xnor UO_1347 (O_1347,N_24133,N_24494);
and UO_1348 (O_1348,N_24110,N_24063);
nand UO_1349 (O_1349,N_24496,N_24361);
nand UO_1350 (O_1350,N_24174,N_24268);
nand UO_1351 (O_1351,N_24214,N_24130);
or UO_1352 (O_1352,N_24998,N_24275);
nand UO_1353 (O_1353,N_24364,N_24365);
xor UO_1354 (O_1354,N_24765,N_24464);
xor UO_1355 (O_1355,N_24621,N_24085);
xnor UO_1356 (O_1356,N_24830,N_24014);
or UO_1357 (O_1357,N_24968,N_24795);
nor UO_1358 (O_1358,N_24030,N_24742);
nor UO_1359 (O_1359,N_24803,N_24590);
nor UO_1360 (O_1360,N_24610,N_24311);
xor UO_1361 (O_1361,N_24347,N_24985);
nor UO_1362 (O_1362,N_24532,N_24354);
nor UO_1363 (O_1363,N_24339,N_24490);
and UO_1364 (O_1364,N_24664,N_24659);
nand UO_1365 (O_1365,N_24895,N_24819);
nand UO_1366 (O_1366,N_24921,N_24149);
nor UO_1367 (O_1367,N_24050,N_24906);
and UO_1368 (O_1368,N_24528,N_24670);
nand UO_1369 (O_1369,N_24892,N_24508);
and UO_1370 (O_1370,N_24070,N_24258);
or UO_1371 (O_1371,N_24920,N_24539);
or UO_1372 (O_1372,N_24509,N_24408);
nand UO_1373 (O_1373,N_24861,N_24752);
xor UO_1374 (O_1374,N_24724,N_24144);
or UO_1375 (O_1375,N_24079,N_24565);
and UO_1376 (O_1376,N_24794,N_24467);
or UO_1377 (O_1377,N_24569,N_24566);
and UO_1378 (O_1378,N_24874,N_24523);
or UO_1379 (O_1379,N_24932,N_24690);
or UO_1380 (O_1380,N_24474,N_24056);
nand UO_1381 (O_1381,N_24055,N_24342);
or UO_1382 (O_1382,N_24420,N_24935);
and UO_1383 (O_1383,N_24280,N_24510);
xnor UO_1384 (O_1384,N_24600,N_24681);
and UO_1385 (O_1385,N_24978,N_24270);
xor UO_1386 (O_1386,N_24449,N_24668);
nand UO_1387 (O_1387,N_24368,N_24046);
nand UO_1388 (O_1388,N_24214,N_24602);
xor UO_1389 (O_1389,N_24731,N_24736);
nor UO_1390 (O_1390,N_24125,N_24259);
and UO_1391 (O_1391,N_24798,N_24732);
nand UO_1392 (O_1392,N_24622,N_24261);
or UO_1393 (O_1393,N_24035,N_24350);
or UO_1394 (O_1394,N_24522,N_24647);
or UO_1395 (O_1395,N_24882,N_24219);
or UO_1396 (O_1396,N_24538,N_24018);
nand UO_1397 (O_1397,N_24803,N_24345);
or UO_1398 (O_1398,N_24674,N_24550);
or UO_1399 (O_1399,N_24401,N_24071);
and UO_1400 (O_1400,N_24838,N_24735);
nor UO_1401 (O_1401,N_24264,N_24711);
or UO_1402 (O_1402,N_24795,N_24100);
xor UO_1403 (O_1403,N_24700,N_24743);
nor UO_1404 (O_1404,N_24728,N_24986);
nor UO_1405 (O_1405,N_24423,N_24526);
and UO_1406 (O_1406,N_24153,N_24995);
xnor UO_1407 (O_1407,N_24231,N_24709);
or UO_1408 (O_1408,N_24817,N_24514);
and UO_1409 (O_1409,N_24149,N_24991);
nor UO_1410 (O_1410,N_24319,N_24327);
nand UO_1411 (O_1411,N_24040,N_24847);
nor UO_1412 (O_1412,N_24331,N_24771);
nor UO_1413 (O_1413,N_24978,N_24735);
nand UO_1414 (O_1414,N_24250,N_24775);
nor UO_1415 (O_1415,N_24460,N_24053);
nand UO_1416 (O_1416,N_24370,N_24767);
nand UO_1417 (O_1417,N_24793,N_24940);
and UO_1418 (O_1418,N_24595,N_24004);
nand UO_1419 (O_1419,N_24803,N_24147);
or UO_1420 (O_1420,N_24426,N_24213);
nor UO_1421 (O_1421,N_24735,N_24185);
xor UO_1422 (O_1422,N_24289,N_24125);
xor UO_1423 (O_1423,N_24523,N_24461);
xnor UO_1424 (O_1424,N_24891,N_24492);
nand UO_1425 (O_1425,N_24872,N_24651);
or UO_1426 (O_1426,N_24549,N_24658);
nor UO_1427 (O_1427,N_24395,N_24442);
xnor UO_1428 (O_1428,N_24502,N_24344);
nand UO_1429 (O_1429,N_24616,N_24155);
xor UO_1430 (O_1430,N_24632,N_24630);
xnor UO_1431 (O_1431,N_24481,N_24938);
xor UO_1432 (O_1432,N_24586,N_24144);
or UO_1433 (O_1433,N_24691,N_24573);
xnor UO_1434 (O_1434,N_24083,N_24214);
or UO_1435 (O_1435,N_24548,N_24089);
nand UO_1436 (O_1436,N_24899,N_24065);
nor UO_1437 (O_1437,N_24692,N_24782);
and UO_1438 (O_1438,N_24575,N_24372);
and UO_1439 (O_1439,N_24114,N_24679);
or UO_1440 (O_1440,N_24758,N_24618);
or UO_1441 (O_1441,N_24867,N_24811);
nand UO_1442 (O_1442,N_24914,N_24132);
nand UO_1443 (O_1443,N_24353,N_24079);
nor UO_1444 (O_1444,N_24038,N_24296);
xnor UO_1445 (O_1445,N_24048,N_24734);
xor UO_1446 (O_1446,N_24053,N_24608);
xor UO_1447 (O_1447,N_24230,N_24995);
and UO_1448 (O_1448,N_24149,N_24241);
and UO_1449 (O_1449,N_24765,N_24554);
and UO_1450 (O_1450,N_24366,N_24848);
nand UO_1451 (O_1451,N_24968,N_24184);
or UO_1452 (O_1452,N_24463,N_24817);
xnor UO_1453 (O_1453,N_24654,N_24008);
or UO_1454 (O_1454,N_24136,N_24727);
xnor UO_1455 (O_1455,N_24604,N_24361);
nor UO_1456 (O_1456,N_24412,N_24952);
xnor UO_1457 (O_1457,N_24030,N_24359);
nand UO_1458 (O_1458,N_24953,N_24078);
and UO_1459 (O_1459,N_24199,N_24395);
nor UO_1460 (O_1460,N_24273,N_24187);
nand UO_1461 (O_1461,N_24871,N_24255);
nand UO_1462 (O_1462,N_24407,N_24539);
and UO_1463 (O_1463,N_24197,N_24077);
nor UO_1464 (O_1464,N_24154,N_24478);
nor UO_1465 (O_1465,N_24866,N_24376);
nand UO_1466 (O_1466,N_24778,N_24755);
xnor UO_1467 (O_1467,N_24077,N_24380);
xnor UO_1468 (O_1468,N_24745,N_24952);
or UO_1469 (O_1469,N_24855,N_24245);
nor UO_1470 (O_1470,N_24857,N_24620);
nand UO_1471 (O_1471,N_24674,N_24197);
xnor UO_1472 (O_1472,N_24039,N_24588);
xnor UO_1473 (O_1473,N_24265,N_24097);
xor UO_1474 (O_1474,N_24350,N_24333);
nand UO_1475 (O_1475,N_24855,N_24820);
nor UO_1476 (O_1476,N_24767,N_24409);
xor UO_1477 (O_1477,N_24589,N_24315);
nor UO_1478 (O_1478,N_24978,N_24288);
nand UO_1479 (O_1479,N_24912,N_24474);
nor UO_1480 (O_1480,N_24239,N_24621);
or UO_1481 (O_1481,N_24417,N_24979);
xnor UO_1482 (O_1482,N_24897,N_24988);
or UO_1483 (O_1483,N_24344,N_24486);
and UO_1484 (O_1484,N_24047,N_24325);
nor UO_1485 (O_1485,N_24936,N_24602);
or UO_1486 (O_1486,N_24231,N_24246);
or UO_1487 (O_1487,N_24472,N_24816);
or UO_1488 (O_1488,N_24655,N_24304);
xor UO_1489 (O_1489,N_24322,N_24268);
and UO_1490 (O_1490,N_24149,N_24458);
nor UO_1491 (O_1491,N_24760,N_24290);
nand UO_1492 (O_1492,N_24610,N_24224);
nor UO_1493 (O_1493,N_24850,N_24832);
nor UO_1494 (O_1494,N_24538,N_24315);
and UO_1495 (O_1495,N_24057,N_24520);
nor UO_1496 (O_1496,N_24584,N_24778);
and UO_1497 (O_1497,N_24864,N_24982);
nor UO_1498 (O_1498,N_24205,N_24624);
nor UO_1499 (O_1499,N_24167,N_24173);
or UO_1500 (O_1500,N_24293,N_24700);
or UO_1501 (O_1501,N_24035,N_24894);
or UO_1502 (O_1502,N_24187,N_24847);
or UO_1503 (O_1503,N_24926,N_24857);
xnor UO_1504 (O_1504,N_24090,N_24527);
and UO_1505 (O_1505,N_24533,N_24820);
and UO_1506 (O_1506,N_24492,N_24331);
nand UO_1507 (O_1507,N_24452,N_24445);
xor UO_1508 (O_1508,N_24957,N_24883);
xor UO_1509 (O_1509,N_24765,N_24933);
and UO_1510 (O_1510,N_24321,N_24674);
xor UO_1511 (O_1511,N_24934,N_24171);
or UO_1512 (O_1512,N_24169,N_24391);
nand UO_1513 (O_1513,N_24188,N_24024);
xor UO_1514 (O_1514,N_24186,N_24694);
nor UO_1515 (O_1515,N_24416,N_24531);
xnor UO_1516 (O_1516,N_24829,N_24212);
or UO_1517 (O_1517,N_24090,N_24962);
xnor UO_1518 (O_1518,N_24677,N_24660);
or UO_1519 (O_1519,N_24475,N_24443);
and UO_1520 (O_1520,N_24833,N_24611);
nor UO_1521 (O_1521,N_24238,N_24404);
nand UO_1522 (O_1522,N_24711,N_24106);
or UO_1523 (O_1523,N_24363,N_24947);
xnor UO_1524 (O_1524,N_24271,N_24091);
xor UO_1525 (O_1525,N_24573,N_24706);
and UO_1526 (O_1526,N_24248,N_24560);
xor UO_1527 (O_1527,N_24129,N_24900);
or UO_1528 (O_1528,N_24437,N_24443);
and UO_1529 (O_1529,N_24063,N_24624);
nand UO_1530 (O_1530,N_24264,N_24194);
and UO_1531 (O_1531,N_24403,N_24193);
and UO_1532 (O_1532,N_24390,N_24633);
xor UO_1533 (O_1533,N_24177,N_24199);
and UO_1534 (O_1534,N_24358,N_24593);
xor UO_1535 (O_1535,N_24894,N_24148);
xor UO_1536 (O_1536,N_24561,N_24459);
nand UO_1537 (O_1537,N_24879,N_24770);
or UO_1538 (O_1538,N_24874,N_24848);
and UO_1539 (O_1539,N_24133,N_24419);
xor UO_1540 (O_1540,N_24743,N_24838);
and UO_1541 (O_1541,N_24070,N_24782);
and UO_1542 (O_1542,N_24190,N_24225);
xnor UO_1543 (O_1543,N_24666,N_24496);
xor UO_1544 (O_1544,N_24081,N_24356);
xor UO_1545 (O_1545,N_24361,N_24407);
and UO_1546 (O_1546,N_24041,N_24102);
nand UO_1547 (O_1547,N_24306,N_24596);
xnor UO_1548 (O_1548,N_24595,N_24235);
and UO_1549 (O_1549,N_24676,N_24386);
and UO_1550 (O_1550,N_24695,N_24703);
and UO_1551 (O_1551,N_24178,N_24938);
and UO_1552 (O_1552,N_24577,N_24311);
or UO_1553 (O_1553,N_24149,N_24902);
or UO_1554 (O_1554,N_24004,N_24056);
xnor UO_1555 (O_1555,N_24829,N_24935);
nand UO_1556 (O_1556,N_24942,N_24408);
or UO_1557 (O_1557,N_24084,N_24071);
or UO_1558 (O_1558,N_24123,N_24556);
or UO_1559 (O_1559,N_24090,N_24569);
xor UO_1560 (O_1560,N_24549,N_24898);
nor UO_1561 (O_1561,N_24587,N_24522);
nor UO_1562 (O_1562,N_24228,N_24369);
xnor UO_1563 (O_1563,N_24918,N_24306);
and UO_1564 (O_1564,N_24035,N_24401);
and UO_1565 (O_1565,N_24660,N_24128);
xor UO_1566 (O_1566,N_24073,N_24923);
nand UO_1567 (O_1567,N_24230,N_24402);
nand UO_1568 (O_1568,N_24227,N_24282);
or UO_1569 (O_1569,N_24837,N_24371);
nand UO_1570 (O_1570,N_24422,N_24584);
xnor UO_1571 (O_1571,N_24798,N_24623);
nor UO_1572 (O_1572,N_24637,N_24611);
or UO_1573 (O_1573,N_24773,N_24700);
nor UO_1574 (O_1574,N_24509,N_24388);
or UO_1575 (O_1575,N_24386,N_24399);
or UO_1576 (O_1576,N_24051,N_24042);
nand UO_1577 (O_1577,N_24698,N_24805);
or UO_1578 (O_1578,N_24319,N_24302);
and UO_1579 (O_1579,N_24405,N_24819);
and UO_1580 (O_1580,N_24263,N_24353);
nor UO_1581 (O_1581,N_24933,N_24065);
and UO_1582 (O_1582,N_24482,N_24781);
or UO_1583 (O_1583,N_24087,N_24870);
nor UO_1584 (O_1584,N_24925,N_24462);
xor UO_1585 (O_1585,N_24065,N_24995);
nand UO_1586 (O_1586,N_24561,N_24038);
or UO_1587 (O_1587,N_24235,N_24462);
and UO_1588 (O_1588,N_24357,N_24964);
nand UO_1589 (O_1589,N_24236,N_24349);
or UO_1590 (O_1590,N_24549,N_24916);
nand UO_1591 (O_1591,N_24296,N_24818);
and UO_1592 (O_1592,N_24097,N_24923);
xor UO_1593 (O_1593,N_24191,N_24507);
nand UO_1594 (O_1594,N_24375,N_24294);
and UO_1595 (O_1595,N_24975,N_24378);
nor UO_1596 (O_1596,N_24935,N_24503);
nand UO_1597 (O_1597,N_24192,N_24261);
xnor UO_1598 (O_1598,N_24320,N_24071);
or UO_1599 (O_1599,N_24274,N_24383);
nand UO_1600 (O_1600,N_24218,N_24403);
nor UO_1601 (O_1601,N_24349,N_24237);
nor UO_1602 (O_1602,N_24368,N_24472);
nand UO_1603 (O_1603,N_24113,N_24489);
and UO_1604 (O_1604,N_24643,N_24070);
nor UO_1605 (O_1605,N_24088,N_24176);
nand UO_1606 (O_1606,N_24737,N_24394);
nor UO_1607 (O_1607,N_24405,N_24937);
nor UO_1608 (O_1608,N_24150,N_24723);
nand UO_1609 (O_1609,N_24475,N_24355);
xor UO_1610 (O_1610,N_24659,N_24863);
or UO_1611 (O_1611,N_24101,N_24647);
nor UO_1612 (O_1612,N_24127,N_24186);
and UO_1613 (O_1613,N_24850,N_24909);
xnor UO_1614 (O_1614,N_24429,N_24620);
or UO_1615 (O_1615,N_24197,N_24588);
or UO_1616 (O_1616,N_24047,N_24128);
nand UO_1617 (O_1617,N_24789,N_24427);
xor UO_1618 (O_1618,N_24302,N_24698);
and UO_1619 (O_1619,N_24308,N_24112);
nand UO_1620 (O_1620,N_24400,N_24181);
or UO_1621 (O_1621,N_24236,N_24951);
xnor UO_1622 (O_1622,N_24125,N_24785);
nor UO_1623 (O_1623,N_24874,N_24072);
xor UO_1624 (O_1624,N_24802,N_24338);
xnor UO_1625 (O_1625,N_24784,N_24883);
and UO_1626 (O_1626,N_24289,N_24587);
or UO_1627 (O_1627,N_24921,N_24962);
and UO_1628 (O_1628,N_24300,N_24996);
and UO_1629 (O_1629,N_24021,N_24731);
or UO_1630 (O_1630,N_24105,N_24972);
xnor UO_1631 (O_1631,N_24600,N_24130);
nor UO_1632 (O_1632,N_24035,N_24356);
nor UO_1633 (O_1633,N_24005,N_24694);
or UO_1634 (O_1634,N_24614,N_24077);
xor UO_1635 (O_1635,N_24942,N_24873);
xnor UO_1636 (O_1636,N_24581,N_24171);
and UO_1637 (O_1637,N_24075,N_24532);
nor UO_1638 (O_1638,N_24095,N_24965);
nor UO_1639 (O_1639,N_24870,N_24432);
xor UO_1640 (O_1640,N_24314,N_24021);
nand UO_1641 (O_1641,N_24402,N_24226);
nand UO_1642 (O_1642,N_24443,N_24912);
or UO_1643 (O_1643,N_24773,N_24244);
or UO_1644 (O_1644,N_24978,N_24785);
nor UO_1645 (O_1645,N_24028,N_24879);
nor UO_1646 (O_1646,N_24021,N_24516);
and UO_1647 (O_1647,N_24049,N_24827);
xnor UO_1648 (O_1648,N_24099,N_24729);
or UO_1649 (O_1649,N_24330,N_24708);
and UO_1650 (O_1650,N_24328,N_24315);
xnor UO_1651 (O_1651,N_24536,N_24487);
xnor UO_1652 (O_1652,N_24421,N_24648);
and UO_1653 (O_1653,N_24129,N_24515);
nor UO_1654 (O_1654,N_24733,N_24074);
and UO_1655 (O_1655,N_24283,N_24275);
nand UO_1656 (O_1656,N_24806,N_24689);
and UO_1657 (O_1657,N_24587,N_24470);
xor UO_1658 (O_1658,N_24670,N_24053);
nand UO_1659 (O_1659,N_24631,N_24082);
xor UO_1660 (O_1660,N_24421,N_24403);
and UO_1661 (O_1661,N_24494,N_24885);
xor UO_1662 (O_1662,N_24301,N_24032);
xor UO_1663 (O_1663,N_24021,N_24245);
nor UO_1664 (O_1664,N_24662,N_24198);
xnor UO_1665 (O_1665,N_24100,N_24653);
xnor UO_1666 (O_1666,N_24126,N_24919);
nor UO_1667 (O_1667,N_24688,N_24318);
nand UO_1668 (O_1668,N_24491,N_24212);
nand UO_1669 (O_1669,N_24844,N_24680);
nor UO_1670 (O_1670,N_24192,N_24644);
or UO_1671 (O_1671,N_24465,N_24452);
nand UO_1672 (O_1672,N_24974,N_24671);
xnor UO_1673 (O_1673,N_24064,N_24212);
nand UO_1674 (O_1674,N_24687,N_24265);
xor UO_1675 (O_1675,N_24986,N_24826);
and UO_1676 (O_1676,N_24796,N_24433);
nor UO_1677 (O_1677,N_24576,N_24534);
nand UO_1678 (O_1678,N_24402,N_24398);
nand UO_1679 (O_1679,N_24403,N_24019);
xor UO_1680 (O_1680,N_24102,N_24247);
xnor UO_1681 (O_1681,N_24211,N_24434);
nand UO_1682 (O_1682,N_24952,N_24030);
nand UO_1683 (O_1683,N_24739,N_24953);
nand UO_1684 (O_1684,N_24022,N_24775);
nand UO_1685 (O_1685,N_24972,N_24500);
nor UO_1686 (O_1686,N_24904,N_24248);
nand UO_1687 (O_1687,N_24430,N_24243);
xnor UO_1688 (O_1688,N_24288,N_24549);
or UO_1689 (O_1689,N_24883,N_24418);
xor UO_1690 (O_1690,N_24038,N_24180);
or UO_1691 (O_1691,N_24012,N_24745);
nand UO_1692 (O_1692,N_24986,N_24432);
and UO_1693 (O_1693,N_24211,N_24622);
nor UO_1694 (O_1694,N_24411,N_24724);
or UO_1695 (O_1695,N_24448,N_24377);
nor UO_1696 (O_1696,N_24813,N_24338);
xor UO_1697 (O_1697,N_24691,N_24663);
or UO_1698 (O_1698,N_24587,N_24182);
nor UO_1699 (O_1699,N_24632,N_24706);
or UO_1700 (O_1700,N_24727,N_24860);
nand UO_1701 (O_1701,N_24519,N_24016);
and UO_1702 (O_1702,N_24739,N_24242);
nand UO_1703 (O_1703,N_24797,N_24055);
nand UO_1704 (O_1704,N_24041,N_24502);
nor UO_1705 (O_1705,N_24497,N_24813);
and UO_1706 (O_1706,N_24901,N_24273);
or UO_1707 (O_1707,N_24101,N_24351);
or UO_1708 (O_1708,N_24004,N_24559);
nand UO_1709 (O_1709,N_24946,N_24837);
or UO_1710 (O_1710,N_24274,N_24819);
or UO_1711 (O_1711,N_24330,N_24415);
and UO_1712 (O_1712,N_24428,N_24684);
and UO_1713 (O_1713,N_24120,N_24519);
nor UO_1714 (O_1714,N_24399,N_24597);
nand UO_1715 (O_1715,N_24809,N_24956);
or UO_1716 (O_1716,N_24171,N_24308);
nor UO_1717 (O_1717,N_24579,N_24993);
and UO_1718 (O_1718,N_24778,N_24421);
and UO_1719 (O_1719,N_24835,N_24415);
nor UO_1720 (O_1720,N_24330,N_24016);
or UO_1721 (O_1721,N_24326,N_24873);
nand UO_1722 (O_1722,N_24991,N_24792);
and UO_1723 (O_1723,N_24221,N_24987);
xor UO_1724 (O_1724,N_24476,N_24293);
nor UO_1725 (O_1725,N_24792,N_24807);
nand UO_1726 (O_1726,N_24220,N_24200);
nor UO_1727 (O_1727,N_24288,N_24222);
nor UO_1728 (O_1728,N_24210,N_24132);
or UO_1729 (O_1729,N_24367,N_24265);
or UO_1730 (O_1730,N_24649,N_24804);
xor UO_1731 (O_1731,N_24097,N_24873);
xor UO_1732 (O_1732,N_24224,N_24909);
xnor UO_1733 (O_1733,N_24108,N_24263);
xnor UO_1734 (O_1734,N_24783,N_24866);
nor UO_1735 (O_1735,N_24545,N_24297);
and UO_1736 (O_1736,N_24454,N_24662);
xor UO_1737 (O_1737,N_24218,N_24596);
and UO_1738 (O_1738,N_24323,N_24509);
nor UO_1739 (O_1739,N_24273,N_24155);
xnor UO_1740 (O_1740,N_24888,N_24598);
xor UO_1741 (O_1741,N_24669,N_24641);
and UO_1742 (O_1742,N_24017,N_24234);
nor UO_1743 (O_1743,N_24614,N_24921);
or UO_1744 (O_1744,N_24905,N_24982);
or UO_1745 (O_1745,N_24463,N_24265);
nand UO_1746 (O_1746,N_24451,N_24468);
nand UO_1747 (O_1747,N_24620,N_24542);
xnor UO_1748 (O_1748,N_24359,N_24632);
nor UO_1749 (O_1749,N_24366,N_24251);
and UO_1750 (O_1750,N_24011,N_24195);
nand UO_1751 (O_1751,N_24697,N_24900);
nor UO_1752 (O_1752,N_24822,N_24889);
xnor UO_1753 (O_1753,N_24118,N_24537);
xnor UO_1754 (O_1754,N_24308,N_24096);
and UO_1755 (O_1755,N_24514,N_24348);
xnor UO_1756 (O_1756,N_24258,N_24344);
xor UO_1757 (O_1757,N_24340,N_24053);
nand UO_1758 (O_1758,N_24450,N_24944);
xnor UO_1759 (O_1759,N_24893,N_24539);
or UO_1760 (O_1760,N_24983,N_24964);
xnor UO_1761 (O_1761,N_24077,N_24081);
or UO_1762 (O_1762,N_24902,N_24198);
and UO_1763 (O_1763,N_24923,N_24160);
and UO_1764 (O_1764,N_24332,N_24242);
xnor UO_1765 (O_1765,N_24991,N_24837);
and UO_1766 (O_1766,N_24651,N_24743);
xor UO_1767 (O_1767,N_24157,N_24252);
xnor UO_1768 (O_1768,N_24864,N_24624);
and UO_1769 (O_1769,N_24981,N_24840);
and UO_1770 (O_1770,N_24675,N_24057);
and UO_1771 (O_1771,N_24076,N_24995);
or UO_1772 (O_1772,N_24630,N_24073);
nor UO_1773 (O_1773,N_24026,N_24901);
nor UO_1774 (O_1774,N_24291,N_24722);
xnor UO_1775 (O_1775,N_24225,N_24517);
nor UO_1776 (O_1776,N_24006,N_24470);
nand UO_1777 (O_1777,N_24735,N_24031);
nand UO_1778 (O_1778,N_24321,N_24886);
nand UO_1779 (O_1779,N_24675,N_24533);
and UO_1780 (O_1780,N_24074,N_24354);
and UO_1781 (O_1781,N_24766,N_24298);
nor UO_1782 (O_1782,N_24961,N_24201);
and UO_1783 (O_1783,N_24217,N_24956);
and UO_1784 (O_1784,N_24330,N_24488);
and UO_1785 (O_1785,N_24124,N_24414);
or UO_1786 (O_1786,N_24273,N_24860);
and UO_1787 (O_1787,N_24883,N_24102);
nor UO_1788 (O_1788,N_24686,N_24010);
and UO_1789 (O_1789,N_24107,N_24544);
nand UO_1790 (O_1790,N_24491,N_24376);
xor UO_1791 (O_1791,N_24969,N_24995);
nand UO_1792 (O_1792,N_24455,N_24136);
xnor UO_1793 (O_1793,N_24872,N_24393);
and UO_1794 (O_1794,N_24637,N_24217);
nand UO_1795 (O_1795,N_24781,N_24817);
and UO_1796 (O_1796,N_24987,N_24243);
or UO_1797 (O_1797,N_24822,N_24384);
xor UO_1798 (O_1798,N_24073,N_24274);
and UO_1799 (O_1799,N_24679,N_24244);
nor UO_1800 (O_1800,N_24144,N_24436);
nand UO_1801 (O_1801,N_24905,N_24162);
nand UO_1802 (O_1802,N_24640,N_24267);
nor UO_1803 (O_1803,N_24330,N_24962);
nor UO_1804 (O_1804,N_24838,N_24787);
nand UO_1805 (O_1805,N_24431,N_24225);
xnor UO_1806 (O_1806,N_24695,N_24563);
nand UO_1807 (O_1807,N_24776,N_24917);
xnor UO_1808 (O_1808,N_24936,N_24585);
xnor UO_1809 (O_1809,N_24360,N_24508);
and UO_1810 (O_1810,N_24998,N_24896);
nor UO_1811 (O_1811,N_24416,N_24331);
nor UO_1812 (O_1812,N_24486,N_24645);
nand UO_1813 (O_1813,N_24486,N_24126);
xor UO_1814 (O_1814,N_24818,N_24812);
or UO_1815 (O_1815,N_24237,N_24665);
or UO_1816 (O_1816,N_24929,N_24329);
xnor UO_1817 (O_1817,N_24719,N_24115);
xor UO_1818 (O_1818,N_24904,N_24648);
xnor UO_1819 (O_1819,N_24913,N_24600);
and UO_1820 (O_1820,N_24697,N_24149);
or UO_1821 (O_1821,N_24473,N_24887);
nor UO_1822 (O_1822,N_24362,N_24102);
or UO_1823 (O_1823,N_24262,N_24247);
nor UO_1824 (O_1824,N_24759,N_24486);
nor UO_1825 (O_1825,N_24199,N_24420);
nand UO_1826 (O_1826,N_24055,N_24231);
nand UO_1827 (O_1827,N_24000,N_24587);
and UO_1828 (O_1828,N_24058,N_24053);
and UO_1829 (O_1829,N_24358,N_24976);
and UO_1830 (O_1830,N_24038,N_24584);
xor UO_1831 (O_1831,N_24674,N_24768);
and UO_1832 (O_1832,N_24514,N_24359);
or UO_1833 (O_1833,N_24416,N_24428);
or UO_1834 (O_1834,N_24744,N_24674);
nand UO_1835 (O_1835,N_24249,N_24352);
and UO_1836 (O_1836,N_24480,N_24108);
nor UO_1837 (O_1837,N_24801,N_24213);
or UO_1838 (O_1838,N_24953,N_24877);
nand UO_1839 (O_1839,N_24248,N_24866);
and UO_1840 (O_1840,N_24522,N_24998);
or UO_1841 (O_1841,N_24749,N_24288);
nand UO_1842 (O_1842,N_24649,N_24364);
and UO_1843 (O_1843,N_24215,N_24810);
and UO_1844 (O_1844,N_24024,N_24350);
nand UO_1845 (O_1845,N_24994,N_24423);
nand UO_1846 (O_1846,N_24105,N_24476);
or UO_1847 (O_1847,N_24248,N_24253);
nand UO_1848 (O_1848,N_24707,N_24268);
xnor UO_1849 (O_1849,N_24746,N_24837);
nand UO_1850 (O_1850,N_24219,N_24837);
nand UO_1851 (O_1851,N_24240,N_24673);
nor UO_1852 (O_1852,N_24111,N_24881);
nor UO_1853 (O_1853,N_24628,N_24701);
xor UO_1854 (O_1854,N_24396,N_24601);
nand UO_1855 (O_1855,N_24701,N_24668);
and UO_1856 (O_1856,N_24673,N_24295);
xor UO_1857 (O_1857,N_24387,N_24003);
nor UO_1858 (O_1858,N_24753,N_24042);
nand UO_1859 (O_1859,N_24681,N_24834);
xnor UO_1860 (O_1860,N_24251,N_24323);
nor UO_1861 (O_1861,N_24095,N_24774);
and UO_1862 (O_1862,N_24657,N_24770);
xnor UO_1863 (O_1863,N_24173,N_24445);
xor UO_1864 (O_1864,N_24216,N_24428);
nor UO_1865 (O_1865,N_24847,N_24149);
and UO_1866 (O_1866,N_24957,N_24917);
and UO_1867 (O_1867,N_24531,N_24764);
xnor UO_1868 (O_1868,N_24003,N_24901);
nand UO_1869 (O_1869,N_24356,N_24704);
nor UO_1870 (O_1870,N_24304,N_24183);
or UO_1871 (O_1871,N_24396,N_24883);
xor UO_1872 (O_1872,N_24582,N_24533);
or UO_1873 (O_1873,N_24749,N_24086);
nor UO_1874 (O_1874,N_24781,N_24670);
or UO_1875 (O_1875,N_24753,N_24427);
nor UO_1876 (O_1876,N_24666,N_24343);
nand UO_1877 (O_1877,N_24920,N_24107);
nor UO_1878 (O_1878,N_24367,N_24553);
or UO_1879 (O_1879,N_24671,N_24233);
or UO_1880 (O_1880,N_24495,N_24880);
and UO_1881 (O_1881,N_24967,N_24416);
or UO_1882 (O_1882,N_24279,N_24704);
or UO_1883 (O_1883,N_24960,N_24469);
xnor UO_1884 (O_1884,N_24657,N_24661);
nor UO_1885 (O_1885,N_24475,N_24895);
and UO_1886 (O_1886,N_24240,N_24788);
nand UO_1887 (O_1887,N_24878,N_24585);
nand UO_1888 (O_1888,N_24559,N_24585);
and UO_1889 (O_1889,N_24911,N_24369);
xor UO_1890 (O_1890,N_24528,N_24676);
nor UO_1891 (O_1891,N_24443,N_24727);
and UO_1892 (O_1892,N_24227,N_24409);
and UO_1893 (O_1893,N_24259,N_24452);
and UO_1894 (O_1894,N_24241,N_24551);
nand UO_1895 (O_1895,N_24136,N_24260);
xnor UO_1896 (O_1896,N_24772,N_24015);
xor UO_1897 (O_1897,N_24974,N_24531);
xnor UO_1898 (O_1898,N_24621,N_24666);
and UO_1899 (O_1899,N_24662,N_24300);
nor UO_1900 (O_1900,N_24956,N_24372);
and UO_1901 (O_1901,N_24761,N_24805);
nand UO_1902 (O_1902,N_24700,N_24299);
nand UO_1903 (O_1903,N_24516,N_24919);
xor UO_1904 (O_1904,N_24358,N_24176);
xor UO_1905 (O_1905,N_24101,N_24837);
or UO_1906 (O_1906,N_24870,N_24710);
and UO_1907 (O_1907,N_24877,N_24322);
nand UO_1908 (O_1908,N_24217,N_24763);
and UO_1909 (O_1909,N_24516,N_24375);
xor UO_1910 (O_1910,N_24695,N_24006);
xnor UO_1911 (O_1911,N_24455,N_24196);
xor UO_1912 (O_1912,N_24226,N_24579);
and UO_1913 (O_1913,N_24957,N_24963);
nand UO_1914 (O_1914,N_24313,N_24098);
nand UO_1915 (O_1915,N_24753,N_24560);
nand UO_1916 (O_1916,N_24753,N_24166);
xnor UO_1917 (O_1917,N_24241,N_24747);
xor UO_1918 (O_1918,N_24108,N_24292);
nand UO_1919 (O_1919,N_24362,N_24133);
nor UO_1920 (O_1920,N_24006,N_24974);
or UO_1921 (O_1921,N_24926,N_24977);
or UO_1922 (O_1922,N_24190,N_24451);
nand UO_1923 (O_1923,N_24231,N_24465);
nor UO_1924 (O_1924,N_24221,N_24292);
nand UO_1925 (O_1925,N_24302,N_24125);
nor UO_1926 (O_1926,N_24594,N_24720);
nand UO_1927 (O_1927,N_24367,N_24617);
nand UO_1928 (O_1928,N_24623,N_24461);
or UO_1929 (O_1929,N_24968,N_24774);
nand UO_1930 (O_1930,N_24089,N_24814);
or UO_1931 (O_1931,N_24009,N_24507);
nand UO_1932 (O_1932,N_24724,N_24669);
xnor UO_1933 (O_1933,N_24688,N_24010);
or UO_1934 (O_1934,N_24204,N_24427);
nor UO_1935 (O_1935,N_24016,N_24832);
or UO_1936 (O_1936,N_24561,N_24207);
and UO_1937 (O_1937,N_24375,N_24114);
and UO_1938 (O_1938,N_24438,N_24677);
xnor UO_1939 (O_1939,N_24385,N_24005);
or UO_1940 (O_1940,N_24408,N_24422);
xnor UO_1941 (O_1941,N_24851,N_24896);
xor UO_1942 (O_1942,N_24882,N_24085);
or UO_1943 (O_1943,N_24342,N_24491);
xnor UO_1944 (O_1944,N_24348,N_24011);
xnor UO_1945 (O_1945,N_24654,N_24773);
and UO_1946 (O_1946,N_24263,N_24472);
nor UO_1947 (O_1947,N_24299,N_24717);
nand UO_1948 (O_1948,N_24944,N_24648);
nor UO_1949 (O_1949,N_24491,N_24802);
and UO_1950 (O_1950,N_24770,N_24956);
or UO_1951 (O_1951,N_24660,N_24364);
nor UO_1952 (O_1952,N_24009,N_24532);
nor UO_1953 (O_1953,N_24218,N_24066);
or UO_1954 (O_1954,N_24320,N_24712);
nor UO_1955 (O_1955,N_24399,N_24482);
nor UO_1956 (O_1956,N_24739,N_24358);
nand UO_1957 (O_1957,N_24960,N_24449);
xor UO_1958 (O_1958,N_24409,N_24988);
xor UO_1959 (O_1959,N_24099,N_24480);
nand UO_1960 (O_1960,N_24995,N_24529);
nor UO_1961 (O_1961,N_24200,N_24313);
nor UO_1962 (O_1962,N_24512,N_24835);
and UO_1963 (O_1963,N_24901,N_24628);
nand UO_1964 (O_1964,N_24531,N_24404);
nor UO_1965 (O_1965,N_24594,N_24814);
or UO_1966 (O_1966,N_24822,N_24589);
nor UO_1967 (O_1967,N_24755,N_24097);
nor UO_1968 (O_1968,N_24054,N_24737);
nor UO_1969 (O_1969,N_24723,N_24292);
nor UO_1970 (O_1970,N_24983,N_24659);
and UO_1971 (O_1971,N_24542,N_24486);
or UO_1972 (O_1972,N_24139,N_24676);
xor UO_1973 (O_1973,N_24270,N_24123);
xnor UO_1974 (O_1974,N_24983,N_24105);
xnor UO_1975 (O_1975,N_24027,N_24986);
nand UO_1976 (O_1976,N_24172,N_24796);
and UO_1977 (O_1977,N_24328,N_24162);
and UO_1978 (O_1978,N_24533,N_24954);
nor UO_1979 (O_1979,N_24733,N_24007);
and UO_1980 (O_1980,N_24517,N_24686);
nor UO_1981 (O_1981,N_24248,N_24021);
nor UO_1982 (O_1982,N_24817,N_24895);
or UO_1983 (O_1983,N_24211,N_24219);
or UO_1984 (O_1984,N_24262,N_24628);
or UO_1985 (O_1985,N_24747,N_24907);
xnor UO_1986 (O_1986,N_24673,N_24290);
nor UO_1987 (O_1987,N_24635,N_24147);
xnor UO_1988 (O_1988,N_24453,N_24082);
or UO_1989 (O_1989,N_24717,N_24364);
xor UO_1990 (O_1990,N_24909,N_24244);
or UO_1991 (O_1991,N_24877,N_24276);
and UO_1992 (O_1992,N_24481,N_24836);
xnor UO_1993 (O_1993,N_24260,N_24544);
nor UO_1994 (O_1994,N_24657,N_24527);
xnor UO_1995 (O_1995,N_24772,N_24572);
nand UO_1996 (O_1996,N_24298,N_24313);
nand UO_1997 (O_1997,N_24997,N_24090);
nor UO_1998 (O_1998,N_24077,N_24954);
nand UO_1999 (O_1999,N_24221,N_24126);
and UO_2000 (O_2000,N_24308,N_24728);
and UO_2001 (O_2001,N_24389,N_24879);
nor UO_2002 (O_2002,N_24120,N_24572);
xnor UO_2003 (O_2003,N_24056,N_24468);
nor UO_2004 (O_2004,N_24572,N_24092);
nor UO_2005 (O_2005,N_24356,N_24017);
or UO_2006 (O_2006,N_24634,N_24269);
nand UO_2007 (O_2007,N_24595,N_24220);
xor UO_2008 (O_2008,N_24961,N_24744);
or UO_2009 (O_2009,N_24274,N_24714);
xor UO_2010 (O_2010,N_24944,N_24490);
nand UO_2011 (O_2011,N_24909,N_24940);
nor UO_2012 (O_2012,N_24426,N_24089);
or UO_2013 (O_2013,N_24613,N_24551);
nor UO_2014 (O_2014,N_24737,N_24779);
nand UO_2015 (O_2015,N_24924,N_24675);
or UO_2016 (O_2016,N_24727,N_24007);
nor UO_2017 (O_2017,N_24698,N_24565);
xnor UO_2018 (O_2018,N_24314,N_24510);
and UO_2019 (O_2019,N_24773,N_24154);
and UO_2020 (O_2020,N_24909,N_24344);
and UO_2021 (O_2021,N_24987,N_24895);
nor UO_2022 (O_2022,N_24097,N_24197);
and UO_2023 (O_2023,N_24620,N_24212);
and UO_2024 (O_2024,N_24413,N_24525);
or UO_2025 (O_2025,N_24428,N_24552);
xor UO_2026 (O_2026,N_24547,N_24038);
and UO_2027 (O_2027,N_24951,N_24896);
or UO_2028 (O_2028,N_24169,N_24432);
and UO_2029 (O_2029,N_24910,N_24637);
and UO_2030 (O_2030,N_24792,N_24317);
or UO_2031 (O_2031,N_24647,N_24137);
nand UO_2032 (O_2032,N_24353,N_24694);
nor UO_2033 (O_2033,N_24368,N_24540);
nor UO_2034 (O_2034,N_24471,N_24675);
or UO_2035 (O_2035,N_24907,N_24384);
and UO_2036 (O_2036,N_24664,N_24543);
nand UO_2037 (O_2037,N_24885,N_24850);
xnor UO_2038 (O_2038,N_24546,N_24251);
and UO_2039 (O_2039,N_24767,N_24754);
xor UO_2040 (O_2040,N_24065,N_24283);
xor UO_2041 (O_2041,N_24413,N_24286);
nand UO_2042 (O_2042,N_24333,N_24897);
nand UO_2043 (O_2043,N_24395,N_24891);
or UO_2044 (O_2044,N_24267,N_24032);
and UO_2045 (O_2045,N_24415,N_24907);
or UO_2046 (O_2046,N_24453,N_24052);
and UO_2047 (O_2047,N_24301,N_24898);
nand UO_2048 (O_2048,N_24978,N_24472);
nand UO_2049 (O_2049,N_24970,N_24500);
nand UO_2050 (O_2050,N_24167,N_24253);
xor UO_2051 (O_2051,N_24193,N_24555);
nor UO_2052 (O_2052,N_24495,N_24196);
and UO_2053 (O_2053,N_24980,N_24867);
xnor UO_2054 (O_2054,N_24982,N_24641);
nand UO_2055 (O_2055,N_24817,N_24679);
xnor UO_2056 (O_2056,N_24698,N_24228);
or UO_2057 (O_2057,N_24536,N_24943);
and UO_2058 (O_2058,N_24345,N_24787);
nand UO_2059 (O_2059,N_24805,N_24726);
or UO_2060 (O_2060,N_24086,N_24421);
nor UO_2061 (O_2061,N_24714,N_24760);
or UO_2062 (O_2062,N_24829,N_24565);
and UO_2063 (O_2063,N_24350,N_24960);
or UO_2064 (O_2064,N_24485,N_24581);
nor UO_2065 (O_2065,N_24634,N_24022);
nor UO_2066 (O_2066,N_24570,N_24163);
or UO_2067 (O_2067,N_24138,N_24671);
nor UO_2068 (O_2068,N_24543,N_24447);
nand UO_2069 (O_2069,N_24325,N_24246);
and UO_2070 (O_2070,N_24451,N_24631);
xnor UO_2071 (O_2071,N_24094,N_24004);
xnor UO_2072 (O_2072,N_24085,N_24501);
and UO_2073 (O_2073,N_24823,N_24317);
nor UO_2074 (O_2074,N_24690,N_24088);
nand UO_2075 (O_2075,N_24411,N_24927);
or UO_2076 (O_2076,N_24057,N_24210);
and UO_2077 (O_2077,N_24927,N_24562);
or UO_2078 (O_2078,N_24669,N_24560);
nand UO_2079 (O_2079,N_24059,N_24297);
or UO_2080 (O_2080,N_24651,N_24738);
nor UO_2081 (O_2081,N_24366,N_24580);
nand UO_2082 (O_2082,N_24342,N_24906);
xor UO_2083 (O_2083,N_24267,N_24011);
xor UO_2084 (O_2084,N_24520,N_24505);
nor UO_2085 (O_2085,N_24037,N_24167);
nor UO_2086 (O_2086,N_24305,N_24492);
or UO_2087 (O_2087,N_24180,N_24857);
and UO_2088 (O_2088,N_24771,N_24662);
and UO_2089 (O_2089,N_24500,N_24152);
xnor UO_2090 (O_2090,N_24797,N_24621);
and UO_2091 (O_2091,N_24590,N_24932);
xnor UO_2092 (O_2092,N_24812,N_24554);
or UO_2093 (O_2093,N_24773,N_24568);
nor UO_2094 (O_2094,N_24084,N_24697);
nor UO_2095 (O_2095,N_24199,N_24702);
nand UO_2096 (O_2096,N_24319,N_24817);
nor UO_2097 (O_2097,N_24547,N_24343);
xor UO_2098 (O_2098,N_24564,N_24257);
xnor UO_2099 (O_2099,N_24382,N_24423);
xor UO_2100 (O_2100,N_24973,N_24130);
nor UO_2101 (O_2101,N_24869,N_24233);
and UO_2102 (O_2102,N_24155,N_24931);
and UO_2103 (O_2103,N_24396,N_24760);
or UO_2104 (O_2104,N_24047,N_24253);
or UO_2105 (O_2105,N_24061,N_24480);
nor UO_2106 (O_2106,N_24907,N_24700);
nand UO_2107 (O_2107,N_24056,N_24336);
nor UO_2108 (O_2108,N_24768,N_24824);
and UO_2109 (O_2109,N_24669,N_24360);
and UO_2110 (O_2110,N_24250,N_24900);
xnor UO_2111 (O_2111,N_24712,N_24285);
or UO_2112 (O_2112,N_24652,N_24934);
or UO_2113 (O_2113,N_24862,N_24433);
nor UO_2114 (O_2114,N_24326,N_24754);
and UO_2115 (O_2115,N_24848,N_24443);
nor UO_2116 (O_2116,N_24821,N_24155);
or UO_2117 (O_2117,N_24052,N_24065);
or UO_2118 (O_2118,N_24195,N_24224);
nor UO_2119 (O_2119,N_24386,N_24286);
and UO_2120 (O_2120,N_24559,N_24466);
and UO_2121 (O_2121,N_24143,N_24551);
nor UO_2122 (O_2122,N_24372,N_24831);
nand UO_2123 (O_2123,N_24310,N_24145);
and UO_2124 (O_2124,N_24900,N_24994);
and UO_2125 (O_2125,N_24152,N_24864);
nor UO_2126 (O_2126,N_24739,N_24094);
nor UO_2127 (O_2127,N_24886,N_24336);
or UO_2128 (O_2128,N_24686,N_24410);
or UO_2129 (O_2129,N_24127,N_24726);
nand UO_2130 (O_2130,N_24182,N_24406);
nand UO_2131 (O_2131,N_24008,N_24943);
or UO_2132 (O_2132,N_24307,N_24336);
and UO_2133 (O_2133,N_24222,N_24720);
or UO_2134 (O_2134,N_24495,N_24548);
or UO_2135 (O_2135,N_24028,N_24714);
and UO_2136 (O_2136,N_24076,N_24063);
nand UO_2137 (O_2137,N_24036,N_24937);
nand UO_2138 (O_2138,N_24504,N_24964);
nand UO_2139 (O_2139,N_24343,N_24331);
nor UO_2140 (O_2140,N_24481,N_24646);
and UO_2141 (O_2141,N_24987,N_24171);
or UO_2142 (O_2142,N_24092,N_24663);
and UO_2143 (O_2143,N_24650,N_24473);
and UO_2144 (O_2144,N_24925,N_24544);
nor UO_2145 (O_2145,N_24059,N_24024);
and UO_2146 (O_2146,N_24814,N_24965);
xor UO_2147 (O_2147,N_24649,N_24284);
and UO_2148 (O_2148,N_24251,N_24742);
nor UO_2149 (O_2149,N_24123,N_24277);
or UO_2150 (O_2150,N_24001,N_24732);
or UO_2151 (O_2151,N_24375,N_24759);
nand UO_2152 (O_2152,N_24855,N_24610);
or UO_2153 (O_2153,N_24844,N_24684);
and UO_2154 (O_2154,N_24868,N_24452);
nor UO_2155 (O_2155,N_24359,N_24209);
xnor UO_2156 (O_2156,N_24661,N_24517);
and UO_2157 (O_2157,N_24840,N_24892);
xor UO_2158 (O_2158,N_24752,N_24214);
nor UO_2159 (O_2159,N_24212,N_24992);
and UO_2160 (O_2160,N_24098,N_24349);
nor UO_2161 (O_2161,N_24413,N_24983);
nand UO_2162 (O_2162,N_24834,N_24450);
nor UO_2163 (O_2163,N_24895,N_24044);
nor UO_2164 (O_2164,N_24397,N_24863);
or UO_2165 (O_2165,N_24236,N_24448);
nor UO_2166 (O_2166,N_24203,N_24123);
nand UO_2167 (O_2167,N_24173,N_24088);
xor UO_2168 (O_2168,N_24915,N_24507);
nor UO_2169 (O_2169,N_24745,N_24388);
or UO_2170 (O_2170,N_24878,N_24649);
and UO_2171 (O_2171,N_24711,N_24583);
nor UO_2172 (O_2172,N_24771,N_24157);
xor UO_2173 (O_2173,N_24436,N_24869);
nand UO_2174 (O_2174,N_24292,N_24841);
and UO_2175 (O_2175,N_24374,N_24834);
and UO_2176 (O_2176,N_24630,N_24352);
nor UO_2177 (O_2177,N_24131,N_24605);
nand UO_2178 (O_2178,N_24349,N_24481);
nor UO_2179 (O_2179,N_24404,N_24120);
xor UO_2180 (O_2180,N_24435,N_24066);
nor UO_2181 (O_2181,N_24979,N_24978);
nand UO_2182 (O_2182,N_24688,N_24741);
nand UO_2183 (O_2183,N_24197,N_24654);
and UO_2184 (O_2184,N_24359,N_24378);
xor UO_2185 (O_2185,N_24022,N_24097);
or UO_2186 (O_2186,N_24352,N_24232);
or UO_2187 (O_2187,N_24914,N_24863);
and UO_2188 (O_2188,N_24910,N_24189);
nor UO_2189 (O_2189,N_24309,N_24093);
nand UO_2190 (O_2190,N_24103,N_24085);
and UO_2191 (O_2191,N_24374,N_24400);
xor UO_2192 (O_2192,N_24733,N_24521);
or UO_2193 (O_2193,N_24528,N_24819);
nand UO_2194 (O_2194,N_24586,N_24610);
xnor UO_2195 (O_2195,N_24210,N_24773);
or UO_2196 (O_2196,N_24963,N_24397);
nor UO_2197 (O_2197,N_24100,N_24433);
and UO_2198 (O_2198,N_24385,N_24187);
or UO_2199 (O_2199,N_24052,N_24061);
and UO_2200 (O_2200,N_24643,N_24777);
or UO_2201 (O_2201,N_24919,N_24250);
nor UO_2202 (O_2202,N_24168,N_24891);
xor UO_2203 (O_2203,N_24483,N_24293);
nand UO_2204 (O_2204,N_24950,N_24458);
and UO_2205 (O_2205,N_24938,N_24421);
and UO_2206 (O_2206,N_24916,N_24147);
xnor UO_2207 (O_2207,N_24714,N_24801);
and UO_2208 (O_2208,N_24912,N_24742);
nor UO_2209 (O_2209,N_24229,N_24815);
xor UO_2210 (O_2210,N_24194,N_24730);
nor UO_2211 (O_2211,N_24374,N_24735);
nor UO_2212 (O_2212,N_24233,N_24506);
nor UO_2213 (O_2213,N_24644,N_24221);
xor UO_2214 (O_2214,N_24632,N_24605);
nor UO_2215 (O_2215,N_24302,N_24276);
or UO_2216 (O_2216,N_24583,N_24411);
or UO_2217 (O_2217,N_24095,N_24685);
nor UO_2218 (O_2218,N_24663,N_24658);
nor UO_2219 (O_2219,N_24002,N_24111);
or UO_2220 (O_2220,N_24674,N_24549);
xor UO_2221 (O_2221,N_24719,N_24132);
nand UO_2222 (O_2222,N_24685,N_24471);
nand UO_2223 (O_2223,N_24488,N_24628);
or UO_2224 (O_2224,N_24506,N_24683);
and UO_2225 (O_2225,N_24366,N_24477);
nor UO_2226 (O_2226,N_24458,N_24400);
xnor UO_2227 (O_2227,N_24929,N_24363);
xnor UO_2228 (O_2228,N_24923,N_24729);
nand UO_2229 (O_2229,N_24458,N_24673);
xnor UO_2230 (O_2230,N_24692,N_24906);
nand UO_2231 (O_2231,N_24884,N_24723);
nand UO_2232 (O_2232,N_24728,N_24644);
and UO_2233 (O_2233,N_24062,N_24872);
and UO_2234 (O_2234,N_24548,N_24410);
or UO_2235 (O_2235,N_24578,N_24610);
nor UO_2236 (O_2236,N_24716,N_24407);
nor UO_2237 (O_2237,N_24135,N_24575);
or UO_2238 (O_2238,N_24519,N_24395);
or UO_2239 (O_2239,N_24891,N_24747);
or UO_2240 (O_2240,N_24810,N_24020);
nand UO_2241 (O_2241,N_24813,N_24540);
nand UO_2242 (O_2242,N_24652,N_24361);
xor UO_2243 (O_2243,N_24867,N_24289);
nand UO_2244 (O_2244,N_24216,N_24504);
nand UO_2245 (O_2245,N_24481,N_24780);
xor UO_2246 (O_2246,N_24784,N_24689);
xor UO_2247 (O_2247,N_24339,N_24504);
nor UO_2248 (O_2248,N_24233,N_24917);
xor UO_2249 (O_2249,N_24527,N_24262);
nor UO_2250 (O_2250,N_24468,N_24018);
nor UO_2251 (O_2251,N_24415,N_24758);
and UO_2252 (O_2252,N_24931,N_24656);
or UO_2253 (O_2253,N_24759,N_24543);
nor UO_2254 (O_2254,N_24307,N_24299);
and UO_2255 (O_2255,N_24035,N_24113);
or UO_2256 (O_2256,N_24087,N_24647);
xnor UO_2257 (O_2257,N_24834,N_24868);
nand UO_2258 (O_2258,N_24560,N_24953);
or UO_2259 (O_2259,N_24849,N_24171);
or UO_2260 (O_2260,N_24071,N_24010);
nor UO_2261 (O_2261,N_24211,N_24713);
and UO_2262 (O_2262,N_24363,N_24823);
or UO_2263 (O_2263,N_24064,N_24388);
xor UO_2264 (O_2264,N_24773,N_24120);
nor UO_2265 (O_2265,N_24099,N_24596);
nor UO_2266 (O_2266,N_24669,N_24486);
and UO_2267 (O_2267,N_24559,N_24903);
or UO_2268 (O_2268,N_24209,N_24801);
nor UO_2269 (O_2269,N_24780,N_24745);
or UO_2270 (O_2270,N_24111,N_24820);
and UO_2271 (O_2271,N_24028,N_24530);
nand UO_2272 (O_2272,N_24570,N_24050);
xor UO_2273 (O_2273,N_24325,N_24034);
or UO_2274 (O_2274,N_24858,N_24246);
nand UO_2275 (O_2275,N_24689,N_24243);
or UO_2276 (O_2276,N_24144,N_24378);
nor UO_2277 (O_2277,N_24977,N_24129);
nor UO_2278 (O_2278,N_24805,N_24493);
nor UO_2279 (O_2279,N_24336,N_24969);
or UO_2280 (O_2280,N_24359,N_24446);
or UO_2281 (O_2281,N_24736,N_24928);
and UO_2282 (O_2282,N_24282,N_24203);
nor UO_2283 (O_2283,N_24157,N_24159);
nand UO_2284 (O_2284,N_24675,N_24341);
or UO_2285 (O_2285,N_24778,N_24598);
nor UO_2286 (O_2286,N_24544,N_24243);
xor UO_2287 (O_2287,N_24100,N_24688);
and UO_2288 (O_2288,N_24474,N_24405);
nor UO_2289 (O_2289,N_24130,N_24657);
nand UO_2290 (O_2290,N_24179,N_24287);
and UO_2291 (O_2291,N_24575,N_24819);
and UO_2292 (O_2292,N_24374,N_24548);
or UO_2293 (O_2293,N_24591,N_24217);
xnor UO_2294 (O_2294,N_24063,N_24056);
nand UO_2295 (O_2295,N_24767,N_24961);
xnor UO_2296 (O_2296,N_24632,N_24374);
and UO_2297 (O_2297,N_24800,N_24825);
nor UO_2298 (O_2298,N_24636,N_24388);
xor UO_2299 (O_2299,N_24794,N_24349);
nand UO_2300 (O_2300,N_24146,N_24809);
nor UO_2301 (O_2301,N_24554,N_24187);
nor UO_2302 (O_2302,N_24411,N_24464);
and UO_2303 (O_2303,N_24580,N_24526);
and UO_2304 (O_2304,N_24168,N_24022);
and UO_2305 (O_2305,N_24531,N_24440);
or UO_2306 (O_2306,N_24491,N_24662);
xor UO_2307 (O_2307,N_24650,N_24350);
xor UO_2308 (O_2308,N_24110,N_24398);
and UO_2309 (O_2309,N_24997,N_24327);
and UO_2310 (O_2310,N_24808,N_24614);
nor UO_2311 (O_2311,N_24758,N_24442);
nor UO_2312 (O_2312,N_24157,N_24352);
or UO_2313 (O_2313,N_24770,N_24409);
nor UO_2314 (O_2314,N_24623,N_24773);
or UO_2315 (O_2315,N_24034,N_24027);
nor UO_2316 (O_2316,N_24837,N_24378);
and UO_2317 (O_2317,N_24883,N_24828);
or UO_2318 (O_2318,N_24018,N_24811);
xor UO_2319 (O_2319,N_24867,N_24325);
or UO_2320 (O_2320,N_24457,N_24191);
and UO_2321 (O_2321,N_24078,N_24682);
or UO_2322 (O_2322,N_24568,N_24823);
nor UO_2323 (O_2323,N_24520,N_24399);
xnor UO_2324 (O_2324,N_24084,N_24430);
or UO_2325 (O_2325,N_24164,N_24765);
xnor UO_2326 (O_2326,N_24639,N_24748);
xor UO_2327 (O_2327,N_24333,N_24385);
and UO_2328 (O_2328,N_24437,N_24426);
or UO_2329 (O_2329,N_24790,N_24634);
xor UO_2330 (O_2330,N_24400,N_24936);
and UO_2331 (O_2331,N_24423,N_24750);
nor UO_2332 (O_2332,N_24933,N_24402);
and UO_2333 (O_2333,N_24415,N_24911);
xnor UO_2334 (O_2334,N_24642,N_24352);
or UO_2335 (O_2335,N_24225,N_24564);
xor UO_2336 (O_2336,N_24407,N_24047);
or UO_2337 (O_2337,N_24632,N_24736);
nand UO_2338 (O_2338,N_24829,N_24184);
and UO_2339 (O_2339,N_24502,N_24590);
and UO_2340 (O_2340,N_24849,N_24952);
or UO_2341 (O_2341,N_24362,N_24233);
nand UO_2342 (O_2342,N_24626,N_24042);
xnor UO_2343 (O_2343,N_24694,N_24002);
nand UO_2344 (O_2344,N_24915,N_24983);
nor UO_2345 (O_2345,N_24403,N_24239);
nand UO_2346 (O_2346,N_24587,N_24901);
xnor UO_2347 (O_2347,N_24359,N_24434);
xor UO_2348 (O_2348,N_24760,N_24498);
nand UO_2349 (O_2349,N_24720,N_24550);
and UO_2350 (O_2350,N_24130,N_24381);
nand UO_2351 (O_2351,N_24217,N_24586);
nor UO_2352 (O_2352,N_24070,N_24762);
xor UO_2353 (O_2353,N_24026,N_24727);
or UO_2354 (O_2354,N_24086,N_24961);
nor UO_2355 (O_2355,N_24008,N_24169);
nor UO_2356 (O_2356,N_24910,N_24710);
xor UO_2357 (O_2357,N_24185,N_24444);
xnor UO_2358 (O_2358,N_24711,N_24545);
nand UO_2359 (O_2359,N_24279,N_24403);
nand UO_2360 (O_2360,N_24741,N_24977);
nor UO_2361 (O_2361,N_24681,N_24175);
xnor UO_2362 (O_2362,N_24337,N_24102);
xnor UO_2363 (O_2363,N_24697,N_24022);
xnor UO_2364 (O_2364,N_24104,N_24907);
nand UO_2365 (O_2365,N_24223,N_24526);
nor UO_2366 (O_2366,N_24115,N_24842);
and UO_2367 (O_2367,N_24106,N_24869);
nand UO_2368 (O_2368,N_24651,N_24474);
or UO_2369 (O_2369,N_24042,N_24465);
xnor UO_2370 (O_2370,N_24072,N_24654);
nand UO_2371 (O_2371,N_24670,N_24954);
or UO_2372 (O_2372,N_24171,N_24660);
and UO_2373 (O_2373,N_24069,N_24776);
xnor UO_2374 (O_2374,N_24169,N_24828);
nor UO_2375 (O_2375,N_24577,N_24735);
and UO_2376 (O_2376,N_24333,N_24319);
or UO_2377 (O_2377,N_24542,N_24766);
or UO_2378 (O_2378,N_24186,N_24775);
nand UO_2379 (O_2379,N_24776,N_24393);
nand UO_2380 (O_2380,N_24998,N_24946);
or UO_2381 (O_2381,N_24551,N_24323);
and UO_2382 (O_2382,N_24005,N_24061);
xor UO_2383 (O_2383,N_24293,N_24875);
xor UO_2384 (O_2384,N_24007,N_24223);
xnor UO_2385 (O_2385,N_24106,N_24150);
or UO_2386 (O_2386,N_24730,N_24168);
or UO_2387 (O_2387,N_24753,N_24553);
or UO_2388 (O_2388,N_24718,N_24901);
nor UO_2389 (O_2389,N_24912,N_24771);
xnor UO_2390 (O_2390,N_24282,N_24762);
nor UO_2391 (O_2391,N_24486,N_24724);
nor UO_2392 (O_2392,N_24136,N_24171);
nand UO_2393 (O_2393,N_24417,N_24760);
nor UO_2394 (O_2394,N_24488,N_24685);
nand UO_2395 (O_2395,N_24566,N_24290);
and UO_2396 (O_2396,N_24260,N_24912);
nor UO_2397 (O_2397,N_24381,N_24869);
xnor UO_2398 (O_2398,N_24572,N_24747);
xor UO_2399 (O_2399,N_24702,N_24248);
nor UO_2400 (O_2400,N_24021,N_24520);
nor UO_2401 (O_2401,N_24466,N_24830);
nand UO_2402 (O_2402,N_24560,N_24700);
nor UO_2403 (O_2403,N_24365,N_24777);
nor UO_2404 (O_2404,N_24218,N_24032);
or UO_2405 (O_2405,N_24354,N_24271);
xor UO_2406 (O_2406,N_24233,N_24649);
nand UO_2407 (O_2407,N_24690,N_24049);
and UO_2408 (O_2408,N_24055,N_24256);
xor UO_2409 (O_2409,N_24173,N_24566);
xor UO_2410 (O_2410,N_24807,N_24031);
nand UO_2411 (O_2411,N_24389,N_24419);
or UO_2412 (O_2412,N_24224,N_24101);
nand UO_2413 (O_2413,N_24604,N_24463);
and UO_2414 (O_2414,N_24759,N_24945);
nor UO_2415 (O_2415,N_24256,N_24493);
nand UO_2416 (O_2416,N_24802,N_24179);
nand UO_2417 (O_2417,N_24351,N_24991);
nor UO_2418 (O_2418,N_24960,N_24825);
and UO_2419 (O_2419,N_24414,N_24162);
xnor UO_2420 (O_2420,N_24584,N_24635);
nor UO_2421 (O_2421,N_24523,N_24083);
xnor UO_2422 (O_2422,N_24706,N_24263);
and UO_2423 (O_2423,N_24914,N_24076);
nor UO_2424 (O_2424,N_24048,N_24313);
and UO_2425 (O_2425,N_24327,N_24698);
xnor UO_2426 (O_2426,N_24327,N_24853);
nor UO_2427 (O_2427,N_24500,N_24740);
or UO_2428 (O_2428,N_24336,N_24219);
or UO_2429 (O_2429,N_24704,N_24437);
and UO_2430 (O_2430,N_24393,N_24300);
nand UO_2431 (O_2431,N_24988,N_24152);
or UO_2432 (O_2432,N_24511,N_24508);
or UO_2433 (O_2433,N_24326,N_24170);
xnor UO_2434 (O_2434,N_24058,N_24518);
xnor UO_2435 (O_2435,N_24343,N_24973);
and UO_2436 (O_2436,N_24721,N_24724);
nor UO_2437 (O_2437,N_24703,N_24842);
nand UO_2438 (O_2438,N_24577,N_24225);
nor UO_2439 (O_2439,N_24016,N_24545);
nor UO_2440 (O_2440,N_24069,N_24790);
nor UO_2441 (O_2441,N_24669,N_24665);
xnor UO_2442 (O_2442,N_24944,N_24387);
nand UO_2443 (O_2443,N_24034,N_24319);
nand UO_2444 (O_2444,N_24253,N_24858);
nor UO_2445 (O_2445,N_24220,N_24251);
or UO_2446 (O_2446,N_24698,N_24039);
nor UO_2447 (O_2447,N_24409,N_24736);
nand UO_2448 (O_2448,N_24831,N_24888);
or UO_2449 (O_2449,N_24745,N_24799);
or UO_2450 (O_2450,N_24235,N_24379);
xnor UO_2451 (O_2451,N_24141,N_24362);
nand UO_2452 (O_2452,N_24900,N_24413);
or UO_2453 (O_2453,N_24050,N_24761);
or UO_2454 (O_2454,N_24725,N_24608);
nor UO_2455 (O_2455,N_24804,N_24926);
or UO_2456 (O_2456,N_24693,N_24175);
or UO_2457 (O_2457,N_24131,N_24452);
nand UO_2458 (O_2458,N_24482,N_24726);
nand UO_2459 (O_2459,N_24061,N_24841);
or UO_2460 (O_2460,N_24140,N_24095);
xnor UO_2461 (O_2461,N_24124,N_24563);
nor UO_2462 (O_2462,N_24842,N_24503);
or UO_2463 (O_2463,N_24084,N_24449);
nand UO_2464 (O_2464,N_24538,N_24833);
nand UO_2465 (O_2465,N_24830,N_24804);
nand UO_2466 (O_2466,N_24082,N_24686);
nand UO_2467 (O_2467,N_24522,N_24788);
xor UO_2468 (O_2468,N_24662,N_24213);
and UO_2469 (O_2469,N_24914,N_24497);
nand UO_2470 (O_2470,N_24878,N_24413);
xor UO_2471 (O_2471,N_24143,N_24685);
or UO_2472 (O_2472,N_24015,N_24397);
and UO_2473 (O_2473,N_24685,N_24541);
and UO_2474 (O_2474,N_24361,N_24941);
and UO_2475 (O_2475,N_24122,N_24707);
and UO_2476 (O_2476,N_24153,N_24277);
and UO_2477 (O_2477,N_24064,N_24513);
nor UO_2478 (O_2478,N_24868,N_24368);
and UO_2479 (O_2479,N_24854,N_24745);
xor UO_2480 (O_2480,N_24450,N_24845);
and UO_2481 (O_2481,N_24629,N_24212);
or UO_2482 (O_2482,N_24286,N_24221);
xnor UO_2483 (O_2483,N_24391,N_24867);
nand UO_2484 (O_2484,N_24413,N_24341);
or UO_2485 (O_2485,N_24445,N_24739);
and UO_2486 (O_2486,N_24773,N_24644);
and UO_2487 (O_2487,N_24472,N_24784);
or UO_2488 (O_2488,N_24164,N_24030);
nor UO_2489 (O_2489,N_24921,N_24698);
and UO_2490 (O_2490,N_24038,N_24752);
or UO_2491 (O_2491,N_24427,N_24077);
or UO_2492 (O_2492,N_24828,N_24306);
xor UO_2493 (O_2493,N_24503,N_24716);
nor UO_2494 (O_2494,N_24550,N_24322);
and UO_2495 (O_2495,N_24645,N_24635);
nor UO_2496 (O_2496,N_24787,N_24818);
or UO_2497 (O_2497,N_24920,N_24495);
nand UO_2498 (O_2498,N_24688,N_24029);
nor UO_2499 (O_2499,N_24746,N_24768);
nor UO_2500 (O_2500,N_24985,N_24174);
nand UO_2501 (O_2501,N_24066,N_24840);
xor UO_2502 (O_2502,N_24326,N_24564);
nand UO_2503 (O_2503,N_24043,N_24870);
nand UO_2504 (O_2504,N_24181,N_24774);
or UO_2505 (O_2505,N_24561,N_24873);
or UO_2506 (O_2506,N_24707,N_24354);
and UO_2507 (O_2507,N_24324,N_24134);
and UO_2508 (O_2508,N_24815,N_24523);
xor UO_2509 (O_2509,N_24789,N_24838);
and UO_2510 (O_2510,N_24101,N_24729);
nor UO_2511 (O_2511,N_24283,N_24294);
and UO_2512 (O_2512,N_24459,N_24828);
nand UO_2513 (O_2513,N_24827,N_24110);
nand UO_2514 (O_2514,N_24556,N_24044);
nand UO_2515 (O_2515,N_24579,N_24920);
xnor UO_2516 (O_2516,N_24627,N_24788);
xnor UO_2517 (O_2517,N_24986,N_24399);
xor UO_2518 (O_2518,N_24002,N_24593);
nand UO_2519 (O_2519,N_24680,N_24724);
nand UO_2520 (O_2520,N_24719,N_24226);
nand UO_2521 (O_2521,N_24028,N_24689);
or UO_2522 (O_2522,N_24970,N_24534);
nor UO_2523 (O_2523,N_24379,N_24072);
xnor UO_2524 (O_2524,N_24485,N_24342);
xnor UO_2525 (O_2525,N_24521,N_24527);
and UO_2526 (O_2526,N_24535,N_24259);
and UO_2527 (O_2527,N_24333,N_24437);
nor UO_2528 (O_2528,N_24389,N_24263);
xor UO_2529 (O_2529,N_24175,N_24882);
nand UO_2530 (O_2530,N_24181,N_24754);
nor UO_2531 (O_2531,N_24346,N_24140);
xnor UO_2532 (O_2532,N_24180,N_24089);
or UO_2533 (O_2533,N_24373,N_24503);
nor UO_2534 (O_2534,N_24180,N_24125);
nand UO_2535 (O_2535,N_24853,N_24811);
nor UO_2536 (O_2536,N_24014,N_24460);
nor UO_2537 (O_2537,N_24484,N_24941);
nor UO_2538 (O_2538,N_24215,N_24889);
nand UO_2539 (O_2539,N_24753,N_24074);
and UO_2540 (O_2540,N_24652,N_24183);
xor UO_2541 (O_2541,N_24003,N_24872);
or UO_2542 (O_2542,N_24351,N_24228);
or UO_2543 (O_2543,N_24800,N_24776);
xor UO_2544 (O_2544,N_24968,N_24263);
or UO_2545 (O_2545,N_24987,N_24935);
xor UO_2546 (O_2546,N_24144,N_24295);
nor UO_2547 (O_2547,N_24213,N_24543);
xnor UO_2548 (O_2548,N_24633,N_24748);
and UO_2549 (O_2549,N_24342,N_24246);
nand UO_2550 (O_2550,N_24230,N_24974);
or UO_2551 (O_2551,N_24296,N_24268);
xor UO_2552 (O_2552,N_24539,N_24478);
nor UO_2553 (O_2553,N_24312,N_24610);
or UO_2554 (O_2554,N_24678,N_24454);
nand UO_2555 (O_2555,N_24028,N_24638);
xnor UO_2556 (O_2556,N_24968,N_24431);
nand UO_2557 (O_2557,N_24926,N_24282);
nand UO_2558 (O_2558,N_24582,N_24938);
and UO_2559 (O_2559,N_24004,N_24891);
nand UO_2560 (O_2560,N_24888,N_24091);
nor UO_2561 (O_2561,N_24710,N_24143);
or UO_2562 (O_2562,N_24954,N_24551);
xor UO_2563 (O_2563,N_24055,N_24753);
nand UO_2564 (O_2564,N_24319,N_24937);
nand UO_2565 (O_2565,N_24931,N_24119);
nor UO_2566 (O_2566,N_24850,N_24876);
and UO_2567 (O_2567,N_24056,N_24692);
or UO_2568 (O_2568,N_24339,N_24867);
nand UO_2569 (O_2569,N_24614,N_24917);
xor UO_2570 (O_2570,N_24000,N_24291);
nand UO_2571 (O_2571,N_24341,N_24596);
or UO_2572 (O_2572,N_24688,N_24960);
or UO_2573 (O_2573,N_24859,N_24675);
xnor UO_2574 (O_2574,N_24455,N_24120);
and UO_2575 (O_2575,N_24941,N_24803);
or UO_2576 (O_2576,N_24596,N_24680);
and UO_2577 (O_2577,N_24811,N_24637);
nand UO_2578 (O_2578,N_24104,N_24438);
and UO_2579 (O_2579,N_24019,N_24281);
nor UO_2580 (O_2580,N_24127,N_24231);
nor UO_2581 (O_2581,N_24160,N_24106);
and UO_2582 (O_2582,N_24337,N_24559);
or UO_2583 (O_2583,N_24268,N_24571);
or UO_2584 (O_2584,N_24220,N_24093);
xor UO_2585 (O_2585,N_24615,N_24974);
xnor UO_2586 (O_2586,N_24002,N_24969);
xor UO_2587 (O_2587,N_24413,N_24848);
or UO_2588 (O_2588,N_24425,N_24848);
or UO_2589 (O_2589,N_24625,N_24504);
and UO_2590 (O_2590,N_24816,N_24095);
nor UO_2591 (O_2591,N_24284,N_24582);
and UO_2592 (O_2592,N_24578,N_24584);
nor UO_2593 (O_2593,N_24350,N_24822);
xor UO_2594 (O_2594,N_24524,N_24934);
xnor UO_2595 (O_2595,N_24076,N_24083);
or UO_2596 (O_2596,N_24126,N_24604);
or UO_2597 (O_2597,N_24898,N_24804);
nand UO_2598 (O_2598,N_24095,N_24280);
and UO_2599 (O_2599,N_24512,N_24545);
or UO_2600 (O_2600,N_24670,N_24813);
nand UO_2601 (O_2601,N_24355,N_24849);
and UO_2602 (O_2602,N_24192,N_24514);
or UO_2603 (O_2603,N_24146,N_24504);
or UO_2604 (O_2604,N_24389,N_24936);
nand UO_2605 (O_2605,N_24893,N_24253);
or UO_2606 (O_2606,N_24779,N_24007);
xnor UO_2607 (O_2607,N_24156,N_24362);
and UO_2608 (O_2608,N_24379,N_24005);
xor UO_2609 (O_2609,N_24450,N_24649);
nor UO_2610 (O_2610,N_24930,N_24709);
and UO_2611 (O_2611,N_24805,N_24613);
nor UO_2612 (O_2612,N_24081,N_24905);
xor UO_2613 (O_2613,N_24150,N_24761);
or UO_2614 (O_2614,N_24334,N_24737);
and UO_2615 (O_2615,N_24000,N_24358);
or UO_2616 (O_2616,N_24861,N_24472);
nor UO_2617 (O_2617,N_24652,N_24915);
nor UO_2618 (O_2618,N_24833,N_24207);
and UO_2619 (O_2619,N_24658,N_24752);
nand UO_2620 (O_2620,N_24981,N_24755);
xnor UO_2621 (O_2621,N_24282,N_24723);
xor UO_2622 (O_2622,N_24343,N_24533);
xor UO_2623 (O_2623,N_24319,N_24050);
or UO_2624 (O_2624,N_24778,N_24104);
xor UO_2625 (O_2625,N_24018,N_24153);
nor UO_2626 (O_2626,N_24243,N_24284);
nand UO_2627 (O_2627,N_24269,N_24970);
nand UO_2628 (O_2628,N_24634,N_24357);
nor UO_2629 (O_2629,N_24695,N_24724);
and UO_2630 (O_2630,N_24844,N_24467);
xnor UO_2631 (O_2631,N_24479,N_24730);
and UO_2632 (O_2632,N_24687,N_24784);
or UO_2633 (O_2633,N_24168,N_24704);
xor UO_2634 (O_2634,N_24073,N_24711);
or UO_2635 (O_2635,N_24138,N_24426);
and UO_2636 (O_2636,N_24220,N_24402);
nor UO_2637 (O_2637,N_24605,N_24584);
or UO_2638 (O_2638,N_24320,N_24090);
or UO_2639 (O_2639,N_24501,N_24859);
and UO_2640 (O_2640,N_24117,N_24462);
nand UO_2641 (O_2641,N_24648,N_24572);
or UO_2642 (O_2642,N_24028,N_24362);
or UO_2643 (O_2643,N_24913,N_24101);
xor UO_2644 (O_2644,N_24931,N_24080);
or UO_2645 (O_2645,N_24757,N_24770);
nor UO_2646 (O_2646,N_24302,N_24460);
or UO_2647 (O_2647,N_24414,N_24302);
nand UO_2648 (O_2648,N_24542,N_24102);
nand UO_2649 (O_2649,N_24635,N_24181);
nor UO_2650 (O_2650,N_24767,N_24165);
nor UO_2651 (O_2651,N_24272,N_24550);
nor UO_2652 (O_2652,N_24316,N_24183);
xor UO_2653 (O_2653,N_24938,N_24968);
nor UO_2654 (O_2654,N_24857,N_24000);
nor UO_2655 (O_2655,N_24471,N_24175);
and UO_2656 (O_2656,N_24581,N_24069);
or UO_2657 (O_2657,N_24243,N_24040);
or UO_2658 (O_2658,N_24348,N_24695);
and UO_2659 (O_2659,N_24489,N_24558);
and UO_2660 (O_2660,N_24818,N_24570);
or UO_2661 (O_2661,N_24613,N_24217);
and UO_2662 (O_2662,N_24567,N_24379);
and UO_2663 (O_2663,N_24931,N_24606);
nand UO_2664 (O_2664,N_24873,N_24934);
nand UO_2665 (O_2665,N_24644,N_24556);
xor UO_2666 (O_2666,N_24352,N_24280);
xor UO_2667 (O_2667,N_24396,N_24476);
nand UO_2668 (O_2668,N_24488,N_24565);
or UO_2669 (O_2669,N_24208,N_24925);
and UO_2670 (O_2670,N_24483,N_24673);
nor UO_2671 (O_2671,N_24938,N_24214);
nand UO_2672 (O_2672,N_24829,N_24408);
nor UO_2673 (O_2673,N_24013,N_24927);
xor UO_2674 (O_2674,N_24578,N_24189);
and UO_2675 (O_2675,N_24365,N_24938);
and UO_2676 (O_2676,N_24469,N_24190);
nor UO_2677 (O_2677,N_24793,N_24410);
nand UO_2678 (O_2678,N_24642,N_24721);
xor UO_2679 (O_2679,N_24535,N_24346);
or UO_2680 (O_2680,N_24044,N_24415);
xor UO_2681 (O_2681,N_24319,N_24070);
nand UO_2682 (O_2682,N_24245,N_24631);
and UO_2683 (O_2683,N_24894,N_24583);
nor UO_2684 (O_2684,N_24887,N_24270);
nand UO_2685 (O_2685,N_24031,N_24174);
nor UO_2686 (O_2686,N_24549,N_24364);
xor UO_2687 (O_2687,N_24292,N_24825);
nor UO_2688 (O_2688,N_24306,N_24998);
nor UO_2689 (O_2689,N_24527,N_24289);
and UO_2690 (O_2690,N_24253,N_24950);
xor UO_2691 (O_2691,N_24033,N_24447);
nand UO_2692 (O_2692,N_24562,N_24145);
nand UO_2693 (O_2693,N_24812,N_24377);
nor UO_2694 (O_2694,N_24833,N_24724);
nand UO_2695 (O_2695,N_24386,N_24515);
or UO_2696 (O_2696,N_24859,N_24299);
and UO_2697 (O_2697,N_24941,N_24402);
xnor UO_2698 (O_2698,N_24150,N_24094);
and UO_2699 (O_2699,N_24888,N_24388);
xor UO_2700 (O_2700,N_24709,N_24425);
or UO_2701 (O_2701,N_24031,N_24944);
nor UO_2702 (O_2702,N_24988,N_24690);
nor UO_2703 (O_2703,N_24176,N_24289);
nor UO_2704 (O_2704,N_24958,N_24194);
xor UO_2705 (O_2705,N_24399,N_24804);
or UO_2706 (O_2706,N_24579,N_24960);
nor UO_2707 (O_2707,N_24598,N_24479);
or UO_2708 (O_2708,N_24823,N_24390);
xnor UO_2709 (O_2709,N_24331,N_24648);
or UO_2710 (O_2710,N_24461,N_24269);
and UO_2711 (O_2711,N_24923,N_24409);
nor UO_2712 (O_2712,N_24431,N_24037);
nor UO_2713 (O_2713,N_24655,N_24882);
nand UO_2714 (O_2714,N_24054,N_24028);
or UO_2715 (O_2715,N_24727,N_24485);
nor UO_2716 (O_2716,N_24890,N_24264);
nand UO_2717 (O_2717,N_24232,N_24992);
or UO_2718 (O_2718,N_24608,N_24042);
and UO_2719 (O_2719,N_24642,N_24583);
nor UO_2720 (O_2720,N_24011,N_24254);
nand UO_2721 (O_2721,N_24614,N_24791);
xnor UO_2722 (O_2722,N_24131,N_24933);
nand UO_2723 (O_2723,N_24620,N_24622);
xnor UO_2724 (O_2724,N_24044,N_24763);
nand UO_2725 (O_2725,N_24059,N_24365);
or UO_2726 (O_2726,N_24628,N_24393);
nand UO_2727 (O_2727,N_24535,N_24268);
or UO_2728 (O_2728,N_24034,N_24916);
and UO_2729 (O_2729,N_24911,N_24667);
xor UO_2730 (O_2730,N_24254,N_24438);
or UO_2731 (O_2731,N_24518,N_24145);
nor UO_2732 (O_2732,N_24390,N_24924);
or UO_2733 (O_2733,N_24392,N_24657);
nand UO_2734 (O_2734,N_24845,N_24084);
nand UO_2735 (O_2735,N_24079,N_24393);
xor UO_2736 (O_2736,N_24851,N_24373);
xnor UO_2737 (O_2737,N_24245,N_24925);
or UO_2738 (O_2738,N_24266,N_24056);
nand UO_2739 (O_2739,N_24389,N_24748);
xnor UO_2740 (O_2740,N_24216,N_24952);
nand UO_2741 (O_2741,N_24346,N_24722);
nand UO_2742 (O_2742,N_24993,N_24879);
or UO_2743 (O_2743,N_24742,N_24082);
and UO_2744 (O_2744,N_24587,N_24307);
nand UO_2745 (O_2745,N_24194,N_24973);
nand UO_2746 (O_2746,N_24181,N_24191);
or UO_2747 (O_2747,N_24383,N_24397);
xor UO_2748 (O_2748,N_24789,N_24912);
or UO_2749 (O_2749,N_24219,N_24263);
and UO_2750 (O_2750,N_24414,N_24125);
xor UO_2751 (O_2751,N_24468,N_24838);
or UO_2752 (O_2752,N_24106,N_24438);
xor UO_2753 (O_2753,N_24146,N_24935);
and UO_2754 (O_2754,N_24986,N_24950);
xor UO_2755 (O_2755,N_24153,N_24081);
or UO_2756 (O_2756,N_24097,N_24415);
xnor UO_2757 (O_2757,N_24272,N_24678);
or UO_2758 (O_2758,N_24916,N_24760);
xor UO_2759 (O_2759,N_24958,N_24019);
and UO_2760 (O_2760,N_24947,N_24632);
and UO_2761 (O_2761,N_24780,N_24766);
nand UO_2762 (O_2762,N_24476,N_24060);
or UO_2763 (O_2763,N_24931,N_24369);
nor UO_2764 (O_2764,N_24642,N_24424);
xnor UO_2765 (O_2765,N_24677,N_24144);
nand UO_2766 (O_2766,N_24542,N_24774);
nand UO_2767 (O_2767,N_24490,N_24432);
xor UO_2768 (O_2768,N_24922,N_24474);
nand UO_2769 (O_2769,N_24291,N_24483);
xor UO_2770 (O_2770,N_24583,N_24833);
xnor UO_2771 (O_2771,N_24578,N_24337);
nand UO_2772 (O_2772,N_24148,N_24912);
or UO_2773 (O_2773,N_24054,N_24300);
or UO_2774 (O_2774,N_24253,N_24734);
nand UO_2775 (O_2775,N_24252,N_24798);
or UO_2776 (O_2776,N_24649,N_24420);
nor UO_2777 (O_2777,N_24895,N_24469);
or UO_2778 (O_2778,N_24761,N_24663);
or UO_2779 (O_2779,N_24010,N_24728);
xnor UO_2780 (O_2780,N_24208,N_24838);
nor UO_2781 (O_2781,N_24596,N_24010);
or UO_2782 (O_2782,N_24421,N_24334);
xnor UO_2783 (O_2783,N_24107,N_24098);
or UO_2784 (O_2784,N_24079,N_24090);
nand UO_2785 (O_2785,N_24509,N_24581);
or UO_2786 (O_2786,N_24962,N_24651);
nor UO_2787 (O_2787,N_24344,N_24767);
xnor UO_2788 (O_2788,N_24070,N_24063);
or UO_2789 (O_2789,N_24358,N_24324);
and UO_2790 (O_2790,N_24682,N_24373);
nor UO_2791 (O_2791,N_24264,N_24284);
and UO_2792 (O_2792,N_24503,N_24962);
nor UO_2793 (O_2793,N_24447,N_24927);
and UO_2794 (O_2794,N_24906,N_24617);
xnor UO_2795 (O_2795,N_24512,N_24093);
nor UO_2796 (O_2796,N_24109,N_24610);
xor UO_2797 (O_2797,N_24332,N_24307);
or UO_2798 (O_2798,N_24821,N_24858);
or UO_2799 (O_2799,N_24988,N_24303);
or UO_2800 (O_2800,N_24686,N_24623);
xor UO_2801 (O_2801,N_24208,N_24730);
xor UO_2802 (O_2802,N_24982,N_24809);
nand UO_2803 (O_2803,N_24437,N_24601);
xor UO_2804 (O_2804,N_24183,N_24887);
or UO_2805 (O_2805,N_24961,N_24125);
nand UO_2806 (O_2806,N_24043,N_24897);
or UO_2807 (O_2807,N_24728,N_24065);
or UO_2808 (O_2808,N_24873,N_24243);
nand UO_2809 (O_2809,N_24529,N_24833);
nand UO_2810 (O_2810,N_24229,N_24416);
nor UO_2811 (O_2811,N_24098,N_24783);
and UO_2812 (O_2812,N_24571,N_24871);
xor UO_2813 (O_2813,N_24159,N_24955);
and UO_2814 (O_2814,N_24556,N_24858);
nand UO_2815 (O_2815,N_24127,N_24403);
nor UO_2816 (O_2816,N_24479,N_24740);
or UO_2817 (O_2817,N_24799,N_24163);
and UO_2818 (O_2818,N_24456,N_24971);
xnor UO_2819 (O_2819,N_24493,N_24743);
or UO_2820 (O_2820,N_24378,N_24976);
and UO_2821 (O_2821,N_24853,N_24585);
nor UO_2822 (O_2822,N_24921,N_24874);
or UO_2823 (O_2823,N_24704,N_24745);
and UO_2824 (O_2824,N_24178,N_24062);
xnor UO_2825 (O_2825,N_24354,N_24338);
or UO_2826 (O_2826,N_24094,N_24462);
and UO_2827 (O_2827,N_24547,N_24238);
xor UO_2828 (O_2828,N_24131,N_24384);
or UO_2829 (O_2829,N_24739,N_24809);
xor UO_2830 (O_2830,N_24647,N_24061);
nor UO_2831 (O_2831,N_24240,N_24693);
or UO_2832 (O_2832,N_24763,N_24375);
nor UO_2833 (O_2833,N_24113,N_24461);
and UO_2834 (O_2834,N_24841,N_24002);
and UO_2835 (O_2835,N_24602,N_24270);
nor UO_2836 (O_2836,N_24035,N_24393);
xnor UO_2837 (O_2837,N_24452,N_24191);
nand UO_2838 (O_2838,N_24313,N_24327);
nand UO_2839 (O_2839,N_24382,N_24053);
nand UO_2840 (O_2840,N_24039,N_24961);
nand UO_2841 (O_2841,N_24020,N_24220);
nand UO_2842 (O_2842,N_24897,N_24073);
nor UO_2843 (O_2843,N_24748,N_24878);
xor UO_2844 (O_2844,N_24547,N_24146);
xnor UO_2845 (O_2845,N_24609,N_24667);
and UO_2846 (O_2846,N_24481,N_24537);
nand UO_2847 (O_2847,N_24661,N_24510);
and UO_2848 (O_2848,N_24059,N_24373);
xnor UO_2849 (O_2849,N_24861,N_24828);
xor UO_2850 (O_2850,N_24592,N_24309);
nand UO_2851 (O_2851,N_24251,N_24435);
xnor UO_2852 (O_2852,N_24354,N_24930);
or UO_2853 (O_2853,N_24978,N_24182);
and UO_2854 (O_2854,N_24263,N_24218);
nand UO_2855 (O_2855,N_24836,N_24716);
nor UO_2856 (O_2856,N_24470,N_24245);
nand UO_2857 (O_2857,N_24043,N_24026);
nand UO_2858 (O_2858,N_24767,N_24826);
and UO_2859 (O_2859,N_24786,N_24763);
or UO_2860 (O_2860,N_24949,N_24204);
xor UO_2861 (O_2861,N_24879,N_24494);
nor UO_2862 (O_2862,N_24010,N_24449);
nand UO_2863 (O_2863,N_24811,N_24622);
nand UO_2864 (O_2864,N_24787,N_24433);
or UO_2865 (O_2865,N_24258,N_24415);
nand UO_2866 (O_2866,N_24882,N_24572);
nand UO_2867 (O_2867,N_24609,N_24548);
nand UO_2868 (O_2868,N_24378,N_24022);
xnor UO_2869 (O_2869,N_24888,N_24874);
nand UO_2870 (O_2870,N_24461,N_24188);
xnor UO_2871 (O_2871,N_24942,N_24169);
and UO_2872 (O_2872,N_24691,N_24930);
nand UO_2873 (O_2873,N_24230,N_24083);
and UO_2874 (O_2874,N_24308,N_24110);
nor UO_2875 (O_2875,N_24231,N_24842);
nor UO_2876 (O_2876,N_24599,N_24034);
nor UO_2877 (O_2877,N_24753,N_24524);
or UO_2878 (O_2878,N_24382,N_24695);
or UO_2879 (O_2879,N_24712,N_24377);
nand UO_2880 (O_2880,N_24502,N_24547);
xnor UO_2881 (O_2881,N_24257,N_24811);
or UO_2882 (O_2882,N_24524,N_24776);
or UO_2883 (O_2883,N_24310,N_24482);
nand UO_2884 (O_2884,N_24201,N_24200);
nor UO_2885 (O_2885,N_24632,N_24936);
or UO_2886 (O_2886,N_24737,N_24940);
xor UO_2887 (O_2887,N_24857,N_24883);
nand UO_2888 (O_2888,N_24883,N_24349);
nor UO_2889 (O_2889,N_24550,N_24834);
nand UO_2890 (O_2890,N_24028,N_24666);
nor UO_2891 (O_2891,N_24294,N_24287);
or UO_2892 (O_2892,N_24828,N_24254);
or UO_2893 (O_2893,N_24762,N_24475);
nand UO_2894 (O_2894,N_24786,N_24356);
xor UO_2895 (O_2895,N_24933,N_24309);
xor UO_2896 (O_2896,N_24750,N_24625);
xnor UO_2897 (O_2897,N_24454,N_24864);
xor UO_2898 (O_2898,N_24449,N_24375);
and UO_2899 (O_2899,N_24044,N_24796);
and UO_2900 (O_2900,N_24752,N_24448);
or UO_2901 (O_2901,N_24392,N_24140);
nand UO_2902 (O_2902,N_24236,N_24116);
or UO_2903 (O_2903,N_24487,N_24753);
or UO_2904 (O_2904,N_24050,N_24781);
nor UO_2905 (O_2905,N_24864,N_24912);
nor UO_2906 (O_2906,N_24609,N_24242);
and UO_2907 (O_2907,N_24502,N_24890);
nor UO_2908 (O_2908,N_24321,N_24351);
and UO_2909 (O_2909,N_24126,N_24007);
and UO_2910 (O_2910,N_24105,N_24039);
nand UO_2911 (O_2911,N_24958,N_24653);
nor UO_2912 (O_2912,N_24362,N_24540);
xnor UO_2913 (O_2913,N_24769,N_24419);
or UO_2914 (O_2914,N_24919,N_24160);
xor UO_2915 (O_2915,N_24800,N_24373);
nand UO_2916 (O_2916,N_24071,N_24830);
nor UO_2917 (O_2917,N_24950,N_24205);
and UO_2918 (O_2918,N_24352,N_24495);
nor UO_2919 (O_2919,N_24688,N_24060);
nor UO_2920 (O_2920,N_24697,N_24830);
xor UO_2921 (O_2921,N_24321,N_24449);
nand UO_2922 (O_2922,N_24431,N_24829);
nor UO_2923 (O_2923,N_24310,N_24662);
or UO_2924 (O_2924,N_24624,N_24766);
or UO_2925 (O_2925,N_24914,N_24657);
and UO_2926 (O_2926,N_24110,N_24080);
nor UO_2927 (O_2927,N_24088,N_24011);
and UO_2928 (O_2928,N_24573,N_24044);
or UO_2929 (O_2929,N_24292,N_24224);
nor UO_2930 (O_2930,N_24374,N_24903);
nand UO_2931 (O_2931,N_24867,N_24233);
nor UO_2932 (O_2932,N_24697,N_24671);
nand UO_2933 (O_2933,N_24673,N_24493);
and UO_2934 (O_2934,N_24972,N_24165);
or UO_2935 (O_2935,N_24737,N_24098);
xnor UO_2936 (O_2936,N_24592,N_24329);
nor UO_2937 (O_2937,N_24923,N_24800);
and UO_2938 (O_2938,N_24761,N_24109);
nor UO_2939 (O_2939,N_24149,N_24752);
and UO_2940 (O_2940,N_24504,N_24973);
xor UO_2941 (O_2941,N_24191,N_24944);
and UO_2942 (O_2942,N_24275,N_24807);
nand UO_2943 (O_2943,N_24264,N_24942);
and UO_2944 (O_2944,N_24751,N_24930);
nor UO_2945 (O_2945,N_24398,N_24926);
xnor UO_2946 (O_2946,N_24440,N_24828);
and UO_2947 (O_2947,N_24392,N_24262);
nor UO_2948 (O_2948,N_24824,N_24949);
xnor UO_2949 (O_2949,N_24664,N_24683);
xor UO_2950 (O_2950,N_24940,N_24045);
or UO_2951 (O_2951,N_24429,N_24894);
or UO_2952 (O_2952,N_24771,N_24096);
nor UO_2953 (O_2953,N_24274,N_24008);
or UO_2954 (O_2954,N_24141,N_24568);
nor UO_2955 (O_2955,N_24362,N_24645);
or UO_2956 (O_2956,N_24837,N_24647);
nor UO_2957 (O_2957,N_24378,N_24926);
xor UO_2958 (O_2958,N_24462,N_24734);
nor UO_2959 (O_2959,N_24998,N_24479);
xor UO_2960 (O_2960,N_24638,N_24831);
nand UO_2961 (O_2961,N_24194,N_24930);
and UO_2962 (O_2962,N_24524,N_24330);
xor UO_2963 (O_2963,N_24603,N_24563);
nand UO_2964 (O_2964,N_24769,N_24223);
and UO_2965 (O_2965,N_24762,N_24668);
nand UO_2966 (O_2966,N_24058,N_24069);
or UO_2967 (O_2967,N_24529,N_24759);
and UO_2968 (O_2968,N_24797,N_24302);
nor UO_2969 (O_2969,N_24183,N_24348);
nor UO_2970 (O_2970,N_24772,N_24305);
nand UO_2971 (O_2971,N_24940,N_24648);
nand UO_2972 (O_2972,N_24454,N_24598);
or UO_2973 (O_2973,N_24604,N_24612);
nor UO_2974 (O_2974,N_24845,N_24840);
xnor UO_2975 (O_2975,N_24690,N_24508);
xor UO_2976 (O_2976,N_24047,N_24815);
xor UO_2977 (O_2977,N_24560,N_24609);
xor UO_2978 (O_2978,N_24668,N_24254);
and UO_2979 (O_2979,N_24714,N_24191);
xnor UO_2980 (O_2980,N_24473,N_24760);
and UO_2981 (O_2981,N_24053,N_24290);
or UO_2982 (O_2982,N_24070,N_24602);
nand UO_2983 (O_2983,N_24499,N_24011);
xor UO_2984 (O_2984,N_24507,N_24737);
and UO_2985 (O_2985,N_24822,N_24268);
or UO_2986 (O_2986,N_24202,N_24148);
and UO_2987 (O_2987,N_24740,N_24972);
xor UO_2988 (O_2988,N_24478,N_24714);
xnor UO_2989 (O_2989,N_24491,N_24640);
or UO_2990 (O_2990,N_24626,N_24321);
nor UO_2991 (O_2991,N_24753,N_24228);
or UO_2992 (O_2992,N_24779,N_24079);
nand UO_2993 (O_2993,N_24934,N_24498);
nand UO_2994 (O_2994,N_24440,N_24360);
nand UO_2995 (O_2995,N_24219,N_24722);
nand UO_2996 (O_2996,N_24235,N_24421);
xnor UO_2997 (O_2997,N_24328,N_24621);
or UO_2998 (O_2998,N_24674,N_24284);
nor UO_2999 (O_2999,N_24471,N_24077);
endmodule