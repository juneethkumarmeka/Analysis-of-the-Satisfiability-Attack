module basic_2500_25000_3000_4_levels_5xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18757,N_18758,N_18759,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18925,N_18926,N_18927,N_18928,N_18929,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18945,N_18946,N_18947,N_18948,N_18949,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19187,N_19188,N_19189,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19456,N_19457,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19628,N_19629,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19651,N_19652,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19669,N_19670,N_19671,N_19672,N_19673,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19731,N_19732,N_19733,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19745,N_19746,N_19747,N_19748,N_19749,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20003,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20021,N_20022,N_20023,N_20024,N_20025,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20323,N_20324,N_20325,N_20326,N_20327,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20594,N_20595,N_20596,N_20599,N_20600,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20745,N_20746,N_20747,N_20748,N_20750,N_20751,N_20752,N_20753,N_20755,N_20756,N_20757,N_20758,N_20759,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20853,N_20854,N_20855,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20946,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21122,N_21123,N_21124,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21157,N_21158,N_21159,N_21160,N_21161,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21378,N_21379,N_21380,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21739,N_21740,N_21741,N_21742,N_21743,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21972,N_21973,N_21974,N_21975,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22119,N_22120,N_22121,N_22122,N_22124,N_22125,N_22126,N_22127,N_22128,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22227,N_22228,N_22229,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22596,N_22597,N_22598,N_22599,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23089,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23115,N_23116,N_23117,N_23118,N_23119,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23226,N_23227,N_23228,N_23229,N_23231,N_23232,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23297,N_23299,N_23300,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23334,N_23335,N_23337,N_23338,N_23339,N_23340,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23352,N_23353,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23675,N_23676,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23991,N_23992,N_23993,N_23994,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24104,N_24105,N_24106,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24225,N_24226,N_24227,N_24228,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24729,N_24730,N_24731,N_24732,N_24733,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24885,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24993,N_24995,N_24996,N_24997,N_24998,N_24999;
nand U0 (N_0,In_289,In_845);
or U1 (N_1,In_306,In_1682);
nor U2 (N_2,In_1164,In_2267);
and U3 (N_3,In_619,In_762);
and U4 (N_4,In_2365,In_2037);
nand U5 (N_5,In_540,In_1013);
nand U6 (N_6,In_2448,In_2409);
and U7 (N_7,In_641,In_1722);
nor U8 (N_8,In_1716,In_668);
or U9 (N_9,In_1436,In_2266);
or U10 (N_10,In_718,In_1049);
nand U11 (N_11,In_2120,In_258);
and U12 (N_12,In_882,In_1751);
nor U13 (N_13,In_1797,In_756);
and U14 (N_14,In_1487,In_935);
and U15 (N_15,In_2455,In_447);
nor U16 (N_16,In_2322,In_1321);
or U17 (N_17,In_623,In_2218);
nor U18 (N_18,In_1654,In_1276);
nand U19 (N_19,In_1069,In_559);
and U20 (N_20,In_596,In_681);
and U21 (N_21,In_1798,In_758);
and U22 (N_22,In_2135,In_989);
or U23 (N_23,In_1620,In_1158);
nor U24 (N_24,In_809,In_1358);
nand U25 (N_25,In_795,In_673);
or U26 (N_26,In_1279,In_1059);
or U27 (N_27,In_1863,In_1005);
nor U28 (N_28,In_235,In_1768);
or U29 (N_29,In_1580,In_2166);
and U30 (N_30,In_2253,In_1033);
nor U31 (N_31,In_671,In_2274);
nor U32 (N_32,In_2466,In_2217);
nor U33 (N_33,In_73,In_1252);
nor U34 (N_34,In_332,In_2432);
and U35 (N_35,In_556,In_2323);
xor U36 (N_36,In_1819,In_483);
and U37 (N_37,In_1366,In_2377);
and U38 (N_38,In_741,In_1198);
or U39 (N_39,In_545,In_1455);
or U40 (N_40,In_320,In_2112);
nand U41 (N_41,In_361,In_807);
xnor U42 (N_42,In_852,In_893);
or U43 (N_43,In_1313,In_755);
and U44 (N_44,In_1216,In_2470);
nand U45 (N_45,In_1893,In_1102);
xor U46 (N_46,In_1979,In_439);
or U47 (N_47,In_2065,In_383);
nor U48 (N_48,In_1532,In_940);
xnor U49 (N_49,In_404,In_2106);
nand U50 (N_50,In_216,In_193);
or U51 (N_51,In_975,In_2092);
nand U52 (N_52,In_1171,In_2304);
nor U53 (N_53,In_660,In_122);
nand U54 (N_54,In_51,In_1361);
xor U55 (N_55,In_244,In_132);
and U56 (N_56,In_1877,In_172);
or U57 (N_57,In_1442,In_1444);
and U58 (N_58,In_1125,In_27);
nor U59 (N_59,In_283,In_2087);
or U60 (N_60,In_980,In_264);
and U61 (N_61,In_1263,In_1464);
and U62 (N_62,In_180,In_1881);
nand U63 (N_63,In_2018,In_1031);
and U64 (N_64,In_2008,In_2183);
nand U65 (N_65,In_1657,In_778);
nand U66 (N_66,In_1937,In_1714);
or U67 (N_67,In_1938,In_1858);
and U68 (N_68,In_1290,In_998);
or U69 (N_69,In_1190,In_1977);
or U70 (N_70,In_1870,In_963);
nand U71 (N_71,In_2070,In_2240);
nor U72 (N_72,In_406,In_611);
and U73 (N_73,In_1367,In_1668);
nor U74 (N_74,In_2172,In_451);
and U75 (N_75,In_1228,In_2096);
xor U76 (N_76,In_2017,In_614);
and U77 (N_77,In_1249,In_1917);
and U78 (N_78,In_2355,In_1450);
nor U79 (N_79,In_1581,In_1909);
or U80 (N_80,In_2440,In_2422);
or U81 (N_81,In_628,In_4);
nand U82 (N_82,In_1619,In_427);
nor U83 (N_83,In_2352,In_2303);
or U84 (N_84,In_584,In_1878);
or U85 (N_85,In_1836,In_1012);
nor U86 (N_86,In_23,In_974);
nor U87 (N_87,In_1422,In_932);
or U88 (N_88,In_835,In_562);
or U89 (N_89,In_663,In_516);
or U90 (N_90,In_651,In_313);
nand U91 (N_91,In_1901,In_2402);
nand U92 (N_92,In_1179,In_1111);
nand U93 (N_93,In_479,In_1117);
nand U94 (N_94,In_1811,In_735);
or U95 (N_95,In_125,In_1478);
and U96 (N_96,In_2149,In_1740);
nor U97 (N_97,In_2156,In_2385);
nand U98 (N_98,In_841,In_914);
nor U99 (N_99,In_1333,In_488);
nor U100 (N_100,In_139,In_515);
and U101 (N_101,In_496,In_2239);
nand U102 (N_102,In_2012,In_714);
and U103 (N_103,In_2427,In_1051);
or U104 (N_104,In_275,In_270);
and U105 (N_105,In_2401,In_1617);
and U106 (N_106,In_357,In_1986);
xnor U107 (N_107,In_1884,In_335);
nor U108 (N_108,In_2250,In_228);
or U109 (N_109,In_2153,In_1411);
nor U110 (N_110,In_1339,In_1502);
or U111 (N_111,In_1500,In_1860);
or U112 (N_112,In_590,In_1952);
nor U113 (N_113,In_195,In_636);
nor U114 (N_114,In_1220,In_911);
and U115 (N_115,In_1058,In_2439);
nand U116 (N_116,In_1443,In_822);
or U117 (N_117,In_676,In_97);
and U118 (N_118,In_1734,In_950);
and U119 (N_119,In_71,In_1757);
nand U120 (N_120,In_2373,In_1570);
xnor U121 (N_121,In_1035,In_2185);
nor U122 (N_122,In_1221,In_1916);
xor U123 (N_123,In_2220,In_1769);
or U124 (N_124,In_269,In_1014);
nor U125 (N_125,In_690,In_1418);
or U126 (N_126,In_2374,In_661);
nand U127 (N_127,In_2223,In_2400);
or U128 (N_128,In_743,In_1155);
xnor U129 (N_129,In_2316,In_494);
nor U130 (N_130,In_246,In_567);
nand U131 (N_131,In_2246,In_492);
nand U132 (N_132,In_2275,In_1868);
or U133 (N_133,In_907,In_50);
or U134 (N_134,In_1785,In_184);
nor U135 (N_135,In_1429,In_182);
and U136 (N_136,In_1146,In_942);
nor U137 (N_137,In_37,In_1783);
xor U138 (N_138,In_521,In_2320);
nor U139 (N_139,In_544,In_2415);
nor U140 (N_140,In_322,In_141);
nor U141 (N_141,In_2372,In_1109);
and U142 (N_142,In_1183,In_2158);
or U143 (N_143,In_9,In_2434);
or U144 (N_144,In_564,In_1618);
nor U145 (N_145,In_2124,In_850);
xnor U146 (N_146,In_644,In_732);
or U147 (N_147,In_236,In_1187);
or U148 (N_148,In_374,In_1037);
nand U149 (N_149,In_2099,In_32);
and U150 (N_150,In_996,In_2359);
and U151 (N_151,In_1498,In_194);
and U152 (N_152,In_314,In_466);
nor U153 (N_153,In_1616,In_210);
or U154 (N_154,In_1627,In_185);
nor U155 (N_155,In_780,In_1650);
or U156 (N_156,In_2035,In_468);
nand U157 (N_157,In_1270,In_298);
nand U158 (N_158,In_2252,In_520);
and U159 (N_159,In_18,In_1019);
xnor U160 (N_160,In_1648,In_1525);
nor U161 (N_161,In_241,In_1862);
and U162 (N_162,In_2358,In_1544);
nor U163 (N_163,In_801,In_819);
xor U164 (N_164,In_2088,In_868);
or U165 (N_165,In_1981,In_1697);
or U166 (N_166,In_1745,In_1001);
and U167 (N_167,In_409,In_165);
nor U168 (N_168,In_666,In_2283);
or U169 (N_169,In_1317,In_2305);
nand U170 (N_170,In_2085,In_616);
nor U171 (N_171,In_1854,In_1805);
nand U172 (N_172,In_371,In_529);
nand U173 (N_173,In_1099,In_465);
or U174 (N_174,In_804,In_2114);
and U175 (N_175,In_1431,In_337);
nand U176 (N_176,In_1390,In_179);
or U177 (N_177,In_1666,In_1482);
nor U178 (N_178,In_1314,In_818);
or U179 (N_179,In_1588,In_338);
and U180 (N_180,In_1073,In_1203);
or U181 (N_181,In_2280,In_1519);
xor U182 (N_182,In_2190,In_2326);
xor U183 (N_183,In_1994,In_1437);
nand U184 (N_184,In_1652,In_1503);
and U185 (N_185,In_426,In_507);
nor U186 (N_186,In_1451,In_978);
and U187 (N_187,In_12,In_2497);
and U188 (N_188,In_171,In_2433);
nor U189 (N_189,In_2136,In_1644);
and U190 (N_190,In_1119,In_669);
and U191 (N_191,In_2339,In_21);
or U192 (N_192,In_1052,In_87);
and U193 (N_193,In_2174,In_1859);
nand U194 (N_194,In_1306,In_2202);
nand U195 (N_195,In_976,In_765);
or U196 (N_196,In_1771,In_1307);
nor U197 (N_197,In_435,In_713);
nand U198 (N_198,In_1828,In_2368);
and U199 (N_199,In_1593,In_2111);
nor U200 (N_200,In_2152,In_464);
or U201 (N_201,In_684,In_467);
xor U202 (N_202,In_1452,In_1839);
or U203 (N_203,In_1621,In_2403);
nand U204 (N_204,In_1910,In_206);
xor U205 (N_205,In_1299,In_829);
nor U206 (N_206,In_2068,In_1707);
and U207 (N_207,In_34,In_568);
and U208 (N_208,In_95,In_2098);
nor U209 (N_209,In_2023,In_1172);
nor U210 (N_210,In_2009,In_2144);
nor U211 (N_211,In_1008,In_393);
nand U212 (N_212,In_149,In_315);
and U213 (N_213,In_1739,In_1492);
nor U214 (N_214,In_821,In_933);
nor U215 (N_215,In_1374,In_1825);
nand U216 (N_216,In_1826,In_929);
or U217 (N_217,In_711,In_473);
nor U218 (N_218,In_1610,In_777);
and U219 (N_219,In_1118,In_2295);
nor U220 (N_220,In_2421,In_1044);
and U221 (N_221,In_757,In_1043);
or U222 (N_222,In_1371,In_1273);
nand U223 (N_223,In_1485,In_1882);
or U224 (N_224,In_284,In_2109);
and U225 (N_225,In_1818,In_891);
or U226 (N_226,In_1505,In_1412);
nor U227 (N_227,In_470,In_2471);
and U228 (N_228,In_1419,In_767);
xnor U229 (N_229,In_2244,In_98);
nand U230 (N_230,In_2454,In_823);
nor U231 (N_231,In_1034,In_952);
nand U232 (N_232,In_2082,In_1346);
nor U233 (N_233,In_2315,In_1733);
nor U234 (N_234,In_2147,In_527);
and U235 (N_235,In_245,In_218);
nor U236 (N_236,In_334,In_700);
and U237 (N_237,In_988,In_396);
xor U238 (N_238,In_1633,In_69);
and U239 (N_239,In_61,In_138);
and U240 (N_240,In_1807,In_2207);
nor U241 (N_241,In_991,In_1082);
nand U242 (N_242,In_670,In_887);
and U243 (N_243,In_930,In_1655);
and U244 (N_244,In_232,In_174);
and U245 (N_245,In_347,In_1914);
and U246 (N_246,In_104,In_1844);
nor U247 (N_247,In_1139,In_2163);
or U248 (N_248,In_1078,In_760);
nor U249 (N_249,In_1085,In_2066);
nor U250 (N_250,In_1792,In_1876);
and U251 (N_251,In_817,In_1106);
nor U252 (N_252,In_548,In_941);
nand U253 (N_253,In_639,In_1754);
xnor U254 (N_254,In_2069,In_1165);
xnor U255 (N_255,In_2363,In_864);
and U256 (N_256,In_2118,In_2298);
or U257 (N_257,In_52,In_220);
and U258 (N_258,In_214,In_2405);
and U259 (N_259,In_2016,In_10);
and U260 (N_260,In_539,In_1223);
or U261 (N_261,In_949,In_634);
nor U262 (N_262,In_2256,In_883);
xor U263 (N_263,In_341,In_311);
and U264 (N_264,In_1706,In_1486);
nor U265 (N_265,In_922,In_606);
nand U266 (N_266,In_746,In_2268);
nor U267 (N_267,In_100,In_1369);
and U268 (N_268,In_415,In_405);
or U269 (N_269,In_505,In_1592);
or U270 (N_270,In_745,In_115);
and U271 (N_271,In_761,In_1202);
nand U272 (N_272,In_1709,In_2321);
or U273 (N_273,In_814,In_1556);
nor U274 (N_274,In_1316,In_412);
and U275 (N_275,In_1022,In_1352);
and U276 (N_276,In_2319,In_792);
nand U277 (N_277,In_1239,In_1027);
nor U278 (N_278,In_2347,In_105);
or U279 (N_279,In_1968,In_1778);
xnor U280 (N_280,In_1423,In_2129);
nand U281 (N_281,In_1267,In_1456);
and U282 (N_282,In_782,In_1721);
nand U283 (N_283,In_798,In_1543);
nor U284 (N_284,In_1238,In_947);
or U285 (N_285,In_1311,In_688);
nand U286 (N_286,In_2429,In_805);
nand U287 (N_287,In_1587,In_323);
xnor U288 (N_288,In_1289,In_1891);
nand U289 (N_289,In_1607,In_885);
nand U290 (N_290,In_912,In_1446);
and U291 (N_291,In_2264,In_1445);
and U292 (N_292,In_1148,In_1218);
or U293 (N_293,In_2182,In_740);
xnor U294 (N_294,In_1736,In_292);
nand U295 (N_295,In_997,In_1808);
or U296 (N_296,In_1056,In_1003);
xor U297 (N_297,In_1935,In_1430);
and U298 (N_298,In_1925,In_155);
and U299 (N_299,In_2067,In_1161);
nand U300 (N_300,In_1386,In_2254);
and U301 (N_301,In_1204,In_2344);
nor U302 (N_302,In_709,In_1883);
nor U303 (N_303,In_2494,In_469);
nand U304 (N_304,In_2450,In_1388);
and U305 (N_305,In_119,In_2044);
nor U306 (N_306,In_1294,In_1920);
nand U307 (N_307,In_1932,In_1300);
and U308 (N_308,In_497,In_2);
xnor U309 (N_309,In_372,In_157);
nor U310 (N_310,In_1775,In_249);
nand U311 (N_311,In_250,In_943);
nor U312 (N_312,In_2195,In_793);
or U313 (N_313,In_2312,In_1061);
nor U314 (N_314,In_2447,In_1115);
or U315 (N_315,In_2128,In_2036);
and U316 (N_316,In_2054,In_2086);
or U317 (N_317,In_580,In_2265);
nand U318 (N_318,In_2030,In_1998);
or U319 (N_319,In_839,In_1961);
nand U320 (N_320,In_621,In_797);
nor U321 (N_321,In_1460,In_589);
nor U322 (N_322,In_13,In_2407);
nand U323 (N_323,In_1271,In_112);
or U324 (N_324,In_2230,In_2313);
nor U325 (N_325,In_1945,In_838);
and U326 (N_326,In_2222,In_475);
or U327 (N_327,In_2213,In_751);
or U328 (N_328,In_788,In_2132);
and U329 (N_329,In_1405,In_2366);
or U330 (N_330,In_860,In_1213);
nand U331 (N_331,In_428,In_1888);
xnor U332 (N_332,In_151,In_456);
nand U333 (N_333,In_188,In_201);
nand U334 (N_334,In_1856,In_1199);
and U335 (N_335,In_1050,In_1800);
nor U336 (N_336,In_1269,In_11);
or U337 (N_337,In_1997,In_909);
or U338 (N_338,In_575,In_2040);
and U339 (N_339,In_1508,In_2333);
and U340 (N_340,In_2110,In_1425);
xnor U341 (N_341,In_847,In_1912);
xor U342 (N_342,In_123,In_1257);
or U343 (N_343,In_2301,In_2042);
or U344 (N_344,In_1334,In_1924);
and U345 (N_345,In_1701,In_1594);
or U346 (N_346,In_2199,In_2367);
nor U347 (N_347,In_855,In_2104);
nand U348 (N_348,In_2210,In_1351);
nor U349 (N_349,In_2105,In_1972);
and U350 (N_350,In_395,In_1934);
nor U351 (N_351,In_716,In_962);
nand U352 (N_352,In_438,In_423);
nand U353 (N_353,In_96,In_1071);
or U354 (N_354,In_1435,In_1195);
nand U355 (N_355,In_1108,In_2272);
nor U356 (N_356,In_225,In_2184);
nor U357 (N_357,In_1156,In_2089);
and U358 (N_358,In_972,In_1853);
xor U359 (N_359,In_14,In_1170);
and U360 (N_360,In_968,In_2376);
nand U361 (N_361,In_1895,In_1140);
xnor U362 (N_362,In_977,In_1393);
xnor U363 (N_363,In_44,In_1735);
and U364 (N_364,In_1340,In_1803);
nor U365 (N_365,In_698,In_531);
or U366 (N_366,In_1599,In_1584);
and U367 (N_367,In_1207,In_2351);
nor U368 (N_368,In_1169,In_2291);
xnor U369 (N_369,In_2318,In_2261);
or U370 (N_370,In_1297,In_422);
and U371 (N_371,In_2251,In_1941);
and U372 (N_372,In_647,In_296);
or U373 (N_373,In_89,In_499);
nand U374 (N_374,In_221,In_461);
or U375 (N_375,In_1522,In_1625);
and U376 (N_376,In_295,In_1950);
or U377 (N_377,In_421,In_1407);
or U378 (N_378,In_2311,In_1766);
nor U379 (N_379,In_2079,In_1890);
and U380 (N_380,In_1394,In_33);
or U381 (N_381,In_1177,In_512);
and U382 (N_382,In_344,In_135);
nor U383 (N_383,In_551,In_2201);
nand U384 (N_384,In_2287,In_731);
nand U385 (N_385,In_457,In_896);
xnor U386 (N_386,In_205,In_1087);
nor U387 (N_387,In_2140,In_1399);
nand U388 (N_388,In_2125,In_1293);
or U389 (N_389,In_152,In_1298);
and U390 (N_390,In_603,In_2233);
or U391 (N_391,In_981,In_1385);
and U392 (N_392,In_1929,In_134);
nand U393 (N_393,In_625,In_2308);
and U394 (N_394,In_2064,In_1142);
nand U395 (N_395,In_74,In_317);
xnor U396 (N_396,In_164,In_343);
nor U397 (N_397,In_695,In_1495);
or U398 (N_398,In_2468,In_2168);
and U399 (N_399,In_523,In_1738);
nand U400 (N_400,In_500,In_2293);
nor U401 (N_401,In_1576,In_476);
nor U402 (N_402,In_1821,In_517);
nand U403 (N_403,In_874,In_747);
nand U404 (N_404,In_1123,In_508);
xnor U405 (N_405,In_859,In_114);
nand U406 (N_406,In_1959,In_1467);
nand U407 (N_407,In_160,In_2097);
nor U408 (N_408,In_316,In_2391);
nor U409 (N_409,In_518,In_199);
or U410 (N_410,In_2478,In_774);
nand U411 (N_411,In_42,In_1404);
and U412 (N_412,In_92,In_953);
nand U413 (N_413,In_1931,In_1824);
nor U414 (N_414,In_2130,In_446);
and U415 (N_415,In_2188,In_1662);
or U416 (N_416,In_858,In_646);
nand U417 (N_417,In_583,In_1903);
and U418 (N_418,In_873,In_2215);
or U419 (N_419,In_1953,In_1806);
nor U420 (N_420,In_552,In_1989);
nor U421 (N_421,In_703,In_305);
nor U422 (N_422,In_1240,In_632);
nor U423 (N_423,In_1215,In_1268);
nand U424 (N_424,In_1749,In_2093);
nor U425 (N_425,In_55,In_274);
and U426 (N_426,In_973,In_1296);
and U427 (N_427,In_120,In_667);
and U428 (N_428,In_1359,In_1206);
and U429 (N_429,In_1678,In_710);
nand U430 (N_430,In_1971,In_878);
nor U431 (N_431,In_1936,In_2050);
or U432 (N_432,In_1174,In_1629);
and U433 (N_433,In_2276,In_2360);
nor U434 (N_434,In_1765,In_1710);
nor U435 (N_435,In_1395,In_2020);
xnor U436 (N_436,In_591,In_2404);
and U437 (N_437,In_1869,In_2115);
or U438 (N_438,In_1250,In_57);
nor U439 (N_439,In_387,In_956);
xnor U440 (N_440,In_1905,In_1951);
xor U441 (N_441,In_40,In_1973);
nand U442 (N_442,In_1605,In_204);
nor U443 (N_443,In_587,In_1597);
xor U444 (N_444,In_1499,In_2340);
or U445 (N_445,In_1135,In_2271);
nand U446 (N_446,In_2495,In_2395);
nor U447 (N_447,In_2383,In_2122);
and U448 (N_448,In_1259,In_1520);
xnor U449 (N_449,In_263,In_2248);
and U450 (N_450,In_678,In_2131);
and U451 (N_451,In_1475,In_720);
nand U452 (N_452,In_166,In_1669);
nand U453 (N_453,In_605,In_1076);
or U454 (N_454,In_2255,In_156);
nor U455 (N_455,In_593,In_547);
nand U456 (N_456,In_524,In_585);
xor U457 (N_457,In_2382,In_178);
nand U458 (N_458,In_794,In_365);
xor U459 (N_459,In_1983,In_1046);
nand U460 (N_460,In_870,In_1055);
nand U461 (N_461,In_916,In_1354);
and U462 (N_462,In_687,In_1687);
nor U463 (N_463,In_1846,In_1992);
nor U464 (N_464,In_253,In_1671);
or U465 (N_465,In_1582,In_853);
or U466 (N_466,In_329,In_1763);
nand U467 (N_467,In_2443,In_1063);
nor U468 (N_468,In_321,In_1718);
nand U469 (N_469,In_2121,In_1674);
and U470 (N_470,In_2225,In_392);
or U471 (N_471,In_356,In_759);
nand U472 (N_472,In_2412,In_1229);
and U473 (N_473,In_2127,In_124);
nor U474 (N_474,In_2080,In_2119);
nor U475 (N_475,In_1466,In_1658);
and U476 (N_476,In_1742,In_1608);
and U477 (N_477,In_2444,In_336);
or U478 (N_478,In_955,In_1070);
nor U479 (N_479,In_693,In_629);
and U480 (N_480,In_433,In_1373);
or U481 (N_481,In_117,In_1673);
or U482 (N_482,In_1965,In_1802);
nand U483 (N_483,In_1384,In_736);
nor U484 (N_484,In_1372,In_187);
nor U485 (N_485,In_1032,In_2282);
nand U486 (N_486,In_328,In_227);
or U487 (N_487,In_2345,In_230);
nand U488 (N_488,In_979,In_1852);
nand U489 (N_489,In_1194,In_620);
nand U490 (N_490,In_2167,In_592);
nand U491 (N_491,In_1801,In_928);
nor U492 (N_492,In_984,In_827);
nand U493 (N_493,In_682,In_2175);
nand U494 (N_494,In_2059,In_482);
nor U495 (N_495,In_108,In_1683);
xor U496 (N_496,In_739,In_487);
and U497 (N_497,In_1360,In_376);
or U498 (N_498,In_1484,In_826);
or U499 (N_499,In_2475,In_712);
nand U500 (N_500,In_203,In_1149);
nand U501 (N_501,In_824,In_432);
and U502 (N_502,In_1681,In_425);
nor U503 (N_503,In_129,In_2489);
nor U504 (N_504,In_1583,In_2033);
or U505 (N_505,In_1157,In_876);
or U506 (N_506,In_1907,In_126);
or U507 (N_507,In_542,In_2187);
or U508 (N_508,In_1089,In_707);
and U509 (N_509,In_1517,In_917);
nor U510 (N_510,In_1676,In_19);
nand U511 (N_511,In_717,In_924);
xnor U512 (N_512,In_1725,In_642);
nor U513 (N_513,In_530,In_708);
nor U514 (N_514,In_1786,In_8);
nor U515 (N_515,In_1023,In_1048);
nand U516 (N_516,In_2456,In_2397);
and U517 (N_517,In_234,In_834);
nor U518 (N_518,In_1141,In_1124);
or U519 (N_519,In_91,In_1006);
xnor U520 (N_520,In_1634,In_675);
nand U521 (N_521,In_2414,In_1133);
nand U522 (N_522,In_566,In_965);
nor U523 (N_523,In_1488,In_2045);
and U524 (N_524,In_202,In_1414);
nor U525 (N_525,In_1128,In_1097);
nand U526 (N_526,In_2235,In_1274);
nand U527 (N_527,In_1472,In_1759);
nand U528 (N_528,In_501,In_888);
or U529 (N_529,In_2231,In_900);
and U530 (N_530,In_176,In_799);
and U531 (N_531,In_2010,In_2257);
or U532 (N_532,In_1086,In_60);
nor U533 (N_533,In_167,In_1966);
and U534 (N_534,In_133,In_2336);
nor U535 (N_535,In_565,In_130);
nand U536 (N_536,In_1840,In_1315);
and U537 (N_537,In_1685,In_1815);
xor U538 (N_538,In_1226,In_1561);
nor U539 (N_539,In_1540,In_2103);
nor U540 (N_540,In_558,In_2179);
nand U541 (N_541,In_1319,In_287);
nor U542 (N_542,In_128,In_24);
xnor U543 (N_543,In_2487,In_1030);
xor U544 (N_544,In_101,In_399);
nor U545 (N_545,In_1723,In_2498);
and U546 (N_546,In_143,In_2461);
or U547 (N_547,In_223,In_1670);
xor U548 (N_548,In_815,In_1477);
or U549 (N_549,In_419,In_471);
nor U550 (N_550,In_1501,In_2356);
nand U551 (N_551,In_1497,In_1962);
nand U552 (N_552,In_577,In_436);
and U553 (N_553,In_1915,In_2162);
nor U554 (N_554,In_595,In_35);
nand U555 (N_555,In_80,In_525);
or U556 (N_556,In_775,In_1378);
nor U557 (N_557,In_102,In_1694);
and U558 (N_558,In_877,In_1160);
or U559 (N_559,In_261,In_2061);
nor U560 (N_560,In_2413,In_2426);
nor U561 (N_561,In_445,In_2476);
xor U562 (N_562,In_1585,In_350);
or U563 (N_563,In_1233,In_1554);
or U564 (N_564,In_1995,In_2260);
or U565 (N_565,In_397,In_463);
xnor U566 (N_566,In_2194,In_1166);
or U567 (N_567,In_607,In_729);
or U568 (N_568,In_382,In_1985);
or U569 (N_569,In_1604,In_1154);
or U570 (N_570,In_1642,In_1295);
xnor U571 (N_571,In_1336,In_535);
nor U572 (N_572,In_1088,In_1667);
and U573 (N_573,In_1506,In_2419);
nor U574 (N_574,In_2200,In_752);
or U575 (N_575,In_1380,In_489);
and U576 (N_576,In_1286,In_1743);
and U577 (N_577,In_1093,In_1849);
or U578 (N_578,In_255,In_672);
and U579 (N_579,In_772,In_2027);
or U580 (N_580,In_262,In_2057);
nor U581 (N_581,In_1062,In_2155);
nand U582 (N_582,In_1980,In_604);
nand U583 (N_583,In_1235,In_291);
nor U584 (N_584,In_1804,In_831);
nor U585 (N_585,In_1323,In_1984);
or U586 (N_586,In_1557,In_889);
xor U587 (N_587,In_840,In_1463);
nand U588 (N_588,In_183,In_2457);
and U589 (N_589,In_526,In_994);
or U590 (N_590,In_763,In_726);
or U591 (N_591,In_2022,In_2191);
nor U592 (N_592,In_1230,In_1251);
and U593 (N_593,In_600,In_2083);
or U594 (N_594,In_598,In_554);
nor U595 (N_595,In_906,In_869);
or U596 (N_596,In_1663,In_2154);
nand U597 (N_597,In_1720,In_1382);
nor U598 (N_598,In_769,In_601);
nor U599 (N_599,In_2134,In_597);
or U600 (N_600,In_683,In_1227);
and U601 (N_601,In_1601,In_948);
nor U602 (N_602,In_2049,In_1025);
nor U603 (N_603,In_1645,In_1098);
xnor U604 (N_604,In_971,In_1782);
nor U605 (N_605,In_538,In_2094);
and U606 (N_606,In_1612,In_1675);
and U607 (N_607,In_1159,In_1162);
or U608 (N_608,In_846,In_1741);
or U609 (N_609,In_2101,In_2410);
nand U610 (N_610,In_790,In_1991);
nor U611 (N_611,In_318,In_1611);
nand U612 (N_612,In_1528,In_413);
or U613 (N_613,In_1153,In_1649);
nand U614 (N_614,In_1489,In_1898);
nand U615 (N_615,In_1563,In_1764);
nand U616 (N_616,In_1827,In_1729);
nand U617 (N_617,In_2445,In_2302);
nand U618 (N_618,In_586,In_2133);
nor U619 (N_619,In_1415,In_1021);
nand U620 (N_620,In_1080,In_2245);
xnor U621 (N_621,In_1090,In_30);
nand U622 (N_622,In_1275,In_1609);
or U623 (N_623,In_1212,In_2000);
nor U624 (N_624,In_39,In_1632);
nand U625 (N_625,In_609,In_502);
nand U626 (N_626,In_1231,In_431);
or U627 (N_627,In_300,In_581);
and U628 (N_628,In_938,In_2227);
and U629 (N_629,In_279,In_2241);
nand U630 (N_630,In_890,In_1304);
nor U631 (N_631,In_1341,In_1122);
nor U632 (N_632,In_1947,In_370);
nand U633 (N_633,In_1075,In_2161);
nand U634 (N_634,In_2141,In_290);
and U635 (N_635,In_1700,In_1281);
nor U636 (N_636,In_1731,In_388);
xor U637 (N_637,In_259,In_2205);
and U638 (N_638,In_2165,In_2453);
nor U639 (N_639,In_816,In_2329);
nand U640 (N_640,In_967,In_1047);
and U641 (N_641,In_1646,In_163);
nor U642 (N_642,In_2203,In_1326);
or U643 (N_643,In_2176,In_1518);
or U644 (N_644,In_1780,In_1103);
nor U645 (N_645,In_925,In_1068);
nor U646 (N_646,In_81,In_408);
and U647 (N_647,In_1322,In_643);
and U648 (N_648,In_553,In_902);
nor U649 (N_649,In_327,In_1175);
or U650 (N_650,In_2212,In_103);
nor U651 (N_651,In_658,In_398);
or U652 (N_652,In_1287,In_1137);
or U653 (N_653,In_161,In_2341);
nand U654 (N_654,In_46,In_2041);
or U655 (N_655,In_207,In_1391);
and U656 (N_656,In_1996,In_113);
nand U657 (N_657,In_2406,In_1922);
or U658 (N_658,In_533,In_1559);
nand U659 (N_659,In_2004,In_842);
or U660 (N_660,In_1232,In_1191);
xor U661 (N_661,In_453,In_1963);
nor U662 (N_662,In_1569,In_2208);
nand U663 (N_663,In_2423,In_1899);
nand U664 (N_664,In_1355,In_2343);
nor U665 (N_665,In_1684,In_648);
nand U666 (N_666,In_67,In_2328);
or U667 (N_667,In_1548,In_1331);
nor U668 (N_668,In_2335,In_1752);
xor U669 (N_669,In_1392,In_662);
nor U670 (N_670,In_1770,In_1236);
nand U671 (N_671,In_339,In_1510);
or U672 (N_672,In_1180,In_1939);
nor U673 (N_673,In_2258,In_1504);
and U674 (N_674,In_753,In_654);
or U675 (N_675,In_2006,In_1698);
nand U676 (N_676,In_1375,In_2332);
or U677 (N_677,In_918,In_2058);
nand U678 (N_678,In_2451,In_1496);
nand U679 (N_679,In_2116,In_2399);
nand U680 (N_680,In_631,In_276);
or U681 (N_681,In_1447,In_2281);
nand U682 (N_682,In_251,In_843);
or U683 (N_683,In_569,In_173);
and U684 (N_684,In_522,In_576);
and U685 (N_685,In_354,In_196);
nand U686 (N_686,In_1779,In_110);
and U687 (N_687,In_1680,In_1784);
nand U688 (N_688,In_534,In_999);
or U689 (N_689,In_2449,In_2073);
xnor U690 (N_690,In_1261,In_653);
or U691 (N_691,In_353,In_1138);
and U692 (N_692,In_1772,In_812);
nand U693 (N_693,In_26,In_1433);
or U694 (N_694,In_1083,In_2075);
nand U695 (N_695,In_175,In_1978);
nor U696 (N_696,In_1831,In_2052);
or U697 (N_697,In_2221,In_2001);
or U698 (N_698,In_181,In_1928);
nand U699 (N_699,In_1222,In_1988);
or U700 (N_700,In_571,In_2394);
or U701 (N_701,In_2024,In_1982);
nor U702 (N_702,In_961,In_1558);
or U703 (N_703,In_2063,In_326);
nor U704 (N_704,In_796,In_514);
and U705 (N_705,In_1579,In_2209);
and U706 (N_706,In_15,In_1449);
nand U707 (N_707,In_281,In_277);
nor U708 (N_708,In_787,In_1930);
or U709 (N_709,In_278,In_458);
and U710 (N_710,In_272,In_191);
or U711 (N_711,In_657,In_411);
and U712 (N_712,In_434,In_699);
nor U713 (N_713,In_1841,In_1458);
nor U714 (N_714,In_1066,In_594);
or U715 (N_715,In_16,In_310);
nor U716 (N_716,In_2032,In_1410);
nand U717 (N_717,In_784,In_2169);
and U718 (N_718,In_1767,In_2148);
xnor U719 (N_719,In_748,In_899);
and U720 (N_720,In_6,In_1483);
or U721 (N_721,In_1441,In_1473);
nand U722 (N_722,In_1084,In_2228);
and U723 (N_723,In_448,In_2047);
nor U724 (N_724,In_2196,In_692);
nor U725 (N_725,In_1578,In_266);
and U726 (N_726,In_1426,In_239);
or U727 (N_727,In_1842,In_1639);
or U728 (N_728,In_420,In_1136);
nand U729 (N_729,In_359,In_866);
and U730 (N_730,In_1549,In_946);
and U731 (N_731,In_1210,In_1516);
and U732 (N_732,In_1555,In_2338);
nor U733 (N_733,In_1699,In_1471);
nand U734 (N_734,In_2357,In_1453);
nand U735 (N_735,In_1531,In_1908);
nor U736 (N_736,In_462,In_1067);
or U737 (N_737,In_513,In_1185);
and U738 (N_738,In_111,In_1328);
nand U739 (N_739,In_1589,In_240);
or U740 (N_740,In_937,In_730);
and U741 (N_741,In_1689,In_1513);
nor U742 (N_742,In_364,In_2013);
and U743 (N_743,In_1911,In_694);
nor U744 (N_744,In_1526,In_1440);
nand U745 (N_745,In_45,In_1541);
nand U746 (N_746,In_1028,In_1291);
xnor U747 (N_747,In_2289,In_1661);
nand U748 (N_748,In_691,In_1552);
nand U749 (N_749,In_2273,In_863);
nand U750 (N_750,In_1241,In_2197);
or U751 (N_751,In_2249,In_2441);
and U752 (N_752,In_2270,In_1246);
and U753 (N_753,In_2430,In_1507);
nor U754 (N_754,In_872,In_2242);
nor U755 (N_755,In_76,In_579);
and U756 (N_756,In_1152,In_1237);
nor U757 (N_757,In_1167,In_2496);
nand U758 (N_758,In_1948,In_146);
or U759 (N_759,In_229,In_1756);
or U760 (N_760,In_1975,In_1774);
nand U761 (N_761,In_894,In_2354);
and U762 (N_762,In_38,In_1283);
nand U763 (N_763,In_954,In_2123);
nand U764 (N_764,In_1002,In_865);
nor U765 (N_765,In_94,In_992);
nor U766 (N_766,In_2039,In_1343);
nand U767 (N_767,In_1688,In_2247);
nor U768 (N_768,In_903,In_455);
and U769 (N_769,In_2198,In_1370);
nor U770 (N_770,In_192,In_2371);
and U771 (N_771,In_1242,In_1760);
or U772 (N_772,In_2408,In_106);
nor U773 (N_773,In_1053,In_2464);
nand U774 (N_774,In_610,In_613);
or U775 (N_775,In_1310,In_2459);
and U776 (N_776,In_1524,In_1857);
nor U777 (N_777,In_1660,In_1095);
or U778 (N_778,In_1398,In_1208);
or U779 (N_779,In_880,In_1260);
nor U780 (N_780,In_2460,In_2084);
nor U781 (N_781,In_511,In_2294);
and U782 (N_782,In_1065,In_2334);
nand U783 (N_783,In_920,In_86);
nor U784 (N_784,In_212,In_783);
nor U785 (N_785,In_1726,In_1253);
xor U786 (N_786,In_944,In_416);
nand U787 (N_787,In_1822,In_1280);
and U788 (N_788,In_1761,In_1960);
and U789 (N_789,In_2139,In_1265);
or U790 (N_790,In_2262,In_1708);
nor U791 (N_791,In_939,In_1817);
and U792 (N_792,In_418,In_352);
nor U793 (N_793,In_503,In_1830);
nand U794 (N_794,In_808,In_504);
or U795 (N_795,In_1356,In_454);
nand U796 (N_796,In_378,In_2028);
or U797 (N_797,In_474,In_340);
nor U798 (N_798,In_1247,In_1182);
nor U799 (N_799,In_2243,In_1598);
and U800 (N_800,In_725,In_1349);
or U801 (N_801,In_983,In_136);
and U802 (N_802,In_247,In_389);
or U803 (N_803,In_252,In_656);
nor U804 (N_804,In_2386,In_381);
nand U805 (N_805,In_1628,In_3);
and U806 (N_806,In_1755,In_1918);
and U807 (N_807,In_982,In_1855);
and U808 (N_808,In_881,In_2237);
nand U809 (N_809,In_375,In_1462);
nor U810 (N_810,In_957,In_85);
nand U811 (N_811,In_1717,In_733);
xor U812 (N_812,In_2046,In_5);
nor U813 (N_813,In_2077,In_2381);
xnor U814 (N_814,In_1732,In_238);
or U815 (N_815,In_1225,In_1077);
and U816 (N_816,In_1461,In_211);
and U817 (N_817,In_2234,In_1186);
or U818 (N_818,In_536,In_1969);
nand U819 (N_819,In_2297,In_685);
or U820 (N_820,In_1192,In_1521);
and U821 (N_821,In_1653,In_2370);
and U822 (N_822,In_1026,In_355);
nor U823 (N_823,In_1596,In_1337);
nand U824 (N_824,In_618,In_2043);
and U825 (N_825,In_875,In_1656);
nand U826 (N_826,In_825,In_2350);
and U827 (N_827,In_1534,In_233);
and U828 (N_828,In_308,In_460);
nand U829 (N_829,In_1214,In_331);
or U830 (N_830,In_2150,In_715);
or U831 (N_831,In_2290,In_951);
nor U832 (N_832,In_1264,In_293);
or U833 (N_833,In_2288,In_1861);
nor U834 (N_834,In_1288,In_2279);
or U835 (N_835,In_848,In_806);
and U836 (N_836,In_704,In_267);
and U837 (N_837,In_150,In_1904);
or U838 (N_838,In_1923,In_2078);
xnor U839 (N_839,In_265,In_612);
or U840 (N_840,In_2307,In_1176);
nand U841 (N_841,In_2226,In_945);
xnor U842 (N_842,In_867,In_960);
or U843 (N_843,In_2436,In_1244);
and U844 (N_844,In_68,In_1746);
xor U845 (N_845,In_2310,In_491);
or U846 (N_846,In_145,In_1416);
and U847 (N_847,In_2390,In_1719);
nand U848 (N_848,In_2126,In_990);
nor U849 (N_849,In_1120,In_2236);
or U850 (N_850,In_1550,In_1637);
nor U851 (N_851,In_1568,In_1000);
nand U852 (N_852,In_2458,In_810);
nor U853 (N_853,In_441,In_987);
or U854 (N_854,In_2113,In_1020);
nand U855 (N_855,In_1514,In_785);
or U856 (N_856,In_495,In_1018);
nand U857 (N_857,In_56,In_2418);
or U858 (N_858,In_1788,In_1809);
nand U859 (N_859,In_1538,In_1560);
and U860 (N_860,In_2337,In_541);
nor U861 (N_861,In_444,In_1638);
and U862 (N_862,In_2482,In_1114);
nand U863 (N_863,In_391,In_1);
and U864 (N_864,In_677,In_1332);
xnor U865 (N_865,In_837,In_1327);
or U866 (N_866,In_555,In_635);
nor U867 (N_867,In_854,In_1009);
xnor U868 (N_868,In_28,In_349);
nor U869 (N_869,In_1427,In_1105);
nor U870 (N_870,In_719,In_1591);
and U871 (N_871,In_2007,In_779);
or U872 (N_872,In_637,In_1094);
nor U873 (N_873,In_2157,In_1643);
nor U874 (N_874,In_1147,In_2011);
and U875 (N_875,In_1234,In_127);
or U876 (N_876,In_1491,In_302);
nand U877 (N_877,In_602,In_510);
or U878 (N_878,In_1567,In_2472);
nand U879 (N_879,In_638,In_271);
or U880 (N_880,In_2138,In_1926);
nand U881 (N_881,In_1955,In_1728);
or U882 (N_882,In_574,In_1562);
nand U883 (N_883,In_904,In_532);
nand U884 (N_884,In_908,In_570);
or U885 (N_885,In_1329,In_7);
nand U886 (N_886,In_170,In_549);
or U887 (N_887,In_2145,In_2296);
and U888 (N_888,In_1603,In_557);
nand U889 (N_889,In_243,In_2181);
or U890 (N_890,In_1515,In_519);
or U891 (N_891,In_36,In_442);
nand U892 (N_892,In_1368,In_385);
nand U893 (N_893,In_1342,In_443);
or U894 (N_894,In_1703,In_1790);
nor U895 (N_895,In_1397,In_1647);
and U896 (N_896,In_879,In_1301);
nor U897 (N_897,In_1168,In_1711);
xor U898 (N_898,In_2211,In_786);
and U899 (N_899,In_2325,In_282);
xnor U900 (N_900,In_1480,In_986);
or U901 (N_901,In_17,In_1602);
or U902 (N_902,In_1173,In_828);
nor U903 (N_903,In_897,In_2029);
nor U904 (N_904,In_2392,In_1837);
or U905 (N_905,In_280,In_330);
and U906 (N_906,In_1181,In_1200);
nor U907 (N_907,In_738,In_1838);
and U908 (N_908,In_2417,In_705);
nand U909 (N_909,In_2331,In_168);
nand U910 (N_910,In_2060,In_2330);
and U911 (N_911,In_1529,In_2189);
xor U912 (N_912,In_781,In_208);
and U913 (N_913,In_1793,In_1737);
or U914 (N_914,In_1303,In_1794);
nand U915 (N_915,In_851,In_472);
or U916 (N_916,In_1921,In_770);
xor U917 (N_917,In_2164,In_297);
nor U918 (N_918,In_1964,In_2100);
xor U919 (N_919,In_177,In_1309);
nor U920 (N_920,In_1163,In_1873);
nor U921 (N_921,In_776,In_1041);
or U922 (N_922,In_2300,In_477);
nor U923 (N_923,In_1403,In_582);
nand U924 (N_924,In_285,In_2317);
and U925 (N_925,In_833,In_1813);
nor U926 (N_926,In_118,In_1396);
nor U927 (N_927,In_1748,In_84);
nand U928 (N_928,In_1586,In_832);
and U929 (N_929,In_198,In_2346);
nand U930 (N_930,In_2277,In_1132);
and U931 (N_931,In_2479,In_1178);
and U932 (N_932,In_1730,In_927);
or U933 (N_933,In_1896,In_362);
xor U934 (N_934,In_1546,In_1064);
and U935 (N_935,In_1545,In_2117);
and U936 (N_936,In_1479,In_2314);
and U937 (N_937,In_49,In_2286);
and U938 (N_938,In_697,In_724);
or U939 (N_939,In_2411,In_2393);
or U940 (N_940,In_2442,In_2015);
or U941 (N_941,In_1409,In_303);
and U942 (N_942,In_72,In_696);
and U943 (N_943,In_1509,In_543);
nor U944 (N_944,In_1566,In_563);
nand U945 (N_945,In_898,In_2369);
nand U946 (N_946,In_728,In_750);
or U947 (N_947,In_1079,In_2428);
xnor U948 (N_948,In_572,In_706);
xnor U949 (N_949,In_1121,In_578);
nor U950 (N_950,In_1535,In_1347);
nor U951 (N_951,In_528,In_2388);
and U952 (N_952,In_1874,In_2463);
nand U953 (N_953,In_78,In_2081);
nand U954 (N_954,In_742,In_377);
nor U955 (N_955,In_1379,In_2269);
xnor U956 (N_956,In_401,In_109);
or U957 (N_957,In_2151,In_1705);
nand U958 (N_958,In_622,In_1193);
or U959 (N_959,In_1913,In_624);
and U960 (N_960,In_2031,In_836);
nand U961 (N_961,In_1713,In_1420);
and U962 (N_962,In_766,In_1695);
or U963 (N_963,In_2467,In_1081);
nor U964 (N_964,In_1245,In_722);
nand U965 (N_965,In_2219,In_1810);
and U966 (N_966,In_608,In_964);
and U967 (N_967,In_800,In_2173);
nor U968 (N_968,In_59,In_1277);
nor U969 (N_969,In_1851,In_913);
and U970 (N_970,In_414,In_1007);
xnor U971 (N_971,In_1595,In_47);
nor U972 (N_972,In_2160,In_1614);
or U973 (N_973,In_506,In_820);
nand U974 (N_974,In_153,In_1151);
nor U975 (N_975,In_1886,In_379);
or U976 (N_976,In_1042,In_1712);
or U977 (N_977,In_1635,In_2170);
and U978 (N_978,In_88,In_1363);
and U979 (N_979,In_301,In_2051);
nor U980 (N_980,In_345,In_926);
nor U981 (N_981,In_2387,In_1272);
nor U982 (N_982,In_915,In_2477);
or U983 (N_983,In_424,In_1432);
or U984 (N_984,In_121,In_2437);
nor U985 (N_985,In_2014,In_573);
nor U986 (N_986,In_65,In_1010);
nand U987 (N_987,In_1747,In_2424);
nand U988 (N_988,In_1974,In_402);
or U989 (N_989,In_1145,In_701);
nand U990 (N_990,In_1335,In_1871);
nand U991 (N_991,In_2048,In_1906);
or U992 (N_992,In_627,In_1211);
or U993 (N_993,In_286,In_2171);
or U994 (N_994,In_1364,In_1640);
and U995 (N_995,In_1919,In_791);
xnor U996 (N_996,In_1577,In_509);
and U997 (N_997,In_363,In_256);
and U998 (N_998,In_368,In_1029);
or U999 (N_999,In_1201,In_1511);
nand U1000 (N_1000,In_1224,In_1308);
nand U1001 (N_1001,In_1434,In_360);
or U1002 (N_1002,In_2396,In_1320);
xor U1003 (N_1003,In_2206,In_1590);
nand U1004 (N_1004,In_1428,In_650);
nor U1005 (N_1005,In_1054,In_2159);
nand U1006 (N_1006,In_1389,In_82);
and U1007 (N_1007,In_1664,In_1820);
xor U1008 (N_1008,In_77,In_1539);
nor U1009 (N_1009,In_1417,In_1045);
nor U1010 (N_1010,In_1787,In_131);
nand U1011 (N_1011,In_390,In_2348);
or U1012 (N_1012,In_1946,In_664);
xor U1013 (N_1013,In_162,In_1624);
or U1014 (N_1014,In_1424,In_744);
xor U1015 (N_1015,In_1016,In_2431);
nor U1016 (N_1016,In_1110,In_1693);
xnor U1017 (N_1017,In_1292,In_1011);
nor U1018 (N_1018,In_1188,In_1057);
nor U1019 (N_1019,In_197,In_1330);
or U1020 (N_1020,In_2216,In_1040);
nor U1021 (N_1021,In_2072,In_99);
and U1022 (N_1022,In_217,In_1127);
nor U1023 (N_1023,In_1565,In_721);
nor U1024 (N_1024,In_1036,In_1957);
nor U1025 (N_1025,In_226,In_2389);
xor U1026 (N_1026,In_1024,In_1864);
or U1027 (N_1027,In_550,In_680);
or U1028 (N_1028,In_1376,In_2002);
or U1029 (N_1029,In_674,In_2438);
nor U1030 (N_1030,In_2481,In_1636);
and U1031 (N_1031,In_1387,In_2285);
and U1032 (N_1032,In_2229,In_231);
nor U1033 (N_1033,In_1381,In_1262);
xor U1034 (N_1034,In_79,In_1150);
nor U1035 (N_1035,In_1812,In_1690);
nand U1036 (N_1036,In_1865,In_386);
nand U1037 (N_1037,In_2143,In_886);
nand U1038 (N_1038,In_1715,In_561);
and U1039 (N_1039,In_2137,In_2292);
xor U1040 (N_1040,In_1527,In_2299);
or U1041 (N_1041,In_209,In_459);
nor U1042 (N_1042,In_1867,In_312);
nand U1043 (N_1043,In_2034,In_1130);
and U1044 (N_1044,In_1457,In_2025);
or U1045 (N_1045,In_811,In_1481);
nand U1046 (N_1046,In_2062,In_1623);
nor U1047 (N_1047,In_856,In_1348);
and U1048 (N_1048,In_2204,In_2485);
nor U1049 (N_1049,In_1400,In_294);
nand U1050 (N_1050,In_1468,In_749);
and U1051 (N_1051,In_394,In_1074);
nand U1052 (N_1052,In_1536,In_2021);
and U1053 (N_1053,In_1902,In_1494);
or U1054 (N_1054,In_2492,In_1875);
xnor U1055 (N_1055,In_346,In_140);
nand U1056 (N_1056,In_1704,In_1547);
nand U1057 (N_1057,In_1551,In_1796);
and U1058 (N_1058,In_649,In_369);
and U1059 (N_1059,In_1615,In_2435);
nand U1060 (N_1060,In_2095,In_789);
nor U1061 (N_1061,In_1872,In_2425);
or U1062 (N_1062,In_1197,In_1104);
xor U1063 (N_1063,In_1574,In_1758);
and U1064 (N_1064,In_2232,In_1015);
or U1065 (N_1065,In_1940,In_2486);
or U1066 (N_1066,In_2353,In_2309);
nor U1067 (N_1067,In_1533,In_2380);
and U1068 (N_1068,In_224,In_1096);
or U1069 (N_1069,In_2055,In_1243);
and U1070 (N_1070,In_1017,In_2026);
or U1071 (N_1071,In_200,In_1184);
nand U1072 (N_1072,In_237,In_633);
nor U1073 (N_1073,In_919,In_367);
nand U1074 (N_1074,In_2142,In_1209);
and U1075 (N_1075,In_1679,In_862);
xnor U1076 (N_1076,In_754,In_333);
and U1077 (N_1077,In_993,In_273);
nor U1078 (N_1078,In_1196,In_921);
nand U1079 (N_1079,In_1887,In_2278);
and U1080 (N_1080,In_248,In_70);
nor U1081 (N_1081,In_1091,In_959);
or U1082 (N_1082,In_1691,In_1324);
nand U1083 (N_1083,In_403,In_450);
and U1084 (N_1084,In_969,In_1958);
nand U1085 (N_1085,In_1776,In_190);
nand U1086 (N_1086,In_83,In_1999);
nand U1087 (N_1087,In_1401,In_366);
or U1088 (N_1088,In_1131,In_686);
nand U1089 (N_1089,In_830,In_58);
xor U1090 (N_1090,In_537,In_546);
or U1091 (N_1091,In_142,In_723);
xnor U1092 (N_1092,In_1448,In_773);
and U1093 (N_1093,In_1266,In_1553);
and U1094 (N_1094,In_485,In_373);
nand U1095 (N_1095,In_1258,In_1248);
xor U1096 (N_1096,In_2090,In_936);
nor U1097 (N_1097,In_1987,In_1564);
nand U1098 (N_1098,In_1383,In_486);
nand U1099 (N_1099,In_1641,In_813);
nand U1100 (N_1100,In_966,In_66);
or U1101 (N_1101,In_25,In_2193);
and U1102 (N_1102,In_1777,In_481);
or U1103 (N_1103,In_1970,In_2108);
nand U1104 (N_1104,In_93,In_1727);
nand U1105 (N_1105,In_1189,In_254);
xnor U1106 (N_1106,In_1490,In_689);
nand U1107 (N_1107,In_351,In_985);
or U1108 (N_1108,In_1512,In_1129);
or U1109 (N_1109,In_737,In_1665);
and U1110 (N_1110,In_1573,In_1692);
and U1111 (N_1111,In_1305,In_144);
and U1112 (N_1112,In_1606,In_1072);
nand U1113 (N_1113,In_1897,In_1835);
nor U1114 (N_1114,In_617,In_560);
and U1115 (N_1115,In_1933,In_53);
nor U1116 (N_1116,In_1060,In_849);
nor U1117 (N_1117,In_1954,In_1469);
and U1118 (N_1118,In_43,In_2488);
and U1119 (N_1119,In_905,In_189);
nand U1120 (N_1120,In_2214,In_2474);
xor U1121 (N_1121,In_1575,In_158);
nand U1122 (N_1122,In_1848,In_1967);
nor U1123 (N_1123,In_1092,In_768);
and U1124 (N_1124,In_1659,In_884);
nand U1125 (N_1125,In_1993,In_2003);
and U1126 (N_1126,In_148,In_348);
nand U1127 (N_1127,In_2342,In_2076);
or U1128 (N_1128,In_1943,In_63);
nor U1129 (N_1129,In_358,In_1949);
and U1130 (N_1130,In_2146,In_958);
and U1131 (N_1131,In_1572,In_1254);
and U1132 (N_1132,In_970,In_2378);
and U1133 (N_1133,In_1144,In_1750);
and U1134 (N_1134,In_1829,In_257);
and U1135 (N_1135,In_288,In_1256);
or U1136 (N_1136,In_309,In_655);
xnor U1137 (N_1137,In_2490,In_679);
nand U1138 (N_1138,In_1672,In_429);
or U1139 (N_1139,In_478,In_2361);
nor U1140 (N_1140,In_480,In_304);
or U1141 (N_1141,In_407,In_1537);
and U1142 (N_1142,In_268,In_186);
xor U1143 (N_1143,In_1762,In_861);
nand U1144 (N_1144,In_1816,In_1312);
nor U1145 (N_1145,In_734,In_1134);
nand U1146 (N_1146,In_1402,In_1470);
nand U1147 (N_1147,In_169,In_2465);
or U1148 (N_1148,In_1613,In_22);
and U1149 (N_1149,In_1791,In_771);
nor U1150 (N_1150,In_1651,In_995);
or U1151 (N_1151,In_892,In_490);
or U1152 (N_1152,In_2259,In_325);
nand U1153 (N_1153,In_1724,In_2473);
or U1154 (N_1154,In_1365,In_626);
and U1155 (N_1155,In_1781,In_645);
or U1156 (N_1156,In_1219,In_1318);
and U1157 (N_1157,In_1823,In_1465);
and U1158 (N_1158,In_1847,In_2102);
or U1159 (N_1159,In_2462,In_659);
and U1160 (N_1160,In_1344,In_1834);
and U1161 (N_1161,In_2107,In_2420);
and U1162 (N_1162,In_159,In_1439);
or U1163 (N_1163,In_2483,In_430);
and U1164 (N_1164,In_2180,In_1696);
nand U1165 (N_1165,In_1476,In_410);
nand U1166 (N_1166,In_342,In_1686);
and U1167 (N_1167,In_1353,In_62);
nor U1168 (N_1168,In_1927,In_324);
xor U1169 (N_1169,In_1302,In_380);
or U1170 (N_1170,In_1631,In_1285);
and U1171 (N_1171,In_1677,In_2452);
and U1172 (N_1172,In_1493,In_1845);
or U1173 (N_1173,In_895,In_1833);
or U1174 (N_1174,In_2491,In_2074);
nor U1175 (N_1175,In_1799,In_1100);
nor U1176 (N_1176,In_1325,In_2263);
or U1177 (N_1177,In_1956,In_484);
xnor U1178 (N_1178,In_803,In_1630);
xor U1179 (N_1179,In_1421,In_213);
xor U1180 (N_1180,In_1866,In_1107);
or U1181 (N_1181,In_2178,In_384);
nand U1182 (N_1182,In_2379,In_727);
or U1183 (N_1183,In_599,In_2306);
and U1184 (N_1184,In_1832,In_154);
nor U1185 (N_1185,In_417,In_652);
nor U1186 (N_1186,In_1892,In_2177);
nor U1187 (N_1187,In_2327,In_1282);
and U1188 (N_1188,In_90,In_1362);
nor U1189 (N_1189,In_0,In_934);
and U1190 (N_1190,In_1345,In_702);
and U1191 (N_1191,In_1413,In_1113);
nor U1192 (N_1192,In_41,In_260);
nor U1193 (N_1193,In_2480,In_2469);
or U1194 (N_1194,In_1879,In_1205);
nand U1195 (N_1195,In_588,In_2398);
nor U1196 (N_1196,In_1702,In_1278);
xor U1197 (N_1197,In_1377,In_931);
or U1198 (N_1198,In_29,In_1004);
nor U1199 (N_1199,In_2499,In_802);
xnor U1200 (N_1200,In_2053,In_2224);
xor U1201 (N_1201,In_665,In_844);
nand U1202 (N_1202,In_31,In_1406);
xor U1203 (N_1203,In_2416,In_1255);
nand U1204 (N_1204,In_48,In_215);
nand U1205 (N_1205,In_449,In_1408);
nand U1206 (N_1206,In_1571,In_1880);
xor U1207 (N_1207,In_437,In_1744);
and U1208 (N_1208,In_1976,In_498);
or U1209 (N_1209,In_1438,In_630);
xnor U1210 (N_1210,In_54,In_1795);
and U1211 (N_1211,In_2091,In_2238);
nor U1212 (N_1212,In_2493,In_107);
and U1213 (N_1213,In_299,In_1942);
or U1214 (N_1214,In_1990,In_2484);
or U1215 (N_1215,In_1284,In_116);
nand U1216 (N_1216,In_1530,In_1523);
nand U1217 (N_1217,In_20,In_1454);
nor U1218 (N_1218,In_64,In_493);
nor U1219 (N_1219,In_1622,In_1038);
or U1220 (N_1220,In_1626,In_923);
and U1221 (N_1221,In_2005,In_2038);
and U1222 (N_1222,In_901,In_764);
and U1223 (N_1223,In_440,In_1542);
or U1224 (N_1224,In_1217,In_2192);
and U1225 (N_1225,In_2362,In_2364);
nor U1226 (N_1226,In_1357,In_2446);
xor U1227 (N_1227,In_1814,In_2056);
nor U1228 (N_1228,In_1944,In_1885);
nand U1229 (N_1229,In_2375,In_75);
nand U1230 (N_1230,In_1889,In_2019);
xnor U1231 (N_1231,In_1773,In_1894);
xor U1232 (N_1232,In_1600,In_1843);
xnor U1233 (N_1233,In_2324,In_319);
xnor U1234 (N_1234,In_2284,In_137);
nor U1235 (N_1235,In_2349,In_400);
nand U1236 (N_1236,In_615,In_222);
nor U1237 (N_1237,In_640,In_307);
or U1238 (N_1238,In_1459,In_910);
nand U1239 (N_1239,In_1039,In_1789);
nor U1240 (N_1240,In_857,In_1101);
nor U1241 (N_1241,In_1753,In_219);
and U1242 (N_1242,In_1116,In_452);
nor U1243 (N_1243,In_2384,In_1350);
and U1244 (N_1244,In_1126,In_1143);
or U1245 (N_1245,In_1900,In_1112);
and U1246 (N_1246,In_1474,In_242);
nor U1247 (N_1247,In_147,In_2071);
nor U1248 (N_1248,In_1850,In_871);
or U1249 (N_1249,In_2186,In_1338);
nand U1250 (N_1250,In_2032,In_1292);
nand U1251 (N_1251,In_1310,In_682);
nand U1252 (N_1252,In_1546,In_1450);
nor U1253 (N_1253,In_1435,In_1896);
or U1254 (N_1254,In_537,In_805);
nor U1255 (N_1255,In_2274,In_937);
nor U1256 (N_1256,In_430,In_1487);
and U1257 (N_1257,In_1012,In_1411);
and U1258 (N_1258,In_1717,In_609);
xor U1259 (N_1259,In_1331,In_1344);
nand U1260 (N_1260,In_1397,In_1534);
or U1261 (N_1261,In_1350,In_1184);
and U1262 (N_1262,In_584,In_1422);
nor U1263 (N_1263,In_2081,In_184);
xnor U1264 (N_1264,In_15,In_710);
or U1265 (N_1265,In_250,In_1975);
nand U1266 (N_1266,In_418,In_856);
and U1267 (N_1267,In_2462,In_1974);
or U1268 (N_1268,In_2067,In_1614);
nor U1269 (N_1269,In_456,In_2360);
or U1270 (N_1270,In_1034,In_628);
and U1271 (N_1271,In_1698,In_1747);
xor U1272 (N_1272,In_1404,In_682);
and U1273 (N_1273,In_545,In_163);
and U1274 (N_1274,In_2330,In_562);
nand U1275 (N_1275,In_2096,In_373);
or U1276 (N_1276,In_28,In_1076);
nand U1277 (N_1277,In_1563,In_850);
xnor U1278 (N_1278,In_2261,In_1210);
nor U1279 (N_1279,In_972,In_1946);
or U1280 (N_1280,In_823,In_2379);
or U1281 (N_1281,In_1909,In_1529);
xnor U1282 (N_1282,In_1860,In_1400);
or U1283 (N_1283,In_2423,In_2043);
or U1284 (N_1284,In_2115,In_1740);
nor U1285 (N_1285,In_1707,In_686);
nor U1286 (N_1286,In_1753,In_723);
or U1287 (N_1287,In_809,In_2440);
xnor U1288 (N_1288,In_1627,In_2042);
nor U1289 (N_1289,In_542,In_1640);
and U1290 (N_1290,In_1286,In_1999);
and U1291 (N_1291,In_1817,In_757);
or U1292 (N_1292,In_1157,In_92);
nor U1293 (N_1293,In_2,In_1950);
and U1294 (N_1294,In_700,In_576);
and U1295 (N_1295,In_1497,In_1476);
and U1296 (N_1296,In_2171,In_1874);
and U1297 (N_1297,In_963,In_86);
xnor U1298 (N_1298,In_1919,In_2487);
nor U1299 (N_1299,In_677,In_2429);
and U1300 (N_1300,In_387,In_1847);
nand U1301 (N_1301,In_1991,In_492);
and U1302 (N_1302,In_1453,In_1939);
or U1303 (N_1303,In_403,In_2048);
or U1304 (N_1304,In_1101,In_1002);
nand U1305 (N_1305,In_665,In_1948);
or U1306 (N_1306,In_1095,In_2011);
xor U1307 (N_1307,In_1924,In_2349);
nor U1308 (N_1308,In_588,In_2476);
or U1309 (N_1309,In_2251,In_2018);
nor U1310 (N_1310,In_1969,In_1150);
and U1311 (N_1311,In_1222,In_776);
nor U1312 (N_1312,In_1408,In_165);
nor U1313 (N_1313,In_23,In_1857);
nor U1314 (N_1314,In_1295,In_234);
or U1315 (N_1315,In_1349,In_252);
or U1316 (N_1316,In_925,In_2178);
or U1317 (N_1317,In_2403,In_2108);
nand U1318 (N_1318,In_435,In_2046);
and U1319 (N_1319,In_135,In_993);
nor U1320 (N_1320,In_172,In_1132);
and U1321 (N_1321,In_22,In_1357);
nor U1322 (N_1322,In_1477,In_1121);
and U1323 (N_1323,In_1365,In_839);
and U1324 (N_1324,In_2368,In_2326);
nand U1325 (N_1325,In_1611,In_1199);
nor U1326 (N_1326,In_226,In_865);
or U1327 (N_1327,In_2461,In_944);
xnor U1328 (N_1328,In_2460,In_1397);
nand U1329 (N_1329,In_23,In_1645);
nor U1330 (N_1330,In_2189,In_2412);
nand U1331 (N_1331,In_536,In_1315);
and U1332 (N_1332,In_1750,In_344);
nand U1333 (N_1333,In_620,In_2199);
nand U1334 (N_1334,In_196,In_2289);
nor U1335 (N_1335,In_1116,In_983);
nor U1336 (N_1336,In_1854,In_1438);
and U1337 (N_1337,In_1138,In_2137);
and U1338 (N_1338,In_2310,In_762);
nand U1339 (N_1339,In_1846,In_656);
and U1340 (N_1340,In_218,In_1371);
or U1341 (N_1341,In_2298,In_2054);
nand U1342 (N_1342,In_1147,In_1445);
and U1343 (N_1343,In_2061,In_1731);
nor U1344 (N_1344,In_815,In_2415);
nor U1345 (N_1345,In_670,In_183);
and U1346 (N_1346,In_1709,In_969);
or U1347 (N_1347,In_1207,In_1332);
and U1348 (N_1348,In_1695,In_274);
nor U1349 (N_1349,In_1047,In_1543);
or U1350 (N_1350,In_865,In_2453);
xor U1351 (N_1351,In_2305,In_2430);
or U1352 (N_1352,In_442,In_456);
and U1353 (N_1353,In_1994,In_602);
and U1354 (N_1354,In_1930,In_2439);
or U1355 (N_1355,In_1195,In_1889);
nand U1356 (N_1356,In_1463,In_221);
or U1357 (N_1357,In_2210,In_158);
and U1358 (N_1358,In_1905,In_1143);
xor U1359 (N_1359,In_1044,In_288);
or U1360 (N_1360,In_2053,In_24);
nand U1361 (N_1361,In_339,In_2266);
nand U1362 (N_1362,In_113,In_530);
and U1363 (N_1363,In_2477,In_85);
or U1364 (N_1364,In_1105,In_1820);
nor U1365 (N_1365,In_205,In_579);
nor U1366 (N_1366,In_2015,In_2331);
nor U1367 (N_1367,In_1909,In_959);
and U1368 (N_1368,In_177,In_1329);
or U1369 (N_1369,In_682,In_1877);
nor U1370 (N_1370,In_379,In_864);
or U1371 (N_1371,In_1758,In_1510);
and U1372 (N_1372,In_732,In_1088);
and U1373 (N_1373,In_629,In_1972);
or U1374 (N_1374,In_2346,In_1049);
and U1375 (N_1375,In_184,In_1403);
or U1376 (N_1376,In_1807,In_1875);
or U1377 (N_1377,In_2448,In_817);
nand U1378 (N_1378,In_464,In_165);
nor U1379 (N_1379,In_2144,In_778);
and U1380 (N_1380,In_2336,In_2159);
nor U1381 (N_1381,In_1728,In_1768);
xor U1382 (N_1382,In_563,In_2275);
nor U1383 (N_1383,In_1070,In_56);
and U1384 (N_1384,In_1841,In_1165);
nand U1385 (N_1385,In_1812,In_629);
and U1386 (N_1386,In_1496,In_1744);
and U1387 (N_1387,In_1353,In_1812);
or U1388 (N_1388,In_644,In_2103);
or U1389 (N_1389,In_40,In_823);
nor U1390 (N_1390,In_472,In_985);
and U1391 (N_1391,In_2442,In_1708);
or U1392 (N_1392,In_915,In_848);
or U1393 (N_1393,In_2371,In_604);
nand U1394 (N_1394,In_461,In_1385);
or U1395 (N_1395,In_2458,In_2290);
xnor U1396 (N_1396,In_823,In_498);
xor U1397 (N_1397,In_550,In_95);
and U1398 (N_1398,In_1666,In_1842);
and U1399 (N_1399,In_2299,In_81);
nor U1400 (N_1400,In_1571,In_155);
nand U1401 (N_1401,In_2307,In_521);
and U1402 (N_1402,In_1052,In_2307);
or U1403 (N_1403,In_30,In_1441);
and U1404 (N_1404,In_1617,In_1286);
and U1405 (N_1405,In_45,In_1947);
nor U1406 (N_1406,In_1601,In_323);
or U1407 (N_1407,In_1039,In_2357);
nand U1408 (N_1408,In_1020,In_1176);
nand U1409 (N_1409,In_653,In_1769);
or U1410 (N_1410,In_759,In_1948);
xnor U1411 (N_1411,In_2415,In_831);
nor U1412 (N_1412,In_2429,In_2090);
and U1413 (N_1413,In_2170,In_563);
and U1414 (N_1414,In_430,In_2044);
nand U1415 (N_1415,In_425,In_1600);
nor U1416 (N_1416,In_605,In_1039);
or U1417 (N_1417,In_1302,In_1585);
and U1418 (N_1418,In_1723,In_2250);
nand U1419 (N_1419,In_2109,In_1882);
nand U1420 (N_1420,In_2172,In_278);
xnor U1421 (N_1421,In_2163,In_1312);
nand U1422 (N_1422,In_1613,In_1534);
nor U1423 (N_1423,In_1851,In_368);
nor U1424 (N_1424,In_1502,In_2005);
nand U1425 (N_1425,In_1014,In_2267);
nor U1426 (N_1426,In_909,In_2468);
nor U1427 (N_1427,In_1748,In_1583);
xnor U1428 (N_1428,In_1186,In_511);
and U1429 (N_1429,In_413,In_1896);
or U1430 (N_1430,In_1322,In_62);
and U1431 (N_1431,In_1612,In_1296);
or U1432 (N_1432,In_754,In_2039);
or U1433 (N_1433,In_665,In_1061);
and U1434 (N_1434,In_335,In_558);
nor U1435 (N_1435,In_743,In_2263);
nor U1436 (N_1436,In_1491,In_1720);
nand U1437 (N_1437,In_99,In_128);
nor U1438 (N_1438,In_1100,In_884);
nand U1439 (N_1439,In_1831,In_628);
or U1440 (N_1440,In_589,In_0);
xnor U1441 (N_1441,In_2067,In_378);
nand U1442 (N_1442,In_325,In_1899);
nand U1443 (N_1443,In_1326,In_1637);
nand U1444 (N_1444,In_1253,In_1398);
nor U1445 (N_1445,In_822,In_211);
nor U1446 (N_1446,In_1608,In_112);
nor U1447 (N_1447,In_260,In_928);
nor U1448 (N_1448,In_2468,In_2055);
and U1449 (N_1449,In_1431,In_671);
and U1450 (N_1450,In_762,In_911);
nor U1451 (N_1451,In_2123,In_1972);
or U1452 (N_1452,In_2007,In_1667);
and U1453 (N_1453,In_1869,In_91);
nor U1454 (N_1454,In_273,In_149);
and U1455 (N_1455,In_227,In_1669);
or U1456 (N_1456,In_852,In_2090);
or U1457 (N_1457,In_1561,In_623);
and U1458 (N_1458,In_880,In_1578);
nand U1459 (N_1459,In_65,In_815);
and U1460 (N_1460,In_471,In_981);
nor U1461 (N_1461,In_909,In_1425);
or U1462 (N_1462,In_1662,In_141);
nand U1463 (N_1463,In_423,In_1340);
nand U1464 (N_1464,In_1284,In_1969);
and U1465 (N_1465,In_883,In_1948);
nand U1466 (N_1466,In_1259,In_1862);
xnor U1467 (N_1467,In_7,In_931);
and U1468 (N_1468,In_2323,In_2123);
nand U1469 (N_1469,In_293,In_537);
xor U1470 (N_1470,In_2173,In_1878);
nand U1471 (N_1471,In_2013,In_71);
nor U1472 (N_1472,In_169,In_1745);
or U1473 (N_1473,In_1524,In_1042);
and U1474 (N_1474,In_66,In_2071);
and U1475 (N_1475,In_1970,In_1433);
and U1476 (N_1476,In_1029,In_413);
xor U1477 (N_1477,In_597,In_1989);
and U1478 (N_1478,In_2381,In_523);
or U1479 (N_1479,In_2049,In_1341);
xor U1480 (N_1480,In_2302,In_858);
and U1481 (N_1481,In_1301,In_2049);
xnor U1482 (N_1482,In_1246,In_2023);
and U1483 (N_1483,In_1822,In_615);
nor U1484 (N_1484,In_2081,In_1137);
or U1485 (N_1485,In_301,In_1032);
nor U1486 (N_1486,In_1194,In_2040);
nand U1487 (N_1487,In_1468,In_1972);
nand U1488 (N_1488,In_1312,In_795);
or U1489 (N_1489,In_297,In_1459);
or U1490 (N_1490,In_813,In_503);
nand U1491 (N_1491,In_1161,In_13);
or U1492 (N_1492,In_1531,In_2152);
or U1493 (N_1493,In_823,In_756);
and U1494 (N_1494,In_642,In_853);
and U1495 (N_1495,In_413,In_2022);
or U1496 (N_1496,In_1724,In_1795);
nand U1497 (N_1497,In_1846,In_2228);
and U1498 (N_1498,In_2469,In_504);
or U1499 (N_1499,In_656,In_2186);
and U1500 (N_1500,In_2381,In_408);
nor U1501 (N_1501,In_262,In_1506);
nand U1502 (N_1502,In_111,In_1376);
or U1503 (N_1503,In_2070,In_2386);
nor U1504 (N_1504,In_600,In_2123);
or U1505 (N_1505,In_1742,In_1073);
nor U1506 (N_1506,In_1710,In_2300);
and U1507 (N_1507,In_1312,In_2437);
or U1508 (N_1508,In_229,In_1207);
xor U1509 (N_1509,In_1881,In_1273);
xnor U1510 (N_1510,In_1857,In_1514);
nor U1511 (N_1511,In_190,In_26);
nand U1512 (N_1512,In_1914,In_463);
or U1513 (N_1513,In_114,In_726);
or U1514 (N_1514,In_1031,In_1315);
or U1515 (N_1515,In_1557,In_669);
and U1516 (N_1516,In_675,In_601);
xor U1517 (N_1517,In_1188,In_1631);
nand U1518 (N_1518,In_1741,In_545);
nor U1519 (N_1519,In_1202,In_1212);
or U1520 (N_1520,In_1415,In_2208);
and U1521 (N_1521,In_981,In_1500);
and U1522 (N_1522,In_2264,In_296);
nor U1523 (N_1523,In_2412,In_496);
nor U1524 (N_1524,In_992,In_1303);
nor U1525 (N_1525,In_1944,In_1252);
nor U1526 (N_1526,In_240,In_1741);
and U1527 (N_1527,In_2097,In_2470);
nor U1528 (N_1528,In_1515,In_1477);
or U1529 (N_1529,In_1213,In_1585);
nor U1530 (N_1530,In_138,In_511);
or U1531 (N_1531,In_473,In_1272);
nor U1532 (N_1532,In_1261,In_1645);
and U1533 (N_1533,In_293,In_1260);
nor U1534 (N_1534,In_111,In_2131);
nand U1535 (N_1535,In_702,In_248);
xor U1536 (N_1536,In_1342,In_1357);
and U1537 (N_1537,In_1973,In_2068);
nor U1538 (N_1538,In_2189,In_193);
and U1539 (N_1539,In_176,In_1790);
nand U1540 (N_1540,In_73,In_375);
or U1541 (N_1541,In_37,In_1850);
xnor U1542 (N_1542,In_440,In_1099);
or U1543 (N_1543,In_463,In_1187);
or U1544 (N_1544,In_1262,In_1531);
xor U1545 (N_1545,In_842,In_905);
xnor U1546 (N_1546,In_1840,In_1722);
or U1547 (N_1547,In_311,In_1134);
nor U1548 (N_1548,In_1224,In_2011);
nor U1549 (N_1549,In_519,In_416);
nand U1550 (N_1550,In_2330,In_2114);
or U1551 (N_1551,In_697,In_1218);
nor U1552 (N_1552,In_754,In_1522);
and U1553 (N_1553,In_920,In_224);
nand U1554 (N_1554,In_203,In_474);
nand U1555 (N_1555,In_2170,In_1439);
and U1556 (N_1556,In_1489,In_368);
or U1557 (N_1557,In_334,In_1433);
and U1558 (N_1558,In_2211,In_2054);
or U1559 (N_1559,In_442,In_1866);
nand U1560 (N_1560,In_624,In_1262);
and U1561 (N_1561,In_1432,In_1544);
nand U1562 (N_1562,In_2429,In_1241);
nor U1563 (N_1563,In_1701,In_711);
nor U1564 (N_1564,In_982,In_1179);
or U1565 (N_1565,In_1839,In_2040);
xor U1566 (N_1566,In_1553,In_1016);
nor U1567 (N_1567,In_1829,In_759);
xor U1568 (N_1568,In_2343,In_527);
and U1569 (N_1569,In_173,In_65);
or U1570 (N_1570,In_2471,In_711);
nor U1571 (N_1571,In_1645,In_882);
or U1572 (N_1572,In_1184,In_242);
nand U1573 (N_1573,In_693,In_1757);
nand U1574 (N_1574,In_1724,In_1744);
and U1575 (N_1575,In_2391,In_932);
nand U1576 (N_1576,In_36,In_1628);
or U1577 (N_1577,In_2058,In_2412);
nor U1578 (N_1578,In_147,In_896);
or U1579 (N_1579,In_2045,In_2280);
and U1580 (N_1580,In_623,In_60);
or U1581 (N_1581,In_739,In_1020);
nor U1582 (N_1582,In_928,In_369);
nor U1583 (N_1583,In_1278,In_165);
or U1584 (N_1584,In_462,In_1861);
xnor U1585 (N_1585,In_1620,In_1877);
nand U1586 (N_1586,In_2276,In_2103);
nor U1587 (N_1587,In_392,In_1529);
nor U1588 (N_1588,In_968,In_772);
nor U1589 (N_1589,In_2460,In_131);
nand U1590 (N_1590,In_2206,In_138);
nand U1591 (N_1591,In_1814,In_1966);
nand U1592 (N_1592,In_464,In_1749);
and U1593 (N_1593,In_1175,In_1487);
and U1594 (N_1594,In_2371,In_10);
nand U1595 (N_1595,In_531,In_2238);
and U1596 (N_1596,In_757,In_1659);
nor U1597 (N_1597,In_548,In_2345);
nand U1598 (N_1598,In_479,In_1296);
xor U1599 (N_1599,In_2343,In_2356);
or U1600 (N_1600,In_445,In_1994);
nor U1601 (N_1601,In_1574,In_1228);
nand U1602 (N_1602,In_2082,In_2378);
and U1603 (N_1603,In_2096,In_2120);
nor U1604 (N_1604,In_667,In_1281);
nor U1605 (N_1605,In_946,In_75);
nor U1606 (N_1606,In_145,In_827);
nor U1607 (N_1607,In_122,In_1826);
nand U1608 (N_1608,In_1812,In_1671);
nor U1609 (N_1609,In_1602,In_413);
nand U1610 (N_1610,In_2190,In_88);
xnor U1611 (N_1611,In_556,In_750);
and U1612 (N_1612,In_414,In_1201);
or U1613 (N_1613,In_291,In_523);
and U1614 (N_1614,In_75,In_1183);
nand U1615 (N_1615,In_1170,In_1253);
nand U1616 (N_1616,In_1273,In_1126);
or U1617 (N_1617,In_1251,In_2267);
or U1618 (N_1618,In_2478,In_1988);
or U1619 (N_1619,In_1082,In_1592);
nor U1620 (N_1620,In_1224,In_292);
xor U1621 (N_1621,In_1987,In_1307);
and U1622 (N_1622,In_1958,In_958);
xnor U1623 (N_1623,In_1112,In_586);
nand U1624 (N_1624,In_104,In_1191);
nand U1625 (N_1625,In_814,In_470);
nand U1626 (N_1626,In_687,In_1362);
and U1627 (N_1627,In_1336,In_1214);
xnor U1628 (N_1628,In_287,In_2267);
nor U1629 (N_1629,In_935,In_259);
or U1630 (N_1630,In_2209,In_1279);
nor U1631 (N_1631,In_866,In_1361);
and U1632 (N_1632,In_288,In_1276);
and U1633 (N_1633,In_929,In_1797);
nand U1634 (N_1634,In_641,In_1874);
and U1635 (N_1635,In_1293,In_288);
nor U1636 (N_1636,In_1774,In_1524);
nand U1637 (N_1637,In_1049,In_2333);
nand U1638 (N_1638,In_1198,In_1156);
or U1639 (N_1639,In_1563,In_191);
and U1640 (N_1640,In_577,In_1669);
nor U1641 (N_1641,In_624,In_1409);
and U1642 (N_1642,In_1596,In_299);
nor U1643 (N_1643,In_290,In_1744);
nor U1644 (N_1644,In_616,In_539);
xnor U1645 (N_1645,In_2255,In_46);
and U1646 (N_1646,In_1233,In_2102);
or U1647 (N_1647,In_1815,In_1682);
nor U1648 (N_1648,In_1163,In_432);
nand U1649 (N_1649,In_1014,In_277);
nor U1650 (N_1650,In_1730,In_1356);
nor U1651 (N_1651,In_783,In_2473);
or U1652 (N_1652,In_431,In_184);
nor U1653 (N_1653,In_1635,In_2384);
nor U1654 (N_1654,In_843,In_924);
and U1655 (N_1655,In_242,In_1868);
and U1656 (N_1656,In_129,In_25);
nor U1657 (N_1657,In_2359,In_2061);
nor U1658 (N_1658,In_1577,In_1914);
nand U1659 (N_1659,In_1201,In_221);
xnor U1660 (N_1660,In_454,In_1134);
or U1661 (N_1661,In_2180,In_1836);
or U1662 (N_1662,In_2317,In_1354);
nor U1663 (N_1663,In_1368,In_2001);
and U1664 (N_1664,In_851,In_2464);
nor U1665 (N_1665,In_504,In_1300);
or U1666 (N_1666,In_1699,In_7);
or U1667 (N_1667,In_63,In_935);
and U1668 (N_1668,In_2387,In_1198);
or U1669 (N_1669,In_1149,In_1146);
xor U1670 (N_1670,In_1423,In_1408);
nand U1671 (N_1671,In_1082,In_2374);
and U1672 (N_1672,In_2168,In_1311);
nor U1673 (N_1673,In_1291,In_1901);
and U1674 (N_1674,In_1898,In_2432);
or U1675 (N_1675,In_1875,In_1939);
nor U1676 (N_1676,In_629,In_120);
nand U1677 (N_1677,In_2322,In_916);
nor U1678 (N_1678,In_2128,In_1001);
or U1679 (N_1679,In_1460,In_656);
nand U1680 (N_1680,In_1666,In_1240);
and U1681 (N_1681,In_1004,In_1997);
and U1682 (N_1682,In_728,In_1823);
or U1683 (N_1683,In_1787,In_803);
nand U1684 (N_1684,In_949,In_33);
xnor U1685 (N_1685,In_758,In_95);
and U1686 (N_1686,In_2489,In_2386);
and U1687 (N_1687,In_730,In_1686);
and U1688 (N_1688,In_1753,In_432);
or U1689 (N_1689,In_179,In_2363);
and U1690 (N_1690,In_1917,In_115);
and U1691 (N_1691,In_280,In_201);
xor U1692 (N_1692,In_1484,In_1570);
xor U1693 (N_1693,In_1997,In_999);
xor U1694 (N_1694,In_524,In_293);
or U1695 (N_1695,In_701,In_228);
and U1696 (N_1696,In_1106,In_441);
nor U1697 (N_1697,In_1261,In_1659);
and U1698 (N_1698,In_1547,In_567);
xor U1699 (N_1699,In_1275,In_293);
or U1700 (N_1700,In_377,In_223);
nand U1701 (N_1701,In_2268,In_2175);
nor U1702 (N_1702,In_2048,In_2213);
nand U1703 (N_1703,In_1419,In_1749);
xor U1704 (N_1704,In_2389,In_221);
nand U1705 (N_1705,In_984,In_1918);
nand U1706 (N_1706,In_1570,In_2181);
nand U1707 (N_1707,In_167,In_441);
nand U1708 (N_1708,In_622,In_1633);
nand U1709 (N_1709,In_1578,In_1623);
nor U1710 (N_1710,In_2042,In_1747);
nor U1711 (N_1711,In_1469,In_2001);
nor U1712 (N_1712,In_364,In_1436);
xor U1713 (N_1713,In_2043,In_960);
nor U1714 (N_1714,In_2105,In_1158);
or U1715 (N_1715,In_2341,In_2163);
or U1716 (N_1716,In_165,In_1814);
or U1717 (N_1717,In_229,In_934);
and U1718 (N_1718,In_889,In_1083);
nor U1719 (N_1719,In_1028,In_1993);
and U1720 (N_1720,In_225,In_1068);
nor U1721 (N_1721,In_113,In_858);
nand U1722 (N_1722,In_151,In_1535);
nor U1723 (N_1723,In_1155,In_1150);
nor U1724 (N_1724,In_2264,In_37);
nor U1725 (N_1725,In_392,In_1793);
and U1726 (N_1726,In_2307,In_43);
and U1727 (N_1727,In_2151,In_530);
nor U1728 (N_1728,In_1031,In_1777);
nor U1729 (N_1729,In_139,In_1760);
nand U1730 (N_1730,In_2467,In_63);
xor U1731 (N_1731,In_1783,In_1644);
or U1732 (N_1732,In_837,In_1000);
and U1733 (N_1733,In_1199,In_348);
xor U1734 (N_1734,In_1411,In_1884);
nor U1735 (N_1735,In_205,In_1717);
and U1736 (N_1736,In_1463,In_276);
or U1737 (N_1737,In_525,In_1527);
nand U1738 (N_1738,In_1160,In_1908);
nand U1739 (N_1739,In_407,In_892);
nand U1740 (N_1740,In_48,In_765);
xor U1741 (N_1741,In_1748,In_1221);
nand U1742 (N_1742,In_1693,In_2069);
or U1743 (N_1743,In_1486,In_1173);
and U1744 (N_1744,In_240,In_311);
or U1745 (N_1745,In_964,In_410);
nand U1746 (N_1746,In_107,In_1846);
or U1747 (N_1747,In_2244,In_372);
nor U1748 (N_1748,In_2190,In_393);
nor U1749 (N_1749,In_2021,In_628);
nand U1750 (N_1750,In_2073,In_2323);
nor U1751 (N_1751,In_2185,In_2468);
nor U1752 (N_1752,In_2419,In_1844);
nor U1753 (N_1753,In_2191,In_868);
or U1754 (N_1754,In_1636,In_2312);
nand U1755 (N_1755,In_790,In_253);
and U1756 (N_1756,In_933,In_875);
nand U1757 (N_1757,In_1549,In_1189);
or U1758 (N_1758,In_1997,In_167);
and U1759 (N_1759,In_1266,In_2497);
nand U1760 (N_1760,In_2490,In_2465);
xnor U1761 (N_1761,In_2100,In_26);
xor U1762 (N_1762,In_1399,In_1190);
or U1763 (N_1763,In_2193,In_1329);
or U1764 (N_1764,In_839,In_1255);
or U1765 (N_1765,In_2077,In_1913);
or U1766 (N_1766,In_2488,In_1537);
nand U1767 (N_1767,In_2407,In_1828);
nor U1768 (N_1768,In_1022,In_1157);
nor U1769 (N_1769,In_705,In_273);
nor U1770 (N_1770,In_170,In_1587);
or U1771 (N_1771,In_1763,In_226);
nor U1772 (N_1772,In_1105,In_1371);
nor U1773 (N_1773,In_394,In_1671);
and U1774 (N_1774,In_2097,In_421);
nand U1775 (N_1775,In_647,In_685);
nor U1776 (N_1776,In_1076,In_1017);
nand U1777 (N_1777,In_1296,In_2168);
nand U1778 (N_1778,In_1125,In_1274);
xnor U1779 (N_1779,In_318,In_180);
and U1780 (N_1780,In_498,In_584);
nor U1781 (N_1781,In_240,In_2050);
nand U1782 (N_1782,In_596,In_946);
xnor U1783 (N_1783,In_357,In_33);
and U1784 (N_1784,In_2041,In_2279);
or U1785 (N_1785,In_584,In_1613);
and U1786 (N_1786,In_1449,In_1443);
and U1787 (N_1787,In_504,In_2200);
nand U1788 (N_1788,In_500,In_1428);
xnor U1789 (N_1789,In_1696,In_2366);
and U1790 (N_1790,In_2470,In_325);
xor U1791 (N_1791,In_414,In_385);
nand U1792 (N_1792,In_2249,In_1233);
or U1793 (N_1793,In_147,In_1992);
xor U1794 (N_1794,In_2020,In_1052);
xor U1795 (N_1795,In_1535,In_920);
nor U1796 (N_1796,In_1744,In_1763);
or U1797 (N_1797,In_2165,In_834);
nand U1798 (N_1798,In_2216,In_132);
nand U1799 (N_1799,In_1146,In_2254);
nor U1800 (N_1800,In_201,In_1092);
and U1801 (N_1801,In_2376,In_1480);
or U1802 (N_1802,In_1520,In_984);
xor U1803 (N_1803,In_2114,In_1888);
nor U1804 (N_1804,In_510,In_1292);
and U1805 (N_1805,In_254,In_1665);
or U1806 (N_1806,In_2277,In_209);
and U1807 (N_1807,In_1358,In_75);
and U1808 (N_1808,In_882,In_241);
or U1809 (N_1809,In_2309,In_527);
or U1810 (N_1810,In_2069,In_258);
nand U1811 (N_1811,In_1171,In_761);
and U1812 (N_1812,In_174,In_1639);
nand U1813 (N_1813,In_1891,In_1157);
nor U1814 (N_1814,In_530,In_2134);
nand U1815 (N_1815,In_271,In_2428);
and U1816 (N_1816,In_1617,In_2252);
and U1817 (N_1817,In_1588,In_1742);
nor U1818 (N_1818,In_1277,In_2226);
and U1819 (N_1819,In_38,In_808);
nand U1820 (N_1820,In_975,In_1695);
or U1821 (N_1821,In_2401,In_234);
or U1822 (N_1822,In_921,In_128);
and U1823 (N_1823,In_688,In_1285);
and U1824 (N_1824,In_304,In_1352);
nand U1825 (N_1825,In_625,In_2326);
and U1826 (N_1826,In_596,In_798);
or U1827 (N_1827,In_1307,In_2343);
and U1828 (N_1828,In_433,In_2407);
and U1829 (N_1829,In_292,In_564);
and U1830 (N_1830,In_1444,In_1550);
nand U1831 (N_1831,In_1888,In_1401);
and U1832 (N_1832,In_2219,In_708);
nor U1833 (N_1833,In_1164,In_1484);
and U1834 (N_1834,In_67,In_1387);
xor U1835 (N_1835,In_2032,In_118);
xor U1836 (N_1836,In_2278,In_573);
nor U1837 (N_1837,In_920,In_761);
xnor U1838 (N_1838,In_383,In_1882);
nand U1839 (N_1839,In_789,In_1106);
or U1840 (N_1840,In_1763,In_1306);
nand U1841 (N_1841,In_146,In_1111);
or U1842 (N_1842,In_1159,In_1904);
and U1843 (N_1843,In_269,In_558);
nor U1844 (N_1844,In_993,In_1328);
nand U1845 (N_1845,In_2041,In_265);
or U1846 (N_1846,In_2113,In_2315);
or U1847 (N_1847,In_2122,In_1964);
and U1848 (N_1848,In_2381,In_1965);
nand U1849 (N_1849,In_1032,In_64);
or U1850 (N_1850,In_424,In_749);
and U1851 (N_1851,In_1328,In_614);
and U1852 (N_1852,In_2411,In_2447);
or U1853 (N_1853,In_34,In_1824);
nor U1854 (N_1854,In_121,In_459);
nor U1855 (N_1855,In_1967,In_1337);
nand U1856 (N_1856,In_729,In_342);
nor U1857 (N_1857,In_1582,In_1208);
and U1858 (N_1858,In_1551,In_1151);
nor U1859 (N_1859,In_2299,In_1966);
nand U1860 (N_1860,In_312,In_499);
nor U1861 (N_1861,In_1452,In_1333);
nand U1862 (N_1862,In_1476,In_938);
xnor U1863 (N_1863,In_1062,In_1088);
nor U1864 (N_1864,In_151,In_2134);
and U1865 (N_1865,In_947,In_1720);
nor U1866 (N_1866,In_886,In_1426);
nand U1867 (N_1867,In_1893,In_2220);
and U1868 (N_1868,In_2353,In_1393);
or U1869 (N_1869,In_933,In_1876);
and U1870 (N_1870,In_650,In_1334);
and U1871 (N_1871,In_96,In_1829);
nor U1872 (N_1872,In_1050,In_865);
xor U1873 (N_1873,In_2057,In_1995);
nor U1874 (N_1874,In_979,In_360);
or U1875 (N_1875,In_1613,In_1460);
nand U1876 (N_1876,In_2301,In_91);
nand U1877 (N_1877,In_259,In_431);
or U1878 (N_1878,In_1224,In_1828);
and U1879 (N_1879,In_1630,In_440);
and U1880 (N_1880,In_2498,In_468);
and U1881 (N_1881,In_379,In_290);
nor U1882 (N_1882,In_845,In_2403);
nor U1883 (N_1883,In_1392,In_933);
nor U1884 (N_1884,In_697,In_1267);
and U1885 (N_1885,In_1343,In_1157);
or U1886 (N_1886,In_1221,In_2442);
or U1887 (N_1887,In_1890,In_941);
or U1888 (N_1888,In_583,In_1539);
or U1889 (N_1889,In_259,In_626);
or U1890 (N_1890,In_508,In_2333);
nand U1891 (N_1891,In_2460,In_1748);
or U1892 (N_1892,In_476,In_1276);
or U1893 (N_1893,In_294,In_2377);
or U1894 (N_1894,In_504,In_1916);
and U1895 (N_1895,In_1578,In_1616);
nand U1896 (N_1896,In_870,In_2242);
or U1897 (N_1897,In_260,In_2161);
nor U1898 (N_1898,In_302,In_2115);
or U1899 (N_1899,In_431,In_44);
or U1900 (N_1900,In_605,In_1879);
nor U1901 (N_1901,In_2193,In_2063);
and U1902 (N_1902,In_1578,In_161);
nor U1903 (N_1903,In_1855,In_2234);
and U1904 (N_1904,In_751,In_1130);
xnor U1905 (N_1905,In_1429,In_582);
and U1906 (N_1906,In_1332,In_822);
or U1907 (N_1907,In_373,In_1836);
nand U1908 (N_1908,In_1682,In_757);
nand U1909 (N_1909,In_1406,In_2028);
and U1910 (N_1910,In_974,In_1888);
nor U1911 (N_1911,In_83,In_784);
xnor U1912 (N_1912,In_1381,In_1899);
and U1913 (N_1913,In_1248,In_1719);
or U1914 (N_1914,In_2289,In_516);
or U1915 (N_1915,In_171,In_994);
nand U1916 (N_1916,In_541,In_198);
xnor U1917 (N_1917,In_2304,In_1408);
or U1918 (N_1918,In_394,In_1002);
nor U1919 (N_1919,In_1772,In_945);
nor U1920 (N_1920,In_1128,In_1708);
nand U1921 (N_1921,In_1930,In_243);
nand U1922 (N_1922,In_1086,In_205);
nand U1923 (N_1923,In_1703,In_1545);
and U1924 (N_1924,In_730,In_1528);
or U1925 (N_1925,In_169,In_1191);
or U1926 (N_1926,In_229,In_2275);
and U1927 (N_1927,In_1410,In_1007);
or U1928 (N_1928,In_1181,In_42);
nand U1929 (N_1929,In_1251,In_1502);
nand U1930 (N_1930,In_782,In_2431);
or U1931 (N_1931,In_1678,In_869);
nand U1932 (N_1932,In_1729,In_2247);
or U1933 (N_1933,In_1775,In_918);
nor U1934 (N_1934,In_1937,In_426);
nor U1935 (N_1935,In_2194,In_2422);
or U1936 (N_1936,In_246,In_1538);
nand U1937 (N_1937,In_2402,In_2259);
nor U1938 (N_1938,In_111,In_442);
or U1939 (N_1939,In_1853,In_1898);
nor U1940 (N_1940,In_1137,In_2447);
and U1941 (N_1941,In_1153,In_513);
nand U1942 (N_1942,In_2444,In_305);
nor U1943 (N_1943,In_2080,In_1425);
and U1944 (N_1944,In_1995,In_1258);
nand U1945 (N_1945,In_1185,In_229);
nor U1946 (N_1946,In_688,In_788);
nor U1947 (N_1947,In_2439,In_1910);
nand U1948 (N_1948,In_1456,In_1821);
nand U1949 (N_1949,In_691,In_1222);
nand U1950 (N_1950,In_2206,In_1879);
xnor U1951 (N_1951,In_702,In_1708);
and U1952 (N_1952,In_1555,In_334);
or U1953 (N_1953,In_1237,In_401);
or U1954 (N_1954,In_2014,In_807);
nor U1955 (N_1955,In_1999,In_2403);
nand U1956 (N_1956,In_272,In_1025);
or U1957 (N_1957,In_747,In_1791);
xnor U1958 (N_1958,In_1503,In_1042);
and U1959 (N_1959,In_2287,In_725);
nor U1960 (N_1960,In_489,In_1640);
nand U1961 (N_1961,In_1938,In_2293);
nor U1962 (N_1962,In_2033,In_491);
nand U1963 (N_1963,In_2378,In_957);
and U1964 (N_1964,In_393,In_2400);
or U1965 (N_1965,In_979,In_406);
nor U1966 (N_1966,In_1750,In_223);
xnor U1967 (N_1967,In_2231,In_411);
nand U1968 (N_1968,In_2049,In_1527);
and U1969 (N_1969,In_860,In_2177);
and U1970 (N_1970,In_1417,In_486);
or U1971 (N_1971,In_2385,In_640);
or U1972 (N_1972,In_280,In_1888);
and U1973 (N_1973,In_1709,In_2269);
and U1974 (N_1974,In_2411,In_1682);
or U1975 (N_1975,In_1041,In_611);
nor U1976 (N_1976,In_1955,In_1504);
xnor U1977 (N_1977,In_1334,In_2451);
nand U1978 (N_1978,In_1962,In_1468);
nor U1979 (N_1979,In_1060,In_2266);
xor U1980 (N_1980,In_1850,In_899);
and U1981 (N_1981,In_1063,In_1502);
nor U1982 (N_1982,In_1118,In_2222);
and U1983 (N_1983,In_163,In_828);
and U1984 (N_1984,In_394,In_455);
nand U1985 (N_1985,In_1628,In_1996);
nand U1986 (N_1986,In_801,In_2338);
and U1987 (N_1987,In_1098,In_2102);
and U1988 (N_1988,In_888,In_103);
or U1989 (N_1989,In_2362,In_1332);
nand U1990 (N_1990,In_1667,In_936);
xor U1991 (N_1991,In_903,In_2353);
nand U1992 (N_1992,In_626,In_1408);
nand U1993 (N_1993,In_2033,In_1156);
xor U1994 (N_1994,In_1479,In_137);
xnor U1995 (N_1995,In_630,In_1049);
or U1996 (N_1996,In_1863,In_458);
or U1997 (N_1997,In_483,In_1740);
or U1998 (N_1998,In_1803,In_294);
nand U1999 (N_1999,In_1514,In_840);
and U2000 (N_2000,In_209,In_697);
nand U2001 (N_2001,In_2270,In_1759);
nand U2002 (N_2002,In_1896,In_1398);
and U2003 (N_2003,In_121,In_1817);
and U2004 (N_2004,In_555,In_1791);
or U2005 (N_2005,In_1559,In_1703);
nor U2006 (N_2006,In_756,In_1595);
and U2007 (N_2007,In_1105,In_110);
and U2008 (N_2008,In_76,In_1784);
nand U2009 (N_2009,In_1377,In_233);
nand U2010 (N_2010,In_2048,In_1521);
nor U2011 (N_2011,In_1771,In_830);
nor U2012 (N_2012,In_662,In_1733);
and U2013 (N_2013,In_1036,In_836);
and U2014 (N_2014,In_1156,In_624);
xnor U2015 (N_2015,In_2037,In_1730);
nor U2016 (N_2016,In_56,In_2254);
and U2017 (N_2017,In_1807,In_2496);
nand U2018 (N_2018,In_2390,In_1850);
xnor U2019 (N_2019,In_2366,In_425);
nor U2020 (N_2020,In_856,In_1616);
and U2021 (N_2021,In_2170,In_427);
nor U2022 (N_2022,In_901,In_1425);
nand U2023 (N_2023,In_2142,In_1197);
nor U2024 (N_2024,In_982,In_783);
and U2025 (N_2025,In_1604,In_2188);
nor U2026 (N_2026,In_926,In_1984);
xor U2027 (N_2027,In_1070,In_2020);
nor U2028 (N_2028,In_1869,In_969);
and U2029 (N_2029,In_2457,In_2146);
nand U2030 (N_2030,In_674,In_1427);
nand U2031 (N_2031,In_1735,In_2277);
and U2032 (N_2032,In_1983,In_695);
nor U2033 (N_2033,In_938,In_2067);
or U2034 (N_2034,In_604,In_276);
and U2035 (N_2035,In_400,In_1014);
or U2036 (N_2036,In_1815,In_2394);
nor U2037 (N_2037,In_723,In_847);
or U2038 (N_2038,In_1202,In_551);
or U2039 (N_2039,In_1760,In_297);
or U2040 (N_2040,In_1142,In_683);
xnor U2041 (N_2041,In_2239,In_1399);
xnor U2042 (N_2042,In_1504,In_1898);
or U2043 (N_2043,In_1966,In_1562);
or U2044 (N_2044,In_411,In_2091);
xnor U2045 (N_2045,In_2007,In_1305);
and U2046 (N_2046,In_1205,In_932);
nand U2047 (N_2047,In_1198,In_19);
xnor U2048 (N_2048,In_2380,In_1630);
and U2049 (N_2049,In_1533,In_226);
xnor U2050 (N_2050,In_2288,In_312);
nand U2051 (N_2051,In_19,In_2151);
nand U2052 (N_2052,In_437,In_941);
nand U2053 (N_2053,In_33,In_1721);
nand U2054 (N_2054,In_434,In_1743);
and U2055 (N_2055,In_1328,In_1945);
or U2056 (N_2056,In_1637,In_267);
and U2057 (N_2057,In_2114,In_363);
nand U2058 (N_2058,In_2199,In_1803);
xor U2059 (N_2059,In_224,In_546);
nand U2060 (N_2060,In_1626,In_1887);
nor U2061 (N_2061,In_1783,In_724);
or U2062 (N_2062,In_1813,In_1516);
nand U2063 (N_2063,In_574,In_2446);
xor U2064 (N_2064,In_1516,In_457);
and U2065 (N_2065,In_41,In_2287);
or U2066 (N_2066,In_1488,In_466);
or U2067 (N_2067,In_2117,In_190);
or U2068 (N_2068,In_1462,In_1816);
nor U2069 (N_2069,In_1179,In_223);
and U2070 (N_2070,In_2205,In_1545);
nand U2071 (N_2071,In_1938,In_221);
or U2072 (N_2072,In_410,In_331);
and U2073 (N_2073,In_2038,In_306);
or U2074 (N_2074,In_1131,In_732);
and U2075 (N_2075,In_893,In_1863);
or U2076 (N_2076,In_367,In_2017);
or U2077 (N_2077,In_1064,In_1180);
and U2078 (N_2078,In_1530,In_1855);
xnor U2079 (N_2079,In_1518,In_244);
xor U2080 (N_2080,In_2392,In_278);
and U2081 (N_2081,In_1586,In_1253);
and U2082 (N_2082,In_1797,In_1716);
nor U2083 (N_2083,In_1758,In_633);
nor U2084 (N_2084,In_1533,In_1022);
nand U2085 (N_2085,In_1423,In_347);
or U2086 (N_2086,In_2303,In_2307);
or U2087 (N_2087,In_508,In_1832);
and U2088 (N_2088,In_983,In_843);
nor U2089 (N_2089,In_1248,In_1418);
xnor U2090 (N_2090,In_2279,In_1780);
nor U2091 (N_2091,In_1074,In_1825);
nand U2092 (N_2092,In_1438,In_1620);
and U2093 (N_2093,In_1572,In_685);
nor U2094 (N_2094,In_2445,In_1399);
or U2095 (N_2095,In_296,In_2029);
or U2096 (N_2096,In_2475,In_2201);
nor U2097 (N_2097,In_1940,In_2463);
and U2098 (N_2098,In_531,In_108);
nand U2099 (N_2099,In_1471,In_1445);
nor U2100 (N_2100,In_2121,In_93);
or U2101 (N_2101,In_839,In_1332);
and U2102 (N_2102,In_742,In_2425);
nor U2103 (N_2103,In_30,In_1081);
or U2104 (N_2104,In_773,In_10);
nand U2105 (N_2105,In_1109,In_1269);
xnor U2106 (N_2106,In_98,In_592);
and U2107 (N_2107,In_1893,In_1900);
nor U2108 (N_2108,In_25,In_2065);
and U2109 (N_2109,In_198,In_2341);
or U2110 (N_2110,In_1750,In_1604);
nand U2111 (N_2111,In_1591,In_2484);
nand U2112 (N_2112,In_1139,In_2176);
and U2113 (N_2113,In_1049,In_272);
xor U2114 (N_2114,In_649,In_403);
or U2115 (N_2115,In_614,In_1943);
and U2116 (N_2116,In_417,In_443);
xor U2117 (N_2117,In_1557,In_635);
nand U2118 (N_2118,In_2080,In_2484);
and U2119 (N_2119,In_2366,In_314);
or U2120 (N_2120,In_1725,In_2265);
or U2121 (N_2121,In_1900,In_1196);
or U2122 (N_2122,In_2418,In_1849);
xor U2123 (N_2123,In_159,In_224);
and U2124 (N_2124,In_409,In_35);
and U2125 (N_2125,In_1204,In_1295);
nor U2126 (N_2126,In_1915,In_806);
or U2127 (N_2127,In_220,In_719);
xor U2128 (N_2128,In_2054,In_1979);
nor U2129 (N_2129,In_1318,In_1868);
or U2130 (N_2130,In_1542,In_1919);
and U2131 (N_2131,In_553,In_779);
nand U2132 (N_2132,In_1630,In_2497);
nand U2133 (N_2133,In_1490,In_223);
nor U2134 (N_2134,In_611,In_794);
and U2135 (N_2135,In_552,In_376);
xor U2136 (N_2136,In_903,In_836);
nand U2137 (N_2137,In_1434,In_1883);
nand U2138 (N_2138,In_1419,In_2118);
nand U2139 (N_2139,In_749,In_1733);
or U2140 (N_2140,In_1358,In_548);
or U2141 (N_2141,In_1872,In_1999);
nand U2142 (N_2142,In_1946,In_1178);
or U2143 (N_2143,In_2121,In_180);
or U2144 (N_2144,In_2265,In_1346);
nand U2145 (N_2145,In_2004,In_545);
xnor U2146 (N_2146,In_1034,In_1833);
or U2147 (N_2147,In_1124,In_2143);
or U2148 (N_2148,In_1809,In_1253);
or U2149 (N_2149,In_2178,In_864);
nor U2150 (N_2150,In_1589,In_2240);
nand U2151 (N_2151,In_571,In_1029);
and U2152 (N_2152,In_1294,In_1921);
or U2153 (N_2153,In_1121,In_2363);
nor U2154 (N_2154,In_638,In_2410);
nand U2155 (N_2155,In_1303,In_1304);
or U2156 (N_2156,In_351,In_162);
nor U2157 (N_2157,In_1305,In_1037);
and U2158 (N_2158,In_1299,In_883);
or U2159 (N_2159,In_371,In_1585);
or U2160 (N_2160,In_519,In_1041);
nand U2161 (N_2161,In_578,In_1156);
nor U2162 (N_2162,In_2128,In_1407);
xor U2163 (N_2163,In_727,In_336);
and U2164 (N_2164,In_1122,In_1214);
and U2165 (N_2165,In_1109,In_1813);
nand U2166 (N_2166,In_1919,In_2346);
nand U2167 (N_2167,In_1932,In_1667);
nand U2168 (N_2168,In_1970,In_58);
and U2169 (N_2169,In_1131,In_729);
xnor U2170 (N_2170,In_420,In_1594);
or U2171 (N_2171,In_2411,In_1571);
xor U2172 (N_2172,In_37,In_631);
or U2173 (N_2173,In_1071,In_888);
nor U2174 (N_2174,In_1242,In_1313);
and U2175 (N_2175,In_1103,In_13);
xor U2176 (N_2176,In_1827,In_1877);
or U2177 (N_2177,In_94,In_2497);
and U2178 (N_2178,In_788,In_491);
nand U2179 (N_2179,In_1397,In_1652);
nand U2180 (N_2180,In_2135,In_914);
nor U2181 (N_2181,In_17,In_2195);
nand U2182 (N_2182,In_2213,In_2364);
nor U2183 (N_2183,In_1775,In_829);
nor U2184 (N_2184,In_403,In_1292);
and U2185 (N_2185,In_932,In_448);
nand U2186 (N_2186,In_1549,In_900);
nand U2187 (N_2187,In_344,In_1235);
or U2188 (N_2188,In_732,In_2194);
or U2189 (N_2189,In_571,In_113);
and U2190 (N_2190,In_2384,In_1010);
or U2191 (N_2191,In_384,In_2335);
and U2192 (N_2192,In_2443,In_17);
xor U2193 (N_2193,In_133,In_918);
or U2194 (N_2194,In_813,In_1925);
nand U2195 (N_2195,In_126,In_615);
nand U2196 (N_2196,In_2287,In_547);
xnor U2197 (N_2197,In_1824,In_1715);
xnor U2198 (N_2198,In_1880,In_1623);
and U2199 (N_2199,In_1644,In_1157);
nand U2200 (N_2200,In_515,In_1176);
nor U2201 (N_2201,In_396,In_2102);
and U2202 (N_2202,In_1403,In_19);
or U2203 (N_2203,In_647,In_2229);
or U2204 (N_2204,In_1961,In_419);
or U2205 (N_2205,In_1049,In_680);
nor U2206 (N_2206,In_363,In_2368);
or U2207 (N_2207,In_352,In_959);
nand U2208 (N_2208,In_1073,In_445);
nand U2209 (N_2209,In_2418,In_23);
nand U2210 (N_2210,In_401,In_1909);
and U2211 (N_2211,In_903,In_898);
xnor U2212 (N_2212,In_1254,In_482);
or U2213 (N_2213,In_850,In_2213);
nor U2214 (N_2214,In_346,In_1846);
nand U2215 (N_2215,In_1231,In_752);
xnor U2216 (N_2216,In_1302,In_1847);
or U2217 (N_2217,In_2326,In_654);
nor U2218 (N_2218,In_953,In_568);
and U2219 (N_2219,In_1622,In_1282);
and U2220 (N_2220,In_1291,In_1898);
or U2221 (N_2221,In_2322,In_1678);
or U2222 (N_2222,In_45,In_2348);
nand U2223 (N_2223,In_1578,In_569);
nand U2224 (N_2224,In_2467,In_30);
nand U2225 (N_2225,In_2092,In_631);
and U2226 (N_2226,In_371,In_1218);
nand U2227 (N_2227,In_1297,In_220);
and U2228 (N_2228,In_1795,In_2324);
and U2229 (N_2229,In_2437,In_1685);
or U2230 (N_2230,In_2176,In_164);
or U2231 (N_2231,In_1378,In_1937);
and U2232 (N_2232,In_1031,In_1612);
nor U2233 (N_2233,In_1398,In_1607);
nand U2234 (N_2234,In_1176,In_462);
and U2235 (N_2235,In_1210,In_1348);
or U2236 (N_2236,In_1050,In_1272);
xor U2237 (N_2237,In_447,In_969);
and U2238 (N_2238,In_135,In_806);
and U2239 (N_2239,In_618,In_430);
or U2240 (N_2240,In_2226,In_1635);
nand U2241 (N_2241,In_577,In_712);
xnor U2242 (N_2242,In_1009,In_85);
nand U2243 (N_2243,In_1045,In_310);
or U2244 (N_2244,In_13,In_1872);
nand U2245 (N_2245,In_776,In_512);
or U2246 (N_2246,In_604,In_1192);
and U2247 (N_2247,In_344,In_1872);
or U2248 (N_2248,In_1721,In_1931);
nand U2249 (N_2249,In_856,In_2206);
nor U2250 (N_2250,In_1499,In_26);
nand U2251 (N_2251,In_895,In_2119);
nand U2252 (N_2252,In_800,In_797);
nand U2253 (N_2253,In_1584,In_684);
or U2254 (N_2254,In_1376,In_420);
nand U2255 (N_2255,In_1507,In_1850);
nand U2256 (N_2256,In_753,In_596);
xnor U2257 (N_2257,In_1008,In_405);
or U2258 (N_2258,In_641,In_1612);
and U2259 (N_2259,In_1005,In_1975);
nor U2260 (N_2260,In_1621,In_2116);
nor U2261 (N_2261,In_1280,In_2046);
nor U2262 (N_2262,In_1743,In_1642);
nand U2263 (N_2263,In_2281,In_1034);
or U2264 (N_2264,In_1418,In_1037);
nor U2265 (N_2265,In_640,In_1558);
nand U2266 (N_2266,In_1692,In_209);
nor U2267 (N_2267,In_1515,In_1152);
xnor U2268 (N_2268,In_1266,In_1063);
nand U2269 (N_2269,In_206,In_454);
nor U2270 (N_2270,In_294,In_150);
nor U2271 (N_2271,In_318,In_127);
nor U2272 (N_2272,In_694,In_1059);
nor U2273 (N_2273,In_1718,In_1447);
xor U2274 (N_2274,In_1811,In_2412);
nand U2275 (N_2275,In_2167,In_318);
nor U2276 (N_2276,In_2385,In_2474);
nand U2277 (N_2277,In_582,In_1761);
or U2278 (N_2278,In_992,In_236);
nor U2279 (N_2279,In_1644,In_440);
or U2280 (N_2280,In_2334,In_1876);
and U2281 (N_2281,In_741,In_412);
nand U2282 (N_2282,In_965,In_736);
nand U2283 (N_2283,In_1500,In_2336);
nand U2284 (N_2284,In_120,In_675);
or U2285 (N_2285,In_823,In_2003);
or U2286 (N_2286,In_1054,In_39);
nor U2287 (N_2287,In_1500,In_750);
and U2288 (N_2288,In_805,In_1232);
or U2289 (N_2289,In_479,In_1806);
or U2290 (N_2290,In_2379,In_590);
nor U2291 (N_2291,In_2436,In_1909);
nor U2292 (N_2292,In_96,In_1795);
and U2293 (N_2293,In_1532,In_2044);
and U2294 (N_2294,In_1556,In_1740);
and U2295 (N_2295,In_578,In_1863);
nand U2296 (N_2296,In_1289,In_544);
nand U2297 (N_2297,In_235,In_1270);
nor U2298 (N_2298,In_503,In_476);
nor U2299 (N_2299,In_602,In_1617);
nor U2300 (N_2300,In_1485,In_534);
or U2301 (N_2301,In_2038,In_809);
nand U2302 (N_2302,In_1719,In_404);
and U2303 (N_2303,In_1659,In_1845);
nor U2304 (N_2304,In_1671,In_2184);
nand U2305 (N_2305,In_314,In_814);
nor U2306 (N_2306,In_1356,In_1958);
nor U2307 (N_2307,In_692,In_667);
nand U2308 (N_2308,In_2220,In_1499);
or U2309 (N_2309,In_933,In_1390);
nand U2310 (N_2310,In_1563,In_1965);
or U2311 (N_2311,In_2079,In_191);
or U2312 (N_2312,In_1891,In_554);
nor U2313 (N_2313,In_838,In_2492);
nor U2314 (N_2314,In_324,In_430);
nand U2315 (N_2315,In_1179,In_1622);
nand U2316 (N_2316,In_52,In_1556);
and U2317 (N_2317,In_1513,In_709);
or U2318 (N_2318,In_281,In_926);
nand U2319 (N_2319,In_270,In_726);
and U2320 (N_2320,In_248,In_2024);
or U2321 (N_2321,In_1871,In_1138);
and U2322 (N_2322,In_2395,In_652);
nand U2323 (N_2323,In_2300,In_1750);
and U2324 (N_2324,In_724,In_797);
or U2325 (N_2325,In_2332,In_455);
or U2326 (N_2326,In_1118,In_2409);
xor U2327 (N_2327,In_317,In_2017);
or U2328 (N_2328,In_272,In_1724);
nor U2329 (N_2329,In_1557,In_2376);
or U2330 (N_2330,In_1627,In_648);
nor U2331 (N_2331,In_699,In_2478);
or U2332 (N_2332,In_2447,In_1422);
xnor U2333 (N_2333,In_871,In_998);
and U2334 (N_2334,In_1068,In_2166);
nor U2335 (N_2335,In_724,In_1545);
and U2336 (N_2336,In_968,In_1780);
nand U2337 (N_2337,In_1677,In_195);
and U2338 (N_2338,In_2457,In_1757);
and U2339 (N_2339,In_901,In_444);
nor U2340 (N_2340,In_583,In_265);
nand U2341 (N_2341,In_1984,In_364);
xor U2342 (N_2342,In_411,In_1148);
nor U2343 (N_2343,In_1075,In_1001);
and U2344 (N_2344,In_174,In_210);
nor U2345 (N_2345,In_1696,In_508);
nor U2346 (N_2346,In_2461,In_1363);
and U2347 (N_2347,In_450,In_1558);
or U2348 (N_2348,In_710,In_806);
nand U2349 (N_2349,In_372,In_2068);
or U2350 (N_2350,In_1853,In_1763);
and U2351 (N_2351,In_1288,In_2149);
or U2352 (N_2352,In_2449,In_737);
nand U2353 (N_2353,In_311,In_1404);
or U2354 (N_2354,In_635,In_1226);
and U2355 (N_2355,In_2353,In_1034);
or U2356 (N_2356,In_1121,In_1713);
nand U2357 (N_2357,In_139,In_912);
nand U2358 (N_2358,In_2002,In_42);
and U2359 (N_2359,In_1888,In_586);
nor U2360 (N_2360,In_2328,In_126);
nand U2361 (N_2361,In_820,In_352);
xor U2362 (N_2362,In_1795,In_1454);
and U2363 (N_2363,In_2390,In_816);
nor U2364 (N_2364,In_1240,In_1063);
or U2365 (N_2365,In_1865,In_2154);
nand U2366 (N_2366,In_1943,In_1855);
xor U2367 (N_2367,In_2023,In_1620);
nand U2368 (N_2368,In_417,In_1533);
or U2369 (N_2369,In_1840,In_779);
nand U2370 (N_2370,In_238,In_1819);
nand U2371 (N_2371,In_1556,In_1320);
or U2372 (N_2372,In_2125,In_1040);
or U2373 (N_2373,In_1511,In_1060);
or U2374 (N_2374,In_1111,In_1718);
and U2375 (N_2375,In_648,In_1312);
and U2376 (N_2376,In_2192,In_2392);
nor U2377 (N_2377,In_94,In_266);
nand U2378 (N_2378,In_390,In_386);
and U2379 (N_2379,In_2496,In_1331);
nand U2380 (N_2380,In_1373,In_1180);
or U2381 (N_2381,In_2314,In_1095);
nand U2382 (N_2382,In_549,In_557);
or U2383 (N_2383,In_2107,In_2098);
or U2384 (N_2384,In_1905,In_760);
nor U2385 (N_2385,In_487,In_1699);
nand U2386 (N_2386,In_2051,In_625);
nand U2387 (N_2387,In_949,In_1163);
nand U2388 (N_2388,In_1959,In_1090);
and U2389 (N_2389,In_383,In_2386);
nor U2390 (N_2390,In_235,In_1569);
nor U2391 (N_2391,In_672,In_1510);
nor U2392 (N_2392,In_89,In_348);
nor U2393 (N_2393,In_2462,In_2187);
nor U2394 (N_2394,In_524,In_1599);
or U2395 (N_2395,In_1235,In_1052);
or U2396 (N_2396,In_1775,In_1270);
nand U2397 (N_2397,In_316,In_1331);
or U2398 (N_2398,In_1427,In_1454);
or U2399 (N_2399,In_639,In_1043);
nor U2400 (N_2400,In_1330,In_576);
or U2401 (N_2401,In_1304,In_992);
nor U2402 (N_2402,In_1647,In_597);
nand U2403 (N_2403,In_2303,In_491);
nor U2404 (N_2404,In_55,In_1896);
nand U2405 (N_2405,In_697,In_1793);
or U2406 (N_2406,In_581,In_348);
xor U2407 (N_2407,In_2168,In_1502);
nand U2408 (N_2408,In_168,In_2098);
xnor U2409 (N_2409,In_855,In_165);
and U2410 (N_2410,In_776,In_1606);
and U2411 (N_2411,In_513,In_1166);
nand U2412 (N_2412,In_180,In_317);
nor U2413 (N_2413,In_859,In_967);
or U2414 (N_2414,In_1611,In_2283);
or U2415 (N_2415,In_1096,In_632);
and U2416 (N_2416,In_1459,In_693);
nor U2417 (N_2417,In_207,In_461);
xor U2418 (N_2418,In_2346,In_1665);
or U2419 (N_2419,In_984,In_286);
or U2420 (N_2420,In_782,In_1726);
and U2421 (N_2421,In_498,In_878);
and U2422 (N_2422,In_1312,In_619);
or U2423 (N_2423,In_1465,In_803);
nand U2424 (N_2424,In_2108,In_2354);
or U2425 (N_2425,In_2149,In_2104);
nand U2426 (N_2426,In_1748,In_131);
nand U2427 (N_2427,In_1433,In_2047);
and U2428 (N_2428,In_222,In_2399);
nor U2429 (N_2429,In_966,In_927);
and U2430 (N_2430,In_2104,In_2182);
and U2431 (N_2431,In_618,In_1977);
nor U2432 (N_2432,In_512,In_533);
nor U2433 (N_2433,In_1924,In_1588);
and U2434 (N_2434,In_329,In_254);
or U2435 (N_2435,In_1104,In_2224);
and U2436 (N_2436,In_2193,In_297);
or U2437 (N_2437,In_1309,In_1540);
or U2438 (N_2438,In_1360,In_1275);
or U2439 (N_2439,In_2219,In_1643);
or U2440 (N_2440,In_2290,In_1476);
and U2441 (N_2441,In_1347,In_1945);
nor U2442 (N_2442,In_1580,In_639);
nand U2443 (N_2443,In_2386,In_768);
nand U2444 (N_2444,In_743,In_475);
nor U2445 (N_2445,In_1281,In_969);
nand U2446 (N_2446,In_867,In_904);
nor U2447 (N_2447,In_1310,In_1598);
nor U2448 (N_2448,In_2070,In_905);
nor U2449 (N_2449,In_1450,In_830);
and U2450 (N_2450,In_2058,In_501);
nand U2451 (N_2451,In_2448,In_1191);
nor U2452 (N_2452,In_2447,In_1234);
and U2453 (N_2453,In_1019,In_1829);
and U2454 (N_2454,In_2268,In_1849);
nor U2455 (N_2455,In_529,In_206);
nor U2456 (N_2456,In_1564,In_319);
nand U2457 (N_2457,In_119,In_312);
nor U2458 (N_2458,In_1500,In_511);
nor U2459 (N_2459,In_1594,In_2142);
or U2460 (N_2460,In_917,In_1095);
nand U2461 (N_2461,In_1944,In_1375);
xor U2462 (N_2462,In_2012,In_410);
and U2463 (N_2463,In_2285,In_1524);
nor U2464 (N_2464,In_2195,In_501);
or U2465 (N_2465,In_358,In_555);
nand U2466 (N_2466,In_727,In_1233);
nor U2467 (N_2467,In_145,In_1314);
or U2468 (N_2468,In_1668,In_112);
nor U2469 (N_2469,In_2265,In_368);
nand U2470 (N_2470,In_2335,In_489);
or U2471 (N_2471,In_2099,In_1159);
or U2472 (N_2472,In_1381,In_1754);
nand U2473 (N_2473,In_2441,In_1848);
nor U2474 (N_2474,In_1929,In_104);
and U2475 (N_2475,In_415,In_2101);
nand U2476 (N_2476,In_2212,In_1149);
and U2477 (N_2477,In_405,In_453);
xor U2478 (N_2478,In_57,In_2208);
and U2479 (N_2479,In_866,In_306);
nand U2480 (N_2480,In_1178,In_2150);
nor U2481 (N_2481,In_1630,In_373);
nand U2482 (N_2482,In_1238,In_1589);
nand U2483 (N_2483,In_1397,In_1493);
and U2484 (N_2484,In_1070,In_118);
or U2485 (N_2485,In_2088,In_2400);
nor U2486 (N_2486,In_128,In_287);
nor U2487 (N_2487,In_1538,In_580);
nand U2488 (N_2488,In_1474,In_171);
or U2489 (N_2489,In_573,In_2378);
nor U2490 (N_2490,In_2130,In_1484);
and U2491 (N_2491,In_31,In_1081);
xnor U2492 (N_2492,In_2160,In_723);
nand U2493 (N_2493,In_2100,In_180);
nand U2494 (N_2494,In_1512,In_66);
nand U2495 (N_2495,In_2050,In_19);
nand U2496 (N_2496,In_2095,In_1041);
and U2497 (N_2497,In_1403,In_1679);
xnor U2498 (N_2498,In_807,In_66);
nor U2499 (N_2499,In_339,In_2153);
xor U2500 (N_2500,In_1547,In_2398);
or U2501 (N_2501,In_1810,In_1995);
nor U2502 (N_2502,In_837,In_472);
nor U2503 (N_2503,In_1724,In_2348);
nor U2504 (N_2504,In_1013,In_2291);
nor U2505 (N_2505,In_990,In_2290);
nor U2506 (N_2506,In_247,In_1167);
xor U2507 (N_2507,In_1439,In_2138);
or U2508 (N_2508,In_2442,In_1097);
nand U2509 (N_2509,In_871,In_2132);
nand U2510 (N_2510,In_1084,In_2389);
or U2511 (N_2511,In_1662,In_214);
or U2512 (N_2512,In_1415,In_1754);
or U2513 (N_2513,In_2177,In_95);
and U2514 (N_2514,In_644,In_865);
nor U2515 (N_2515,In_169,In_776);
nand U2516 (N_2516,In_1975,In_2473);
or U2517 (N_2517,In_703,In_1239);
and U2518 (N_2518,In_1763,In_701);
nand U2519 (N_2519,In_609,In_1101);
or U2520 (N_2520,In_1179,In_1094);
nor U2521 (N_2521,In_259,In_1680);
xnor U2522 (N_2522,In_1190,In_2086);
and U2523 (N_2523,In_370,In_1792);
xor U2524 (N_2524,In_926,In_1376);
nor U2525 (N_2525,In_453,In_125);
nand U2526 (N_2526,In_1783,In_274);
nor U2527 (N_2527,In_574,In_2183);
nor U2528 (N_2528,In_215,In_1499);
nor U2529 (N_2529,In_1398,In_1823);
and U2530 (N_2530,In_2414,In_2198);
nand U2531 (N_2531,In_1779,In_1967);
nand U2532 (N_2532,In_1857,In_1746);
or U2533 (N_2533,In_2327,In_1420);
xor U2534 (N_2534,In_2355,In_1261);
nand U2535 (N_2535,In_1078,In_1100);
or U2536 (N_2536,In_2114,In_1035);
nand U2537 (N_2537,In_1437,In_1993);
nor U2538 (N_2538,In_1588,In_2057);
nor U2539 (N_2539,In_1967,In_948);
or U2540 (N_2540,In_438,In_2014);
nor U2541 (N_2541,In_1676,In_1337);
or U2542 (N_2542,In_2470,In_1189);
nor U2543 (N_2543,In_634,In_1219);
xnor U2544 (N_2544,In_627,In_199);
nor U2545 (N_2545,In_2034,In_1914);
nand U2546 (N_2546,In_1023,In_1087);
nor U2547 (N_2547,In_164,In_1499);
and U2548 (N_2548,In_2166,In_1626);
nand U2549 (N_2549,In_199,In_206);
nor U2550 (N_2550,In_1980,In_1772);
or U2551 (N_2551,In_1131,In_1343);
or U2552 (N_2552,In_2345,In_1287);
or U2553 (N_2553,In_1355,In_952);
xnor U2554 (N_2554,In_363,In_1796);
and U2555 (N_2555,In_2396,In_1896);
xnor U2556 (N_2556,In_135,In_2219);
or U2557 (N_2557,In_349,In_1503);
or U2558 (N_2558,In_274,In_2487);
or U2559 (N_2559,In_602,In_710);
nor U2560 (N_2560,In_492,In_1561);
or U2561 (N_2561,In_1234,In_1646);
xor U2562 (N_2562,In_1253,In_1436);
nand U2563 (N_2563,In_355,In_240);
and U2564 (N_2564,In_1573,In_504);
or U2565 (N_2565,In_646,In_1818);
nor U2566 (N_2566,In_37,In_2292);
or U2567 (N_2567,In_581,In_1075);
nand U2568 (N_2568,In_1278,In_247);
nand U2569 (N_2569,In_337,In_1293);
xor U2570 (N_2570,In_438,In_1847);
and U2571 (N_2571,In_251,In_1233);
nand U2572 (N_2572,In_2031,In_2454);
nand U2573 (N_2573,In_1601,In_614);
or U2574 (N_2574,In_2180,In_1782);
xor U2575 (N_2575,In_564,In_42);
nor U2576 (N_2576,In_520,In_468);
and U2577 (N_2577,In_384,In_1071);
nand U2578 (N_2578,In_512,In_919);
and U2579 (N_2579,In_2373,In_2429);
xnor U2580 (N_2580,In_1525,In_1171);
and U2581 (N_2581,In_812,In_1123);
and U2582 (N_2582,In_599,In_1146);
nand U2583 (N_2583,In_1389,In_1797);
or U2584 (N_2584,In_1124,In_1396);
nor U2585 (N_2585,In_998,In_1511);
nand U2586 (N_2586,In_1970,In_849);
and U2587 (N_2587,In_105,In_64);
or U2588 (N_2588,In_1113,In_2006);
and U2589 (N_2589,In_419,In_326);
or U2590 (N_2590,In_22,In_874);
nand U2591 (N_2591,In_1348,In_38);
or U2592 (N_2592,In_892,In_2185);
nand U2593 (N_2593,In_1270,In_581);
nand U2594 (N_2594,In_1836,In_1705);
or U2595 (N_2595,In_1641,In_1544);
or U2596 (N_2596,In_956,In_1487);
or U2597 (N_2597,In_1483,In_1773);
or U2598 (N_2598,In_58,In_2388);
or U2599 (N_2599,In_1897,In_885);
nand U2600 (N_2600,In_1948,In_1739);
and U2601 (N_2601,In_1968,In_1460);
or U2602 (N_2602,In_1652,In_228);
nor U2603 (N_2603,In_1493,In_713);
and U2604 (N_2604,In_898,In_1725);
and U2605 (N_2605,In_594,In_1656);
and U2606 (N_2606,In_769,In_425);
or U2607 (N_2607,In_1301,In_290);
or U2608 (N_2608,In_1471,In_74);
xor U2609 (N_2609,In_1851,In_165);
and U2610 (N_2610,In_2412,In_2382);
and U2611 (N_2611,In_575,In_2308);
and U2612 (N_2612,In_1343,In_144);
and U2613 (N_2613,In_567,In_1382);
and U2614 (N_2614,In_759,In_1531);
nand U2615 (N_2615,In_768,In_1285);
nor U2616 (N_2616,In_1204,In_1297);
or U2617 (N_2617,In_1665,In_268);
nand U2618 (N_2618,In_462,In_1649);
nand U2619 (N_2619,In_1926,In_244);
and U2620 (N_2620,In_700,In_1985);
xnor U2621 (N_2621,In_413,In_567);
and U2622 (N_2622,In_1501,In_7);
nor U2623 (N_2623,In_157,In_1373);
and U2624 (N_2624,In_1431,In_1450);
and U2625 (N_2625,In_53,In_696);
and U2626 (N_2626,In_1431,In_275);
and U2627 (N_2627,In_298,In_2093);
and U2628 (N_2628,In_2367,In_882);
or U2629 (N_2629,In_1898,In_1060);
or U2630 (N_2630,In_1751,In_1690);
nor U2631 (N_2631,In_1840,In_2167);
xnor U2632 (N_2632,In_1085,In_1347);
or U2633 (N_2633,In_1974,In_1391);
or U2634 (N_2634,In_2079,In_2242);
and U2635 (N_2635,In_1456,In_1249);
nor U2636 (N_2636,In_2151,In_854);
or U2637 (N_2637,In_1576,In_2018);
nor U2638 (N_2638,In_1377,In_1967);
nor U2639 (N_2639,In_1486,In_147);
or U2640 (N_2640,In_1245,In_2483);
and U2641 (N_2641,In_645,In_2291);
and U2642 (N_2642,In_2454,In_1873);
or U2643 (N_2643,In_2116,In_2241);
nand U2644 (N_2644,In_1723,In_1795);
and U2645 (N_2645,In_2298,In_419);
or U2646 (N_2646,In_1058,In_501);
nand U2647 (N_2647,In_1059,In_2347);
nand U2648 (N_2648,In_1779,In_44);
and U2649 (N_2649,In_2344,In_1317);
nor U2650 (N_2650,In_381,In_145);
and U2651 (N_2651,In_2019,In_626);
nand U2652 (N_2652,In_1905,In_530);
and U2653 (N_2653,In_146,In_1451);
nand U2654 (N_2654,In_1713,In_497);
nor U2655 (N_2655,In_1444,In_596);
nor U2656 (N_2656,In_959,In_2024);
and U2657 (N_2657,In_127,In_1713);
xor U2658 (N_2658,In_659,In_2033);
nor U2659 (N_2659,In_1362,In_1488);
nand U2660 (N_2660,In_2400,In_2162);
xor U2661 (N_2661,In_804,In_379);
nor U2662 (N_2662,In_1202,In_2424);
or U2663 (N_2663,In_2299,In_924);
or U2664 (N_2664,In_645,In_2005);
nand U2665 (N_2665,In_2306,In_1428);
nor U2666 (N_2666,In_195,In_2384);
xnor U2667 (N_2667,In_416,In_2473);
or U2668 (N_2668,In_247,In_1486);
nand U2669 (N_2669,In_339,In_1508);
nor U2670 (N_2670,In_830,In_779);
xor U2671 (N_2671,In_112,In_760);
nor U2672 (N_2672,In_2069,In_1882);
nand U2673 (N_2673,In_1061,In_916);
nor U2674 (N_2674,In_1553,In_2224);
or U2675 (N_2675,In_1285,In_938);
nand U2676 (N_2676,In_2362,In_154);
nand U2677 (N_2677,In_1919,In_1129);
nand U2678 (N_2678,In_720,In_1725);
xor U2679 (N_2679,In_2324,In_750);
and U2680 (N_2680,In_1559,In_1256);
nand U2681 (N_2681,In_818,In_1122);
xnor U2682 (N_2682,In_2019,In_1401);
xnor U2683 (N_2683,In_2306,In_576);
nand U2684 (N_2684,In_1498,In_1697);
nand U2685 (N_2685,In_131,In_597);
nor U2686 (N_2686,In_2257,In_1123);
and U2687 (N_2687,In_2238,In_1804);
xnor U2688 (N_2688,In_2448,In_319);
or U2689 (N_2689,In_813,In_1171);
and U2690 (N_2690,In_823,In_739);
nand U2691 (N_2691,In_1394,In_186);
and U2692 (N_2692,In_1392,In_888);
nand U2693 (N_2693,In_1916,In_577);
nor U2694 (N_2694,In_1050,In_445);
or U2695 (N_2695,In_10,In_1398);
and U2696 (N_2696,In_585,In_403);
or U2697 (N_2697,In_2485,In_54);
and U2698 (N_2698,In_2289,In_913);
nand U2699 (N_2699,In_2182,In_614);
nor U2700 (N_2700,In_2488,In_2457);
and U2701 (N_2701,In_1322,In_1406);
and U2702 (N_2702,In_1364,In_2419);
or U2703 (N_2703,In_2026,In_888);
xnor U2704 (N_2704,In_929,In_2297);
nor U2705 (N_2705,In_1713,In_1374);
nand U2706 (N_2706,In_2347,In_1508);
nand U2707 (N_2707,In_1364,In_361);
and U2708 (N_2708,In_413,In_36);
nor U2709 (N_2709,In_1319,In_95);
nand U2710 (N_2710,In_1085,In_1288);
nand U2711 (N_2711,In_2294,In_66);
nand U2712 (N_2712,In_2452,In_1805);
nor U2713 (N_2713,In_2246,In_2014);
nor U2714 (N_2714,In_1895,In_352);
nor U2715 (N_2715,In_1373,In_782);
nand U2716 (N_2716,In_479,In_1535);
or U2717 (N_2717,In_1695,In_1183);
nor U2718 (N_2718,In_1237,In_445);
nand U2719 (N_2719,In_920,In_335);
nand U2720 (N_2720,In_1798,In_1138);
nand U2721 (N_2721,In_1825,In_2195);
xnor U2722 (N_2722,In_1313,In_393);
or U2723 (N_2723,In_612,In_337);
nand U2724 (N_2724,In_166,In_763);
nand U2725 (N_2725,In_1526,In_2458);
nor U2726 (N_2726,In_1610,In_1687);
nand U2727 (N_2727,In_2220,In_700);
or U2728 (N_2728,In_2334,In_53);
or U2729 (N_2729,In_1720,In_1445);
nor U2730 (N_2730,In_479,In_1456);
nand U2731 (N_2731,In_497,In_1439);
or U2732 (N_2732,In_1106,In_972);
or U2733 (N_2733,In_1662,In_1172);
xnor U2734 (N_2734,In_824,In_209);
or U2735 (N_2735,In_90,In_1283);
nand U2736 (N_2736,In_633,In_342);
nand U2737 (N_2737,In_1680,In_1687);
and U2738 (N_2738,In_173,In_1437);
nand U2739 (N_2739,In_1641,In_675);
nor U2740 (N_2740,In_2412,In_1144);
nor U2741 (N_2741,In_171,In_550);
xnor U2742 (N_2742,In_2074,In_20);
nor U2743 (N_2743,In_244,In_1495);
and U2744 (N_2744,In_1790,In_2234);
nor U2745 (N_2745,In_1366,In_787);
nand U2746 (N_2746,In_588,In_1896);
nor U2747 (N_2747,In_2263,In_1274);
nand U2748 (N_2748,In_52,In_325);
nand U2749 (N_2749,In_294,In_1766);
xnor U2750 (N_2750,In_1909,In_1614);
or U2751 (N_2751,In_983,In_166);
nor U2752 (N_2752,In_712,In_1010);
nand U2753 (N_2753,In_293,In_2192);
or U2754 (N_2754,In_1699,In_901);
nand U2755 (N_2755,In_345,In_517);
nand U2756 (N_2756,In_2477,In_1309);
and U2757 (N_2757,In_770,In_1684);
nand U2758 (N_2758,In_424,In_2027);
or U2759 (N_2759,In_2047,In_2234);
nor U2760 (N_2760,In_1355,In_544);
nor U2761 (N_2761,In_1026,In_762);
nand U2762 (N_2762,In_1703,In_1423);
and U2763 (N_2763,In_539,In_1609);
or U2764 (N_2764,In_2060,In_282);
nor U2765 (N_2765,In_2025,In_1195);
nand U2766 (N_2766,In_1326,In_1588);
nor U2767 (N_2767,In_2486,In_1641);
nor U2768 (N_2768,In_1567,In_308);
and U2769 (N_2769,In_246,In_1634);
or U2770 (N_2770,In_487,In_765);
or U2771 (N_2771,In_1850,In_1729);
or U2772 (N_2772,In_1283,In_273);
nor U2773 (N_2773,In_111,In_2421);
nand U2774 (N_2774,In_289,In_702);
nand U2775 (N_2775,In_1997,In_1381);
or U2776 (N_2776,In_447,In_1450);
and U2777 (N_2777,In_2286,In_1047);
nor U2778 (N_2778,In_187,In_1792);
and U2779 (N_2779,In_1614,In_1541);
and U2780 (N_2780,In_1731,In_2291);
nand U2781 (N_2781,In_1380,In_146);
nor U2782 (N_2782,In_1247,In_1184);
and U2783 (N_2783,In_356,In_151);
or U2784 (N_2784,In_435,In_276);
and U2785 (N_2785,In_1243,In_2348);
nand U2786 (N_2786,In_319,In_1100);
and U2787 (N_2787,In_1800,In_39);
or U2788 (N_2788,In_1932,In_706);
nor U2789 (N_2789,In_478,In_1686);
or U2790 (N_2790,In_2272,In_360);
or U2791 (N_2791,In_1243,In_519);
nand U2792 (N_2792,In_1052,In_1185);
nor U2793 (N_2793,In_66,In_1262);
or U2794 (N_2794,In_876,In_1242);
nand U2795 (N_2795,In_457,In_1482);
and U2796 (N_2796,In_1924,In_706);
or U2797 (N_2797,In_166,In_796);
nand U2798 (N_2798,In_2097,In_1342);
nand U2799 (N_2799,In_827,In_972);
nand U2800 (N_2800,In_467,In_1738);
nor U2801 (N_2801,In_454,In_1943);
and U2802 (N_2802,In_1269,In_247);
and U2803 (N_2803,In_1493,In_2270);
nor U2804 (N_2804,In_2029,In_1383);
nor U2805 (N_2805,In_1447,In_1023);
and U2806 (N_2806,In_1324,In_806);
and U2807 (N_2807,In_713,In_951);
or U2808 (N_2808,In_653,In_25);
and U2809 (N_2809,In_2147,In_117);
xnor U2810 (N_2810,In_1893,In_1434);
nor U2811 (N_2811,In_1510,In_980);
and U2812 (N_2812,In_1361,In_1664);
nand U2813 (N_2813,In_2499,In_986);
nor U2814 (N_2814,In_986,In_1645);
or U2815 (N_2815,In_920,In_66);
nand U2816 (N_2816,In_2021,In_2203);
nor U2817 (N_2817,In_247,In_293);
and U2818 (N_2818,In_461,In_2113);
or U2819 (N_2819,In_1020,In_2156);
nand U2820 (N_2820,In_148,In_94);
or U2821 (N_2821,In_525,In_1307);
nor U2822 (N_2822,In_887,In_2265);
nand U2823 (N_2823,In_720,In_2);
or U2824 (N_2824,In_547,In_1575);
nand U2825 (N_2825,In_2248,In_2164);
or U2826 (N_2826,In_2423,In_1450);
nand U2827 (N_2827,In_730,In_765);
or U2828 (N_2828,In_2099,In_1560);
or U2829 (N_2829,In_120,In_1046);
or U2830 (N_2830,In_1149,In_69);
or U2831 (N_2831,In_1330,In_1361);
nor U2832 (N_2832,In_697,In_94);
and U2833 (N_2833,In_2177,In_1300);
and U2834 (N_2834,In_202,In_98);
and U2835 (N_2835,In_434,In_349);
nor U2836 (N_2836,In_955,In_1843);
and U2837 (N_2837,In_2042,In_671);
nor U2838 (N_2838,In_1839,In_186);
nor U2839 (N_2839,In_1744,In_2169);
and U2840 (N_2840,In_2272,In_1535);
nor U2841 (N_2841,In_893,In_2103);
and U2842 (N_2842,In_1836,In_77);
and U2843 (N_2843,In_1423,In_2064);
and U2844 (N_2844,In_1201,In_1245);
nor U2845 (N_2845,In_854,In_1066);
and U2846 (N_2846,In_438,In_618);
or U2847 (N_2847,In_1557,In_1468);
and U2848 (N_2848,In_424,In_2262);
nor U2849 (N_2849,In_2498,In_32);
xnor U2850 (N_2850,In_2425,In_975);
xnor U2851 (N_2851,In_2297,In_976);
xnor U2852 (N_2852,In_1248,In_392);
nor U2853 (N_2853,In_1807,In_1585);
nand U2854 (N_2854,In_1388,In_2182);
or U2855 (N_2855,In_994,In_2138);
nor U2856 (N_2856,In_2357,In_112);
nand U2857 (N_2857,In_2433,In_1614);
xor U2858 (N_2858,In_1271,In_1558);
nand U2859 (N_2859,In_547,In_1472);
nand U2860 (N_2860,In_855,In_2419);
nand U2861 (N_2861,In_2086,In_1001);
or U2862 (N_2862,In_383,In_1230);
nand U2863 (N_2863,In_2046,In_822);
nand U2864 (N_2864,In_1626,In_2202);
and U2865 (N_2865,In_987,In_2493);
nor U2866 (N_2866,In_1922,In_1255);
and U2867 (N_2867,In_675,In_1596);
and U2868 (N_2868,In_1361,In_1095);
nor U2869 (N_2869,In_1655,In_2016);
or U2870 (N_2870,In_911,In_2289);
and U2871 (N_2871,In_585,In_416);
nand U2872 (N_2872,In_1550,In_1290);
nand U2873 (N_2873,In_740,In_2136);
nor U2874 (N_2874,In_874,In_2309);
or U2875 (N_2875,In_2029,In_2261);
and U2876 (N_2876,In_613,In_706);
nor U2877 (N_2877,In_1403,In_375);
or U2878 (N_2878,In_1481,In_465);
nand U2879 (N_2879,In_1605,In_1417);
xor U2880 (N_2880,In_1832,In_442);
and U2881 (N_2881,In_471,In_1548);
nor U2882 (N_2882,In_1893,In_1757);
nor U2883 (N_2883,In_1702,In_1915);
xor U2884 (N_2884,In_856,In_1316);
nor U2885 (N_2885,In_466,In_2305);
and U2886 (N_2886,In_559,In_179);
or U2887 (N_2887,In_779,In_1902);
nor U2888 (N_2888,In_1037,In_729);
nand U2889 (N_2889,In_2329,In_1929);
nand U2890 (N_2890,In_506,In_2060);
nor U2891 (N_2891,In_1538,In_1490);
and U2892 (N_2892,In_1410,In_1988);
and U2893 (N_2893,In_378,In_1591);
or U2894 (N_2894,In_188,In_2096);
nand U2895 (N_2895,In_1218,In_250);
and U2896 (N_2896,In_2193,In_2383);
nand U2897 (N_2897,In_481,In_175);
nand U2898 (N_2898,In_898,In_2370);
and U2899 (N_2899,In_455,In_1270);
nor U2900 (N_2900,In_401,In_1128);
nor U2901 (N_2901,In_1726,In_1761);
nor U2902 (N_2902,In_2099,In_503);
nand U2903 (N_2903,In_2117,In_1457);
or U2904 (N_2904,In_1017,In_1685);
or U2905 (N_2905,In_938,In_1192);
nand U2906 (N_2906,In_110,In_1081);
and U2907 (N_2907,In_2347,In_721);
and U2908 (N_2908,In_193,In_1709);
or U2909 (N_2909,In_802,In_1259);
nand U2910 (N_2910,In_128,In_2156);
nand U2911 (N_2911,In_230,In_2151);
nor U2912 (N_2912,In_2095,In_2105);
or U2913 (N_2913,In_570,In_1682);
xnor U2914 (N_2914,In_814,In_1330);
and U2915 (N_2915,In_1388,In_1091);
or U2916 (N_2916,In_1001,In_975);
nand U2917 (N_2917,In_1971,In_646);
nor U2918 (N_2918,In_208,In_576);
nor U2919 (N_2919,In_73,In_768);
nand U2920 (N_2920,In_1076,In_2108);
and U2921 (N_2921,In_2316,In_1626);
or U2922 (N_2922,In_300,In_272);
nor U2923 (N_2923,In_1303,In_283);
and U2924 (N_2924,In_994,In_2390);
or U2925 (N_2925,In_907,In_1640);
and U2926 (N_2926,In_1992,In_2454);
xor U2927 (N_2927,In_456,In_353);
nor U2928 (N_2928,In_43,In_2346);
nand U2929 (N_2929,In_2222,In_1093);
and U2930 (N_2930,In_1911,In_904);
nor U2931 (N_2931,In_1527,In_484);
and U2932 (N_2932,In_2124,In_296);
and U2933 (N_2933,In_1066,In_180);
nand U2934 (N_2934,In_479,In_1115);
and U2935 (N_2935,In_2209,In_2415);
nor U2936 (N_2936,In_2131,In_1838);
and U2937 (N_2937,In_649,In_1958);
or U2938 (N_2938,In_1653,In_180);
or U2939 (N_2939,In_348,In_1279);
nand U2940 (N_2940,In_1129,In_299);
nand U2941 (N_2941,In_1739,In_1879);
nand U2942 (N_2942,In_520,In_1000);
xor U2943 (N_2943,In_1386,In_2395);
nand U2944 (N_2944,In_839,In_1231);
and U2945 (N_2945,In_2007,In_1639);
nand U2946 (N_2946,In_258,In_2409);
and U2947 (N_2947,In_1581,In_1001);
nor U2948 (N_2948,In_55,In_1219);
nand U2949 (N_2949,In_2449,In_1522);
nand U2950 (N_2950,In_624,In_1587);
xnor U2951 (N_2951,In_876,In_825);
or U2952 (N_2952,In_998,In_1513);
nand U2953 (N_2953,In_1034,In_207);
or U2954 (N_2954,In_746,In_2101);
nor U2955 (N_2955,In_1977,In_1970);
and U2956 (N_2956,In_1984,In_2055);
or U2957 (N_2957,In_21,In_1879);
or U2958 (N_2958,In_1600,In_1514);
nor U2959 (N_2959,In_1222,In_581);
or U2960 (N_2960,In_662,In_2359);
or U2961 (N_2961,In_2442,In_90);
nor U2962 (N_2962,In_2186,In_1858);
nor U2963 (N_2963,In_1541,In_1873);
xor U2964 (N_2964,In_783,In_2396);
xor U2965 (N_2965,In_1595,In_994);
or U2966 (N_2966,In_694,In_2395);
nand U2967 (N_2967,In_1832,In_47);
or U2968 (N_2968,In_1717,In_2271);
and U2969 (N_2969,In_2115,In_2395);
nand U2970 (N_2970,In_1819,In_2077);
or U2971 (N_2971,In_1331,In_380);
or U2972 (N_2972,In_493,In_651);
xor U2973 (N_2973,In_950,In_1527);
nand U2974 (N_2974,In_253,In_2110);
nor U2975 (N_2975,In_1504,In_197);
nand U2976 (N_2976,In_1246,In_1214);
and U2977 (N_2977,In_1914,In_477);
and U2978 (N_2978,In_425,In_296);
or U2979 (N_2979,In_2382,In_2185);
and U2980 (N_2980,In_2491,In_327);
nor U2981 (N_2981,In_1524,In_603);
and U2982 (N_2982,In_540,In_642);
nor U2983 (N_2983,In_1553,In_1629);
and U2984 (N_2984,In_1939,In_552);
and U2985 (N_2985,In_2464,In_446);
or U2986 (N_2986,In_1084,In_81);
nand U2987 (N_2987,In_2105,In_1496);
nor U2988 (N_2988,In_1795,In_1290);
and U2989 (N_2989,In_1320,In_735);
nor U2990 (N_2990,In_951,In_789);
xor U2991 (N_2991,In_1542,In_97);
or U2992 (N_2992,In_899,In_740);
nand U2993 (N_2993,In_302,In_2130);
and U2994 (N_2994,In_1722,In_2030);
nand U2995 (N_2995,In_1761,In_2027);
or U2996 (N_2996,In_2210,In_212);
nor U2997 (N_2997,In_445,In_1748);
nor U2998 (N_2998,In_125,In_1103);
nor U2999 (N_2999,In_1159,In_2429);
nand U3000 (N_3000,In_1137,In_2239);
or U3001 (N_3001,In_2050,In_2055);
nand U3002 (N_3002,In_1856,In_1499);
nand U3003 (N_3003,In_767,In_2125);
xnor U3004 (N_3004,In_249,In_1352);
and U3005 (N_3005,In_841,In_996);
or U3006 (N_3006,In_1275,In_857);
or U3007 (N_3007,In_745,In_353);
nand U3008 (N_3008,In_505,In_1156);
nor U3009 (N_3009,In_2031,In_1720);
nor U3010 (N_3010,In_90,In_609);
nor U3011 (N_3011,In_1919,In_982);
nor U3012 (N_3012,In_600,In_262);
nor U3013 (N_3013,In_356,In_930);
nand U3014 (N_3014,In_71,In_1949);
and U3015 (N_3015,In_1473,In_454);
xor U3016 (N_3016,In_92,In_1190);
nor U3017 (N_3017,In_2219,In_1507);
and U3018 (N_3018,In_2208,In_2246);
nor U3019 (N_3019,In_1787,In_558);
xnor U3020 (N_3020,In_399,In_665);
nor U3021 (N_3021,In_40,In_145);
or U3022 (N_3022,In_892,In_2056);
and U3023 (N_3023,In_1598,In_1826);
nor U3024 (N_3024,In_126,In_1117);
nor U3025 (N_3025,In_539,In_2075);
and U3026 (N_3026,In_1495,In_583);
nand U3027 (N_3027,In_270,In_1315);
nor U3028 (N_3028,In_1924,In_2281);
nor U3029 (N_3029,In_719,In_1253);
or U3030 (N_3030,In_1581,In_1168);
and U3031 (N_3031,In_159,In_1036);
xnor U3032 (N_3032,In_1789,In_1715);
nor U3033 (N_3033,In_2359,In_788);
or U3034 (N_3034,In_2430,In_2482);
or U3035 (N_3035,In_1414,In_2106);
nor U3036 (N_3036,In_2170,In_2473);
nor U3037 (N_3037,In_311,In_1599);
and U3038 (N_3038,In_1765,In_1725);
and U3039 (N_3039,In_341,In_519);
or U3040 (N_3040,In_2480,In_2378);
nor U3041 (N_3041,In_848,In_432);
and U3042 (N_3042,In_569,In_172);
or U3043 (N_3043,In_1093,In_2220);
nor U3044 (N_3044,In_1157,In_2360);
nand U3045 (N_3045,In_1149,In_1851);
or U3046 (N_3046,In_1982,In_1820);
and U3047 (N_3047,In_2205,In_2379);
nor U3048 (N_3048,In_248,In_657);
nor U3049 (N_3049,In_2324,In_1488);
nand U3050 (N_3050,In_1610,In_991);
nand U3051 (N_3051,In_1249,In_740);
and U3052 (N_3052,In_1097,In_1778);
xnor U3053 (N_3053,In_1470,In_2372);
or U3054 (N_3054,In_1700,In_470);
or U3055 (N_3055,In_420,In_1439);
xor U3056 (N_3056,In_2163,In_1664);
nor U3057 (N_3057,In_1876,In_819);
nand U3058 (N_3058,In_2326,In_2257);
nor U3059 (N_3059,In_414,In_2020);
and U3060 (N_3060,In_182,In_223);
or U3061 (N_3061,In_414,In_1154);
nor U3062 (N_3062,In_485,In_1141);
and U3063 (N_3063,In_1017,In_2394);
and U3064 (N_3064,In_2146,In_1098);
nor U3065 (N_3065,In_2082,In_1701);
nand U3066 (N_3066,In_2351,In_183);
nor U3067 (N_3067,In_176,In_242);
and U3068 (N_3068,In_211,In_2436);
nor U3069 (N_3069,In_764,In_2039);
nand U3070 (N_3070,In_748,In_1799);
or U3071 (N_3071,In_261,In_1151);
or U3072 (N_3072,In_920,In_2213);
or U3073 (N_3073,In_966,In_1908);
xor U3074 (N_3074,In_828,In_1578);
and U3075 (N_3075,In_1915,In_47);
xnor U3076 (N_3076,In_2327,In_126);
and U3077 (N_3077,In_2344,In_2267);
xor U3078 (N_3078,In_673,In_563);
or U3079 (N_3079,In_539,In_25);
nand U3080 (N_3080,In_2202,In_1718);
nor U3081 (N_3081,In_1226,In_1403);
and U3082 (N_3082,In_46,In_441);
and U3083 (N_3083,In_1626,In_2011);
xnor U3084 (N_3084,In_564,In_1508);
and U3085 (N_3085,In_887,In_547);
and U3086 (N_3086,In_556,In_2025);
nor U3087 (N_3087,In_85,In_2073);
nand U3088 (N_3088,In_1599,In_1151);
or U3089 (N_3089,In_201,In_647);
nand U3090 (N_3090,In_378,In_1221);
and U3091 (N_3091,In_1510,In_1645);
or U3092 (N_3092,In_995,In_1187);
xnor U3093 (N_3093,In_1213,In_478);
or U3094 (N_3094,In_985,In_2053);
nand U3095 (N_3095,In_2361,In_1657);
or U3096 (N_3096,In_1412,In_1732);
and U3097 (N_3097,In_504,In_2422);
nand U3098 (N_3098,In_32,In_303);
xor U3099 (N_3099,In_1780,In_2222);
xor U3100 (N_3100,In_2112,In_2380);
xnor U3101 (N_3101,In_1895,In_467);
or U3102 (N_3102,In_615,In_724);
xor U3103 (N_3103,In_2089,In_50);
nand U3104 (N_3104,In_1499,In_1287);
or U3105 (N_3105,In_999,In_114);
nand U3106 (N_3106,In_2332,In_806);
or U3107 (N_3107,In_234,In_169);
and U3108 (N_3108,In_1808,In_2359);
and U3109 (N_3109,In_1820,In_2142);
nor U3110 (N_3110,In_1724,In_1667);
nand U3111 (N_3111,In_708,In_2456);
nor U3112 (N_3112,In_352,In_1890);
or U3113 (N_3113,In_696,In_1924);
and U3114 (N_3114,In_314,In_83);
nor U3115 (N_3115,In_1907,In_195);
nor U3116 (N_3116,In_1079,In_1210);
or U3117 (N_3117,In_1217,In_196);
or U3118 (N_3118,In_787,In_1452);
or U3119 (N_3119,In_756,In_1236);
nand U3120 (N_3120,In_973,In_2480);
and U3121 (N_3121,In_1300,In_1033);
or U3122 (N_3122,In_880,In_969);
and U3123 (N_3123,In_745,In_872);
nor U3124 (N_3124,In_323,In_1757);
nand U3125 (N_3125,In_677,In_418);
nand U3126 (N_3126,In_1151,In_286);
nor U3127 (N_3127,In_14,In_2344);
nor U3128 (N_3128,In_796,In_1991);
and U3129 (N_3129,In_2173,In_2452);
xor U3130 (N_3130,In_1970,In_414);
nor U3131 (N_3131,In_871,In_402);
nand U3132 (N_3132,In_58,In_1257);
nor U3133 (N_3133,In_1994,In_1500);
nor U3134 (N_3134,In_1467,In_444);
or U3135 (N_3135,In_1770,In_1466);
nor U3136 (N_3136,In_1151,In_2494);
nor U3137 (N_3137,In_1989,In_1061);
and U3138 (N_3138,In_501,In_1403);
and U3139 (N_3139,In_944,In_1994);
or U3140 (N_3140,In_2382,In_159);
and U3141 (N_3141,In_1417,In_2218);
nand U3142 (N_3142,In_739,In_295);
nor U3143 (N_3143,In_1251,In_1413);
nor U3144 (N_3144,In_942,In_825);
nor U3145 (N_3145,In_1585,In_1984);
or U3146 (N_3146,In_1818,In_802);
and U3147 (N_3147,In_1158,In_802);
nor U3148 (N_3148,In_745,In_1844);
nor U3149 (N_3149,In_1313,In_2140);
and U3150 (N_3150,In_296,In_1638);
nor U3151 (N_3151,In_398,In_1902);
nand U3152 (N_3152,In_1584,In_1105);
nand U3153 (N_3153,In_103,In_25);
nor U3154 (N_3154,In_1959,In_1821);
nor U3155 (N_3155,In_1331,In_2095);
nor U3156 (N_3156,In_929,In_1406);
nand U3157 (N_3157,In_65,In_2453);
or U3158 (N_3158,In_1650,In_211);
and U3159 (N_3159,In_642,In_1167);
nand U3160 (N_3160,In_808,In_1492);
and U3161 (N_3161,In_1732,In_2303);
and U3162 (N_3162,In_2117,In_1152);
and U3163 (N_3163,In_235,In_462);
xor U3164 (N_3164,In_1968,In_532);
or U3165 (N_3165,In_1227,In_1985);
and U3166 (N_3166,In_2175,In_757);
and U3167 (N_3167,In_1420,In_425);
or U3168 (N_3168,In_2498,In_323);
or U3169 (N_3169,In_554,In_918);
or U3170 (N_3170,In_944,In_718);
xor U3171 (N_3171,In_1273,In_831);
and U3172 (N_3172,In_2366,In_2104);
nor U3173 (N_3173,In_503,In_1933);
or U3174 (N_3174,In_3,In_115);
xor U3175 (N_3175,In_382,In_474);
nor U3176 (N_3176,In_512,In_158);
nor U3177 (N_3177,In_2024,In_174);
xnor U3178 (N_3178,In_378,In_207);
nand U3179 (N_3179,In_902,In_406);
nor U3180 (N_3180,In_1263,In_2363);
xnor U3181 (N_3181,In_2468,In_945);
or U3182 (N_3182,In_648,In_2361);
nor U3183 (N_3183,In_666,In_2395);
nor U3184 (N_3184,In_1677,In_456);
nand U3185 (N_3185,In_1873,In_1105);
or U3186 (N_3186,In_1302,In_2344);
nand U3187 (N_3187,In_827,In_749);
nor U3188 (N_3188,In_1803,In_1760);
and U3189 (N_3189,In_2388,In_397);
nand U3190 (N_3190,In_97,In_668);
and U3191 (N_3191,In_502,In_464);
or U3192 (N_3192,In_1855,In_1287);
nor U3193 (N_3193,In_1963,In_2463);
nor U3194 (N_3194,In_1770,In_2424);
nand U3195 (N_3195,In_972,In_1131);
and U3196 (N_3196,In_677,In_504);
nand U3197 (N_3197,In_2298,In_1949);
nand U3198 (N_3198,In_2125,In_1333);
and U3199 (N_3199,In_967,In_2295);
and U3200 (N_3200,In_121,In_96);
nor U3201 (N_3201,In_1415,In_2189);
nand U3202 (N_3202,In_1633,In_1947);
and U3203 (N_3203,In_1991,In_576);
nand U3204 (N_3204,In_1541,In_916);
or U3205 (N_3205,In_1615,In_668);
xnor U3206 (N_3206,In_1178,In_1415);
and U3207 (N_3207,In_2216,In_2107);
nand U3208 (N_3208,In_194,In_1326);
and U3209 (N_3209,In_2181,In_443);
nor U3210 (N_3210,In_140,In_157);
and U3211 (N_3211,In_940,In_1623);
nand U3212 (N_3212,In_789,In_2289);
and U3213 (N_3213,In_2214,In_695);
or U3214 (N_3214,In_2099,In_1026);
nor U3215 (N_3215,In_1260,In_2257);
xnor U3216 (N_3216,In_689,In_2302);
and U3217 (N_3217,In_307,In_1625);
or U3218 (N_3218,In_1647,In_232);
and U3219 (N_3219,In_1203,In_796);
and U3220 (N_3220,In_584,In_1911);
nand U3221 (N_3221,In_1959,In_1951);
nand U3222 (N_3222,In_590,In_582);
or U3223 (N_3223,In_76,In_1336);
nor U3224 (N_3224,In_1207,In_1160);
and U3225 (N_3225,In_1587,In_1143);
or U3226 (N_3226,In_2043,In_1163);
or U3227 (N_3227,In_2141,In_1971);
and U3228 (N_3228,In_646,In_148);
nand U3229 (N_3229,In_2049,In_153);
and U3230 (N_3230,In_2148,In_2477);
and U3231 (N_3231,In_2048,In_1982);
nor U3232 (N_3232,In_1315,In_1933);
xor U3233 (N_3233,In_684,In_17);
and U3234 (N_3234,In_1567,In_2142);
nor U3235 (N_3235,In_772,In_1982);
nand U3236 (N_3236,In_1916,In_1402);
nor U3237 (N_3237,In_909,In_1649);
nand U3238 (N_3238,In_148,In_1957);
xor U3239 (N_3239,In_1019,In_485);
nor U3240 (N_3240,In_859,In_140);
and U3241 (N_3241,In_1534,In_182);
nor U3242 (N_3242,In_1587,In_2451);
nor U3243 (N_3243,In_968,In_333);
and U3244 (N_3244,In_1469,In_1350);
and U3245 (N_3245,In_2405,In_2410);
nor U3246 (N_3246,In_262,In_565);
nor U3247 (N_3247,In_2493,In_1002);
or U3248 (N_3248,In_1879,In_1893);
nand U3249 (N_3249,In_1370,In_1972);
nor U3250 (N_3250,In_1515,In_2062);
and U3251 (N_3251,In_1731,In_605);
or U3252 (N_3252,In_858,In_529);
nand U3253 (N_3253,In_1415,In_1796);
and U3254 (N_3254,In_2388,In_264);
nand U3255 (N_3255,In_722,In_1687);
or U3256 (N_3256,In_2260,In_561);
and U3257 (N_3257,In_2222,In_797);
nand U3258 (N_3258,In_120,In_462);
and U3259 (N_3259,In_28,In_1559);
and U3260 (N_3260,In_1446,In_1529);
nand U3261 (N_3261,In_56,In_2119);
and U3262 (N_3262,In_408,In_2331);
and U3263 (N_3263,In_438,In_2475);
and U3264 (N_3264,In_1387,In_233);
or U3265 (N_3265,In_444,In_1842);
and U3266 (N_3266,In_813,In_1274);
nor U3267 (N_3267,In_112,In_1328);
and U3268 (N_3268,In_2063,In_1417);
nor U3269 (N_3269,In_1180,In_1670);
nor U3270 (N_3270,In_1915,In_1786);
nand U3271 (N_3271,In_872,In_1868);
nor U3272 (N_3272,In_1077,In_1086);
nand U3273 (N_3273,In_2073,In_746);
and U3274 (N_3274,In_394,In_1577);
nand U3275 (N_3275,In_1242,In_1290);
and U3276 (N_3276,In_787,In_2456);
nand U3277 (N_3277,In_1530,In_550);
nor U3278 (N_3278,In_1087,In_16);
or U3279 (N_3279,In_713,In_278);
nand U3280 (N_3280,In_1436,In_2498);
nand U3281 (N_3281,In_1213,In_2109);
or U3282 (N_3282,In_438,In_1061);
nor U3283 (N_3283,In_1533,In_1306);
and U3284 (N_3284,In_82,In_793);
nor U3285 (N_3285,In_943,In_1365);
or U3286 (N_3286,In_994,In_1243);
nor U3287 (N_3287,In_1041,In_1460);
nor U3288 (N_3288,In_250,In_297);
xnor U3289 (N_3289,In_2106,In_1598);
and U3290 (N_3290,In_1217,In_1762);
nor U3291 (N_3291,In_2058,In_142);
or U3292 (N_3292,In_2316,In_2074);
and U3293 (N_3293,In_877,In_2272);
nor U3294 (N_3294,In_1425,In_1822);
nor U3295 (N_3295,In_960,In_2293);
and U3296 (N_3296,In_254,In_1798);
and U3297 (N_3297,In_2031,In_2310);
or U3298 (N_3298,In_1371,In_397);
or U3299 (N_3299,In_2189,In_688);
or U3300 (N_3300,In_2450,In_1941);
or U3301 (N_3301,In_2075,In_1817);
or U3302 (N_3302,In_172,In_2419);
and U3303 (N_3303,In_1936,In_1573);
and U3304 (N_3304,In_889,In_201);
or U3305 (N_3305,In_847,In_1662);
nand U3306 (N_3306,In_277,In_317);
and U3307 (N_3307,In_2392,In_409);
xnor U3308 (N_3308,In_2344,In_525);
nor U3309 (N_3309,In_705,In_2230);
and U3310 (N_3310,In_289,In_1577);
or U3311 (N_3311,In_435,In_680);
nand U3312 (N_3312,In_1258,In_915);
nand U3313 (N_3313,In_1226,In_2197);
or U3314 (N_3314,In_32,In_1604);
or U3315 (N_3315,In_70,In_1466);
and U3316 (N_3316,In_1783,In_311);
nand U3317 (N_3317,In_2277,In_1381);
nand U3318 (N_3318,In_2307,In_2357);
nor U3319 (N_3319,In_1205,In_208);
and U3320 (N_3320,In_429,In_44);
and U3321 (N_3321,In_688,In_2363);
nor U3322 (N_3322,In_1910,In_2288);
nand U3323 (N_3323,In_1568,In_2344);
nor U3324 (N_3324,In_2393,In_1209);
and U3325 (N_3325,In_1589,In_275);
xnor U3326 (N_3326,In_2064,In_2008);
xor U3327 (N_3327,In_2450,In_824);
nand U3328 (N_3328,In_925,In_1067);
nor U3329 (N_3329,In_600,In_1934);
nand U3330 (N_3330,In_2276,In_0);
nor U3331 (N_3331,In_379,In_2358);
nor U3332 (N_3332,In_330,In_818);
nand U3333 (N_3333,In_1015,In_882);
and U3334 (N_3334,In_1908,In_1629);
or U3335 (N_3335,In_441,In_2256);
nor U3336 (N_3336,In_1530,In_2133);
nor U3337 (N_3337,In_2307,In_1446);
nor U3338 (N_3338,In_311,In_579);
nand U3339 (N_3339,In_2323,In_753);
or U3340 (N_3340,In_1434,In_2224);
xor U3341 (N_3341,In_1600,In_957);
and U3342 (N_3342,In_1522,In_480);
and U3343 (N_3343,In_1100,In_1384);
nor U3344 (N_3344,In_1419,In_1161);
nand U3345 (N_3345,In_2073,In_1387);
and U3346 (N_3346,In_1870,In_1672);
and U3347 (N_3347,In_46,In_43);
nand U3348 (N_3348,In_2060,In_1074);
or U3349 (N_3349,In_627,In_1302);
nand U3350 (N_3350,In_1384,In_2268);
nand U3351 (N_3351,In_1261,In_2258);
nand U3352 (N_3352,In_882,In_614);
nor U3353 (N_3353,In_818,In_110);
and U3354 (N_3354,In_1588,In_2467);
nand U3355 (N_3355,In_100,In_1504);
and U3356 (N_3356,In_1639,In_1082);
nand U3357 (N_3357,In_511,In_1557);
nand U3358 (N_3358,In_1505,In_1624);
and U3359 (N_3359,In_100,In_1521);
nor U3360 (N_3360,In_2113,In_2384);
nand U3361 (N_3361,In_345,In_697);
nor U3362 (N_3362,In_557,In_216);
nor U3363 (N_3363,In_1899,In_1096);
or U3364 (N_3364,In_1286,In_2321);
and U3365 (N_3365,In_414,In_1190);
or U3366 (N_3366,In_714,In_1005);
nor U3367 (N_3367,In_141,In_1956);
and U3368 (N_3368,In_1670,In_1790);
nor U3369 (N_3369,In_888,In_1915);
xor U3370 (N_3370,In_98,In_574);
xor U3371 (N_3371,In_1358,In_1075);
or U3372 (N_3372,In_2169,In_642);
nor U3373 (N_3373,In_2274,In_1834);
and U3374 (N_3374,In_1952,In_1616);
nand U3375 (N_3375,In_594,In_2361);
or U3376 (N_3376,In_1735,In_534);
or U3377 (N_3377,In_2249,In_2495);
or U3378 (N_3378,In_445,In_1379);
or U3379 (N_3379,In_2398,In_2265);
and U3380 (N_3380,In_1386,In_865);
or U3381 (N_3381,In_1082,In_954);
nor U3382 (N_3382,In_1145,In_1809);
nand U3383 (N_3383,In_100,In_958);
and U3384 (N_3384,In_2039,In_1953);
xnor U3385 (N_3385,In_460,In_490);
and U3386 (N_3386,In_80,In_1378);
nor U3387 (N_3387,In_2257,In_854);
and U3388 (N_3388,In_2463,In_2353);
nand U3389 (N_3389,In_313,In_876);
nor U3390 (N_3390,In_1105,In_1116);
or U3391 (N_3391,In_901,In_2076);
or U3392 (N_3392,In_1989,In_1639);
xnor U3393 (N_3393,In_74,In_881);
or U3394 (N_3394,In_2058,In_1237);
nor U3395 (N_3395,In_1997,In_258);
nand U3396 (N_3396,In_1756,In_1102);
and U3397 (N_3397,In_183,In_1138);
nor U3398 (N_3398,In_245,In_2218);
nand U3399 (N_3399,In_1785,In_2460);
nand U3400 (N_3400,In_2294,In_583);
or U3401 (N_3401,In_2215,In_1758);
nand U3402 (N_3402,In_1517,In_122);
or U3403 (N_3403,In_553,In_1303);
and U3404 (N_3404,In_2243,In_1784);
and U3405 (N_3405,In_2289,In_2172);
and U3406 (N_3406,In_90,In_1144);
or U3407 (N_3407,In_2443,In_1854);
xnor U3408 (N_3408,In_916,In_1831);
nor U3409 (N_3409,In_579,In_2147);
or U3410 (N_3410,In_2400,In_43);
or U3411 (N_3411,In_34,In_2431);
nor U3412 (N_3412,In_1754,In_615);
nor U3413 (N_3413,In_14,In_82);
or U3414 (N_3414,In_1867,In_1334);
or U3415 (N_3415,In_1331,In_2399);
nor U3416 (N_3416,In_2374,In_196);
nand U3417 (N_3417,In_451,In_1548);
or U3418 (N_3418,In_1840,In_241);
or U3419 (N_3419,In_1267,In_1526);
and U3420 (N_3420,In_847,In_2178);
xor U3421 (N_3421,In_1871,In_1164);
and U3422 (N_3422,In_292,In_956);
nand U3423 (N_3423,In_1127,In_876);
nand U3424 (N_3424,In_990,In_757);
or U3425 (N_3425,In_1901,In_540);
nand U3426 (N_3426,In_1366,In_2184);
and U3427 (N_3427,In_301,In_799);
and U3428 (N_3428,In_1044,In_2332);
nand U3429 (N_3429,In_1092,In_538);
and U3430 (N_3430,In_1066,In_312);
nand U3431 (N_3431,In_1619,In_2149);
or U3432 (N_3432,In_2192,In_22);
or U3433 (N_3433,In_174,In_1287);
or U3434 (N_3434,In_870,In_1050);
or U3435 (N_3435,In_984,In_254);
nand U3436 (N_3436,In_2411,In_543);
nand U3437 (N_3437,In_1834,In_100);
xnor U3438 (N_3438,In_1790,In_1692);
nand U3439 (N_3439,In_1926,In_2232);
nor U3440 (N_3440,In_729,In_2406);
or U3441 (N_3441,In_1292,In_74);
nor U3442 (N_3442,In_2039,In_369);
and U3443 (N_3443,In_2019,In_2276);
nor U3444 (N_3444,In_2135,In_1086);
and U3445 (N_3445,In_1442,In_2372);
nor U3446 (N_3446,In_23,In_932);
nor U3447 (N_3447,In_720,In_430);
nor U3448 (N_3448,In_2292,In_2165);
nor U3449 (N_3449,In_663,In_172);
and U3450 (N_3450,In_1723,In_900);
or U3451 (N_3451,In_189,In_322);
nand U3452 (N_3452,In_1836,In_2050);
or U3453 (N_3453,In_1126,In_1899);
or U3454 (N_3454,In_507,In_817);
and U3455 (N_3455,In_654,In_508);
and U3456 (N_3456,In_1489,In_1506);
nand U3457 (N_3457,In_692,In_171);
nor U3458 (N_3458,In_2355,In_1483);
and U3459 (N_3459,In_534,In_723);
or U3460 (N_3460,In_2380,In_452);
xnor U3461 (N_3461,In_49,In_1166);
and U3462 (N_3462,In_1342,In_767);
xnor U3463 (N_3463,In_2309,In_1818);
and U3464 (N_3464,In_2307,In_1517);
nand U3465 (N_3465,In_1024,In_2378);
nor U3466 (N_3466,In_418,In_1027);
and U3467 (N_3467,In_1215,In_367);
and U3468 (N_3468,In_1536,In_650);
or U3469 (N_3469,In_2388,In_415);
nand U3470 (N_3470,In_304,In_379);
or U3471 (N_3471,In_688,In_2219);
nand U3472 (N_3472,In_739,In_377);
and U3473 (N_3473,In_1490,In_2493);
nor U3474 (N_3474,In_410,In_1769);
xnor U3475 (N_3475,In_2461,In_307);
nand U3476 (N_3476,In_2337,In_79);
or U3477 (N_3477,In_1277,In_484);
or U3478 (N_3478,In_221,In_1574);
and U3479 (N_3479,In_521,In_1911);
and U3480 (N_3480,In_363,In_236);
nand U3481 (N_3481,In_760,In_21);
or U3482 (N_3482,In_2053,In_130);
and U3483 (N_3483,In_574,In_1117);
nor U3484 (N_3484,In_528,In_900);
xnor U3485 (N_3485,In_171,In_1759);
xor U3486 (N_3486,In_1007,In_104);
or U3487 (N_3487,In_659,In_714);
nand U3488 (N_3488,In_492,In_841);
nand U3489 (N_3489,In_843,In_1568);
nor U3490 (N_3490,In_1396,In_1523);
and U3491 (N_3491,In_422,In_681);
and U3492 (N_3492,In_2281,In_2309);
nor U3493 (N_3493,In_1387,In_2253);
and U3494 (N_3494,In_113,In_1692);
and U3495 (N_3495,In_1548,In_1482);
nand U3496 (N_3496,In_1099,In_11);
nand U3497 (N_3497,In_1185,In_2376);
or U3498 (N_3498,In_749,In_971);
xnor U3499 (N_3499,In_2226,In_501);
xor U3500 (N_3500,In_1289,In_1346);
nand U3501 (N_3501,In_1042,In_2410);
nor U3502 (N_3502,In_2225,In_523);
or U3503 (N_3503,In_297,In_2064);
and U3504 (N_3504,In_1969,In_2370);
and U3505 (N_3505,In_364,In_1267);
nor U3506 (N_3506,In_1679,In_2420);
and U3507 (N_3507,In_2495,In_391);
and U3508 (N_3508,In_69,In_2133);
nand U3509 (N_3509,In_1847,In_701);
and U3510 (N_3510,In_1120,In_1286);
nor U3511 (N_3511,In_1938,In_1819);
nor U3512 (N_3512,In_2100,In_2136);
nor U3513 (N_3513,In_723,In_726);
nand U3514 (N_3514,In_848,In_2037);
or U3515 (N_3515,In_874,In_907);
nor U3516 (N_3516,In_2496,In_670);
and U3517 (N_3517,In_1420,In_1464);
and U3518 (N_3518,In_45,In_492);
nand U3519 (N_3519,In_1747,In_2142);
xor U3520 (N_3520,In_399,In_1279);
or U3521 (N_3521,In_302,In_1336);
nor U3522 (N_3522,In_866,In_27);
and U3523 (N_3523,In_185,In_637);
nor U3524 (N_3524,In_1747,In_1251);
nand U3525 (N_3525,In_880,In_564);
xor U3526 (N_3526,In_2028,In_1566);
nand U3527 (N_3527,In_40,In_214);
xnor U3528 (N_3528,In_1068,In_40);
or U3529 (N_3529,In_1825,In_1190);
nand U3530 (N_3530,In_193,In_166);
and U3531 (N_3531,In_2228,In_1133);
nor U3532 (N_3532,In_1274,In_12);
and U3533 (N_3533,In_1082,In_508);
or U3534 (N_3534,In_2433,In_2198);
nand U3535 (N_3535,In_1760,In_1298);
and U3536 (N_3536,In_657,In_280);
nor U3537 (N_3537,In_1042,In_2304);
and U3538 (N_3538,In_255,In_472);
xnor U3539 (N_3539,In_923,In_2139);
nand U3540 (N_3540,In_2047,In_1199);
nor U3541 (N_3541,In_1119,In_1000);
and U3542 (N_3542,In_872,In_1130);
nor U3543 (N_3543,In_236,In_1098);
nand U3544 (N_3544,In_135,In_2009);
nor U3545 (N_3545,In_96,In_2020);
and U3546 (N_3546,In_2412,In_1577);
and U3547 (N_3547,In_2356,In_16);
nor U3548 (N_3548,In_2093,In_1457);
and U3549 (N_3549,In_583,In_2033);
or U3550 (N_3550,In_1445,In_1940);
nor U3551 (N_3551,In_1092,In_1383);
and U3552 (N_3552,In_2418,In_270);
nand U3553 (N_3553,In_1232,In_913);
xnor U3554 (N_3554,In_432,In_2069);
nor U3555 (N_3555,In_1311,In_200);
nand U3556 (N_3556,In_2339,In_945);
nand U3557 (N_3557,In_464,In_1337);
nand U3558 (N_3558,In_36,In_365);
or U3559 (N_3559,In_2494,In_347);
and U3560 (N_3560,In_2274,In_1645);
nand U3561 (N_3561,In_98,In_289);
nand U3562 (N_3562,In_540,In_438);
or U3563 (N_3563,In_372,In_2497);
nor U3564 (N_3564,In_1364,In_113);
and U3565 (N_3565,In_1207,In_1169);
and U3566 (N_3566,In_1384,In_1298);
and U3567 (N_3567,In_1102,In_2092);
and U3568 (N_3568,In_1397,In_299);
nand U3569 (N_3569,In_2194,In_105);
nand U3570 (N_3570,In_570,In_1925);
and U3571 (N_3571,In_493,In_1153);
nand U3572 (N_3572,In_2420,In_1869);
or U3573 (N_3573,In_527,In_1664);
xnor U3574 (N_3574,In_2288,In_681);
and U3575 (N_3575,In_1767,In_2248);
nor U3576 (N_3576,In_800,In_1409);
nor U3577 (N_3577,In_1473,In_448);
or U3578 (N_3578,In_1720,In_1368);
nor U3579 (N_3579,In_390,In_525);
and U3580 (N_3580,In_2356,In_2018);
and U3581 (N_3581,In_2280,In_2132);
nor U3582 (N_3582,In_2469,In_2084);
and U3583 (N_3583,In_2266,In_1049);
xor U3584 (N_3584,In_205,In_266);
or U3585 (N_3585,In_1302,In_1723);
nand U3586 (N_3586,In_2411,In_1936);
nand U3587 (N_3587,In_640,In_815);
nand U3588 (N_3588,In_40,In_126);
nand U3589 (N_3589,In_1220,In_1335);
xor U3590 (N_3590,In_128,In_1238);
and U3591 (N_3591,In_1619,In_1544);
nand U3592 (N_3592,In_2126,In_369);
and U3593 (N_3593,In_1012,In_1801);
or U3594 (N_3594,In_452,In_1300);
or U3595 (N_3595,In_1569,In_1116);
and U3596 (N_3596,In_1968,In_333);
and U3597 (N_3597,In_2228,In_0);
nand U3598 (N_3598,In_1577,In_973);
nand U3599 (N_3599,In_51,In_906);
nor U3600 (N_3600,In_1028,In_2185);
or U3601 (N_3601,In_2245,In_432);
or U3602 (N_3602,In_14,In_691);
and U3603 (N_3603,In_1581,In_1429);
nand U3604 (N_3604,In_781,In_1345);
or U3605 (N_3605,In_2337,In_2195);
or U3606 (N_3606,In_1789,In_1988);
xnor U3607 (N_3607,In_745,In_1486);
or U3608 (N_3608,In_1982,In_1697);
or U3609 (N_3609,In_426,In_130);
nor U3610 (N_3610,In_1797,In_1769);
nor U3611 (N_3611,In_1971,In_806);
and U3612 (N_3612,In_1663,In_1664);
nor U3613 (N_3613,In_192,In_1750);
nand U3614 (N_3614,In_2385,In_578);
nor U3615 (N_3615,In_1778,In_1372);
or U3616 (N_3616,In_489,In_1438);
xnor U3617 (N_3617,In_1655,In_1746);
xor U3618 (N_3618,In_1235,In_2359);
and U3619 (N_3619,In_1953,In_2376);
nor U3620 (N_3620,In_274,In_927);
xnor U3621 (N_3621,In_2226,In_47);
or U3622 (N_3622,In_838,In_872);
xnor U3623 (N_3623,In_305,In_2081);
and U3624 (N_3624,In_1769,In_413);
and U3625 (N_3625,In_1873,In_502);
nand U3626 (N_3626,In_1962,In_1823);
or U3627 (N_3627,In_2070,In_2287);
nand U3628 (N_3628,In_1519,In_1806);
nand U3629 (N_3629,In_993,In_106);
xnor U3630 (N_3630,In_933,In_727);
and U3631 (N_3631,In_2316,In_2151);
and U3632 (N_3632,In_1841,In_258);
nor U3633 (N_3633,In_1113,In_1608);
or U3634 (N_3634,In_1637,In_2257);
or U3635 (N_3635,In_295,In_1995);
nor U3636 (N_3636,In_1021,In_638);
and U3637 (N_3637,In_2343,In_1471);
nor U3638 (N_3638,In_1567,In_17);
nand U3639 (N_3639,In_2384,In_2093);
or U3640 (N_3640,In_166,In_1858);
nand U3641 (N_3641,In_1288,In_380);
and U3642 (N_3642,In_2427,In_2407);
nor U3643 (N_3643,In_1741,In_99);
or U3644 (N_3644,In_1422,In_2313);
nand U3645 (N_3645,In_246,In_1405);
nand U3646 (N_3646,In_895,In_2467);
nor U3647 (N_3647,In_1311,In_2030);
xor U3648 (N_3648,In_2261,In_1585);
and U3649 (N_3649,In_564,In_2406);
xor U3650 (N_3650,In_1106,In_1165);
nor U3651 (N_3651,In_291,In_2018);
nand U3652 (N_3652,In_453,In_2220);
nand U3653 (N_3653,In_665,In_432);
nor U3654 (N_3654,In_1657,In_1149);
nor U3655 (N_3655,In_952,In_1212);
nand U3656 (N_3656,In_1621,In_91);
nor U3657 (N_3657,In_1141,In_2310);
xnor U3658 (N_3658,In_1912,In_266);
xor U3659 (N_3659,In_1085,In_414);
or U3660 (N_3660,In_1247,In_1750);
nand U3661 (N_3661,In_580,In_818);
or U3662 (N_3662,In_2030,In_2281);
nand U3663 (N_3663,In_802,In_1350);
nand U3664 (N_3664,In_1355,In_1920);
or U3665 (N_3665,In_2370,In_1901);
nand U3666 (N_3666,In_1285,In_926);
xnor U3667 (N_3667,In_355,In_33);
or U3668 (N_3668,In_1679,In_633);
nand U3669 (N_3669,In_1310,In_219);
or U3670 (N_3670,In_2296,In_79);
or U3671 (N_3671,In_2487,In_273);
and U3672 (N_3672,In_30,In_684);
or U3673 (N_3673,In_633,In_2446);
and U3674 (N_3674,In_2081,In_1321);
nand U3675 (N_3675,In_822,In_169);
and U3676 (N_3676,In_1872,In_952);
xor U3677 (N_3677,In_1427,In_890);
or U3678 (N_3678,In_1392,In_1193);
or U3679 (N_3679,In_1017,In_2240);
and U3680 (N_3680,In_529,In_1077);
or U3681 (N_3681,In_1546,In_983);
and U3682 (N_3682,In_964,In_265);
and U3683 (N_3683,In_1218,In_397);
nor U3684 (N_3684,In_2261,In_1009);
and U3685 (N_3685,In_1547,In_1313);
xor U3686 (N_3686,In_1862,In_2389);
and U3687 (N_3687,In_1187,In_1697);
and U3688 (N_3688,In_175,In_1567);
nand U3689 (N_3689,In_2019,In_133);
nor U3690 (N_3690,In_2378,In_2210);
or U3691 (N_3691,In_1485,In_1813);
and U3692 (N_3692,In_1027,In_1016);
or U3693 (N_3693,In_1707,In_1288);
nand U3694 (N_3694,In_1032,In_555);
and U3695 (N_3695,In_949,In_2191);
or U3696 (N_3696,In_698,In_124);
nand U3697 (N_3697,In_83,In_2082);
or U3698 (N_3698,In_1375,In_197);
nand U3699 (N_3699,In_2131,In_486);
nand U3700 (N_3700,In_2040,In_397);
or U3701 (N_3701,In_1229,In_984);
nand U3702 (N_3702,In_1540,In_393);
nand U3703 (N_3703,In_1744,In_2110);
or U3704 (N_3704,In_1564,In_2323);
nand U3705 (N_3705,In_2163,In_2005);
or U3706 (N_3706,In_1595,In_1189);
and U3707 (N_3707,In_1621,In_1057);
or U3708 (N_3708,In_1388,In_181);
and U3709 (N_3709,In_1094,In_269);
nor U3710 (N_3710,In_1202,In_2454);
or U3711 (N_3711,In_820,In_248);
or U3712 (N_3712,In_969,In_1460);
nand U3713 (N_3713,In_2449,In_2426);
or U3714 (N_3714,In_2399,In_2190);
nand U3715 (N_3715,In_501,In_1341);
nand U3716 (N_3716,In_16,In_1025);
and U3717 (N_3717,In_1316,In_1324);
nand U3718 (N_3718,In_2146,In_107);
nor U3719 (N_3719,In_617,In_92);
and U3720 (N_3720,In_1072,In_1224);
nor U3721 (N_3721,In_1090,In_437);
nor U3722 (N_3722,In_593,In_1178);
and U3723 (N_3723,In_1609,In_1460);
nor U3724 (N_3724,In_732,In_1278);
or U3725 (N_3725,In_1886,In_1197);
nor U3726 (N_3726,In_49,In_1586);
nand U3727 (N_3727,In_2393,In_414);
nand U3728 (N_3728,In_847,In_1345);
xor U3729 (N_3729,In_1938,In_1971);
nor U3730 (N_3730,In_467,In_2268);
or U3731 (N_3731,In_737,In_864);
nor U3732 (N_3732,In_1726,In_1226);
nor U3733 (N_3733,In_2327,In_64);
or U3734 (N_3734,In_71,In_2173);
nor U3735 (N_3735,In_654,In_358);
nand U3736 (N_3736,In_1354,In_357);
and U3737 (N_3737,In_1245,In_1269);
and U3738 (N_3738,In_1876,In_2293);
nand U3739 (N_3739,In_2104,In_1209);
nand U3740 (N_3740,In_2130,In_2132);
nor U3741 (N_3741,In_33,In_637);
and U3742 (N_3742,In_888,In_1417);
nor U3743 (N_3743,In_754,In_332);
nand U3744 (N_3744,In_564,In_2063);
or U3745 (N_3745,In_1079,In_1169);
and U3746 (N_3746,In_962,In_1410);
xor U3747 (N_3747,In_888,In_717);
nor U3748 (N_3748,In_490,In_1959);
nor U3749 (N_3749,In_2250,In_1213);
and U3750 (N_3750,In_2181,In_1659);
nand U3751 (N_3751,In_2262,In_174);
nor U3752 (N_3752,In_272,In_2382);
and U3753 (N_3753,In_1072,In_1354);
nand U3754 (N_3754,In_1642,In_1289);
and U3755 (N_3755,In_1984,In_1817);
nand U3756 (N_3756,In_2060,In_693);
and U3757 (N_3757,In_1476,In_1271);
or U3758 (N_3758,In_1148,In_1528);
nand U3759 (N_3759,In_680,In_698);
or U3760 (N_3760,In_2418,In_1537);
and U3761 (N_3761,In_803,In_2377);
nand U3762 (N_3762,In_1227,In_373);
or U3763 (N_3763,In_1714,In_387);
nand U3764 (N_3764,In_876,In_1993);
nor U3765 (N_3765,In_1459,In_31);
nor U3766 (N_3766,In_139,In_1133);
and U3767 (N_3767,In_411,In_1092);
and U3768 (N_3768,In_1588,In_2442);
xnor U3769 (N_3769,In_509,In_2152);
nor U3770 (N_3770,In_1227,In_1192);
and U3771 (N_3771,In_2272,In_1491);
or U3772 (N_3772,In_344,In_977);
nor U3773 (N_3773,In_369,In_2255);
and U3774 (N_3774,In_139,In_1272);
nor U3775 (N_3775,In_2219,In_801);
nor U3776 (N_3776,In_1269,In_2367);
or U3777 (N_3777,In_1528,In_277);
nor U3778 (N_3778,In_1439,In_260);
or U3779 (N_3779,In_1143,In_2250);
nand U3780 (N_3780,In_2201,In_1058);
nand U3781 (N_3781,In_1307,In_2031);
or U3782 (N_3782,In_968,In_809);
nand U3783 (N_3783,In_1918,In_2061);
nor U3784 (N_3784,In_983,In_801);
nand U3785 (N_3785,In_2377,In_2487);
nand U3786 (N_3786,In_2133,In_199);
nand U3787 (N_3787,In_432,In_1628);
nor U3788 (N_3788,In_518,In_533);
and U3789 (N_3789,In_794,In_1563);
or U3790 (N_3790,In_242,In_1889);
nor U3791 (N_3791,In_1471,In_243);
nand U3792 (N_3792,In_2466,In_2463);
nand U3793 (N_3793,In_2250,In_49);
and U3794 (N_3794,In_1949,In_1034);
nor U3795 (N_3795,In_1936,In_309);
and U3796 (N_3796,In_1342,In_937);
nor U3797 (N_3797,In_1351,In_215);
nand U3798 (N_3798,In_755,In_568);
and U3799 (N_3799,In_890,In_1138);
nor U3800 (N_3800,In_2173,In_2045);
nand U3801 (N_3801,In_937,In_2116);
and U3802 (N_3802,In_1878,In_223);
and U3803 (N_3803,In_1059,In_560);
nand U3804 (N_3804,In_1672,In_1299);
or U3805 (N_3805,In_1095,In_711);
nand U3806 (N_3806,In_1652,In_2475);
and U3807 (N_3807,In_1166,In_1747);
and U3808 (N_3808,In_1844,In_1270);
or U3809 (N_3809,In_54,In_672);
nand U3810 (N_3810,In_955,In_6);
nor U3811 (N_3811,In_557,In_361);
nand U3812 (N_3812,In_350,In_1958);
nand U3813 (N_3813,In_598,In_2271);
or U3814 (N_3814,In_2422,In_2333);
or U3815 (N_3815,In_537,In_2483);
nand U3816 (N_3816,In_669,In_586);
or U3817 (N_3817,In_1542,In_388);
nor U3818 (N_3818,In_1950,In_228);
nand U3819 (N_3819,In_2326,In_359);
and U3820 (N_3820,In_2465,In_1563);
xnor U3821 (N_3821,In_79,In_599);
and U3822 (N_3822,In_763,In_138);
and U3823 (N_3823,In_2004,In_521);
nor U3824 (N_3824,In_131,In_1555);
nand U3825 (N_3825,In_2261,In_503);
xnor U3826 (N_3826,In_1021,In_2092);
nor U3827 (N_3827,In_99,In_1560);
and U3828 (N_3828,In_1318,In_2107);
nor U3829 (N_3829,In_1294,In_1544);
or U3830 (N_3830,In_2157,In_201);
xor U3831 (N_3831,In_1448,In_944);
nor U3832 (N_3832,In_944,In_353);
nand U3833 (N_3833,In_276,In_87);
and U3834 (N_3834,In_1364,In_470);
and U3835 (N_3835,In_2065,In_695);
nor U3836 (N_3836,In_505,In_1211);
nand U3837 (N_3837,In_1140,In_1458);
or U3838 (N_3838,In_2048,In_1004);
nor U3839 (N_3839,In_1559,In_634);
nand U3840 (N_3840,In_659,In_1629);
or U3841 (N_3841,In_1361,In_1057);
or U3842 (N_3842,In_358,In_344);
xor U3843 (N_3843,In_1461,In_67);
nand U3844 (N_3844,In_910,In_1896);
xnor U3845 (N_3845,In_1509,In_2344);
nand U3846 (N_3846,In_2477,In_416);
nor U3847 (N_3847,In_2353,In_1408);
or U3848 (N_3848,In_1854,In_1314);
or U3849 (N_3849,In_2027,In_153);
or U3850 (N_3850,In_1598,In_1660);
nand U3851 (N_3851,In_1050,In_2392);
nand U3852 (N_3852,In_1239,In_2131);
or U3853 (N_3853,In_919,In_813);
and U3854 (N_3854,In_1782,In_692);
and U3855 (N_3855,In_2111,In_1479);
or U3856 (N_3856,In_778,In_66);
xnor U3857 (N_3857,In_1533,In_1044);
or U3858 (N_3858,In_99,In_1660);
nand U3859 (N_3859,In_1420,In_1605);
nor U3860 (N_3860,In_91,In_2010);
nand U3861 (N_3861,In_2211,In_1633);
or U3862 (N_3862,In_1759,In_1434);
nand U3863 (N_3863,In_1626,In_825);
or U3864 (N_3864,In_1766,In_1212);
nand U3865 (N_3865,In_336,In_203);
nand U3866 (N_3866,In_2380,In_161);
and U3867 (N_3867,In_782,In_1330);
or U3868 (N_3868,In_425,In_1153);
and U3869 (N_3869,In_244,In_2427);
or U3870 (N_3870,In_1252,In_1148);
or U3871 (N_3871,In_2235,In_2061);
or U3872 (N_3872,In_2247,In_1816);
or U3873 (N_3873,In_1308,In_1320);
nor U3874 (N_3874,In_648,In_2462);
nand U3875 (N_3875,In_2084,In_548);
and U3876 (N_3876,In_994,In_2354);
xnor U3877 (N_3877,In_1006,In_1230);
nor U3878 (N_3878,In_2020,In_1844);
nand U3879 (N_3879,In_1534,In_1074);
nor U3880 (N_3880,In_2382,In_1540);
nor U3881 (N_3881,In_1603,In_1526);
nor U3882 (N_3882,In_1280,In_484);
xnor U3883 (N_3883,In_1633,In_412);
and U3884 (N_3884,In_2426,In_31);
and U3885 (N_3885,In_1551,In_326);
nand U3886 (N_3886,In_404,In_770);
or U3887 (N_3887,In_2133,In_1485);
nand U3888 (N_3888,In_2180,In_1632);
and U3889 (N_3889,In_845,In_1174);
nor U3890 (N_3890,In_2440,In_2263);
nor U3891 (N_3891,In_1200,In_490);
or U3892 (N_3892,In_1815,In_988);
nand U3893 (N_3893,In_594,In_848);
xnor U3894 (N_3894,In_2133,In_494);
xor U3895 (N_3895,In_2172,In_454);
or U3896 (N_3896,In_419,In_169);
nand U3897 (N_3897,In_2218,In_485);
or U3898 (N_3898,In_1417,In_753);
or U3899 (N_3899,In_1914,In_606);
nand U3900 (N_3900,In_1239,In_1139);
or U3901 (N_3901,In_1504,In_2052);
or U3902 (N_3902,In_702,In_786);
nor U3903 (N_3903,In_1752,In_202);
nor U3904 (N_3904,In_2328,In_529);
and U3905 (N_3905,In_308,In_659);
and U3906 (N_3906,In_524,In_299);
nand U3907 (N_3907,In_1270,In_1078);
and U3908 (N_3908,In_332,In_911);
nand U3909 (N_3909,In_1975,In_1713);
nand U3910 (N_3910,In_755,In_718);
nand U3911 (N_3911,In_827,In_2084);
and U3912 (N_3912,In_1743,In_335);
nor U3913 (N_3913,In_695,In_1202);
or U3914 (N_3914,In_1478,In_1425);
xnor U3915 (N_3915,In_152,In_766);
or U3916 (N_3916,In_967,In_2153);
xnor U3917 (N_3917,In_378,In_1809);
nor U3918 (N_3918,In_5,In_285);
and U3919 (N_3919,In_552,In_2357);
and U3920 (N_3920,In_2116,In_2334);
and U3921 (N_3921,In_2306,In_691);
and U3922 (N_3922,In_1644,In_2286);
nand U3923 (N_3923,In_1708,In_2286);
and U3924 (N_3924,In_1935,In_748);
or U3925 (N_3925,In_1468,In_1441);
or U3926 (N_3926,In_1449,In_1820);
or U3927 (N_3927,In_2001,In_1134);
and U3928 (N_3928,In_1460,In_1449);
or U3929 (N_3929,In_2187,In_840);
or U3930 (N_3930,In_657,In_2329);
nor U3931 (N_3931,In_318,In_1173);
nor U3932 (N_3932,In_1402,In_887);
nor U3933 (N_3933,In_232,In_2272);
nor U3934 (N_3934,In_564,In_1840);
and U3935 (N_3935,In_718,In_2149);
nand U3936 (N_3936,In_606,In_1486);
nor U3937 (N_3937,In_1441,In_3);
nor U3938 (N_3938,In_2001,In_672);
and U3939 (N_3939,In_843,In_2277);
or U3940 (N_3940,In_1757,In_139);
nor U3941 (N_3941,In_1154,In_868);
nand U3942 (N_3942,In_2331,In_178);
nor U3943 (N_3943,In_1272,In_61);
or U3944 (N_3944,In_1542,In_588);
and U3945 (N_3945,In_2046,In_530);
nand U3946 (N_3946,In_1975,In_1531);
or U3947 (N_3947,In_1178,In_418);
nor U3948 (N_3948,In_71,In_1268);
and U3949 (N_3949,In_1410,In_1897);
or U3950 (N_3950,In_1876,In_179);
and U3951 (N_3951,In_946,In_150);
xor U3952 (N_3952,In_2336,In_426);
nor U3953 (N_3953,In_192,In_50);
nor U3954 (N_3954,In_918,In_1657);
nand U3955 (N_3955,In_62,In_1314);
and U3956 (N_3956,In_1891,In_423);
and U3957 (N_3957,In_129,In_495);
xnor U3958 (N_3958,In_369,In_1567);
nand U3959 (N_3959,In_1878,In_226);
or U3960 (N_3960,In_1035,In_131);
or U3961 (N_3961,In_1217,In_1038);
nand U3962 (N_3962,In_483,In_238);
nor U3963 (N_3963,In_591,In_763);
xnor U3964 (N_3964,In_121,In_1402);
and U3965 (N_3965,In_2209,In_558);
and U3966 (N_3966,In_2044,In_643);
nand U3967 (N_3967,In_783,In_1308);
or U3968 (N_3968,In_435,In_1574);
nand U3969 (N_3969,In_505,In_743);
nand U3970 (N_3970,In_2098,In_334);
xor U3971 (N_3971,In_988,In_435);
and U3972 (N_3972,In_828,In_225);
nand U3973 (N_3973,In_2161,In_1183);
nor U3974 (N_3974,In_64,In_2453);
nor U3975 (N_3975,In_928,In_1019);
and U3976 (N_3976,In_2094,In_779);
nor U3977 (N_3977,In_1550,In_1746);
nand U3978 (N_3978,In_344,In_639);
nand U3979 (N_3979,In_2066,In_2033);
nor U3980 (N_3980,In_486,In_419);
xor U3981 (N_3981,In_1343,In_93);
nand U3982 (N_3982,In_963,In_1116);
nor U3983 (N_3983,In_1510,In_51);
or U3984 (N_3984,In_1972,In_1723);
nand U3985 (N_3985,In_250,In_1581);
or U3986 (N_3986,In_183,In_503);
and U3987 (N_3987,In_2485,In_992);
and U3988 (N_3988,In_2407,In_1046);
nand U3989 (N_3989,In_456,In_1090);
nand U3990 (N_3990,In_2420,In_264);
or U3991 (N_3991,In_40,In_1941);
and U3992 (N_3992,In_2287,In_318);
nor U3993 (N_3993,In_2315,In_250);
nand U3994 (N_3994,In_2316,In_2341);
nand U3995 (N_3995,In_1928,In_2272);
and U3996 (N_3996,In_849,In_1525);
or U3997 (N_3997,In_571,In_2164);
nand U3998 (N_3998,In_326,In_1949);
nor U3999 (N_3999,In_647,In_2475);
nand U4000 (N_4000,In_241,In_1189);
nand U4001 (N_4001,In_262,In_1436);
nor U4002 (N_4002,In_1055,In_1902);
nand U4003 (N_4003,In_139,In_1047);
or U4004 (N_4004,In_2342,In_2314);
nor U4005 (N_4005,In_2090,In_804);
or U4006 (N_4006,In_1585,In_1084);
and U4007 (N_4007,In_476,In_2285);
and U4008 (N_4008,In_2151,In_281);
and U4009 (N_4009,In_331,In_1754);
nand U4010 (N_4010,In_2255,In_1511);
and U4011 (N_4011,In_30,In_2392);
and U4012 (N_4012,In_155,In_370);
and U4013 (N_4013,In_858,In_2266);
or U4014 (N_4014,In_1602,In_1871);
and U4015 (N_4015,In_1943,In_447);
and U4016 (N_4016,In_1213,In_903);
nor U4017 (N_4017,In_885,In_1424);
and U4018 (N_4018,In_82,In_812);
and U4019 (N_4019,In_196,In_2378);
nand U4020 (N_4020,In_1598,In_44);
and U4021 (N_4021,In_1172,In_2259);
and U4022 (N_4022,In_137,In_2365);
nand U4023 (N_4023,In_1997,In_1531);
nand U4024 (N_4024,In_157,In_1110);
nand U4025 (N_4025,In_1790,In_2054);
and U4026 (N_4026,In_911,In_178);
nand U4027 (N_4027,In_2375,In_720);
and U4028 (N_4028,In_2176,In_40);
xnor U4029 (N_4029,In_843,In_1283);
nor U4030 (N_4030,In_933,In_2443);
nor U4031 (N_4031,In_458,In_2299);
nand U4032 (N_4032,In_1740,In_1894);
or U4033 (N_4033,In_52,In_733);
or U4034 (N_4034,In_1343,In_805);
and U4035 (N_4035,In_1597,In_366);
nor U4036 (N_4036,In_732,In_2222);
or U4037 (N_4037,In_1652,In_480);
nand U4038 (N_4038,In_363,In_2335);
and U4039 (N_4039,In_33,In_657);
nand U4040 (N_4040,In_185,In_2088);
nor U4041 (N_4041,In_235,In_428);
nand U4042 (N_4042,In_1895,In_1669);
or U4043 (N_4043,In_464,In_888);
or U4044 (N_4044,In_677,In_2030);
nand U4045 (N_4045,In_57,In_1020);
and U4046 (N_4046,In_536,In_1568);
and U4047 (N_4047,In_1106,In_1082);
nand U4048 (N_4048,In_1007,In_2060);
or U4049 (N_4049,In_1651,In_1461);
xnor U4050 (N_4050,In_616,In_1130);
and U4051 (N_4051,In_2175,In_1047);
nand U4052 (N_4052,In_1377,In_732);
or U4053 (N_4053,In_1579,In_2121);
or U4054 (N_4054,In_1558,In_950);
xor U4055 (N_4055,In_1303,In_771);
and U4056 (N_4056,In_739,In_2239);
xnor U4057 (N_4057,In_1224,In_1982);
nand U4058 (N_4058,In_1640,In_2195);
nor U4059 (N_4059,In_1779,In_113);
or U4060 (N_4060,In_1655,In_51);
or U4061 (N_4061,In_1525,In_1784);
nand U4062 (N_4062,In_78,In_1791);
nand U4063 (N_4063,In_1912,In_1303);
or U4064 (N_4064,In_427,In_2176);
nor U4065 (N_4065,In_1966,In_1647);
and U4066 (N_4066,In_788,In_377);
and U4067 (N_4067,In_615,In_1952);
nor U4068 (N_4068,In_659,In_2414);
nor U4069 (N_4069,In_778,In_1095);
nand U4070 (N_4070,In_1092,In_2327);
nor U4071 (N_4071,In_253,In_2468);
nand U4072 (N_4072,In_2211,In_1364);
nor U4073 (N_4073,In_222,In_1338);
xor U4074 (N_4074,In_100,In_1288);
or U4075 (N_4075,In_1329,In_1663);
nand U4076 (N_4076,In_1163,In_983);
nor U4077 (N_4077,In_957,In_2327);
nand U4078 (N_4078,In_1413,In_962);
and U4079 (N_4079,In_1993,In_117);
nand U4080 (N_4080,In_712,In_324);
xnor U4081 (N_4081,In_1171,In_923);
and U4082 (N_4082,In_263,In_262);
or U4083 (N_4083,In_2133,In_634);
nand U4084 (N_4084,In_1225,In_924);
nand U4085 (N_4085,In_133,In_49);
nand U4086 (N_4086,In_1034,In_1415);
xnor U4087 (N_4087,In_1040,In_2053);
nor U4088 (N_4088,In_152,In_270);
xnor U4089 (N_4089,In_439,In_351);
or U4090 (N_4090,In_1051,In_2251);
nor U4091 (N_4091,In_1168,In_676);
xor U4092 (N_4092,In_1419,In_708);
nand U4093 (N_4093,In_2270,In_7);
nor U4094 (N_4094,In_1627,In_122);
nor U4095 (N_4095,In_864,In_1367);
and U4096 (N_4096,In_197,In_1323);
xnor U4097 (N_4097,In_655,In_1434);
or U4098 (N_4098,In_735,In_146);
nor U4099 (N_4099,In_1970,In_1088);
nand U4100 (N_4100,In_425,In_1474);
nor U4101 (N_4101,In_2343,In_450);
nor U4102 (N_4102,In_1944,In_1325);
or U4103 (N_4103,In_1111,In_1674);
or U4104 (N_4104,In_1422,In_154);
nand U4105 (N_4105,In_1204,In_2105);
or U4106 (N_4106,In_482,In_855);
and U4107 (N_4107,In_2232,In_190);
nand U4108 (N_4108,In_50,In_248);
and U4109 (N_4109,In_2353,In_1512);
and U4110 (N_4110,In_1944,In_1560);
nand U4111 (N_4111,In_1601,In_590);
nand U4112 (N_4112,In_175,In_1558);
and U4113 (N_4113,In_2018,In_1820);
nand U4114 (N_4114,In_41,In_1885);
nor U4115 (N_4115,In_1741,In_2229);
and U4116 (N_4116,In_1621,In_1194);
or U4117 (N_4117,In_2227,In_55);
nand U4118 (N_4118,In_1496,In_819);
or U4119 (N_4119,In_657,In_1403);
nor U4120 (N_4120,In_921,In_1292);
or U4121 (N_4121,In_948,In_1197);
or U4122 (N_4122,In_795,In_2460);
nor U4123 (N_4123,In_2268,In_853);
and U4124 (N_4124,In_2413,In_228);
nor U4125 (N_4125,In_448,In_2214);
or U4126 (N_4126,In_1279,In_1311);
nor U4127 (N_4127,In_887,In_27);
nor U4128 (N_4128,In_512,In_1148);
and U4129 (N_4129,In_623,In_339);
nand U4130 (N_4130,In_173,In_2161);
nor U4131 (N_4131,In_2235,In_892);
or U4132 (N_4132,In_1007,In_1611);
nor U4133 (N_4133,In_2351,In_905);
and U4134 (N_4134,In_1639,In_2181);
nand U4135 (N_4135,In_1038,In_432);
nand U4136 (N_4136,In_1288,In_2468);
nor U4137 (N_4137,In_1416,In_369);
and U4138 (N_4138,In_470,In_2002);
xnor U4139 (N_4139,In_332,In_1483);
and U4140 (N_4140,In_62,In_1545);
or U4141 (N_4141,In_1533,In_1832);
xor U4142 (N_4142,In_320,In_1738);
and U4143 (N_4143,In_1403,In_742);
nand U4144 (N_4144,In_164,In_1386);
nor U4145 (N_4145,In_1554,In_2044);
nand U4146 (N_4146,In_374,In_71);
or U4147 (N_4147,In_416,In_859);
nor U4148 (N_4148,In_18,In_1060);
and U4149 (N_4149,In_1077,In_1462);
nor U4150 (N_4150,In_1947,In_968);
or U4151 (N_4151,In_1509,In_2389);
xnor U4152 (N_4152,In_471,In_1689);
and U4153 (N_4153,In_401,In_1987);
nand U4154 (N_4154,In_2397,In_1340);
nor U4155 (N_4155,In_2128,In_1661);
nor U4156 (N_4156,In_13,In_1070);
nor U4157 (N_4157,In_457,In_776);
or U4158 (N_4158,In_625,In_527);
nor U4159 (N_4159,In_778,In_175);
and U4160 (N_4160,In_1566,In_80);
nand U4161 (N_4161,In_946,In_2103);
xor U4162 (N_4162,In_728,In_941);
and U4163 (N_4163,In_593,In_2086);
and U4164 (N_4164,In_538,In_1545);
nand U4165 (N_4165,In_1819,In_20);
xor U4166 (N_4166,In_1111,In_2065);
nor U4167 (N_4167,In_2444,In_1277);
nand U4168 (N_4168,In_640,In_1765);
xor U4169 (N_4169,In_1683,In_333);
xnor U4170 (N_4170,In_752,In_1639);
and U4171 (N_4171,In_1391,In_2105);
nand U4172 (N_4172,In_2457,In_1503);
nand U4173 (N_4173,In_1318,In_390);
and U4174 (N_4174,In_475,In_1673);
nand U4175 (N_4175,In_299,In_1709);
nand U4176 (N_4176,In_563,In_644);
nor U4177 (N_4177,In_2304,In_1835);
and U4178 (N_4178,In_585,In_2054);
nand U4179 (N_4179,In_1769,In_674);
xnor U4180 (N_4180,In_2497,In_740);
xnor U4181 (N_4181,In_1078,In_294);
nor U4182 (N_4182,In_705,In_1302);
xor U4183 (N_4183,In_501,In_1977);
nand U4184 (N_4184,In_524,In_2105);
nand U4185 (N_4185,In_680,In_1271);
nand U4186 (N_4186,In_931,In_1640);
nand U4187 (N_4187,In_1230,In_291);
and U4188 (N_4188,In_597,In_1327);
nor U4189 (N_4189,In_1696,In_499);
or U4190 (N_4190,In_2181,In_1656);
nand U4191 (N_4191,In_435,In_882);
nand U4192 (N_4192,In_439,In_2267);
nand U4193 (N_4193,In_2293,In_1824);
nor U4194 (N_4194,In_2138,In_1176);
or U4195 (N_4195,In_1163,In_707);
or U4196 (N_4196,In_1163,In_1488);
nor U4197 (N_4197,In_1765,In_1149);
or U4198 (N_4198,In_818,In_1585);
nand U4199 (N_4199,In_1234,In_307);
nand U4200 (N_4200,In_271,In_519);
xnor U4201 (N_4201,In_1581,In_527);
and U4202 (N_4202,In_1240,In_1406);
and U4203 (N_4203,In_1351,In_2017);
nor U4204 (N_4204,In_1259,In_557);
nor U4205 (N_4205,In_2420,In_1173);
or U4206 (N_4206,In_324,In_983);
nand U4207 (N_4207,In_622,In_1217);
nor U4208 (N_4208,In_2313,In_2104);
or U4209 (N_4209,In_2350,In_1695);
or U4210 (N_4210,In_789,In_29);
nor U4211 (N_4211,In_186,In_692);
nor U4212 (N_4212,In_1955,In_802);
and U4213 (N_4213,In_830,In_2192);
and U4214 (N_4214,In_940,In_2033);
nor U4215 (N_4215,In_1017,In_443);
nor U4216 (N_4216,In_1396,In_2009);
nand U4217 (N_4217,In_38,In_291);
nor U4218 (N_4218,In_2196,In_25);
and U4219 (N_4219,In_1504,In_324);
xnor U4220 (N_4220,In_1450,In_1064);
nand U4221 (N_4221,In_1224,In_1330);
and U4222 (N_4222,In_822,In_814);
and U4223 (N_4223,In_1788,In_13);
nor U4224 (N_4224,In_295,In_2155);
nor U4225 (N_4225,In_813,In_1770);
nand U4226 (N_4226,In_2467,In_440);
and U4227 (N_4227,In_977,In_680);
and U4228 (N_4228,In_1363,In_1867);
or U4229 (N_4229,In_2133,In_335);
nor U4230 (N_4230,In_627,In_2333);
and U4231 (N_4231,In_506,In_2070);
and U4232 (N_4232,In_472,In_1403);
nand U4233 (N_4233,In_2177,In_2330);
nand U4234 (N_4234,In_742,In_1184);
nor U4235 (N_4235,In_2140,In_1721);
or U4236 (N_4236,In_605,In_1606);
xnor U4237 (N_4237,In_785,In_2047);
nand U4238 (N_4238,In_2052,In_60);
nor U4239 (N_4239,In_2243,In_2114);
nor U4240 (N_4240,In_1070,In_555);
or U4241 (N_4241,In_923,In_1028);
nand U4242 (N_4242,In_2,In_2382);
nand U4243 (N_4243,In_856,In_2019);
xor U4244 (N_4244,In_34,In_2125);
and U4245 (N_4245,In_2383,In_391);
and U4246 (N_4246,In_441,In_1539);
xor U4247 (N_4247,In_437,In_322);
or U4248 (N_4248,In_1076,In_2053);
or U4249 (N_4249,In_2107,In_1505);
nor U4250 (N_4250,In_1540,In_1707);
nand U4251 (N_4251,In_295,In_1838);
and U4252 (N_4252,In_2055,In_1592);
and U4253 (N_4253,In_837,In_1788);
or U4254 (N_4254,In_221,In_1623);
or U4255 (N_4255,In_1178,In_965);
nand U4256 (N_4256,In_2186,In_737);
and U4257 (N_4257,In_1593,In_880);
nand U4258 (N_4258,In_1012,In_2308);
and U4259 (N_4259,In_1991,In_563);
or U4260 (N_4260,In_1126,In_284);
or U4261 (N_4261,In_204,In_2286);
or U4262 (N_4262,In_2040,In_2250);
nor U4263 (N_4263,In_2041,In_1290);
nor U4264 (N_4264,In_641,In_2251);
nand U4265 (N_4265,In_1583,In_1088);
nor U4266 (N_4266,In_1213,In_2499);
nor U4267 (N_4267,In_1719,In_1747);
nor U4268 (N_4268,In_1354,In_527);
or U4269 (N_4269,In_933,In_423);
nor U4270 (N_4270,In_2158,In_2412);
and U4271 (N_4271,In_142,In_2281);
or U4272 (N_4272,In_116,In_12);
or U4273 (N_4273,In_231,In_494);
nand U4274 (N_4274,In_600,In_852);
or U4275 (N_4275,In_2401,In_1680);
nor U4276 (N_4276,In_1019,In_2392);
nor U4277 (N_4277,In_91,In_2028);
or U4278 (N_4278,In_556,In_1854);
nor U4279 (N_4279,In_1807,In_685);
or U4280 (N_4280,In_1664,In_128);
nand U4281 (N_4281,In_2402,In_2131);
nor U4282 (N_4282,In_212,In_1025);
nand U4283 (N_4283,In_541,In_2177);
and U4284 (N_4284,In_1245,In_1324);
xor U4285 (N_4285,In_1113,In_2053);
xor U4286 (N_4286,In_1686,In_1662);
nand U4287 (N_4287,In_1723,In_676);
nand U4288 (N_4288,In_543,In_2006);
nand U4289 (N_4289,In_34,In_1707);
and U4290 (N_4290,In_1079,In_658);
nor U4291 (N_4291,In_2332,In_1455);
or U4292 (N_4292,In_519,In_55);
or U4293 (N_4293,In_1485,In_1994);
or U4294 (N_4294,In_1099,In_1726);
or U4295 (N_4295,In_269,In_2432);
nand U4296 (N_4296,In_1396,In_1818);
nor U4297 (N_4297,In_139,In_893);
and U4298 (N_4298,In_1003,In_1667);
and U4299 (N_4299,In_2316,In_835);
and U4300 (N_4300,In_885,In_2023);
and U4301 (N_4301,In_2372,In_1088);
nand U4302 (N_4302,In_1122,In_621);
and U4303 (N_4303,In_1048,In_1940);
xor U4304 (N_4304,In_1476,In_2387);
xor U4305 (N_4305,In_1023,In_1281);
nor U4306 (N_4306,In_1780,In_396);
and U4307 (N_4307,In_1490,In_1938);
and U4308 (N_4308,In_1568,In_633);
nor U4309 (N_4309,In_831,In_2346);
or U4310 (N_4310,In_2180,In_125);
nand U4311 (N_4311,In_1020,In_1652);
nor U4312 (N_4312,In_1365,In_1603);
and U4313 (N_4313,In_1099,In_565);
xnor U4314 (N_4314,In_1334,In_59);
and U4315 (N_4315,In_724,In_2429);
or U4316 (N_4316,In_2049,In_2291);
nand U4317 (N_4317,In_1380,In_482);
or U4318 (N_4318,In_1004,In_39);
nand U4319 (N_4319,In_2436,In_2373);
nor U4320 (N_4320,In_1714,In_1448);
nor U4321 (N_4321,In_2059,In_2047);
and U4322 (N_4322,In_327,In_1644);
or U4323 (N_4323,In_1957,In_1307);
and U4324 (N_4324,In_1986,In_1054);
nand U4325 (N_4325,In_1028,In_357);
and U4326 (N_4326,In_1993,In_1011);
nand U4327 (N_4327,In_2356,In_2133);
nor U4328 (N_4328,In_481,In_2366);
or U4329 (N_4329,In_1730,In_920);
xnor U4330 (N_4330,In_324,In_2428);
and U4331 (N_4331,In_96,In_629);
xnor U4332 (N_4332,In_811,In_1871);
or U4333 (N_4333,In_1660,In_1747);
or U4334 (N_4334,In_1096,In_1602);
or U4335 (N_4335,In_411,In_1976);
and U4336 (N_4336,In_1942,In_608);
or U4337 (N_4337,In_569,In_2466);
nor U4338 (N_4338,In_1361,In_698);
nor U4339 (N_4339,In_1726,In_1500);
nor U4340 (N_4340,In_1082,In_2074);
nand U4341 (N_4341,In_2408,In_2100);
nor U4342 (N_4342,In_39,In_102);
or U4343 (N_4343,In_1422,In_149);
nand U4344 (N_4344,In_2150,In_1582);
nor U4345 (N_4345,In_1964,In_1264);
or U4346 (N_4346,In_1015,In_1635);
or U4347 (N_4347,In_1135,In_1980);
nand U4348 (N_4348,In_798,In_2393);
xnor U4349 (N_4349,In_541,In_550);
or U4350 (N_4350,In_1942,In_1913);
nor U4351 (N_4351,In_76,In_215);
nand U4352 (N_4352,In_1738,In_339);
xor U4353 (N_4353,In_1821,In_15);
nor U4354 (N_4354,In_622,In_2176);
nand U4355 (N_4355,In_563,In_635);
or U4356 (N_4356,In_1987,In_414);
xnor U4357 (N_4357,In_973,In_432);
xnor U4358 (N_4358,In_1074,In_2370);
nand U4359 (N_4359,In_2089,In_1877);
nor U4360 (N_4360,In_1324,In_872);
or U4361 (N_4361,In_1927,In_2150);
nand U4362 (N_4362,In_91,In_1115);
and U4363 (N_4363,In_1135,In_1697);
and U4364 (N_4364,In_2478,In_460);
and U4365 (N_4365,In_369,In_121);
nand U4366 (N_4366,In_1728,In_2010);
or U4367 (N_4367,In_2014,In_52);
and U4368 (N_4368,In_2121,In_209);
nor U4369 (N_4369,In_362,In_1334);
xnor U4370 (N_4370,In_2178,In_2324);
nor U4371 (N_4371,In_2106,In_2386);
or U4372 (N_4372,In_1400,In_1858);
nand U4373 (N_4373,In_2478,In_113);
or U4374 (N_4374,In_435,In_42);
nand U4375 (N_4375,In_1075,In_2335);
nor U4376 (N_4376,In_1742,In_1380);
xor U4377 (N_4377,In_1310,In_1114);
nand U4378 (N_4378,In_345,In_367);
nand U4379 (N_4379,In_75,In_2180);
nor U4380 (N_4380,In_2036,In_26);
and U4381 (N_4381,In_20,In_1212);
nand U4382 (N_4382,In_610,In_1903);
and U4383 (N_4383,In_96,In_1312);
and U4384 (N_4384,In_1359,In_2163);
nand U4385 (N_4385,In_1725,In_839);
and U4386 (N_4386,In_65,In_407);
nor U4387 (N_4387,In_1428,In_1845);
xnor U4388 (N_4388,In_573,In_807);
nor U4389 (N_4389,In_436,In_864);
nand U4390 (N_4390,In_1213,In_1618);
nor U4391 (N_4391,In_1568,In_1453);
or U4392 (N_4392,In_421,In_1779);
xor U4393 (N_4393,In_2086,In_352);
nor U4394 (N_4394,In_1689,In_1548);
or U4395 (N_4395,In_747,In_2177);
or U4396 (N_4396,In_2170,In_2350);
or U4397 (N_4397,In_1791,In_1429);
and U4398 (N_4398,In_1163,In_80);
nand U4399 (N_4399,In_539,In_1889);
xnor U4400 (N_4400,In_1198,In_1265);
nand U4401 (N_4401,In_462,In_11);
nor U4402 (N_4402,In_693,In_64);
nor U4403 (N_4403,In_79,In_2211);
or U4404 (N_4404,In_252,In_245);
or U4405 (N_4405,In_28,In_695);
nor U4406 (N_4406,In_2141,In_1748);
nand U4407 (N_4407,In_2023,In_1512);
and U4408 (N_4408,In_1863,In_1101);
nand U4409 (N_4409,In_1820,In_1790);
nor U4410 (N_4410,In_1469,In_1642);
and U4411 (N_4411,In_2086,In_1280);
and U4412 (N_4412,In_2189,In_1065);
nor U4413 (N_4413,In_1505,In_2487);
and U4414 (N_4414,In_69,In_2373);
or U4415 (N_4415,In_432,In_734);
nor U4416 (N_4416,In_196,In_1140);
or U4417 (N_4417,In_1746,In_724);
nand U4418 (N_4418,In_1535,In_951);
xnor U4419 (N_4419,In_2065,In_1452);
xor U4420 (N_4420,In_1844,In_873);
nand U4421 (N_4421,In_457,In_1175);
or U4422 (N_4422,In_2376,In_1710);
or U4423 (N_4423,In_1978,In_854);
and U4424 (N_4424,In_1919,In_1024);
nand U4425 (N_4425,In_1516,In_1292);
and U4426 (N_4426,In_1672,In_2380);
nand U4427 (N_4427,In_1288,In_532);
or U4428 (N_4428,In_1637,In_500);
xnor U4429 (N_4429,In_2479,In_463);
or U4430 (N_4430,In_552,In_1814);
nor U4431 (N_4431,In_2426,In_1865);
nor U4432 (N_4432,In_996,In_754);
and U4433 (N_4433,In_1107,In_2154);
and U4434 (N_4434,In_659,In_453);
nand U4435 (N_4435,In_1007,In_1789);
nor U4436 (N_4436,In_11,In_1097);
nor U4437 (N_4437,In_1587,In_8);
and U4438 (N_4438,In_114,In_961);
nor U4439 (N_4439,In_401,In_1870);
nor U4440 (N_4440,In_2364,In_1662);
nand U4441 (N_4441,In_984,In_175);
nand U4442 (N_4442,In_2032,In_1050);
xnor U4443 (N_4443,In_332,In_1347);
and U4444 (N_4444,In_2147,In_403);
nand U4445 (N_4445,In_922,In_710);
and U4446 (N_4446,In_1319,In_919);
nand U4447 (N_4447,In_2434,In_2318);
and U4448 (N_4448,In_2001,In_1209);
or U4449 (N_4449,In_1494,In_224);
or U4450 (N_4450,In_410,In_1467);
nor U4451 (N_4451,In_979,In_444);
and U4452 (N_4452,In_1358,In_326);
or U4453 (N_4453,In_1227,In_127);
nor U4454 (N_4454,In_1456,In_1908);
nand U4455 (N_4455,In_1347,In_2329);
and U4456 (N_4456,In_2153,In_2227);
nor U4457 (N_4457,In_1471,In_870);
and U4458 (N_4458,In_138,In_488);
nor U4459 (N_4459,In_2137,In_1755);
nand U4460 (N_4460,In_70,In_28);
xnor U4461 (N_4461,In_2114,In_1319);
nor U4462 (N_4462,In_194,In_608);
nor U4463 (N_4463,In_2477,In_663);
nor U4464 (N_4464,In_2078,In_551);
and U4465 (N_4465,In_1192,In_1041);
nor U4466 (N_4466,In_1525,In_1546);
xnor U4467 (N_4467,In_434,In_1173);
nand U4468 (N_4468,In_1298,In_1498);
xnor U4469 (N_4469,In_1195,In_291);
and U4470 (N_4470,In_1764,In_1003);
and U4471 (N_4471,In_2280,In_453);
nor U4472 (N_4472,In_1497,In_700);
nor U4473 (N_4473,In_873,In_333);
nand U4474 (N_4474,In_1895,In_1913);
nor U4475 (N_4475,In_1897,In_979);
and U4476 (N_4476,In_839,In_2239);
nor U4477 (N_4477,In_2122,In_1021);
and U4478 (N_4478,In_604,In_742);
xor U4479 (N_4479,In_1178,In_2434);
and U4480 (N_4480,In_2163,In_2043);
xor U4481 (N_4481,In_72,In_2415);
and U4482 (N_4482,In_1400,In_603);
nand U4483 (N_4483,In_205,In_570);
or U4484 (N_4484,In_549,In_991);
xnor U4485 (N_4485,In_1443,In_1006);
and U4486 (N_4486,In_856,In_566);
nand U4487 (N_4487,In_2157,In_1275);
nor U4488 (N_4488,In_482,In_1009);
nand U4489 (N_4489,In_752,In_271);
or U4490 (N_4490,In_1364,In_1805);
or U4491 (N_4491,In_225,In_139);
and U4492 (N_4492,In_1126,In_1404);
nand U4493 (N_4493,In_462,In_1622);
or U4494 (N_4494,In_699,In_1166);
or U4495 (N_4495,In_1706,In_128);
nor U4496 (N_4496,In_61,In_938);
xor U4497 (N_4497,In_1860,In_124);
nor U4498 (N_4498,In_308,In_993);
and U4499 (N_4499,In_1026,In_1023);
or U4500 (N_4500,In_2081,In_801);
nand U4501 (N_4501,In_2216,In_2266);
nor U4502 (N_4502,In_360,In_930);
or U4503 (N_4503,In_2001,In_922);
or U4504 (N_4504,In_143,In_69);
or U4505 (N_4505,In_2444,In_1680);
nand U4506 (N_4506,In_2080,In_2288);
nand U4507 (N_4507,In_2037,In_1265);
xnor U4508 (N_4508,In_1807,In_2276);
and U4509 (N_4509,In_1874,In_495);
and U4510 (N_4510,In_2108,In_26);
nor U4511 (N_4511,In_183,In_48);
nor U4512 (N_4512,In_836,In_804);
and U4513 (N_4513,In_457,In_2460);
nand U4514 (N_4514,In_365,In_704);
nand U4515 (N_4515,In_692,In_2383);
nand U4516 (N_4516,In_1503,In_1380);
nand U4517 (N_4517,In_909,In_755);
and U4518 (N_4518,In_1826,In_923);
or U4519 (N_4519,In_1222,In_2248);
nand U4520 (N_4520,In_991,In_1471);
nand U4521 (N_4521,In_2343,In_587);
xnor U4522 (N_4522,In_147,In_1315);
nand U4523 (N_4523,In_1776,In_2469);
nor U4524 (N_4524,In_2386,In_2045);
nand U4525 (N_4525,In_894,In_2309);
nor U4526 (N_4526,In_2077,In_1779);
or U4527 (N_4527,In_445,In_1399);
nand U4528 (N_4528,In_1146,In_121);
and U4529 (N_4529,In_2141,In_1228);
and U4530 (N_4530,In_895,In_938);
or U4531 (N_4531,In_1654,In_2187);
xnor U4532 (N_4532,In_779,In_1832);
or U4533 (N_4533,In_1139,In_1835);
and U4534 (N_4534,In_2232,In_2280);
and U4535 (N_4535,In_1881,In_2298);
or U4536 (N_4536,In_756,In_1370);
nand U4537 (N_4537,In_984,In_2265);
and U4538 (N_4538,In_1770,In_1832);
nor U4539 (N_4539,In_783,In_1339);
and U4540 (N_4540,In_2396,In_2453);
nor U4541 (N_4541,In_578,In_1752);
nand U4542 (N_4542,In_579,In_1838);
nor U4543 (N_4543,In_2038,In_1);
and U4544 (N_4544,In_364,In_1538);
nor U4545 (N_4545,In_1020,In_854);
and U4546 (N_4546,In_647,In_155);
nor U4547 (N_4547,In_484,In_1403);
and U4548 (N_4548,In_114,In_2085);
or U4549 (N_4549,In_2053,In_397);
or U4550 (N_4550,In_2479,In_2028);
nor U4551 (N_4551,In_1623,In_1751);
xnor U4552 (N_4552,In_134,In_1132);
and U4553 (N_4553,In_1878,In_28);
or U4554 (N_4554,In_871,In_2156);
nor U4555 (N_4555,In_482,In_1382);
or U4556 (N_4556,In_999,In_950);
nand U4557 (N_4557,In_626,In_993);
nand U4558 (N_4558,In_2432,In_1966);
nor U4559 (N_4559,In_1108,In_249);
or U4560 (N_4560,In_1159,In_959);
nor U4561 (N_4561,In_1975,In_116);
and U4562 (N_4562,In_1424,In_1806);
or U4563 (N_4563,In_1075,In_1100);
xnor U4564 (N_4564,In_2415,In_267);
and U4565 (N_4565,In_1316,In_1857);
nor U4566 (N_4566,In_2405,In_812);
xor U4567 (N_4567,In_782,In_629);
nand U4568 (N_4568,In_1680,In_1858);
or U4569 (N_4569,In_304,In_2363);
or U4570 (N_4570,In_891,In_214);
or U4571 (N_4571,In_1708,In_2302);
nor U4572 (N_4572,In_880,In_194);
nand U4573 (N_4573,In_2351,In_2271);
nand U4574 (N_4574,In_965,In_2189);
nor U4575 (N_4575,In_887,In_1158);
nor U4576 (N_4576,In_1374,In_1596);
nor U4577 (N_4577,In_434,In_2233);
or U4578 (N_4578,In_2483,In_2023);
or U4579 (N_4579,In_2400,In_738);
or U4580 (N_4580,In_1529,In_2333);
xnor U4581 (N_4581,In_1299,In_1552);
and U4582 (N_4582,In_1906,In_353);
xnor U4583 (N_4583,In_599,In_1731);
or U4584 (N_4584,In_161,In_52);
nand U4585 (N_4585,In_2302,In_1382);
nand U4586 (N_4586,In_2158,In_1668);
or U4587 (N_4587,In_1737,In_975);
nand U4588 (N_4588,In_1475,In_882);
nand U4589 (N_4589,In_1777,In_1711);
and U4590 (N_4590,In_45,In_1808);
nor U4591 (N_4591,In_371,In_675);
nor U4592 (N_4592,In_24,In_1997);
and U4593 (N_4593,In_1418,In_558);
and U4594 (N_4594,In_1870,In_2495);
xor U4595 (N_4595,In_291,In_1992);
nor U4596 (N_4596,In_2124,In_1206);
xnor U4597 (N_4597,In_1403,In_647);
nor U4598 (N_4598,In_887,In_1362);
or U4599 (N_4599,In_87,In_1082);
and U4600 (N_4600,In_1959,In_1516);
and U4601 (N_4601,In_1208,In_1388);
nor U4602 (N_4602,In_1160,In_1384);
and U4603 (N_4603,In_123,In_1601);
nor U4604 (N_4604,In_2376,In_385);
xnor U4605 (N_4605,In_763,In_880);
nor U4606 (N_4606,In_1726,In_1094);
or U4607 (N_4607,In_385,In_1569);
nand U4608 (N_4608,In_2248,In_987);
and U4609 (N_4609,In_1673,In_1963);
nor U4610 (N_4610,In_568,In_1631);
and U4611 (N_4611,In_1327,In_2051);
nor U4612 (N_4612,In_1259,In_1329);
and U4613 (N_4613,In_789,In_1618);
or U4614 (N_4614,In_1453,In_895);
nor U4615 (N_4615,In_80,In_1247);
and U4616 (N_4616,In_1120,In_385);
or U4617 (N_4617,In_2263,In_1561);
or U4618 (N_4618,In_890,In_1880);
or U4619 (N_4619,In_387,In_1723);
nor U4620 (N_4620,In_2450,In_1136);
nand U4621 (N_4621,In_683,In_1730);
nor U4622 (N_4622,In_1936,In_2122);
nor U4623 (N_4623,In_257,In_577);
nand U4624 (N_4624,In_1439,In_101);
nand U4625 (N_4625,In_1770,In_2196);
nand U4626 (N_4626,In_647,In_1383);
or U4627 (N_4627,In_1892,In_1706);
and U4628 (N_4628,In_987,In_1489);
or U4629 (N_4629,In_528,In_1532);
nand U4630 (N_4630,In_1970,In_1759);
or U4631 (N_4631,In_1795,In_630);
and U4632 (N_4632,In_326,In_2306);
xor U4633 (N_4633,In_2114,In_423);
nor U4634 (N_4634,In_1554,In_1668);
nor U4635 (N_4635,In_2343,In_291);
xnor U4636 (N_4636,In_774,In_1344);
or U4637 (N_4637,In_894,In_1836);
and U4638 (N_4638,In_875,In_988);
and U4639 (N_4639,In_264,In_1565);
or U4640 (N_4640,In_1441,In_1755);
or U4641 (N_4641,In_1318,In_1435);
or U4642 (N_4642,In_34,In_2028);
and U4643 (N_4643,In_1946,In_636);
and U4644 (N_4644,In_2213,In_1795);
and U4645 (N_4645,In_390,In_2428);
and U4646 (N_4646,In_1641,In_1627);
nor U4647 (N_4647,In_1082,In_2142);
nor U4648 (N_4648,In_1089,In_2360);
or U4649 (N_4649,In_1244,In_448);
nand U4650 (N_4650,In_1582,In_410);
nor U4651 (N_4651,In_1629,In_1794);
nor U4652 (N_4652,In_1196,In_402);
nor U4653 (N_4653,In_1295,In_1849);
nand U4654 (N_4654,In_1123,In_2429);
xnor U4655 (N_4655,In_2468,In_2498);
or U4656 (N_4656,In_1686,In_173);
nor U4657 (N_4657,In_624,In_1102);
and U4658 (N_4658,In_1800,In_1062);
and U4659 (N_4659,In_1771,In_1993);
or U4660 (N_4660,In_1821,In_1950);
and U4661 (N_4661,In_939,In_1);
nor U4662 (N_4662,In_261,In_2342);
xor U4663 (N_4663,In_2098,In_1120);
xnor U4664 (N_4664,In_1526,In_2368);
or U4665 (N_4665,In_803,In_1280);
nand U4666 (N_4666,In_1365,In_750);
xor U4667 (N_4667,In_1239,In_1878);
nand U4668 (N_4668,In_248,In_576);
and U4669 (N_4669,In_1410,In_285);
nor U4670 (N_4670,In_141,In_2420);
xnor U4671 (N_4671,In_426,In_842);
nor U4672 (N_4672,In_131,In_208);
and U4673 (N_4673,In_1326,In_2016);
nor U4674 (N_4674,In_587,In_1537);
nor U4675 (N_4675,In_2123,In_1638);
and U4676 (N_4676,In_1374,In_1842);
or U4677 (N_4677,In_351,In_357);
nor U4678 (N_4678,In_1420,In_196);
nand U4679 (N_4679,In_2278,In_2109);
nand U4680 (N_4680,In_1699,In_77);
nand U4681 (N_4681,In_1323,In_2121);
xor U4682 (N_4682,In_2313,In_1796);
nand U4683 (N_4683,In_2396,In_1368);
or U4684 (N_4684,In_814,In_873);
nand U4685 (N_4685,In_2327,In_156);
nor U4686 (N_4686,In_860,In_714);
or U4687 (N_4687,In_1733,In_1462);
nor U4688 (N_4688,In_1724,In_986);
nor U4689 (N_4689,In_1307,In_1278);
nand U4690 (N_4690,In_2468,In_2411);
nor U4691 (N_4691,In_2391,In_2237);
nor U4692 (N_4692,In_23,In_689);
or U4693 (N_4693,In_691,In_1893);
or U4694 (N_4694,In_1293,In_43);
and U4695 (N_4695,In_1210,In_970);
or U4696 (N_4696,In_926,In_81);
and U4697 (N_4697,In_1907,In_71);
nor U4698 (N_4698,In_2459,In_62);
or U4699 (N_4699,In_473,In_498);
nor U4700 (N_4700,In_1719,In_811);
and U4701 (N_4701,In_2047,In_366);
or U4702 (N_4702,In_174,In_603);
nor U4703 (N_4703,In_1868,In_783);
nor U4704 (N_4704,In_513,In_2137);
and U4705 (N_4705,In_238,In_1392);
nor U4706 (N_4706,In_644,In_83);
and U4707 (N_4707,In_2278,In_1491);
nand U4708 (N_4708,In_752,In_433);
and U4709 (N_4709,In_1390,In_717);
nor U4710 (N_4710,In_2419,In_1327);
nand U4711 (N_4711,In_1339,In_1538);
nand U4712 (N_4712,In_2398,In_795);
and U4713 (N_4713,In_1557,In_1370);
nor U4714 (N_4714,In_1215,In_953);
xor U4715 (N_4715,In_83,In_1892);
nand U4716 (N_4716,In_683,In_2000);
xor U4717 (N_4717,In_861,In_2104);
or U4718 (N_4718,In_922,In_408);
nand U4719 (N_4719,In_641,In_149);
nand U4720 (N_4720,In_1787,In_2404);
nor U4721 (N_4721,In_1096,In_1802);
or U4722 (N_4722,In_752,In_292);
xnor U4723 (N_4723,In_43,In_401);
and U4724 (N_4724,In_577,In_2121);
nand U4725 (N_4725,In_469,In_1789);
and U4726 (N_4726,In_581,In_1922);
and U4727 (N_4727,In_1061,In_1452);
nand U4728 (N_4728,In_1948,In_476);
or U4729 (N_4729,In_122,In_1942);
nor U4730 (N_4730,In_2163,In_2423);
or U4731 (N_4731,In_1970,In_232);
or U4732 (N_4732,In_528,In_438);
or U4733 (N_4733,In_1589,In_1366);
nor U4734 (N_4734,In_1694,In_149);
nand U4735 (N_4735,In_238,In_249);
and U4736 (N_4736,In_1261,In_2434);
nor U4737 (N_4737,In_758,In_2488);
or U4738 (N_4738,In_780,In_759);
nand U4739 (N_4739,In_1871,In_1929);
or U4740 (N_4740,In_58,In_2448);
and U4741 (N_4741,In_382,In_461);
and U4742 (N_4742,In_2092,In_175);
nor U4743 (N_4743,In_239,In_1431);
nor U4744 (N_4744,In_1680,In_1078);
and U4745 (N_4745,In_1377,In_2124);
nand U4746 (N_4746,In_392,In_2234);
nand U4747 (N_4747,In_912,In_1132);
nor U4748 (N_4748,In_1020,In_887);
nand U4749 (N_4749,In_1036,In_2341);
nand U4750 (N_4750,In_1149,In_264);
xnor U4751 (N_4751,In_1851,In_1847);
nand U4752 (N_4752,In_1053,In_2142);
nand U4753 (N_4753,In_465,In_76);
nor U4754 (N_4754,In_412,In_1666);
nand U4755 (N_4755,In_1226,In_2257);
and U4756 (N_4756,In_1852,In_1781);
and U4757 (N_4757,In_1519,In_706);
nor U4758 (N_4758,In_2089,In_2152);
or U4759 (N_4759,In_1633,In_626);
nor U4760 (N_4760,In_918,In_859);
nand U4761 (N_4761,In_32,In_576);
and U4762 (N_4762,In_520,In_355);
nor U4763 (N_4763,In_2118,In_1753);
nand U4764 (N_4764,In_1145,In_317);
nand U4765 (N_4765,In_324,In_634);
nor U4766 (N_4766,In_1679,In_2390);
nor U4767 (N_4767,In_2410,In_1059);
nand U4768 (N_4768,In_1636,In_966);
or U4769 (N_4769,In_1260,In_1826);
nand U4770 (N_4770,In_282,In_1139);
and U4771 (N_4771,In_1601,In_1037);
nor U4772 (N_4772,In_777,In_1577);
or U4773 (N_4773,In_328,In_1125);
or U4774 (N_4774,In_1582,In_1237);
and U4775 (N_4775,In_1505,In_75);
nor U4776 (N_4776,In_1230,In_1217);
nor U4777 (N_4777,In_263,In_1729);
nand U4778 (N_4778,In_1994,In_544);
nor U4779 (N_4779,In_269,In_204);
nor U4780 (N_4780,In_649,In_584);
and U4781 (N_4781,In_688,In_1834);
nor U4782 (N_4782,In_806,In_173);
nor U4783 (N_4783,In_1330,In_2221);
nand U4784 (N_4784,In_1884,In_2217);
and U4785 (N_4785,In_2369,In_1700);
xor U4786 (N_4786,In_2083,In_1804);
nor U4787 (N_4787,In_499,In_949);
nor U4788 (N_4788,In_1794,In_97);
nor U4789 (N_4789,In_424,In_859);
nand U4790 (N_4790,In_1439,In_1328);
xor U4791 (N_4791,In_1038,In_731);
nand U4792 (N_4792,In_1941,In_411);
nand U4793 (N_4793,In_2157,In_1273);
xnor U4794 (N_4794,In_1827,In_1853);
or U4795 (N_4795,In_1351,In_1307);
nor U4796 (N_4796,In_1784,In_2150);
nor U4797 (N_4797,In_191,In_1154);
nand U4798 (N_4798,In_508,In_1492);
nand U4799 (N_4799,In_1901,In_1298);
nand U4800 (N_4800,In_1073,In_1260);
xor U4801 (N_4801,In_1243,In_1274);
nor U4802 (N_4802,In_1660,In_62);
and U4803 (N_4803,In_605,In_1787);
nand U4804 (N_4804,In_1246,In_712);
nor U4805 (N_4805,In_1352,In_797);
nand U4806 (N_4806,In_140,In_1600);
xnor U4807 (N_4807,In_1816,In_790);
or U4808 (N_4808,In_293,In_1436);
or U4809 (N_4809,In_163,In_697);
nand U4810 (N_4810,In_2324,In_119);
nor U4811 (N_4811,In_202,In_360);
and U4812 (N_4812,In_1625,In_2114);
and U4813 (N_4813,In_1235,In_249);
nand U4814 (N_4814,In_1437,In_1967);
and U4815 (N_4815,In_2490,In_202);
nand U4816 (N_4816,In_26,In_1088);
nor U4817 (N_4817,In_1826,In_261);
nand U4818 (N_4818,In_1907,In_268);
xnor U4819 (N_4819,In_673,In_2126);
or U4820 (N_4820,In_1087,In_539);
or U4821 (N_4821,In_1542,In_1960);
nor U4822 (N_4822,In_1687,In_2488);
and U4823 (N_4823,In_1956,In_1334);
nand U4824 (N_4824,In_121,In_2015);
nor U4825 (N_4825,In_936,In_219);
nand U4826 (N_4826,In_1776,In_1052);
xor U4827 (N_4827,In_1702,In_341);
xnor U4828 (N_4828,In_1096,In_1855);
nor U4829 (N_4829,In_1384,In_2131);
and U4830 (N_4830,In_1025,In_1999);
xor U4831 (N_4831,In_518,In_1638);
or U4832 (N_4832,In_2217,In_1631);
and U4833 (N_4833,In_1742,In_106);
or U4834 (N_4834,In_35,In_977);
xor U4835 (N_4835,In_2306,In_2134);
and U4836 (N_4836,In_963,In_92);
and U4837 (N_4837,In_1240,In_370);
or U4838 (N_4838,In_738,In_1208);
or U4839 (N_4839,In_1848,In_875);
or U4840 (N_4840,In_2086,In_1583);
nor U4841 (N_4841,In_1025,In_1651);
nor U4842 (N_4842,In_2040,In_1782);
or U4843 (N_4843,In_1116,In_1424);
or U4844 (N_4844,In_391,In_1940);
nand U4845 (N_4845,In_1920,In_2438);
and U4846 (N_4846,In_2274,In_1357);
and U4847 (N_4847,In_549,In_2486);
xnor U4848 (N_4848,In_1212,In_2488);
xor U4849 (N_4849,In_187,In_480);
xor U4850 (N_4850,In_1999,In_1837);
nand U4851 (N_4851,In_1219,In_329);
nor U4852 (N_4852,In_1825,In_2409);
nand U4853 (N_4853,In_905,In_1937);
or U4854 (N_4854,In_766,In_1913);
nor U4855 (N_4855,In_1630,In_519);
nor U4856 (N_4856,In_2464,In_1894);
xor U4857 (N_4857,In_1044,In_617);
nor U4858 (N_4858,In_777,In_152);
nand U4859 (N_4859,In_2057,In_857);
xnor U4860 (N_4860,In_1903,In_1146);
nor U4861 (N_4861,In_1538,In_2382);
and U4862 (N_4862,In_2182,In_2228);
and U4863 (N_4863,In_499,In_682);
nor U4864 (N_4864,In_719,In_171);
nand U4865 (N_4865,In_918,In_829);
and U4866 (N_4866,In_2258,In_1485);
nor U4867 (N_4867,In_535,In_1175);
and U4868 (N_4868,In_545,In_1787);
or U4869 (N_4869,In_375,In_729);
nand U4870 (N_4870,In_1590,In_1172);
nand U4871 (N_4871,In_2313,In_1690);
nor U4872 (N_4872,In_1936,In_2429);
and U4873 (N_4873,In_568,In_2395);
and U4874 (N_4874,In_378,In_1847);
nor U4875 (N_4875,In_2039,In_1588);
nand U4876 (N_4876,In_1195,In_1210);
xor U4877 (N_4877,In_1199,In_174);
nand U4878 (N_4878,In_1040,In_2341);
nor U4879 (N_4879,In_1871,In_662);
and U4880 (N_4880,In_2486,In_451);
or U4881 (N_4881,In_1296,In_1471);
and U4882 (N_4882,In_2231,In_1867);
xnor U4883 (N_4883,In_627,In_260);
nor U4884 (N_4884,In_2350,In_167);
nor U4885 (N_4885,In_1452,In_1149);
xnor U4886 (N_4886,In_604,In_129);
or U4887 (N_4887,In_868,In_1138);
or U4888 (N_4888,In_1371,In_1844);
xor U4889 (N_4889,In_570,In_1562);
xor U4890 (N_4890,In_977,In_1976);
nand U4891 (N_4891,In_1132,In_2157);
nor U4892 (N_4892,In_862,In_899);
and U4893 (N_4893,In_112,In_1874);
nand U4894 (N_4894,In_621,In_684);
and U4895 (N_4895,In_1469,In_1229);
xnor U4896 (N_4896,In_1033,In_252);
and U4897 (N_4897,In_838,In_1381);
or U4898 (N_4898,In_1051,In_509);
nand U4899 (N_4899,In_654,In_1227);
xor U4900 (N_4900,In_2089,In_281);
and U4901 (N_4901,In_2170,In_2004);
and U4902 (N_4902,In_2394,In_203);
or U4903 (N_4903,In_1368,In_91);
and U4904 (N_4904,In_1597,In_135);
and U4905 (N_4905,In_592,In_120);
xnor U4906 (N_4906,In_20,In_1553);
nor U4907 (N_4907,In_2059,In_661);
or U4908 (N_4908,In_2149,In_1451);
or U4909 (N_4909,In_1384,In_1425);
or U4910 (N_4910,In_327,In_308);
and U4911 (N_4911,In_496,In_1663);
and U4912 (N_4912,In_1972,In_1715);
and U4913 (N_4913,In_870,In_2186);
and U4914 (N_4914,In_2464,In_2051);
xnor U4915 (N_4915,In_450,In_1540);
nand U4916 (N_4916,In_222,In_1067);
nand U4917 (N_4917,In_2419,In_2168);
xnor U4918 (N_4918,In_891,In_1612);
or U4919 (N_4919,In_363,In_2380);
nor U4920 (N_4920,In_2426,In_1989);
and U4921 (N_4921,In_93,In_2215);
nor U4922 (N_4922,In_2200,In_2273);
nand U4923 (N_4923,In_1409,In_1955);
or U4924 (N_4924,In_1708,In_1616);
xnor U4925 (N_4925,In_241,In_2043);
or U4926 (N_4926,In_2367,In_2093);
or U4927 (N_4927,In_1463,In_1301);
and U4928 (N_4928,In_2233,In_2499);
or U4929 (N_4929,In_2423,In_777);
or U4930 (N_4930,In_1538,In_1785);
nand U4931 (N_4931,In_410,In_1047);
and U4932 (N_4932,In_1285,In_2495);
xnor U4933 (N_4933,In_1119,In_412);
and U4934 (N_4934,In_1275,In_2398);
or U4935 (N_4935,In_1840,In_902);
nor U4936 (N_4936,In_2271,In_2218);
nand U4937 (N_4937,In_2237,In_1914);
nor U4938 (N_4938,In_1667,In_1761);
nand U4939 (N_4939,In_1158,In_602);
and U4940 (N_4940,In_1913,In_556);
and U4941 (N_4941,In_1949,In_2376);
nand U4942 (N_4942,In_1406,In_484);
nor U4943 (N_4943,In_1030,In_777);
nand U4944 (N_4944,In_1675,In_2279);
xor U4945 (N_4945,In_1763,In_672);
nand U4946 (N_4946,In_514,In_376);
nor U4947 (N_4947,In_1191,In_1045);
nor U4948 (N_4948,In_239,In_884);
nand U4949 (N_4949,In_419,In_129);
and U4950 (N_4950,In_1099,In_2159);
or U4951 (N_4951,In_2322,In_1775);
and U4952 (N_4952,In_1136,In_436);
and U4953 (N_4953,In_742,In_550);
nand U4954 (N_4954,In_530,In_2475);
and U4955 (N_4955,In_1057,In_466);
and U4956 (N_4956,In_1632,In_228);
or U4957 (N_4957,In_1142,In_2485);
xnor U4958 (N_4958,In_90,In_862);
nor U4959 (N_4959,In_1206,In_226);
nor U4960 (N_4960,In_863,In_1927);
nand U4961 (N_4961,In_1797,In_2117);
and U4962 (N_4962,In_457,In_2115);
and U4963 (N_4963,In_972,In_177);
nand U4964 (N_4964,In_1722,In_1719);
xnor U4965 (N_4965,In_2102,In_1777);
nand U4966 (N_4966,In_88,In_2221);
xnor U4967 (N_4967,In_1273,In_2209);
nand U4968 (N_4968,In_2005,In_494);
nor U4969 (N_4969,In_1932,In_1851);
and U4970 (N_4970,In_575,In_647);
nor U4971 (N_4971,In_731,In_1385);
nor U4972 (N_4972,In_2016,In_2192);
nor U4973 (N_4973,In_1825,In_1700);
or U4974 (N_4974,In_924,In_363);
nand U4975 (N_4975,In_679,In_2097);
nand U4976 (N_4976,In_2093,In_2114);
or U4977 (N_4977,In_1785,In_91);
nand U4978 (N_4978,In_1987,In_911);
nor U4979 (N_4979,In_1343,In_315);
and U4980 (N_4980,In_2111,In_243);
xnor U4981 (N_4981,In_2394,In_473);
or U4982 (N_4982,In_2082,In_1473);
or U4983 (N_4983,In_1262,In_1529);
and U4984 (N_4984,In_1625,In_425);
xor U4985 (N_4985,In_1955,In_2342);
xor U4986 (N_4986,In_694,In_951);
and U4987 (N_4987,In_628,In_1830);
nand U4988 (N_4988,In_399,In_1028);
nor U4989 (N_4989,In_2057,In_431);
and U4990 (N_4990,In_1830,In_1078);
nand U4991 (N_4991,In_590,In_571);
or U4992 (N_4992,In_2171,In_1561);
nor U4993 (N_4993,In_1262,In_1462);
xor U4994 (N_4994,In_1444,In_59);
xor U4995 (N_4995,In_395,In_175);
nand U4996 (N_4996,In_2484,In_2427);
and U4997 (N_4997,In_908,In_806);
nand U4998 (N_4998,In_2321,In_1893);
and U4999 (N_4999,In_825,In_931);
and U5000 (N_5000,In_2428,In_1895);
nand U5001 (N_5001,In_2298,In_1080);
nor U5002 (N_5002,In_1263,In_2210);
nor U5003 (N_5003,In_402,In_376);
nand U5004 (N_5004,In_136,In_2277);
nor U5005 (N_5005,In_1120,In_950);
xor U5006 (N_5006,In_2095,In_1621);
or U5007 (N_5007,In_351,In_733);
or U5008 (N_5008,In_2284,In_1736);
nand U5009 (N_5009,In_1972,In_140);
or U5010 (N_5010,In_1007,In_1313);
nor U5011 (N_5011,In_2332,In_1822);
or U5012 (N_5012,In_1132,In_2194);
xor U5013 (N_5013,In_153,In_119);
or U5014 (N_5014,In_2471,In_202);
or U5015 (N_5015,In_1059,In_1643);
or U5016 (N_5016,In_75,In_1749);
and U5017 (N_5017,In_736,In_1210);
or U5018 (N_5018,In_104,In_2275);
nor U5019 (N_5019,In_181,In_2185);
nand U5020 (N_5020,In_869,In_563);
and U5021 (N_5021,In_2440,In_1807);
nand U5022 (N_5022,In_690,In_2337);
nand U5023 (N_5023,In_2150,In_1244);
and U5024 (N_5024,In_2493,In_616);
nor U5025 (N_5025,In_185,In_1890);
xnor U5026 (N_5026,In_1539,In_956);
and U5027 (N_5027,In_1524,In_1650);
or U5028 (N_5028,In_1211,In_2272);
nor U5029 (N_5029,In_1641,In_2096);
or U5030 (N_5030,In_1232,In_1443);
and U5031 (N_5031,In_2495,In_2027);
and U5032 (N_5032,In_1203,In_2427);
and U5033 (N_5033,In_90,In_1753);
or U5034 (N_5034,In_1342,In_415);
xnor U5035 (N_5035,In_12,In_1373);
nand U5036 (N_5036,In_413,In_760);
nand U5037 (N_5037,In_1746,In_2106);
or U5038 (N_5038,In_1136,In_187);
nor U5039 (N_5039,In_2307,In_35);
and U5040 (N_5040,In_947,In_945);
and U5041 (N_5041,In_2432,In_1594);
nand U5042 (N_5042,In_905,In_1954);
or U5043 (N_5043,In_2392,In_1215);
nor U5044 (N_5044,In_1902,In_611);
nor U5045 (N_5045,In_40,In_1468);
or U5046 (N_5046,In_608,In_554);
or U5047 (N_5047,In_1452,In_2481);
and U5048 (N_5048,In_2086,In_913);
xor U5049 (N_5049,In_1696,In_1290);
or U5050 (N_5050,In_2385,In_1365);
nor U5051 (N_5051,In_1839,In_2329);
or U5052 (N_5052,In_31,In_2434);
nand U5053 (N_5053,In_125,In_118);
xnor U5054 (N_5054,In_1233,In_1958);
and U5055 (N_5055,In_2366,In_1340);
xnor U5056 (N_5056,In_1770,In_2067);
nand U5057 (N_5057,In_1086,In_861);
nand U5058 (N_5058,In_352,In_246);
and U5059 (N_5059,In_235,In_319);
nand U5060 (N_5060,In_2020,In_146);
nor U5061 (N_5061,In_1806,In_2137);
and U5062 (N_5062,In_1545,In_1419);
nor U5063 (N_5063,In_162,In_576);
nor U5064 (N_5064,In_1060,In_941);
nand U5065 (N_5065,In_120,In_268);
xnor U5066 (N_5066,In_1185,In_45);
and U5067 (N_5067,In_37,In_9);
or U5068 (N_5068,In_268,In_536);
or U5069 (N_5069,In_190,In_1115);
or U5070 (N_5070,In_1941,In_1775);
nor U5071 (N_5071,In_1698,In_940);
and U5072 (N_5072,In_1136,In_2406);
or U5073 (N_5073,In_192,In_2051);
or U5074 (N_5074,In_493,In_1660);
xor U5075 (N_5075,In_844,In_2270);
nand U5076 (N_5076,In_2477,In_840);
and U5077 (N_5077,In_1662,In_1988);
nor U5078 (N_5078,In_1476,In_579);
and U5079 (N_5079,In_2333,In_1023);
nand U5080 (N_5080,In_2306,In_1841);
nand U5081 (N_5081,In_1443,In_1193);
or U5082 (N_5082,In_1202,In_2484);
nand U5083 (N_5083,In_290,In_1831);
nor U5084 (N_5084,In_1169,In_42);
or U5085 (N_5085,In_1347,In_2399);
and U5086 (N_5086,In_177,In_1756);
nor U5087 (N_5087,In_202,In_1010);
nand U5088 (N_5088,In_683,In_160);
nand U5089 (N_5089,In_2113,In_1297);
and U5090 (N_5090,In_2160,In_1527);
or U5091 (N_5091,In_1233,In_451);
or U5092 (N_5092,In_140,In_2489);
or U5093 (N_5093,In_1143,In_1512);
or U5094 (N_5094,In_155,In_168);
or U5095 (N_5095,In_510,In_1208);
nor U5096 (N_5096,In_1288,In_1701);
nor U5097 (N_5097,In_2360,In_586);
xor U5098 (N_5098,In_1890,In_696);
and U5099 (N_5099,In_655,In_2465);
or U5100 (N_5100,In_613,In_983);
or U5101 (N_5101,In_668,In_314);
nor U5102 (N_5102,In_874,In_619);
nor U5103 (N_5103,In_1466,In_786);
or U5104 (N_5104,In_2293,In_1231);
nor U5105 (N_5105,In_154,In_1505);
and U5106 (N_5106,In_1730,In_375);
nor U5107 (N_5107,In_1009,In_873);
nand U5108 (N_5108,In_2318,In_648);
nor U5109 (N_5109,In_918,In_948);
nor U5110 (N_5110,In_1726,In_1433);
nor U5111 (N_5111,In_1221,In_37);
nand U5112 (N_5112,In_719,In_2259);
nor U5113 (N_5113,In_803,In_239);
nand U5114 (N_5114,In_613,In_1902);
or U5115 (N_5115,In_466,In_219);
and U5116 (N_5116,In_1278,In_705);
or U5117 (N_5117,In_1030,In_1811);
or U5118 (N_5118,In_1135,In_447);
and U5119 (N_5119,In_555,In_1485);
nand U5120 (N_5120,In_1139,In_388);
nand U5121 (N_5121,In_474,In_1390);
nor U5122 (N_5122,In_480,In_1230);
nor U5123 (N_5123,In_1552,In_2393);
or U5124 (N_5124,In_1662,In_2469);
or U5125 (N_5125,In_2403,In_220);
or U5126 (N_5126,In_1003,In_2294);
nand U5127 (N_5127,In_841,In_2021);
nor U5128 (N_5128,In_2279,In_2154);
or U5129 (N_5129,In_1803,In_540);
nor U5130 (N_5130,In_249,In_1943);
xor U5131 (N_5131,In_1517,In_1460);
nand U5132 (N_5132,In_1424,In_1824);
nor U5133 (N_5133,In_1703,In_111);
nor U5134 (N_5134,In_30,In_2150);
nand U5135 (N_5135,In_24,In_1675);
and U5136 (N_5136,In_510,In_1147);
nand U5137 (N_5137,In_391,In_90);
or U5138 (N_5138,In_1583,In_1928);
and U5139 (N_5139,In_1538,In_498);
and U5140 (N_5140,In_1006,In_1310);
and U5141 (N_5141,In_1637,In_2131);
nor U5142 (N_5142,In_2409,In_363);
and U5143 (N_5143,In_503,In_123);
or U5144 (N_5144,In_1412,In_1693);
nand U5145 (N_5145,In_771,In_1217);
or U5146 (N_5146,In_2141,In_2334);
nor U5147 (N_5147,In_1118,In_961);
or U5148 (N_5148,In_1230,In_2323);
or U5149 (N_5149,In_783,In_2341);
xnor U5150 (N_5150,In_1972,In_1385);
and U5151 (N_5151,In_1615,In_1875);
or U5152 (N_5152,In_1142,In_736);
xor U5153 (N_5153,In_1758,In_871);
xor U5154 (N_5154,In_117,In_1667);
nor U5155 (N_5155,In_855,In_32);
and U5156 (N_5156,In_1425,In_1405);
and U5157 (N_5157,In_1184,In_845);
and U5158 (N_5158,In_732,In_1442);
nor U5159 (N_5159,In_420,In_1336);
nor U5160 (N_5160,In_199,In_1044);
nor U5161 (N_5161,In_2107,In_475);
nor U5162 (N_5162,In_504,In_744);
and U5163 (N_5163,In_1680,In_457);
nor U5164 (N_5164,In_314,In_839);
nand U5165 (N_5165,In_2057,In_257);
and U5166 (N_5166,In_389,In_1235);
and U5167 (N_5167,In_2107,In_529);
or U5168 (N_5168,In_1865,In_1714);
and U5169 (N_5169,In_2280,In_1879);
and U5170 (N_5170,In_1812,In_444);
and U5171 (N_5171,In_2328,In_1715);
or U5172 (N_5172,In_1087,In_981);
xor U5173 (N_5173,In_2002,In_2280);
nor U5174 (N_5174,In_2088,In_1742);
nand U5175 (N_5175,In_155,In_2362);
nand U5176 (N_5176,In_2027,In_1120);
or U5177 (N_5177,In_716,In_430);
nor U5178 (N_5178,In_1671,In_653);
or U5179 (N_5179,In_38,In_1663);
nand U5180 (N_5180,In_1437,In_1817);
or U5181 (N_5181,In_960,In_1798);
nand U5182 (N_5182,In_1655,In_1013);
nand U5183 (N_5183,In_572,In_143);
xor U5184 (N_5184,In_2069,In_185);
nand U5185 (N_5185,In_1396,In_1914);
or U5186 (N_5186,In_357,In_1080);
or U5187 (N_5187,In_1457,In_634);
nor U5188 (N_5188,In_2208,In_831);
or U5189 (N_5189,In_1723,In_1605);
nand U5190 (N_5190,In_1512,In_713);
and U5191 (N_5191,In_353,In_2407);
nand U5192 (N_5192,In_618,In_598);
and U5193 (N_5193,In_575,In_233);
xor U5194 (N_5194,In_1198,In_1000);
nor U5195 (N_5195,In_1995,In_377);
or U5196 (N_5196,In_811,In_1244);
nor U5197 (N_5197,In_1735,In_1427);
nor U5198 (N_5198,In_1507,In_951);
and U5199 (N_5199,In_1298,In_1843);
or U5200 (N_5200,In_2150,In_1884);
nand U5201 (N_5201,In_1976,In_1305);
nor U5202 (N_5202,In_1554,In_356);
and U5203 (N_5203,In_1015,In_2399);
and U5204 (N_5204,In_180,In_590);
and U5205 (N_5205,In_1268,In_224);
nand U5206 (N_5206,In_1251,In_2383);
nor U5207 (N_5207,In_297,In_923);
nand U5208 (N_5208,In_1893,In_1268);
nand U5209 (N_5209,In_885,In_1129);
or U5210 (N_5210,In_2181,In_1250);
and U5211 (N_5211,In_200,In_1897);
and U5212 (N_5212,In_2473,In_334);
xor U5213 (N_5213,In_1899,In_1577);
or U5214 (N_5214,In_896,In_653);
and U5215 (N_5215,In_1732,In_1674);
xnor U5216 (N_5216,In_1519,In_2264);
and U5217 (N_5217,In_1837,In_2447);
nand U5218 (N_5218,In_2067,In_1197);
or U5219 (N_5219,In_655,In_1277);
nand U5220 (N_5220,In_1392,In_331);
nand U5221 (N_5221,In_1497,In_1114);
xnor U5222 (N_5222,In_361,In_83);
xnor U5223 (N_5223,In_2426,In_216);
nand U5224 (N_5224,In_1282,In_1566);
and U5225 (N_5225,In_1667,In_1743);
and U5226 (N_5226,In_1877,In_1209);
nor U5227 (N_5227,In_2130,In_20);
and U5228 (N_5228,In_835,In_1540);
nand U5229 (N_5229,In_1737,In_2083);
xor U5230 (N_5230,In_1939,In_2095);
nor U5231 (N_5231,In_91,In_21);
nor U5232 (N_5232,In_1187,In_2078);
nand U5233 (N_5233,In_1859,In_477);
and U5234 (N_5234,In_2209,In_1016);
or U5235 (N_5235,In_238,In_1021);
nor U5236 (N_5236,In_84,In_619);
and U5237 (N_5237,In_2446,In_1640);
nand U5238 (N_5238,In_1988,In_914);
nor U5239 (N_5239,In_2193,In_2203);
nor U5240 (N_5240,In_1573,In_2368);
or U5241 (N_5241,In_2371,In_526);
and U5242 (N_5242,In_92,In_70);
and U5243 (N_5243,In_1081,In_132);
nand U5244 (N_5244,In_1509,In_670);
and U5245 (N_5245,In_1932,In_659);
and U5246 (N_5246,In_1371,In_2216);
nand U5247 (N_5247,In_2277,In_1276);
nand U5248 (N_5248,In_2321,In_1259);
or U5249 (N_5249,In_731,In_2115);
and U5250 (N_5250,In_1377,In_926);
nor U5251 (N_5251,In_680,In_1436);
nand U5252 (N_5252,In_444,In_1961);
or U5253 (N_5253,In_1649,In_1051);
and U5254 (N_5254,In_2045,In_161);
nand U5255 (N_5255,In_1261,In_545);
and U5256 (N_5256,In_610,In_1835);
xnor U5257 (N_5257,In_2134,In_619);
nand U5258 (N_5258,In_1838,In_337);
nor U5259 (N_5259,In_135,In_2255);
and U5260 (N_5260,In_1749,In_2271);
or U5261 (N_5261,In_419,In_1148);
and U5262 (N_5262,In_1561,In_558);
and U5263 (N_5263,In_2210,In_1935);
xor U5264 (N_5264,In_1291,In_1545);
and U5265 (N_5265,In_786,In_491);
nand U5266 (N_5266,In_96,In_2481);
nand U5267 (N_5267,In_2440,In_2398);
or U5268 (N_5268,In_2438,In_1668);
nand U5269 (N_5269,In_1465,In_1616);
and U5270 (N_5270,In_2239,In_1866);
or U5271 (N_5271,In_2351,In_547);
and U5272 (N_5272,In_339,In_1676);
nor U5273 (N_5273,In_1851,In_1924);
xor U5274 (N_5274,In_533,In_487);
nand U5275 (N_5275,In_2005,In_284);
xnor U5276 (N_5276,In_4,In_2192);
nand U5277 (N_5277,In_2106,In_1200);
nand U5278 (N_5278,In_706,In_644);
nand U5279 (N_5279,In_2176,In_34);
nor U5280 (N_5280,In_477,In_453);
nand U5281 (N_5281,In_627,In_204);
or U5282 (N_5282,In_1207,In_1692);
nor U5283 (N_5283,In_637,In_2357);
nand U5284 (N_5284,In_439,In_2294);
or U5285 (N_5285,In_77,In_1262);
and U5286 (N_5286,In_974,In_1827);
and U5287 (N_5287,In_1751,In_2390);
and U5288 (N_5288,In_1999,In_1672);
nand U5289 (N_5289,In_2286,In_1114);
nor U5290 (N_5290,In_522,In_1375);
and U5291 (N_5291,In_1648,In_426);
or U5292 (N_5292,In_1073,In_1351);
nor U5293 (N_5293,In_826,In_2042);
nand U5294 (N_5294,In_1061,In_1773);
nor U5295 (N_5295,In_1556,In_1046);
xor U5296 (N_5296,In_2293,In_2410);
or U5297 (N_5297,In_864,In_2263);
nand U5298 (N_5298,In_1597,In_1252);
nor U5299 (N_5299,In_1132,In_1423);
or U5300 (N_5300,In_1855,In_2486);
xor U5301 (N_5301,In_134,In_2032);
or U5302 (N_5302,In_1768,In_251);
nand U5303 (N_5303,In_1299,In_2289);
nor U5304 (N_5304,In_739,In_126);
and U5305 (N_5305,In_2081,In_2293);
nor U5306 (N_5306,In_1667,In_475);
or U5307 (N_5307,In_1646,In_1115);
xnor U5308 (N_5308,In_1967,In_1890);
and U5309 (N_5309,In_1659,In_217);
xor U5310 (N_5310,In_323,In_1037);
or U5311 (N_5311,In_645,In_1443);
nor U5312 (N_5312,In_913,In_1481);
and U5313 (N_5313,In_300,In_2093);
nor U5314 (N_5314,In_1624,In_2098);
nor U5315 (N_5315,In_1716,In_1545);
xor U5316 (N_5316,In_2094,In_2467);
nand U5317 (N_5317,In_644,In_641);
nor U5318 (N_5318,In_1320,In_715);
nor U5319 (N_5319,In_2000,In_550);
xnor U5320 (N_5320,In_1450,In_1242);
nor U5321 (N_5321,In_1722,In_661);
nand U5322 (N_5322,In_2043,In_1287);
and U5323 (N_5323,In_1839,In_931);
or U5324 (N_5324,In_39,In_2128);
nand U5325 (N_5325,In_2204,In_1727);
xor U5326 (N_5326,In_320,In_1465);
or U5327 (N_5327,In_93,In_2268);
nor U5328 (N_5328,In_726,In_724);
nor U5329 (N_5329,In_955,In_76);
nand U5330 (N_5330,In_291,In_1224);
and U5331 (N_5331,In_1383,In_2407);
or U5332 (N_5332,In_1458,In_2208);
nand U5333 (N_5333,In_2212,In_2241);
nor U5334 (N_5334,In_730,In_1696);
and U5335 (N_5335,In_466,In_1202);
nand U5336 (N_5336,In_1881,In_18);
nor U5337 (N_5337,In_1731,In_495);
nand U5338 (N_5338,In_232,In_1491);
or U5339 (N_5339,In_1163,In_2157);
nand U5340 (N_5340,In_500,In_498);
and U5341 (N_5341,In_926,In_2421);
nor U5342 (N_5342,In_1340,In_285);
xnor U5343 (N_5343,In_1687,In_1817);
and U5344 (N_5344,In_845,In_1170);
or U5345 (N_5345,In_88,In_195);
nor U5346 (N_5346,In_1399,In_2059);
nor U5347 (N_5347,In_1214,In_2474);
nor U5348 (N_5348,In_574,In_937);
or U5349 (N_5349,In_1889,In_1988);
xnor U5350 (N_5350,In_68,In_2442);
or U5351 (N_5351,In_1269,In_2057);
or U5352 (N_5352,In_1496,In_34);
and U5353 (N_5353,In_793,In_90);
xnor U5354 (N_5354,In_928,In_1709);
nor U5355 (N_5355,In_845,In_2451);
nor U5356 (N_5356,In_404,In_1977);
and U5357 (N_5357,In_983,In_1840);
or U5358 (N_5358,In_470,In_1678);
or U5359 (N_5359,In_1637,In_1795);
and U5360 (N_5360,In_384,In_2359);
xor U5361 (N_5361,In_1270,In_2421);
nand U5362 (N_5362,In_2069,In_1069);
or U5363 (N_5363,In_2322,In_2147);
or U5364 (N_5364,In_2139,In_1542);
or U5365 (N_5365,In_1310,In_797);
xnor U5366 (N_5366,In_1954,In_106);
nor U5367 (N_5367,In_1094,In_2226);
or U5368 (N_5368,In_1438,In_1335);
and U5369 (N_5369,In_1887,In_2224);
nor U5370 (N_5370,In_610,In_185);
and U5371 (N_5371,In_775,In_1905);
nand U5372 (N_5372,In_836,In_464);
nand U5373 (N_5373,In_1710,In_2182);
or U5374 (N_5374,In_595,In_1442);
xor U5375 (N_5375,In_1271,In_2160);
or U5376 (N_5376,In_543,In_609);
and U5377 (N_5377,In_1679,In_1889);
or U5378 (N_5378,In_2440,In_191);
nor U5379 (N_5379,In_261,In_2135);
or U5380 (N_5380,In_1880,In_1635);
nand U5381 (N_5381,In_399,In_1655);
nor U5382 (N_5382,In_1212,In_270);
nand U5383 (N_5383,In_1193,In_529);
xor U5384 (N_5384,In_211,In_818);
and U5385 (N_5385,In_704,In_2155);
or U5386 (N_5386,In_1010,In_349);
nand U5387 (N_5387,In_1333,In_2079);
nor U5388 (N_5388,In_106,In_324);
or U5389 (N_5389,In_1664,In_1657);
and U5390 (N_5390,In_733,In_514);
nand U5391 (N_5391,In_2373,In_2496);
nor U5392 (N_5392,In_821,In_1460);
or U5393 (N_5393,In_2067,In_1445);
xor U5394 (N_5394,In_464,In_576);
or U5395 (N_5395,In_732,In_1569);
nor U5396 (N_5396,In_617,In_1649);
nor U5397 (N_5397,In_77,In_2015);
or U5398 (N_5398,In_1707,In_1977);
xnor U5399 (N_5399,In_1985,In_236);
and U5400 (N_5400,In_292,In_191);
nand U5401 (N_5401,In_248,In_1469);
nand U5402 (N_5402,In_2198,In_1540);
nor U5403 (N_5403,In_2119,In_1210);
or U5404 (N_5404,In_1611,In_308);
and U5405 (N_5405,In_186,In_2142);
nor U5406 (N_5406,In_1125,In_910);
or U5407 (N_5407,In_2091,In_1403);
and U5408 (N_5408,In_95,In_1252);
nand U5409 (N_5409,In_2475,In_586);
nand U5410 (N_5410,In_328,In_1905);
nand U5411 (N_5411,In_800,In_493);
nor U5412 (N_5412,In_1,In_2069);
nand U5413 (N_5413,In_22,In_1757);
or U5414 (N_5414,In_1676,In_1574);
or U5415 (N_5415,In_1021,In_209);
nor U5416 (N_5416,In_1563,In_315);
or U5417 (N_5417,In_1522,In_937);
nor U5418 (N_5418,In_1164,In_390);
and U5419 (N_5419,In_1473,In_1568);
and U5420 (N_5420,In_689,In_2285);
nor U5421 (N_5421,In_379,In_394);
or U5422 (N_5422,In_1637,In_447);
nand U5423 (N_5423,In_2126,In_615);
or U5424 (N_5424,In_953,In_1620);
or U5425 (N_5425,In_114,In_1140);
and U5426 (N_5426,In_1734,In_2080);
or U5427 (N_5427,In_2226,In_1582);
nand U5428 (N_5428,In_469,In_781);
and U5429 (N_5429,In_2472,In_26);
xor U5430 (N_5430,In_2356,In_484);
and U5431 (N_5431,In_24,In_155);
nand U5432 (N_5432,In_1259,In_712);
and U5433 (N_5433,In_1804,In_1613);
nand U5434 (N_5434,In_507,In_200);
nor U5435 (N_5435,In_95,In_1593);
and U5436 (N_5436,In_726,In_18);
nand U5437 (N_5437,In_87,In_789);
or U5438 (N_5438,In_292,In_1815);
or U5439 (N_5439,In_1157,In_1837);
nand U5440 (N_5440,In_469,In_2031);
nor U5441 (N_5441,In_1227,In_888);
and U5442 (N_5442,In_331,In_294);
and U5443 (N_5443,In_2302,In_632);
or U5444 (N_5444,In_327,In_1357);
and U5445 (N_5445,In_172,In_1585);
and U5446 (N_5446,In_1602,In_173);
nor U5447 (N_5447,In_68,In_927);
and U5448 (N_5448,In_1765,In_1617);
nand U5449 (N_5449,In_17,In_1861);
or U5450 (N_5450,In_949,In_275);
and U5451 (N_5451,In_2404,In_686);
nand U5452 (N_5452,In_288,In_862);
and U5453 (N_5453,In_243,In_67);
or U5454 (N_5454,In_763,In_1896);
nor U5455 (N_5455,In_655,In_2202);
nor U5456 (N_5456,In_91,In_1787);
or U5457 (N_5457,In_1729,In_408);
or U5458 (N_5458,In_2113,In_1852);
xor U5459 (N_5459,In_1978,In_782);
nor U5460 (N_5460,In_631,In_1521);
nand U5461 (N_5461,In_825,In_139);
and U5462 (N_5462,In_24,In_2394);
or U5463 (N_5463,In_1560,In_963);
nor U5464 (N_5464,In_177,In_1859);
or U5465 (N_5465,In_1675,In_455);
and U5466 (N_5466,In_650,In_1389);
nand U5467 (N_5467,In_526,In_897);
nor U5468 (N_5468,In_2275,In_986);
or U5469 (N_5469,In_1568,In_882);
nand U5470 (N_5470,In_2103,In_78);
and U5471 (N_5471,In_2091,In_1644);
nor U5472 (N_5472,In_2485,In_2009);
or U5473 (N_5473,In_1231,In_197);
and U5474 (N_5474,In_1883,In_799);
nor U5475 (N_5475,In_2027,In_1087);
xor U5476 (N_5476,In_2355,In_177);
or U5477 (N_5477,In_285,In_690);
nand U5478 (N_5478,In_2456,In_1940);
and U5479 (N_5479,In_1563,In_1931);
xor U5480 (N_5480,In_1063,In_2310);
and U5481 (N_5481,In_1245,In_1808);
nand U5482 (N_5482,In_292,In_324);
and U5483 (N_5483,In_835,In_1905);
nand U5484 (N_5484,In_733,In_678);
and U5485 (N_5485,In_665,In_1117);
xnor U5486 (N_5486,In_2092,In_329);
or U5487 (N_5487,In_71,In_1553);
and U5488 (N_5488,In_1550,In_1790);
and U5489 (N_5489,In_2162,In_2449);
and U5490 (N_5490,In_2397,In_319);
or U5491 (N_5491,In_1478,In_139);
nand U5492 (N_5492,In_1925,In_1501);
nor U5493 (N_5493,In_1190,In_2068);
nor U5494 (N_5494,In_1582,In_1538);
or U5495 (N_5495,In_781,In_1584);
and U5496 (N_5496,In_1064,In_1383);
and U5497 (N_5497,In_525,In_947);
and U5498 (N_5498,In_2336,In_2144);
nand U5499 (N_5499,In_1340,In_881);
nand U5500 (N_5500,In_1837,In_1515);
nor U5501 (N_5501,In_723,In_654);
and U5502 (N_5502,In_1727,In_489);
nand U5503 (N_5503,In_1992,In_1868);
and U5504 (N_5504,In_9,In_10);
nand U5505 (N_5505,In_1372,In_1109);
nand U5506 (N_5506,In_1076,In_1009);
and U5507 (N_5507,In_381,In_1911);
or U5508 (N_5508,In_1122,In_519);
or U5509 (N_5509,In_869,In_2311);
nor U5510 (N_5510,In_408,In_1857);
nor U5511 (N_5511,In_902,In_730);
nor U5512 (N_5512,In_2160,In_783);
nand U5513 (N_5513,In_2097,In_208);
or U5514 (N_5514,In_2390,In_2107);
nor U5515 (N_5515,In_654,In_422);
nand U5516 (N_5516,In_448,In_420);
nor U5517 (N_5517,In_2118,In_1575);
or U5518 (N_5518,In_1173,In_2337);
nor U5519 (N_5519,In_2086,In_362);
nor U5520 (N_5520,In_1951,In_2079);
or U5521 (N_5521,In_2115,In_1499);
nand U5522 (N_5522,In_809,In_2383);
nor U5523 (N_5523,In_2030,In_1583);
or U5524 (N_5524,In_1481,In_1666);
and U5525 (N_5525,In_30,In_1929);
nor U5526 (N_5526,In_953,In_450);
nand U5527 (N_5527,In_2487,In_1217);
xnor U5528 (N_5528,In_2410,In_1728);
or U5529 (N_5529,In_1697,In_412);
xor U5530 (N_5530,In_1537,In_1503);
nand U5531 (N_5531,In_497,In_1110);
or U5532 (N_5532,In_2162,In_2144);
nor U5533 (N_5533,In_219,In_1034);
xor U5534 (N_5534,In_2071,In_806);
nand U5535 (N_5535,In_1007,In_993);
or U5536 (N_5536,In_1863,In_1887);
and U5537 (N_5537,In_701,In_971);
nand U5538 (N_5538,In_1535,In_1686);
or U5539 (N_5539,In_377,In_901);
nand U5540 (N_5540,In_1734,In_110);
nor U5541 (N_5541,In_164,In_336);
or U5542 (N_5542,In_2200,In_1572);
nor U5543 (N_5543,In_804,In_2099);
and U5544 (N_5544,In_2284,In_212);
nand U5545 (N_5545,In_319,In_35);
nor U5546 (N_5546,In_735,In_1627);
or U5547 (N_5547,In_1955,In_251);
and U5548 (N_5548,In_315,In_1973);
nor U5549 (N_5549,In_759,In_303);
nand U5550 (N_5550,In_947,In_1851);
or U5551 (N_5551,In_33,In_263);
nor U5552 (N_5552,In_1083,In_1328);
or U5553 (N_5553,In_651,In_339);
nand U5554 (N_5554,In_923,In_2110);
nand U5555 (N_5555,In_881,In_1711);
nand U5556 (N_5556,In_1378,In_27);
nand U5557 (N_5557,In_1876,In_1363);
or U5558 (N_5558,In_1939,In_1797);
nor U5559 (N_5559,In_2006,In_1297);
and U5560 (N_5560,In_2325,In_2191);
nand U5561 (N_5561,In_1073,In_1005);
and U5562 (N_5562,In_2302,In_1787);
and U5563 (N_5563,In_379,In_1328);
or U5564 (N_5564,In_1600,In_2309);
nand U5565 (N_5565,In_1725,In_1853);
xor U5566 (N_5566,In_1737,In_1715);
and U5567 (N_5567,In_1827,In_1804);
nor U5568 (N_5568,In_2286,In_1538);
xor U5569 (N_5569,In_2002,In_1513);
and U5570 (N_5570,In_2086,In_732);
or U5571 (N_5571,In_1293,In_126);
and U5572 (N_5572,In_482,In_1802);
xor U5573 (N_5573,In_2078,In_1348);
nand U5574 (N_5574,In_286,In_75);
nand U5575 (N_5575,In_120,In_3);
nand U5576 (N_5576,In_2112,In_1960);
or U5577 (N_5577,In_1289,In_1174);
xor U5578 (N_5578,In_612,In_1522);
nor U5579 (N_5579,In_1250,In_1082);
nand U5580 (N_5580,In_599,In_1344);
and U5581 (N_5581,In_384,In_1267);
and U5582 (N_5582,In_2459,In_1319);
nand U5583 (N_5583,In_81,In_92);
xnor U5584 (N_5584,In_1606,In_1630);
or U5585 (N_5585,In_2381,In_1448);
nand U5586 (N_5586,In_2203,In_1985);
nand U5587 (N_5587,In_1419,In_745);
and U5588 (N_5588,In_1863,In_736);
nand U5589 (N_5589,In_1875,In_1873);
nor U5590 (N_5590,In_1567,In_96);
nor U5591 (N_5591,In_567,In_2447);
or U5592 (N_5592,In_1160,In_1490);
nor U5593 (N_5593,In_1311,In_2183);
or U5594 (N_5594,In_838,In_556);
and U5595 (N_5595,In_644,In_1493);
and U5596 (N_5596,In_746,In_335);
or U5597 (N_5597,In_1576,In_1555);
and U5598 (N_5598,In_1207,In_1982);
nor U5599 (N_5599,In_1020,In_418);
nor U5600 (N_5600,In_2154,In_340);
nand U5601 (N_5601,In_2065,In_336);
or U5602 (N_5602,In_733,In_557);
xor U5603 (N_5603,In_1986,In_1305);
or U5604 (N_5604,In_1209,In_999);
and U5605 (N_5605,In_2145,In_2117);
nor U5606 (N_5606,In_964,In_1070);
nor U5607 (N_5607,In_222,In_2059);
nand U5608 (N_5608,In_1041,In_1848);
nor U5609 (N_5609,In_2106,In_25);
nor U5610 (N_5610,In_1116,In_2215);
nor U5611 (N_5611,In_67,In_694);
nor U5612 (N_5612,In_312,In_1970);
and U5613 (N_5613,In_1136,In_1781);
and U5614 (N_5614,In_1832,In_1638);
or U5615 (N_5615,In_219,In_260);
nand U5616 (N_5616,In_434,In_508);
or U5617 (N_5617,In_2031,In_1349);
and U5618 (N_5618,In_701,In_1841);
xor U5619 (N_5619,In_2256,In_1216);
nor U5620 (N_5620,In_2481,In_1986);
nand U5621 (N_5621,In_411,In_1821);
and U5622 (N_5622,In_2257,In_1591);
and U5623 (N_5623,In_922,In_424);
xnor U5624 (N_5624,In_414,In_2356);
nor U5625 (N_5625,In_2280,In_483);
nor U5626 (N_5626,In_1272,In_820);
and U5627 (N_5627,In_2404,In_253);
nand U5628 (N_5628,In_501,In_325);
nor U5629 (N_5629,In_1555,In_12);
nor U5630 (N_5630,In_224,In_1131);
or U5631 (N_5631,In_558,In_2077);
or U5632 (N_5632,In_1492,In_311);
or U5633 (N_5633,In_1709,In_1887);
nor U5634 (N_5634,In_912,In_1843);
nor U5635 (N_5635,In_229,In_448);
or U5636 (N_5636,In_2065,In_96);
or U5637 (N_5637,In_627,In_704);
or U5638 (N_5638,In_1736,In_2109);
nand U5639 (N_5639,In_1428,In_283);
nand U5640 (N_5640,In_2149,In_1710);
or U5641 (N_5641,In_635,In_605);
nand U5642 (N_5642,In_1009,In_2300);
nor U5643 (N_5643,In_1191,In_1488);
xor U5644 (N_5644,In_69,In_834);
nand U5645 (N_5645,In_1494,In_521);
and U5646 (N_5646,In_471,In_1053);
nor U5647 (N_5647,In_1458,In_2044);
nor U5648 (N_5648,In_2439,In_202);
nand U5649 (N_5649,In_679,In_1914);
or U5650 (N_5650,In_1314,In_2038);
and U5651 (N_5651,In_213,In_507);
nor U5652 (N_5652,In_1556,In_1142);
and U5653 (N_5653,In_301,In_1193);
nor U5654 (N_5654,In_1903,In_1907);
or U5655 (N_5655,In_150,In_812);
or U5656 (N_5656,In_1222,In_62);
or U5657 (N_5657,In_2165,In_258);
and U5658 (N_5658,In_1906,In_1940);
and U5659 (N_5659,In_930,In_62);
nand U5660 (N_5660,In_1552,In_844);
nand U5661 (N_5661,In_1533,In_535);
xnor U5662 (N_5662,In_852,In_1028);
and U5663 (N_5663,In_1508,In_2219);
nand U5664 (N_5664,In_518,In_2014);
and U5665 (N_5665,In_1826,In_791);
xnor U5666 (N_5666,In_1684,In_1874);
nand U5667 (N_5667,In_2226,In_1026);
and U5668 (N_5668,In_1847,In_1529);
xnor U5669 (N_5669,In_758,In_472);
nor U5670 (N_5670,In_2197,In_725);
and U5671 (N_5671,In_2207,In_323);
or U5672 (N_5672,In_1500,In_1951);
nand U5673 (N_5673,In_1327,In_2196);
and U5674 (N_5674,In_2266,In_1987);
and U5675 (N_5675,In_1738,In_1455);
or U5676 (N_5676,In_1662,In_1640);
and U5677 (N_5677,In_2406,In_1675);
and U5678 (N_5678,In_156,In_217);
or U5679 (N_5679,In_198,In_2445);
xor U5680 (N_5680,In_628,In_113);
nor U5681 (N_5681,In_402,In_2307);
nand U5682 (N_5682,In_561,In_818);
nor U5683 (N_5683,In_2017,In_672);
nand U5684 (N_5684,In_675,In_1965);
and U5685 (N_5685,In_2487,In_1668);
nand U5686 (N_5686,In_567,In_1708);
nand U5687 (N_5687,In_876,In_798);
nor U5688 (N_5688,In_2131,In_1274);
or U5689 (N_5689,In_31,In_2123);
nor U5690 (N_5690,In_498,In_2079);
and U5691 (N_5691,In_653,In_1996);
nor U5692 (N_5692,In_2115,In_2279);
and U5693 (N_5693,In_2029,In_1494);
or U5694 (N_5694,In_2116,In_1905);
and U5695 (N_5695,In_1758,In_2380);
and U5696 (N_5696,In_1778,In_898);
nor U5697 (N_5697,In_1009,In_196);
or U5698 (N_5698,In_18,In_1155);
or U5699 (N_5699,In_314,In_622);
and U5700 (N_5700,In_2152,In_742);
nor U5701 (N_5701,In_1885,In_264);
and U5702 (N_5702,In_1052,In_2173);
nand U5703 (N_5703,In_1583,In_2341);
or U5704 (N_5704,In_1652,In_174);
nor U5705 (N_5705,In_367,In_1689);
nor U5706 (N_5706,In_1575,In_1851);
nand U5707 (N_5707,In_304,In_467);
or U5708 (N_5708,In_1404,In_1923);
nand U5709 (N_5709,In_1082,In_2172);
nand U5710 (N_5710,In_697,In_1761);
nor U5711 (N_5711,In_1684,In_874);
and U5712 (N_5712,In_577,In_335);
nor U5713 (N_5713,In_519,In_787);
nand U5714 (N_5714,In_1144,In_982);
or U5715 (N_5715,In_1202,In_1497);
and U5716 (N_5716,In_440,In_1470);
xnor U5717 (N_5717,In_2334,In_2499);
nand U5718 (N_5718,In_563,In_1685);
xor U5719 (N_5719,In_1534,In_720);
xnor U5720 (N_5720,In_418,In_366);
xnor U5721 (N_5721,In_683,In_114);
nor U5722 (N_5722,In_907,In_1748);
nor U5723 (N_5723,In_1201,In_1238);
nor U5724 (N_5724,In_402,In_2096);
and U5725 (N_5725,In_1550,In_1465);
nand U5726 (N_5726,In_419,In_361);
nor U5727 (N_5727,In_760,In_301);
nand U5728 (N_5728,In_2035,In_22);
or U5729 (N_5729,In_2328,In_2469);
and U5730 (N_5730,In_336,In_354);
nor U5731 (N_5731,In_962,In_1232);
and U5732 (N_5732,In_641,In_1637);
and U5733 (N_5733,In_1060,In_171);
nand U5734 (N_5734,In_1227,In_2447);
and U5735 (N_5735,In_1417,In_2258);
or U5736 (N_5736,In_1139,In_123);
xor U5737 (N_5737,In_863,In_1991);
nand U5738 (N_5738,In_815,In_1980);
or U5739 (N_5739,In_950,In_1840);
or U5740 (N_5740,In_604,In_1072);
nand U5741 (N_5741,In_824,In_2365);
or U5742 (N_5742,In_1844,In_859);
nor U5743 (N_5743,In_1002,In_2016);
or U5744 (N_5744,In_1613,In_1797);
nor U5745 (N_5745,In_980,In_1637);
nor U5746 (N_5746,In_911,In_1813);
and U5747 (N_5747,In_1867,In_1002);
xnor U5748 (N_5748,In_1696,In_2378);
and U5749 (N_5749,In_44,In_404);
and U5750 (N_5750,In_1493,In_1737);
and U5751 (N_5751,In_2258,In_1342);
nor U5752 (N_5752,In_1056,In_1877);
nand U5753 (N_5753,In_1124,In_1871);
xnor U5754 (N_5754,In_896,In_1762);
and U5755 (N_5755,In_1890,In_773);
and U5756 (N_5756,In_1201,In_1536);
nor U5757 (N_5757,In_1548,In_270);
or U5758 (N_5758,In_2385,In_813);
nand U5759 (N_5759,In_2469,In_2033);
or U5760 (N_5760,In_1521,In_2000);
nand U5761 (N_5761,In_14,In_2391);
or U5762 (N_5762,In_2428,In_1794);
and U5763 (N_5763,In_785,In_445);
xnor U5764 (N_5764,In_2242,In_687);
nand U5765 (N_5765,In_826,In_1538);
and U5766 (N_5766,In_569,In_1945);
nand U5767 (N_5767,In_1649,In_1662);
nor U5768 (N_5768,In_560,In_1904);
and U5769 (N_5769,In_1001,In_1551);
or U5770 (N_5770,In_1129,In_685);
or U5771 (N_5771,In_2475,In_60);
and U5772 (N_5772,In_834,In_1500);
nor U5773 (N_5773,In_2470,In_1165);
nand U5774 (N_5774,In_1777,In_431);
or U5775 (N_5775,In_354,In_2248);
nor U5776 (N_5776,In_1279,In_2231);
or U5777 (N_5777,In_521,In_2111);
and U5778 (N_5778,In_1456,In_1086);
xor U5779 (N_5779,In_1095,In_638);
or U5780 (N_5780,In_1946,In_556);
xor U5781 (N_5781,In_1106,In_2439);
and U5782 (N_5782,In_2399,In_1950);
xor U5783 (N_5783,In_91,In_1769);
or U5784 (N_5784,In_177,In_1669);
nand U5785 (N_5785,In_2388,In_1219);
nand U5786 (N_5786,In_1944,In_976);
nand U5787 (N_5787,In_1267,In_1331);
nand U5788 (N_5788,In_1447,In_2116);
nand U5789 (N_5789,In_1753,In_1885);
xnor U5790 (N_5790,In_1457,In_883);
nand U5791 (N_5791,In_1731,In_1200);
or U5792 (N_5792,In_1454,In_2040);
and U5793 (N_5793,In_711,In_1976);
xnor U5794 (N_5794,In_42,In_1071);
nand U5795 (N_5795,In_1025,In_1251);
nand U5796 (N_5796,In_14,In_1335);
nand U5797 (N_5797,In_1376,In_2285);
nand U5798 (N_5798,In_917,In_1059);
or U5799 (N_5799,In_894,In_1460);
or U5800 (N_5800,In_2119,In_1228);
and U5801 (N_5801,In_1118,In_1453);
nand U5802 (N_5802,In_2410,In_1854);
xor U5803 (N_5803,In_1916,In_91);
and U5804 (N_5804,In_398,In_2195);
and U5805 (N_5805,In_1732,In_1030);
xor U5806 (N_5806,In_956,In_427);
xor U5807 (N_5807,In_2147,In_1622);
nor U5808 (N_5808,In_631,In_972);
nand U5809 (N_5809,In_1945,In_865);
and U5810 (N_5810,In_784,In_705);
or U5811 (N_5811,In_165,In_793);
and U5812 (N_5812,In_1924,In_2421);
nor U5813 (N_5813,In_797,In_1378);
xor U5814 (N_5814,In_1919,In_1881);
or U5815 (N_5815,In_2268,In_498);
and U5816 (N_5816,In_888,In_176);
nor U5817 (N_5817,In_2186,In_22);
nand U5818 (N_5818,In_1341,In_1739);
nand U5819 (N_5819,In_682,In_2398);
or U5820 (N_5820,In_2405,In_1258);
nand U5821 (N_5821,In_2268,In_2147);
nand U5822 (N_5822,In_590,In_2446);
or U5823 (N_5823,In_2433,In_2263);
nor U5824 (N_5824,In_1629,In_1245);
or U5825 (N_5825,In_1395,In_937);
nand U5826 (N_5826,In_664,In_1140);
and U5827 (N_5827,In_1226,In_306);
nand U5828 (N_5828,In_1140,In_2441);
nor U5829 (N_5829,In_1815,In_1515);
nand U5830 (N_5830,In_1485,In_1107);
nor U5831 (N_5831,In_1343,In_2317);
or U5832 (N_5832,In_932,In_1718);
nor U5833 (N_5833,In_952,In_874);
and U5834 (N_5834,In_1660,In_2166);
xnor U5835 (N_5835,In_1047,In_2369);
xor U5836 (N_5836,In_1466,In_2458);
nand U5837 (N_5837,In_2091,In_1512);
or U5838 (N_5838,In_2449,In_2218);
and U5839 (N_5839,In_1850,In_407);
nand U5840 (N_5840,In_37,In_1736);
nand U5841 (N_5841,In_2109,In_1439);
nand U5842 (N_5842,In_2113,In_719);
nand U5843 (N_5843,In_407,In_1300);
nand U5844 (N_5844,In_844,In_698);
nor U5845 (N_5845,In_882,In_1916);
or U5846 (N_5846,In_2417,In_531);
and U5847 (N_5847,In_2306,In_2045);
nor U5848 (N_5848,In_1537,In_762);
and U5849 (N_5849,In_219,In_893);
xor U5850 (N_5850,In_2337,In_640);
nand U5851 (N_5851,In_52,In_2089);
xnor U5852 (N_5852,In_1636,In_2114);
nor U5853 (N_5853,In_2039,In_1075);
nor U5854 (N_5854,In_2296,In_128);
nor U5855 (N_5855,In_1155,In_974);
xnor U5856 (N_5856,In_1175,In_1210);
and U5857 (N_5857,In_225,In_779);
or U5858 (N_5858,In_2097,In_1344);
or U5859 (N_5859,In_2036,In_1887);
xnor U5860 (N_5860,In_2347,In_5);
or U5861 (N_5861,In_2291,In_1730);
and U5862 (N_5862,In_973,In_620);
xnor U5863 (N_5863,In_178,In_1418);
or U5864 (N_5864,In_1478,In_1950);
nand U5865 (N_5865,In_2156,In_1625);
and U5866 (N_5866,In_819,In_1549);
nand U5867 (N_5867,In_1299,In_2222);
or U5868 (N_5868,In_415,In_1816);
nor U5869 (N_5869,In_1405,In_34);
xor U5870 (N_5870,In_509,In_2439);
nor U5871 (N_5871,In_922,In_1763);
xor U5872 (N_5872,In_3,In_2308);
nor U5873 (N_5873,In_1811,In_78);
or U5874 (N_5874,In_2498,In_524);
nor U5875 (N_5875,In_1339,In_2385);
or U5876 (N_5876,In_1867,In_582);
nor U5877 (N_5877,In_2263,In_2365);
nand U5878 (N_5878,In_1656,In_55);
nand U5879 (N_5879,In_1542,In_1554);
or U5880 (N_5880,In_1622,In_1300);
nand U5881 (N_5881,In_369,In_2477);
or U5882 (N_5882,In_1181,In_854);
nand U5883 (N_5883,In_2205,In_1034);
xnor U5884 (N_5884,In_310,In_2041);
and U5885 (N_5885,In_770,In_943);
nand U5886 (N_5886,In_75,In_986);
or U5887 (N_5887,In_891,In_378);
nand U5888 (N_5888,In_261,In_2327);
nor U5889 (N_5889,In_267,In_2394);
nand U5890 (N_5890,In_1412,In_283);
and U5891 (N_5891,In_645,In_291);
nor U5892 (N_5892,In_116,In_1072);
and U5893 (N_5893,In_381,In_1741);
nand U5894 (N_5894,In_1906,In_940);
or U5895 (N_5895,In_2294,In_281);
or U5896 (N_5896,In_1151,In_1515);
or U5897 (N_5897,In_1729,In_486);
or U5898 (N_5898,In_1120,In_820);
xnor U5899 (N_5899,In_2350,In_813);
and U5900 (N_5900,In_2468,In_1940);
nor U5901 (N_5901,In_1030,In_1007);
nor U5902 (N_5902,In_1542,In_205);
and U5903 (N_5903,In_832,In_1679);
nor U5904 (N_5904,In_1281,In_1712);
nor U5905 (N_5905,In_276,In_1853);
and U5906 (N_5906,In_223,In_80);
nand U5907 (N_5907,In_1078,In_2207);
or U5908 (N_5908,In_984,In_988);
nor U5909 (N_5909,In_1959,In_1546);
and U5910 (N_5910,In_1793,In_1996);
xnor U5911 (N_5911,In_760,In_1723);
or U5912 (N_5912,In_1791,In_1513);
nand U5913 (N_5913,In_449,In_1500);
or U5914 (N_5914,In_2327,In_2207);
xnor U5915 (N_5915,In_2477,In_2499);
nand U5916 (N_5916,In_398,In_1626);
nor U5917 (N_5917,In_1554,In_1883);
or U5918 (N_5918,In_570,In_1278);
and U5919 (N_5919,In_2066,In_1327);
and U5920 (N_5920,In_209,In_168);
nand U5921 (N_5921,In_1641,In_1663);
nand U5922 (N_5922,In_1127,In_1932);
nand U5923 (N_5923,In_457,In_2100);
xnor U5924 (N_5924,In_1881,In_2368);
or U5925 (N_5925,In_350,In_1100);
or U5926 (N_5926,In_1734,In_2181);
or U5927 (N_5927,In_184,In_2223);
xor U5928 (N_5928,In_1838,In_2273);
nand U5929 (N_5929,In_1919,In_177);
and U5930 (N_5930,In_1706,In_469);
and U5931 (N_5931,In_2079,In_1446);
nand U5932 (N_5932,In_2124,In_1059);
nand U5933 (N_5933,In_53,In_1719);
and U5934 (N_5934,In_1738,In_1751);
nand U5935 (N_5935,In_780,In_1205);
nor U5936 (N_5936,In_2046,In_1536);
and U5937 (N_5937,In_2137,In_1253);
or U5938 (N_5938,In_2292,In_310);
or U5939 (N_5939,In_1935,In_1698);
or U5940 (N_5940,In_1977,In_1257);
or U5941 (N_5941,In_655,In_253);
nand U5942 (N_5942,In_2406,In_711);
or U5943 (N_5943,In_2208,In_2084);
and U5944 (N_5944,In_994,In_742);
nand U5945 (N_5945,In_865,In_2162);
or U5946 (N_5946,In_747,In_186);
nand U5947 (N_5947,In_834,In_1850);
or U5948 (N_5948,In_679,In_941);
and U5949 (N_5949,In_660,In_550);
xor U5950 (N_5950,In_711,In_2245);
nor U5951 (N_5951,In_1029,In_2339);
and U5952 (N_5952,In_2319,In_188);
nor U5953 (N_5953,In_2491,In_535);
xor U5954 (N_5954,In_1660,In_2435);
nor U5955 (N_5955,In_2433,In_2092);
or U5956 (N_5956,In_55,In_1187);
or U5957 (N_5957,In_2162,In_1321);
nand U5958 (N_5958,In_801,In_1942);
nor U5959 (N_5959,In_493,In_2454);
nand U5960 (N_5960,In_1686,In_2235);
nand U5961 (N_5961,In_1657,In_774);
xor U5962 (N_5962,In_1673,In_1495);
and U5963 (N_5963,In_1929,In_2019);
nor U5964 (N_5964,In_851,In_1773);
nor U5965 (N_5965,In_76,In_841);
or U5966 (N_5966,In_763,In_2233);
xnor U5967 (N_5967,In_2369,In_2311);
xnor U5968 (N_5968,In_1271,In_1990);
nand U5969 (N_5969,In_297,In_352);
and U5970 (N_5970,In_1580,In_2369);
nand U5971 (N_5971,In_180,In_749);
xnor U5972 (N_5972,In_1509,In_1585);
nand U5973 (N_5973,In_100,In_46);
and U5974 (N_5974,In_547,In_565);
nor U5975 (N_5975,In_1426,In_1455);
xor U5976 (N_5976,In_35,In_25);
nor U5977 (N_5977,In_2269,In_384);
and U5978 (N_5978,In_688,In_698);
and U5979 (N_5979,In_1903,In_1797);
nor U5980 (N_5980,In_2365,In_1490);
nor U5981 (N_5981,In_249,In_479);
or U5982 (N_5982,In_51,In_1705);
nand U5983 (N_5983,In_1985,In_2424);
nand U5984 (N_5984,In_1524,In_636);
or U5985 (N_5985,In_945,In_1334);
nand U5986 (N_5986,In_1138,In_1756);
or U5987 (N_5987,In_1024,In_1939);
or U5988 (N_5988,In_1959,In_1106);
and U5989 (N_5989,In_979,In_982);
nor U5990 (N_5990,In_1174,In_109);
and U5991 (N_5991,In_1204,In_138);
nand U5992 (N_5992,In_1209,In_2004);
nand U5993 (N_5993,In_1501,In_792);
or U5994 (N_5994,In_1136,In_949);
nor U5995 (N_5995,In_1837,In_461);
and U5996 (N_5996,In_1948,In_1938);
and U5997 (N_5997,In_327,In_1386);
nor U5998 (N_5998,In_1081,In_2430);
and U5999 (N_5999,In_1977,In_1655);
or U6000 (N_6000,In_1825,In_1387);
nand U6001 (N_6001,In_1696,In_505);
nor U6002 (N_6002,In_992,In_1393);
or U6003 (N_6003,In_1442,In_181);
and U6004 (N_6004,In_250,In_2311);
nor U6005 (N_6005,In_148,In_106);
nor U6006 (N_6006,In_934,In_1289);
or U6007 (N_6007,In_982,In_1173);
and U6008 (N_6008,In_1064,In_2044);
nor U6009 (N_6009,In_1725,In_1923);
nand U6010 (N_6010,In_1880,In_1446);
or U6011 (N_6011,In_160,In_1294);
nor U6012 (N_6012,In_539,In_23);
or U6013 (N_6013,In_999,In_1176);
and U6014 (N_6014,In_2215,In_298);
xor U6015 (N_6015,In_279,In_2474);
or U6016 (N_6016,In_1109,In_1151);
nand U6017 (N_6017,In_2109,In_2306);
nand U6018 (N_6018,In_1110,In_2467);
nor U6019 (N_6019,In_940,In_1990);
or U6020 (N_6020,In_2090,In_1028);
nand U6021 (N_6021,In_1469,In_1075);
or U6022 (N_6022,In_397,In_1435);
and U6023 (N_6023,In_1814,In_800);
nor U6024 (N_6024,In_2321,In_1511);
or U6025 (N_6025,In_1956,In_502);
nand U6026 (N_6026,In_47,In_555);
or U6027 (N_6027,In_1744,In_275);
and U6028 (N_6028,In_1753,In_1839);
and U6029 (N_6029,In_2008,In_2443);
or U6030 (N_6030,In_1270,In_1227);
and U6031 (N_6031,In_2104,In_1659);
xnor U6032 (N_6032,In_1769,In_1875);
or U6033 (N_6033,In_610,In_92);
and U6034 (N_6034,In_395,In_1342);
nor U6035 (N_6035,In_506,In_476);
and U6036 (N_6036,In_339,In_33);
and U6037 (N_6037,In_594,In_608);
nor U6038 (N_6038,In_774,In_92);
or U6039 (N_6039,In_1163,In_1244);
or U6040 (N_6040,In_138,In_2124);
and U6041 (N_6041,In_1749,In_1833);
or U6042 (N_6042,In_2007,In_2132);
nand U6043 (N_6043,In_350,In_1614);
nor U6044 (N_6044,In_1672,In_1373);
nor U6045 (N_6045,In_624,In_2056);
and U6046 (N_6046,In_298,In_2113);
xnor U6047 (N_6047,In_2075,In_487);
and U6048 (N_6048,In_1322,In_216);
and U6049 (N_6049,In_386,In_1450);
nor U6050 (N_6050,In_445,In_1160);
and U6051 (N_6051,In_99,In_1508);
nor U6052 (N_6052,In_219,In_1869);
nor U6053 (N_6053,In_996,In_489);
nand U6054 (N_6054,In_594,In_101);
or U6055 (N_6055,In_1263,In_447);
or U6056 (N_6056,In_493,In_2429);
and U6057 (N_6057,In_198,In_1301);
or U6058 (N_6058,In_109,In_1748);
or U6059 (N_6059,In_520,In_2352);
nor U6060 (N_6060,In_2344,In_1872);
or U6061 (N_6061,In_835,In_256);
nor U6062 (N_6062,In_1797,In_466);
nand U6063 (N_6063,In_212,In_416);
nand U6064 (N_6064,In_2274,In_2443);
or U6065 (N_6065,In_2384,In_1276);
nor U6066 (N_6066,In_1850,In_551);
xnor U6067 (N_6067,In_1604,In_1818);
xnor U6068 (N_6068,In_1366,In_2161);
nand U6069 (N_6069,In_1805,In_584);
or U6070 (N_6070,In_1624,In_2286);
nor U6071 (N_6071,In_2443,In_155);
nor U6072 (N_6072,In_653,In_146);
and U6073 (N_6073,In_1930,In_1375);
nor U6074 (N_6074,In_2315,In_296);
and U6075 (N_6075,In_1582,In_674);
or U6076 (N_6076,In_697,In_1116);
and U6077 (N_6077,In_750,In_1843);
nor U6078 (N_6078,In_252,In_903);
xor U6079 (N_6079,In_548,In_1070);
xnor U6080 (N_6080,In_1254,In_2259);
nand U6081 (N_6081,In_2010,In_1376);
xnor U6082 (N_6082,In_2101,In_1501);
and U6083 (N_6083,In_1119,In_1966);
or U6084 (N_6084,In_2175,In_304);
nor U6085 (N_6085,In_981,In_665);
and U6086 (N_6086,In_1806,In_6);
or U6087 (N_6087,In_2402,In_271);
nor U6088 (N_6088,In_1162,In_2461);
or U6089 (N_6089,In_1355,In_1614);
nand U6090 (N_6090,In_1782,In_2309);
nand U6091 (N_6091,In_2394,In_2376);
nand U6092 (N_6092,In_718,In_359);
nor U6093 (N_6093,In_494,In_1797);
nor U6094 (N_6094,In_283,In_1664);
nor U6095 (N_6095,In_215,In_1504);
or U6096 (N_6096,In_1506,In_875);
or U6097 (N_6097,In_1213,In_885);
nor U6098 (N_6098,In_1949,In_2001);
or U6099 (N_6099,In_1476,In_51);
and U6100 (N_6100,In_1819,In_2299);
and U6101 (N_6101,In_578,In_2348);
and U6102 (N_6102,In_915,In_291);
nand U6103 (N_6103,In_2215,In_249);
nor U6104 (N_6104,In_1598,In_2200);
or U6105 (N_6105,In_1699,In_591);
nand U6106 (N_6106,In_625,In_2332);
and U6107 (N_6107,In_2107,In_2099);
nor U6108 (N_6108,In_1201,In_2056);
and U6109 (N_6109,In_1694,In_1219);
nor U6110 (N_6110,In_2242,In_1160);
and U6111 (N_6111,In_2305,In_1482);
or U6112 (N_6112,In_927,In_228);
nor U6113 (N_6113,In_356,In_1085);
xor U6114 (N_6114,In_1692,In_1701);
or U6115 (N_6115,In_619,In_658);
nor U6116 (N_6116,In_2071,In_659);
nand U6117 (N_6117,In_1583,In_2068);
or U6118 (N_6118,In_1951,In_569);
nor U6119 (N_6119,In_2166,In_1789);
or U6120 (N_6120,In_1395,In_840);
nor U6121 (N_6121,In_1890,In_1952);
xnor U6122 (N_6122,In_2444,In_899);
nor U6123 (N_6123,In_263,In_765);
nand U6124 (N_6124,In_1416,In_2143);
nor U6125 (N_6125,In_900,In_2355);
xor U6126 (N_6126,In_579,In_1112);
and U6127 (N_6127,In_2181,In_1967);
or U6128 (N_6128,In_1858,In_759);
and U6129 (N_6129,In_812,In_2363);
or U6130 (N_6130,In_77,In_881);
nand U6131 (N_6131,In_1123,In_1431);
nand U6132 (N_6132,In_2471,In_67);
nor U6133 (N_6133,In_1606,In_1177);
nand U6134 (N_6134,In_898,In_2062);
nand U6135 (N_6135,In_707,In_2306);
xor U6136 (N_6136,In_2003,In_1919);
and U6137 (N_6137,In_1689,In_517);
and U6138 (N_6138,In_2322,In_513);
nand U6139 (N_6139,In_2128,In_1234);
or U6140 (N_6140,In_1312,In_167);
or U6141 (N_6141,In_804,In_1929);
or U6142 (N_6142,In_1333,In_2237);
or U6143 (N_6143,In_1246,In_1787);
nor U6144 (N_6144,In_1716,In_920);
nand U6145 (N_6145,In_11,In_208);
nor U6146 (N_6146,In_805,In_2025);
nand U6147 (N_6147,In_528,In_2285);
and U6148 (N_6148,In_1085,In_1283);
or U6149 (N_6149,In_158,In_805);
nand U6150 (N_6150,In_785,In_2309);
and U6151 (N_6151,In_1896,In_356);
nand U6152 (N_6152,In_576,In_513);
nor U6153 (N_6153,In_2022,In_380);
and U6154 (N_6154,In_2321,In_1676);
nand U6155 (N_6155,In_1324,In_1727);
xor U6156 (N_6156,In_1426,In_1796);
xor U6157 (N_6157,In_1707,In_374);
nand U6158 (N_6158,In_52,In_1726);
or U6159 (N_6159,In_570,In_524);
or U6160 (N_6160,In_690,In_2123);
or U6161 (N_6161,In_2003,In_2151);
nor U6162 (N_6162,In_2231,In_486);
nand U6163 (N_6163,In_751,In_2262);
nand U6164 (N_6164,In_979,In_680);
xnor U6165 (N_6165,In_822,In_136);
or U6166 (N_6166,In_1077,In_204);
or U6167 (N_6167,In_1466,In_426);
xor U6168 (N_6168,In_774,In_1102);
or U6169 (N_6169,In_800,In_738);
nand U6170 (N_6170,In_1634,In_761);
and U6171 (N_6171,In_1664,In_394);
or U6172 (N_6172,In_2394,In_1840);
xor U6173 (N_6173,In_1924,In_2148);
xnor U6174 (N_6174,In_1452,In_567);
nand U6175 (N_6175,In_931,In_1465);
nand U6176 (N_6176,In_186,In_1334);
nor U6177 (N_6177,In_2031,In_1377);
nand U6178 (N_6178,In_420,In_680);
nor U6179 (N_6179,In_1665,In_533);
or U6180 (N_6180,In_1700,In_729);
or U6181 (N_6181,In_2341,In_1682);
and U6182 (N_6182,In_2095,In_41);
or U6183 (N_6183,In_890,In_525);
or U6184 (N_6184,In_2217,In_2);
nand U6185 (N_6185,In_507,In_941);
or U6186 (N_6186,In_1433,In_204);
nor U6187 (N_6187,In_1526,In_44);
xor U6188 (N_6188,In_2206,In_888);
nand U6189 (N_6189,In_913,In_948);
or U6190 (N_6190,In_880,In_396);
and U6191 (N_6191,In_1719,In_1345);
nand U6192 (N_6192,In_182,In_570);
or U6193 (N_6193,In_1562,In_2063);
xnor U6194 (N_6194,In_370,In_1230);
or U6195 (N_6195,In_369,In_1568);
and U6196 (N_6196,In_2164,In_1837);
xnor U6197 (N_6197,In_1576,In_1091);
and U6198 (N_6198,In_1203,In_2228);
and U6199 (N_6199,In_444,In_2415);
xnor U6200 (N_6200,In_1673,In_1712);
and U6201 (N_6201,In_2242,In_666);
nand U6202 (N_6202,In_1684,In_575);
nor U6203 (N_6203,In_973,In_1246);
xor U6204 (N_6204,In_509,In_1925);
or U6205 (N_6205,In_2145,In_1462);
and U6206 (N_6206,In_644,In_1448);
nand U6207 (N_6207,In_2300,In_1718);
or U6208 (N_6208,In_1516,In_279);
or U6209 (N_6209,In_420,In_443);
and U6210 (N_6210,In_1583,In_2184);
and U6211 (N_6211,In_801,In_2147);
nand U6212 (N_6212,In_1830,In_1501);
nand U6213 (N_6213,In_108,In_1641);
or U6214 (N_6214,In_1870,In_1540);
nand U6215 (N_6215,In_2095,In_1661);
and U6216 (N_6216,In_2331,In_2363);
nor U6217 (N_6217,In_509,In_523);
nor U6218 (N_6218,In_150,In_742);
and U6219 (N_6219,In_250,In_2322);
or U6220 (N_6220,In_2213,In_2325);
or U6221 (N_6221,In_114,In_1634);
nor U6222 (N_6222,In_438,In_1711);
and U6223 (N_6223,In_2472,In_504);
nand U6224 (N_6224,In_1807,In_1115);
and U6225 (N_6225,In_2129,In_1580);
or U6226 (N_6226,In_1328,In_1050);
nand U6227 (N_6227,In_1034,In_605);
nor U6228 (N_6228,In_1140,In_925);
nand U6229 (N_6229,In_2283,In_19);
nor U6230 (N_6230,In_1279,In_316);
and U6231 (N_6231,In_1978,In_179);
or U6232 (N_6232,In_522,In_1585);
or U6233 (N_6233,In_925,In_1783);
or U6234 (N_6234,In_715,In_958);
or U6235 (N_6235,In_1672,In_509);
and U6236 (N_6236,In_2469,In_409);
nor U6237 (N_6237,In_381,In_1335);
nand U6238 (N_6238,In_97,In_1629);
and U6239 (N_6239,In_1382,In_634);
nand U6240 (N_6240,In_913,In_1239);
or U6241 (N_6241,In_1580,In_1419);
nand U6242 (N_6242,In_1599,In_1909);
nor U6243 (N_6243,In_355,In_61);
and U6244 (N_6244,In_357,In_1903);
nor U6245 (N_6245,In_2306,In_865);
nand U6246 (N_6246,In_2057,In_2240);
nand U6247 (N_6247,In_2462,In_1868);
and U6248 (N_6248,In_1610,In_908);
nand U6249 (N_6249,In_1238,In_485);
nor U6250 (N_6250,N_4397,N_660);
or U6251 (N_6251,N_4794,N_4432);
or U6252 (N_6252,N_2179,N_5470);
nor U6253 (N_6253,N_3051,N_3745);
nand U6254 (N_6254,N_12,N_2169);
xor U6255 (N_6255,N_1374,N_4467);
nor U6256 (N_6256,N_5877,N_5241);
nor U6257 (N_6257,N_5252,N_2384);
nand U6258 (N_6258,N_1084,N_6017);
and U6259 (N_6259,N_5993,N_2688);
xnor U6260 (N_6260,N_2087,N_767);
or U6261 (N_6261,N_353,N_1465);
nor U6262 (N_6262,N_1083,N_192);
or U6263 (N_6263,N_987,N_6031);
and U6264 (N_6264,N_2332,N_5208);
nor U6265 (N_6265,N_5537,N_59);
and U6266 (N_6266,N_5750,N_2427);
or U6267 (N_6267,N_4192,N_1421);
nand U6268 (N_6268,N_2155,N_3289);
and U6269 (N_6269,N_2206,N_982);
or U6270 (N_6270,N_5076,N_340);
nor U6271 (N_6271,N_6000,N_2767);
xnor U6272 (N_6272,N_3275,N_5826);
or U6273 (N_6273,N_1672,N_4279);
nor U6274 (N_6274,N_2006,N_222);
and U6275 (N_6275,N_3415,N_28);
or U6276 (N_6276,N_3291,N_1329);
and U6277 (N_6277,N_1483,N_1489);
or U6278 (N_6278,N_27,N_1363);
nand U6279 (N_6279,N_4350,N_1664);
nand U6280 (N_6280,N_675,N_422);
nand U6281 (N_6281,N_4946,N_5060);
nor U6282 (N_6282,N_5142,N_3206);
or U6283 (N_6283,N_3121,N_1395);
nor U6284 (N_6284,N_4578,N_5866);
and U6285 (N_6285,N_5668,N_6235);
or U6286 (N_6286,N_1979,N_609);
nand U6287 (N_6287,N_5068,N_4155);
and U6288 (N_6288,N_4511,N_5871);
and U6289 (N_6289,N_4713,N_605);
nor U6290 (N_6290,N_2758,N_1713);
nand U6291 (N_6291,N_5564,N_3537);
and U6292 (N_6292,N_2947,N_4071);
nor U6293 (N_6293,N_4124,N_3615);
or U6294 (N_6294,N_3429,N_2553);
nor U6295 (N_6295,N_4743,N_3073);
nand U6296 (N_6296,N_5897,N_5628);
and U6297 (N_6297,N_3678,N_846);
nor U6298 (N_6298,N_131,N_4342);
nor U6299 (N_6299,N_410,N_397);
nand U6300 (N_6300,N_5495,N_3979);
nand U6301 (N_6301,N_5723,N_5304);
or U6302 (N_6302,N_302,N_3440);
nor U6303 (N_6303,N_4662,N_4327);
nor U6304 (N_6304,N_2345,N_2451);
and U6305 (N_6305,N_3027,N_306);
xnor U6306 (N_6306,N_1457,N_2189);
and U6307 (N_6307,N_3556,N_4533);
nor U6308 (N_6308,N_3817,N_25);
nand U6309 (N_6309,N_5693,N_2662);
and U6310 (N_6310,N_907,N_2673);
and U6311 (N_6311,N_2964,N_78);
or U6312 (N_6312,N_2356,N_2483);
nor U6313 (N_6313,N_4005,N_2791);
nor U6314 (N_6314,N_369,N_1358);
nand U6315 (N_6315,N_2055,N_511);
xnor U6316 (N_6316,N_273,N_4276);
nand U6317 (N_6317,N_4750,N_6116);
or U6318 (N_6318,N_4621,N_447);
or U6319 (N_6319,N_6143,N_1637);
nand U6320 (N_6320,N_2918,N_2242);
nand U6321 (N_6321,N_2629,N_4484);
or U6322 (N_6322,N_5019,N_4730);
nand U6323 (N_6323,N_4336,N_3428);
or U6324 (N_6324,N_3956,N_2834);
or U6325 (N_6325,N_2637,N_5057);
nand U6326 (N_6326,N_739,N_3792);
xor U6327 (N_6327,N_4892,N_6187);
and U6328 (N_6328,N_4692,N_2812);
and U6329 (N_6329,N_1812,N_5480);
and U6330 (N_6330,N_4772,N_5383);
xnor U6331 (N_6331,N_2591,N_5914);
xnor U6332 (N_6332,N_5545,N_3744);
nor U6333 (N_6333,N_769,N_3198);
xor U6334 (N_6334,N_4244,N_2174);
nor U6335 (N_6335,N_1028,N_3418);
nand U6336 (N_6336,N_1272,N_2742);
xor U6337 (N_6337,N_1779,N_3990);
and U6338 (N_6338,N_3007,N_5679);
or U6339 (N_6339,N_3046,N_1256);
nor U6340 (N_6340,N_2073,N_3177);
nand U6341 (N_6341,N_2221,N_2154);
and U6342 (N_6342,N_470,N_3168);
nor U6343 (N_6343,N_2140,N_1828);
and U6344 (N_6344,N_2121,N_957);
nand U6345 (N_6345,N_5376,N_2912);
nor U6346 (N_6346,N_2255,N_4359);
or U6347 (N_6347,N_1703,N_3855);
nor U6348 (N_6348,N_5539,N_3759);
or U6349 (N_6349,N_5810,N_4115);
nand U6350 (N_6350,N_129,N_459);
nand U6351 (N_6351,N_2922,N_4473);
and U6352 (N_6352,N_5793,N_978);
nor U6353 (N_6353,N_2103,N_3783);
nand U6354 (N_6354,N_1924,N_2645);
and U6355 (N_6355,N_1230,N_4275);
nand U6356 (N_6356,N_291,N_5682);
nand U6357 (N_6357,N_2752,N_2233);
nand U6358 (N_6358,N_2899,N_5748);
or U6359 (N_6359,N_5279,N_4616);
nand U6360 (N_6360,N_2884,N_5104);
nand U6361 (N_6361,N_655,N_3774);
nand U6362 (N_6362,N_4067,N_3015);
or U6363 (N_6363,N_2753,N_4482);
and U6364 (N_6364,N_3715,N_3589);
or U6365 (N_6365,N_1052,N_159);
and U6366 (N_6366,N_2850,N_489);
and U6367 (N_6367,N_1579,N_5603);
and U6368 (N_6368,N_5811,N_689);
and U6369 (N_6369,N_3602,N_5116);
or U6370 (N_6370,N_218,N_5642);
and U6371 (N_6371,N_2247,N_3521);
nor U6372 (N_6372,N_2407,N_2901);
nor U6373 (N_6373,N_4537,N_4838);
and U6374 (N_6374,N_1134,N_2041);
nor U6375 (N_6375,N_3565,N_0);
and U6376 (N_6376,N_3607,N_2487);
nand U6377 (N_6377,N_3323,N_4615);
xnor U6378 (N_6378,N_6041,N_5059);
nor U6379 (N_6379,N_4294,N_2913);
and U6380 (N_6380,N_455,N_5342);
nand U6381 (N_6381,N_5360,N_2231);
nand U6382 (N_6382,N_1627,N_3445);
and U6383 (N_6383,N_3184,N_4219);
or U6384 (N_6384,N_3501,N_4626);
nor U6385 (N_6385,N_4898,N_4924);
or U6386 (N_6386,N_2663,N_4221);
xnor U6387 (N_6387,N_797,N_3626);
xor U6388 (N_6388,N_3224,N_1001);
nor U6389 (N_6389,N_731,N_5952);
and U6390 (N_6390,N_1033,N_2605);
nand U6391 (N_6391,N_3298,N_2581);
nor U6392 (N_6392,N_3303,N_5751);
nand U6393 (N_6393,N_755,N_1614);
nand U6394 (N_6394,N_436,N_5168);
nor U6395 (N_6395,N_4056,N_5688);
or U6396 (N_6396,N_96,N_5233);
and U6397 (N_6397,N_1138,N_5187);
or U6398 (N_6398,N_3236,N_6006);
nor U6399 (N_6399,N_2872,N_4521);
nand U6400 (N_6400,N_5198,N_2720);
nor U6401 (N_6401,N_2162,N_5542);
nor U6402 (N_6402,N_5906,N_2107);
nand U6403 (N_6403,N_2744,N_6182);
and U6404 (N_6404,N_3373,N_2430);
or U6405 (N_6405,N_6170,N_1195);
nor U6406 (N_6406,N_5591,N_3505);
xnor U6407 (N_6407,N_5113,N_4760);
nor U6408 (N_6408,N_5126,N_2725);
and U6409 (N_6409,N_2439,N_5053);
or U6410 (N_6410,N_3125,N_3735);
or U6411 (N_6411,N_5441,N_1660);
and U6412 (N_6412,N_1181,N_1311);
nand U6413 (N_6413,N_5246,N_2965);
xor U6414 (N_6414,N_4877,N_3919);
or U6415 (N_6415,N_5926,N_1042);
nand U6416 (N_6416,N_3689,N_2651);
and U6417 (N_6417,N_814,N_3761);
nor U6418 (N_6418,N_2788,N_1902);
nand U6419 (N_6419,N_6191,N_1620);
nor U6420 (N_6420,N_2340,N_2484);
nor U6421 (N_6421,N_64,N_5734);
or U6422 (N_6422,N_5247,N_631);
nand U6423 (N_6423,N_4190,N_3773);
nor U6424 (N_6424,N_3378,N_5715);
nor U6425 (N_6425,N_624,N_6236);
and U6426 (N_6426,N_238,N_1456);
and U6427 (N_6427,N_475,N_3999);
nand U6428 (N_6428,N_493,N_1989);
or U6429 (N_6429,N_4801,N_4901);
nand U6430 (N_6430,N_2690,N_5692);
or U6431 (N_6431,N_4462,N_231);
or U6432 (N_6432,N_5499,N_5838);
and U6433 (N_6433,N_1549,N_5128);
nand U6434 (N_6434,N_4265,N_2153);
or U6435 (N_6435,N_191,N_4287);
nand U6436 (N_6436,N_2759,N_1861);
nor U6437 (N_6437,N_2893,N_4572);
xor U6438 (N_6438,N_2448,N_4790);
nor U6439 (N_6439,N_1510,N_5489);
or U6440 (N_6440,N_1880,N_5590);
or U6441 (N_6441,N_3695,N_1727);
and U6442 (N_6442,N_3880,N_6022);
xnor U6443 (N_6443,N_1332,N_3078);
nand U6444 (N_6444,N_2717,N_2074);
and U6445 (N_6445,N_1190,N_709);
nor U6446 (N_6446,N_1261,N_3476);
or U6447 (N_6447,N_666,N_5308);
nor U6448 (N_6448,N_5686,N_3732);
nor U6449 (N_6449,N_4514,N_1977);
xnor U6450 (N_6450,N_3606,N_522);
nand U6451 (N_6451,N_3708,N_3424);
or U6452 (N_6452,N_3686,N_2318);
nor U6453 (N_6453,N_2403,N_4340);
nand U6454 (N_6454,N_2787,N_5042);
or U6455 (N_6455,N_3662,N_760);
or U6456 (N_6456,N_2226,N_6240);
nand U6457 (N_6457,N_4673,N_1937);
and U6458 (N_6458,N_5905,N_305);
nand U6459 (N_6459,N_4003,N_3392);
and U6460 (N_6460,N_498,N_5690);
or U6461 (N_6461,N_714,N_4856);
nand U6462 (N_6462,N_6192,N_3642);
nor U6463 (N_6463,N_3684,N_2931);
or U6464 (N_6464,N_2993,N_1928);
and U6465 (N_6465,N_5959,N_5791);
and U6466 (N_6466,N_4367,N_5215);
and U6467 (N_6467,N_2832,N_2590);
or U6468 (N_6468,N_5784,N_2096);
or U6469 (N_6469,N_4025,N_2889);
nand U6470 (N_6470,N_1952,N_546);
and U6471 (N_6471,N_398,N_5164);
or U6472 (N_6472,N_3203,N_3118);
and U6473 (N_6473,N_2664,N_2846);
nand U6474 (N_6474,N_2997,N_1189);
or U6475 (N_6475,N_1923,N_325);
or U6476 (N_6476,N_4288,N_1273);
and U6477 (N_6477,N_3232,N_1246);
or U6478 (N_6478,N_2296,N_3713);
xnor U6479 (N_6479,N_1583,N_3605);
nand U6480 (N_6480,N_4303,N_4365);
nand U6481 (N_6481,N_2186,N_124);
or U6482 (N_6482,N_2995,N_827);
nor U6483 (N_6483,N_719,N_501);
or U6484 (N_6484,N_5744,N_5435);
nand U6485 (N_6485,N_5795,N_2792);
nor U6486 (N_6486,N_2397,N_2085);
nand U6487 (N_6487,N_258,N_2566);
or U6488 (N_6488,N_632,N_2953);
or U6489 (N_6489,N_621,N_3658);
xnor U6490 (N_6490,N_1499,N_1161);
nand U6491 (N_6491,N_5722,N_2497);
and U6492 (N_6492,N_3912,N_463);
nor U6493 (N_6493,N_6066,N_516);
and U6494 (N_6494,N_1663,N_920);
and U6495 (N_6495,N_4836,N_2774);
or U6496 (N_6496,N_5765,N_4550);
xnor U6497 (N_6497,N_1178,N_2277);
and U6498 (N_6498,N_3044,N_134);
nor U6499 (N_6499,N_4,N_5989);
or U6500 (N_6500,N_4420,N_2502);
and U6501 (N_6501,N_1903,N_2088);
nand U6502 (N_6502,N_5641,N_2279);
nand U6503 (N_6503,N_5622,N_5779);
or U6504 (N_6504,N_999,N_1142);
nor U6505 (N_6505,N_861,N_4180);
xnor U6506 (N_6506,N_5630,N_1186);
nor U6507 (N_6507,N_2385,N_2926);
nor U6508 (N_6508,N_4110,N_3472);
xor U6509 (N_6509,N_5340,N_2676);
xnor U6510 (N_6510,N_2429,N_806);
or U6511 (N_6511,N_4907,N_2090);
xnor U6512 (N_6512,N_454,N_6168);
nand U6513 (N_6513,N_2544,N_6058);
nand U6514 (N_6514,N_4001,N_2089);
nor U6515 (N_6515,N_2881,N_610);
or U6516 (N_6516,N_3871,N_2500);
nand U6517 (N_6517,N_771,N_2008);
nor U6518 (N_6518,N_3274,N_989);
nor U6519 (N_6519,N_5970,N_2132);
nand U6520 (N_6520,N_1648,N_5217);
nand U6521 (N_6521,N_5865,N_5423);
xor U6522 (N_6522,N_3398,N_6220);
or U6523 (N_6523,N_5892,N_1055);
or U6524 (N_6524,N_5592,N_2421);
or U6525 (N_6525,N_2921,N_132);
nand U6526 (N_6526,N_418,N_4900);
or U6527 (N_6527,N_5052,N_1742);
and U6528 (N_6528,N_245,N_1316);
nor U6529 (N_6529,N_4218,N_4169);
nand U6530 (N_6530,N_2061,N_2498);
nand U6531 (N_6531,N_2406,N_4940);
nor U6532 (N_6532,N_5106,N_2895);
and U6533 (N_6533,N_3486,N_721);
and U6534 (N_6534,N_429,N_6205);
nand U6535 (N_6535,N_4771,N_5260);
or U6536 (N_6536,N_3857,N_3115);
or U6537 (N_6537,N_2391,N_4691);
or U6538 (N_6538,N_2026,N_394);
nand U6539 (N_6539,N_2422,N_1407);
or U6540 (N_6540,N_5492,N_4006);
or U6541 (N_6541,N_3220,N_3191);
or U6542 (N_6542,N_5139,N_3267);
or U6543 (N_6543,N_4595,N_5840);
xnor U6544 (N_6544,N_770,N_5913);
and U6545 (N_6545,N_2288,N_1623);
and U6546 (N_6546,N_2256,N_5268);
nand U6547 (N_6547,N_5929,N_2811);
and U6548 (N_6548,N_2178,N_1271);
or U6549 (N_6549,N_693,N_6027);
and U6550 (N_6550,N_4752,N_2719);
or U6551 (N_6551,N_5685,N_3535);
nor U6552 (N_6552,N_4463,N_1757);
and U6553 (N_6553,N_168,N_4422);
xnor U6554 (N_6554,N_6070,N_4131);
nor U6555 (N_6555,N_2253,N_1211);
nor U6556 (N_6556,N_5928,N_3601);
and U6557 (N_6557,N_4126,N_4822);
nand U6558 (N_6558,N_3213,N_4748);
nor U6559 (N_6559,N_1561,N_1177);
nor U6560 (N_6560,N_1452,N_3076);
nand U6561 (N_6561,N_3229,N_5829);
and U6562 (N_6562,N_5498,N_1964);
nor U6563 (N_6563,N_870,N_4008);
and U6564 (N_6564,N_4204,N_3622);
nor U6565 (N_6565,N_4174,N_5798);
or U6566 (N_6566,N_5200,N_1864);
nand U6567 (N_6567,N_836,N_3061);
nor U6568 (N_6568,N_5796,N_2749);
and U6569 (N_6569,N_3139,N_1221);
or U6570 (N_6570,N_2799,N_4364);
nor U6571 (N_6571,N_3681,N_2819);
and U6572 (N_6572,N_4609,N_311);
and U6573 (N_6573,N_1149,N_1080);
nand U6574 (N_6574,N_2489,N_164);
nor U6575 (N_6575,N_1507,N_3780);
nand U6576 (N_6576,N_1064,N_691);
or U6577 (N_6577,N_3557,N_3109);
and U6578 (N_6578,N_443,N_3301);
and U6579 (N_6579,N_648,N_788);
and U6580 (N_6580,N_5302,N_2337);
nand U6581 (N_6581,N_6232,N_5319);
and U6582 (N_6582,N_662,N_4850);
nor U6583 (N_6583,N_5061,N_653);
and U6584 (N_6584,N_2207,N_1093);
nor U6585 (N_6585,N_3748,N_1790);
or U6586 (N_6586,N_3087,N_3442);
or U6587 (N_6587,N_6131,N_3820);
and U6588 (N_6588,N_3917,N_469);
nand U6589 (N_6589,N_2547,N_3515);
nor U6590 (N_6590,N_1689,N_3936);
and U6591 (N_6591,N_3964,N_521);
or U6592 (N_6592,N_101,N_3733);
nand U6593 (N_6593,N_4164,N_365);
or U6594 (N_6594,N_3562,N_2350);
nor U6595 (N_6595,N_3215,N_4886);
xnor U6596 (N_6596,N_5957,N_5945);
nand U6597 (N_6597,N_2550,N_1766);
nor U6598 (N_6598,N_6098,N_4992);
and U6599 (N_6599,N_888,N_5131);
nor U6600 (N_6600,N_4211,N_3370);
nor U6601 (N_6601,N_4459,N_1558);
or U6602 (N_6602,N_6044,N_1108);
nor U6603 (N_6603,N_5743,N_3927);
xor U6604 (N_6604,N_5420,N_3390);
or U6605 (N_6605,N_4077,N_3103);
or U6606 (N_6606,N_1262,N_565);
nor U6607 (N_6607,N_4251,N_6062);
or U6608 (N_6608,N_2761,N_5310);
or U6609 (N_6609,N_4358,N_2348);
and U6610 (N_6610,N_1213,N_2560);
nand U6611 (N_6611,N_2248,N_1225);
or U6612 (N_6612,N_528,N_4338);
and U6613 (N_6613,N_5875,N_223);
and U6614 (N_6614,N_4304,N_5226);
nand U6615 (N_6615,N_3063,N_4208);
xnor U6616 (N_6616,N_5396,N_4542);
or U6617 (N_6617,N_5493,N_3402);
and U6618 (N_6618,N_1845,N_3978);
or U6619 (N_6619,N_5457,N_2038);
and U6620 (N_6620,N_4577,N_3039);
nand U6621 (N_6621,N_2595,N_5065);
and U6622 (N_6622,N_6053,N_308);
and U6623 (N_6623,N_4929,N_2685);
nand U6624 (N_6624,N_5017,N_4347);
nand U6625 (N_6625,N_4425,N_5083);
or U6626 (N_6626,N_3644,N_5465);
xor U6627 (N_6627,N_2769,N_3668);
or U6628 (N_6628,N_5425,N_6206);
and U6629 (N_6629,N_2567,N_5315);
or U6630 (N_6630,N_1053,N_3721);
nand U6631 (N_6631,N_1085,N_1473);
and U6632 (N_6632,N_160,N_5801);
nand U6633 (N_6633,N_2346,N_3954);
xnor U6634 (N_6634,N_1884,N_3040);
or U6635 (N_6635,N_5123,N_2488);
and U6636 (N_6636,N_4402,N_3105);
nand U6637 (N_6637,N_4674,N_4627);
or U6638 (N_6638,N_883,N_3838);
or U6639 (N_6639,N_4150,N_787);
nand U6640 (N_6640,N_381,N_188);
nand U6641 (N_6641,N_4400,N_6169);
or U6642 (N_6642,N_3908,N_4483);
xor U6643 (N_6643,N_4580,N_2493);
and U6644 (N_6644,N_525,N_4060);
xor U6645 (N_6645,N_3434,N_4575);
or U6646 (N_6646,N_3102,N_1811);
nor U6647 (N_6647,N_951,N_2149);
nand U6648 (N_6648,N_3878,N_1467);
or U6649 (N_6649,N_2815,N_5627);
xor U6650 (N_6650,N_2896,N_2113);
nor U6651 (N_6651,N_1240,N_4464);
and U6652 (N_6652,N_3348,N_1393);
nor U6653 (N_6653,N_765,N_2275);
nand U6654 (N_6654,N_3849,N_83);
nand U6655 (N_6655,N_3764,N_2444);
and U6656 (N_6656,N_3423,N_5011);
xor U6657 (N_6657,N_2521,N_5063);
nand U6658 (N_6658,N_1842,N_5588);
or U6659 (N_6659,N_1597,N_1799);
nand U6660 (N_6660,N_321,N_2136);
nand U6661 (N_6661,N_530,N_3380);
nor U6662 (N_6662,N_2798,N_5277);
xnor U6663 (N_6663,N_2943,N_2830);
nand U6664 (N_6664,N_1258,N_3329);
or U6665 (N_6665,N_5307,N_4374);
xnor U6666 (N_6666,N_3616,N_1062);
nor U6667 (N_6667,N_819,N_562);
or U6668 (N_6668,N_4032,N_1185);
nor U6669 (N_6669,N_4096,N_2682);
nand U6670 (N_6670,N_6184,N_2092);
nor U6671 (N_6671,N_1744,N_1763);
nor U6672 (N_6672,N_917,N_1343);
or U6673 (N_6673,N_1012,N_98);
and U6674 (N_6674,N_1450,N_4565);
nand U6675 (N_6675,N_4243,N_4234);
nor U6676 (N_6676,N_3057,N_3197);
or U6677 (N_6677,N_3987,N_3794);
nand U6678 (N_6678,N_2644,N_3116);
or U6679 (N_6679,N_684,N_3711);
and U6680 (N_6680,N_3969,N_4184);
and U6681 (N_6681,N_5047,N_563);
xnor U6682 (N_6682,N_3189,N_6189);
nor U6683 (N_6683,N_4997,N_2621);
nand U6684 (N_6684,N_4270,N_3459);
and U6685 (N_6685,N_3417,N_2050);
and U6686 (N_6686,N_3186,N_4369);
nand U6687 (N_6687,N_342,N_294);
and U6688 (N_6688,N_442,N_3050);
nor U6689 (N_6689,N_4194,N_389);
nor U6690 (N_6690,N_4848,N_4883);
and U6691 (N_6691,N_1982,N_4751);
nand U6692 (N_6692,N_1530,N_3330);
or U6693 (N_6693,N_2710,N_2083);
or U6694 (N_6694,N_3547,N_4593);
nand U6695 (N_6695,N_6198,N_1596);
or U6696 (N_6696,N_5931,N_5280);
and U6697 (N_6697,N_1398,N_3974);
nor U6698 (N_6698,N_5256,N_1600);
nor U6699 (N_6699,N_2857,N_217);
nand U6700 (N_6700,N_207,N_5884);
and U6701 (N_6701,N_3464,N_933);
and U6702 (N_6702,N_3079,N_5180);
nor U6703 (N_6703,N_1708,N_3449);
or U6704 (N_6704,N_3122,N_3584);
nand U6705 (N_6705,N_4398,N_1518);
and U6706 (N_6706,N_569,N_1775);
or U6707 (N_6707,N_3381,N_5272);
nor U6708 (N_6708,N_3988,N_5450);
and U6709 (N_6709,N_3159,N_1544);
and U6710 (N_6710,N_5717,N_6081);
nor U6711 (N_6711,N_4535,N_5559);
nor U6712 (N_6712,N_1961,N_3003);
or U6713 (N_6713,N_2698,N_3344);
or U6714 (N_6714,N_5817,N_4185);
nor U6715 (N_6715,N_5286,N_2920);
nor U6716 (N_6716,N_3368,N_5570);
nand U6717 (N_6717,N_1575,N_3130);
xor U6718 (N_6718,N_3529,N_3829);
or U6719 (N_6719,N_5610,N_3870);
nor U6720 (N_6720,N_6229,N_829);
and U6721 (N_6721,N_1797,N_2104);
nand U6722 (N_6722,N_4817,N_3929);
nand U6723 (N_6723,N_2152,N_3045);
and U6724 (N_6724,N_5954,N_5626);
and U6725 (N_6725,N_2184,N_4293);
nor U6726 (N_6726,N_2196,N_4503);
nand U6727 (N_6727,N_479,N_3913);
or U6728 (N_6728,N_2908,N_4348);
or U6729 (N_6729,N_5872,N_816);
nor U6730 (N_6730,N_2115,N_3327);
or U6731 (N_6731,N_3004,N_4882);
nand U6732 (N_6732,N_2400,N_1014);
nand U6733 (N_6733,N_5469,N_40);
nand U6734 (N_6734,N_4305,N_3725);
and U6735 (N_6735,N_2613,N_5548);
nand U6736 (N_6736,N_2584,N_5546);
or U6737 (N_6737,N_3724,N_1427);
and U6738 (N_6738,N_4183,N_1586);
nor U6739 (N_6739,N_4754,N_5400);
nand U6740 (N_6740,N_3798,N_1434);
nand U6741 (N_6741,N_6149,N_4529);
nor U6742 (N_6742,N_2843,N_3570);
and U6743 (N_6743,N_1346,N_4435);
nor U6744 (N_6744,N_5073,N_108);
or U6745 (N_6745,N_4939,N_1022);
nand U6746 (N_6746,N_2431,N_1432);
and U6747 (N_6747,N_636,N_2582);
nor U6748 (N_6748,N_4443,N_5703);
nand U6749 (N_6749,N_6175,N_5012);
and U6750 (N_6750,N_1041,N_3238);
and U6751 (N_6751,N_4741,N_5834);
or U6752 (N_6752,N_5245,N_3770);
or U6753 (N_6753,N_3207,N_1141);
xnor U6754 (N_6754,N_2696,N_2117);
or U6755 (N_6755,N_1255,N_4870);
or U6756 (N_6756,N_668,N_1043);
and U6757 (N_6757,N_3223,N_6241);
and U6758 (N_6758,N_4745,N_5809);
and U6759 (N_6759,N_3270,N_2963);
or U6760 (N_6760,N_3135,N_3875);
nand U6761 (N_6761,N_681,N_1382);
nand U6762 (N_6762,N_5852,N_558);
xnor U6763 (N_6763,N_1418,N_264);
or U6764 (N_6764,N_4372,N_3740);
and U6765 (N_6765,N_4531,N_5443);
and U6766 (N_6766,N_4203,N_5941);
nor U6767 (N_6767,N_5220,N_4442);
nor U6768 (N_6768,N_4547,N_437);
nor U6769 (N_6769,N_537,N_5389);
nor U6770 (N_6770,N_3884,N_2370);
nand U6771 (N_6771,N_6215,N_2699);
and U6772 (N_6772,N_665,N_4157);
nand U6773 (N_6773,N_5500,N_1194);
and U6774 (N_6774,N_155,N_3636);
nand U6775 (N_6775,N_1249,N_975);
and U6776 (N_6776,N_4371,N_4023);
nand U6777 (N_6777,N_6012,N_2765);
and U6778 (N_6778,N_4798,N_3852);
nand U6779 (N_6779,N_5384,N_3613);
nor U6780 (N_6780,N_1698,N_5481);
nor U6781 (N_6781,N_2986,N_2093);
and U6782 (N_6782,N_6005,N_1445);
nor U6783 (N_6783,N_6172,N_4661);
and U6784 (N_6784,N_4642,N_2777);
nand U6785 (N_6785,N_1686,N_598);
nand U6786 (N_6786,N_2649,N_439);
xor U6787 (N_6787,N_5419,N_1867);
nand U6788 (N_6788,N_2924,N_4292);
or U6789 (N_6789,N_1943,N_41);
and U6790 (N_6790,N_4705,N_3036);
or U6791 (N_6791,N_4281,N_984);
or U6792 (N_6792,N_2326,N_4970);
and U6793 (N_6793,N_1389,N_4624);
xor U6794 (N_6794,N_1006,N_5681);
nand U6795 (N_6795,N_4853,N_5487);
or U6796 (N_6796,N_768,N_3660);
nor U6797 (N_6797,N_5949,N_67);
and U6798 (N_6798,N_3996,N_146);
or U6799 (N_6799,N_2951,N_574);
and U6800 (N_6800,N_5265,N_4197);
and U6801 (N_6801,N_1061,N_3782);
and U6802 (N_6802,N_2958,N_2883);
or U6803 (N_6803,N_1949,N_117);
or U6804 (N_6804,N_3552,N_4935);
nand U6805 (N_6805,N_4296,N_5696);
nor U6806 (N_6806,N_2928,N_6114);
or U6807 (N_6807,N_2261,N_4914);
and U6808 (N_6808,N_5231,N_3172);
or U6809 (N_6809,N_4306,N_5074);
nor U6810 (N_6810,N_3819,N_3810);
and U6811 (N_6811,N_3287,N_5090);
or U6812 (N_6812,N_3372,N_1191);
and U6813 (N_6813,N_2005,N_1859);
nand U6814 (N_6814,N_2658,N_3856);
and U6815 (N_6815,N_1426,N_5109);
or U6816 (N_6816,N_348,N_5413);
or U6817 (N_6817,N_4048,N_3179);
nand U6818 (N_6818,N_918,N_2244);
nor U6819 (N_6819,N_4544,N_1980);
xnor U6820 (N_6820,N_5386,N_541);
and U6821 (N_6821,N_5115,N_1215);
nand U6822 (N_6822,N_2434,N_2873);
or U6823 (N_6823,N_3253,N_402);
nor U6824 (N_6824,N_3869,N_2564);
or U6825 (N_6825,N_4796,N_4522);
nand U6826 (N_6826,N_5214,N_5602);
or U6827 (N_6827,N_2210,N_6217);
or U6828 (N_6828,N_3407,N_2833);
xnor U6829 (N_6829,N_5510,N_1865);
and U6830 (N_6830,N_2723,N_5740);
or U6831 (N_6831,N_555,N_3261);
nand U6832 (N_6832,N_4002,N_2329);
nand U6833 (N_6833,N_2655,N_3347);
nand U6834 (N_6834,N_589,N_1403);
xor U6835 (N_6835,N_3574,N_2372);
xnor U6836 (N_6836,N_4539,N_5161);
nand U6837 (N_6837,N_6124,N_1264);
and U6838 (N_6838,N_3337,N_3032);
nand U6839 (N_6839,N_4816,N_2029);
nor U6840 (N_6840,N_1863,N_2976);
nand U6841 (N_6841,N_3243,N_1328);
nor U6842 (N_6842,N_3395,N_412);
and U6843 (N_6843,N_128,N_2627);
or U6844 (N_6844,N_4598,N_4659);
or U6845 (N_6845,N_5025,N_1585);
xor U6846 (N_6846,N_519,N_3316);
nor U6847 (N_6847,N_1163,N_1210);
nor U6848 (N_6848,N_3359,N_4682);
xor U6849 (N_6849,N_496,N_4740);
nand U6850 (N_6850,N_2084,N_1103);
and U6851 (N_6851,N_5656,N_1617);
and U6852 (N_6852,N_858,N_5325);
nor U6853 (N_6853,N_2359,N_3541);
nand U6854 (N_6854,N_5985,N_409);
and U6855 (N_6855,N_2606,N_5759);
and U6856 (N_6856,N_1184,N_1926);
or U6857 (N_6857,N_3382,N_341);
and U6858 (N_6858,N_4507,N_6025);
or U6859 (N_6859,N_4102,N_5221);
nor U6860 (N_6860,N_4317,N_529);
nor U6861 (N_6861,N_6065,N_3800);
xnor U6862 (N_6862,N_2894,N_3144);
and U6863 (N_6863,N_6171,N_3893);
nor U6864 (N_6864,N_5756,N_6033);
or U6865 (N_6865,N_2257,N_2365);
or U6866 (N_6866,N_5111,N_2570);
and U6867 (N_6867,N_5196,N_727);
and U6868 (N_6868,N_659,N_5758);
nand U6869 (N_6869,N_1645,N_6127);
nor U6870 (N_6870,N_1629,N_2989);
nor U6871 (N_6871,N_6129,N_4264);
or U6872 (N_6872,N_2527,N_5227);
nor U6873 (N_6873,N_3767,N_5009);
and U6874 (N_6874,N_4241,N_332);
and U6875 (N_6875,N_5399,N_2433);
and U6876 (N_6876,N_1688,N_5034);
and U6877 (N_6877,N_1187,N_1063);
or U6878 (N_6878,N_2079,N_3384);
and U6879 (N_6879,N_1071,N_3910);
and U6880 (N_6880,N_5624,N_3221);
or U6881 (N_6881,N_316,N_901);
nor U6882 (N_6882,N_2373,N_5857);
and U6883 (N_6883,N_3731,N_1312);
and U6884 (N_6884,N_4592,N_2646);
xor U6885 (N_6885,N_200,N_2063);
and U6886 (N_6886,N_1453,N_105);
nor U6887 (N_6887,N_3319,N_427);
nor U6888 (N_6888,N_5364,N_3414);
nand U6889 (N_6889,N_2598,N_315);
xor U6890 (N_6890,N_4829,N_4053);
and U6891 (N_6891,N_5851,N_2888);
and U6892 (N_6892,N_6023,N_4468);
nand U6893 (N_6893,N_3518,N_2124);
and U6894 (N_6894,N_5922,N_650);
xor U6895 (N_6895,N_2990,N_3190);
nand U6896 (N_6896,N_80,N_4323);
and U6897 (N_6897,N_6145,N_6218);
nor U6898 (N_6898,N_4825,N_2094);
xor U6899 (N_6899,N_4384,N_4387);
and U6900 (N_6900,N_1634,N_5427);
nand U6901 (N_6901,N_6030,N_3980);
nand U6902 (N_6902,N_4007,N_3802);
and U6903 (N_6903,N_2474,N_937);
xnor U6904 (N_6904,N_5710,N_4827);
xor U6905 (N_6905,N_540,N_3690);
nor U6906 (N_6906,N_60,N_254);
nand U6907 (N_6907,N_3193,N_891);
nor U6908 (N_6908,N_3548,N_1833);
nand U6909 (N_6909,N_2344,N_490);
or U6910 (N_6910,N_5638,N_3113);
or U6911 (N_6911,N_5547,N_5752);
nor U6912 (N_6912,N_3655,N_5655);
or U6913 (N_6913,N_1386,N_3504);
or U6914 (N_6914,N_375,N_3482);
and U6915 (N_6915,N_1628,N_5856);
and U6916 (N_6916,N_5040,N_3326);
or U6917 (N_6917,N_266,N_1994);
nor U6918 (N_6918,N_18,N_4637);
xnor U6919 (N_6919,N_3095,N_3132);
or U6920 (N_6920,N_3700,N_5071);
nand U6921 (N_6921,N_2361,N_5295);
and U6922 (N_6922,N_890,N_4638);
nor U6923 (N_6923,N_3072,N_6102);
nand U6924 (N_6924,N_1564,N_2935);
and U6925 (N_6925,N_2035,N_4412);
nor U6926 (N_6926,N_3332,N_6176);
nand U6927 (N_6927,N_3961,N_1168);
or U6928 (N_6928,N_970,N_1515);
or U6929 (N_6929,N_784,N_4461);
nor U6930 (N_6930,N_87,N_5640);
nand U6931 (N_6931,N_1260,N_2848);
or U6932 (N_6932,N_35,N_4087);
or U6933 (N_6933,N_4114,N_2401);
nand U6934 (N_6934,N_1953,N_1337);
and U6935 (N_6935,N_1218,N_3101);
or U6936 (N_6936,N_3091,N_4132);
and U6937 (N_6937,N_3951,N_1487);
or U6938 (N_6938,N_5583,N_4207);
nand U6939 (N_6939,N_687,N_4749);
nand U6940 (N_6940,N_3020,N_5863);
and U6941 (N_6941,N_5978,N_945);
nand U6942 (N_6942,N_643,N_4910);
and U6943 (N_6943,N_695,N_1622);
nor U6944 (N_6944,N_4497,N_1731);
nand U6945 (N_6945,N_4681,N_4041);
and U6946 (N_6946,N_4653,N_1874);
nand U6947 (N_6947,N_4499,N_4538);
nor U6948 (N_6948,N_1069,N_1543);
xnor U6949 (N_6949,N_6103,N_2838);
or U6950 (N_6950,N_652,N_6136);
nand U6951 (N_6951,N_467,N_3981);
nand U6952 (N_6952,N_710,N_4298);
nor U6953 (N_6953,N_664,N_5428);
nor U6954 (N_6954,N_2985,N_362);
and U6955 (N_6955,N_3208,N_1245);
nand U6956 (N_6956,N_2071,N_1746);
nand U6957 (N_6957,N_5720,N_5550);
and U6958 (N_6958,N_766,N_4419);
nand U6959 (N_6959,N_2371,N_3010);
xor U6960 (N_6960,N_5097,N_5648);
nor U6961 (N_6961,N_5484,N_4187);
or U6962 (N_6962,N_3409,N_2106);
nand U6963 (N_6963,N_1931,N_1661);
or U6964 (N_6964,N_1409,N_161);
nor U6965 (N_6965,N_2641,N_502);
nand U6966 (N_6966,N_6135,N_2782);
or U6967 (N_6967,N_5297,N_6222);
nand U6968 (N_6968,N_1472,N_5845);
xnor U6969 (N_6969,N_3768,N_3771);
and U6970 (N_6970,N_2158,N_110);
or U6971 (N_6971,N_2300,N_3062);
nand U6972 (N_6972,N_505,N_3466);
and U6973 (N_6973,N_1986,N_5658);
and U6974 (N_6974,N_2501,N_1758);
and U6975 (N_6975,N_1146,N_2952);
or U6976 (N_6976,N_869,N_4927);
or U6977 (N_6977,N_4396,N_3047);
and U6978 (N_6978,N_5424,N_899);
or U6979 (N_6979,N_1153,N_4065);
or U6980 (N_6980,N_488,N_980);
xnor U6981 (N_6981,N_567,N_355);
and U6982 (N_6982,N_4971,N_3833);
nor U6983 (N_6983,N_3879,N_3357);
nor U6984 (N_6984,N_5899,N_6100);
or U6985 (N_6985,N_4236,N_446);
or U6986 (N_6986,N_724,N_5939);
nand U6987 (N_6987,N_4302,N_5725);
nor U6988 (N_6988,N_5653,N_374);
nor U6989 (N_6989,N_4328,N_1878);
or U6990 (N_6990,N_805,N_4788);
or U6991 (N_6991,N_4502,N_1886);
or U6992 (N_6992,N_4523,N_3592);
nand U6993 (N_6993,N_3456,N_5584);
nor U6994 (N_6994,N_5924,N_5527);
nor U6995 (N_6995,N_2388,N_1370);
nor U6996 (N_6996,N_3022,N_4330);
and U6997 (N_6997,N_3926,N_3006);
and U6998 (N_6998,N_1339,N_3753);
or U6999 (N_6999,N_376,N_2416);
or U7000 (N_7000,N_3104,N_1765);
and U7001 (N_7001,N_2554,N_5918);
nand U7002 (N_7002,N_4668,N_6076);
and U7003 (N_7003,N_1520,N_3614);
and U7004 (N_7004,N_2659,N_6163);
or U7005 (N_7005,N_889,N_2054);
or U7006 (N_7006,N_904,N_4310);
and U7007 (N_7007,N_5405,N_3000);
nand U7008 (N_7008,N_6173,N_3450);
and U7009 (N_7009,N_1201,N_1723);
or U7010 (N_7010,N_2847,N_3830);
xor U7011 (N_7011,N_5543,N_1545);
or U7012 (N_7012,N_5329,N_599);
nand U7013 (N_7013,N_74,N_4257);
or U7014 (N_7014,N_4408,N_1718);
nand U7015 (N_7015,N_4278,N_1947);
or U7016 (N_7016,N_4012,N_841);
nand U7017 (N_7017,N_3968,N_4307);
nand U7018 (N_7018,N_3314,N_840);
or U7019 (N_7019,N_2171,N_5431);
or U7020 (N_7020,N_4256,N_5596);
nand U7021 (N_7021,N_1443,N_4839);
and U7022 (N_7022,N_4489,N_4647);
or U7023 (N_7023,N_4163,N_391);
nand U7024 (N_7024,N_343,N_756);
xor U7025 (N_7025,N_2642,N_1428);
nor U7026 (N_7026,N_4201,N_3488);
and U7027 (N_7027,N_5996,N_2841);
nor U7028 (N_7028,N_301,N_5770);
or U7029 (N_7029,N_4631,N_3310);
and U7030 (N_7030,N_2380,N_4118);
and U7031 (N_7031,N_5379,N_1344);
and U7032 (N_7032,N_5045,N_965);
and U7033 (N_7033,N_6115,N_13);
or U7034 (N_7034,N_5575,N_1078);
xor U7035 (N_7035,N_2375,N_5771);
nor U7036 (N_7036,N_1956,N_837);
xor U7037 (N_7037,N_6207,N_5948);
and U7038 (N_7038,N_6133,N_6085);
and U7039 (N_7039,N_276,N_5582);
or U7040 (N_7040,N_4312,N_1322);
nor U7041 (N_7041,N_1948,N_5299);
xor U7042 (N_7042,N_4113,N_5745);
nand U7043 (N_7043,N_189,N_431);
or U7044 (N_7044,N_5967,N_5615);
and U7045 (N_7045,N_425,N_3608);
nand U7046 (N_7046,N_4506,N_364);
nor U7047 (N_7047,N_54,N_4229);
xor U7048 (N_7048,N_4120,N_5084);
xor U7049 (N_7049,N_5485,N_1335);
nand U7050 (N_7050,N_2389,N_617);
or U7051 (N_7051,N_5205,N_5154);
and U7052 (N_7052,N_6050,N_3300);
xnor U7053 (N_7053,N_5563,N_3264);
nand U7054 (N_7054,N_2491,N_5446);
xor U7055 (N_7055,N_3550,N_3824);
nand U7056 (N_7056,N_3728,N_5188);
xnor U7057 (N_7057,N_651,N_1590);
nor U7058 (N_7058,N_1820,N_3339);
xnor U7059 (N_7059,N_3242,N_5651);
nor U7060 (N_7060,N_1008,N_3140);
or U7061 (N_7061,N_1853,N_845);
and U7062 (N_7062,N_4460,N_4979);
xnor U7063 (N_7063,N_2764,N_3473);
and U7064 (N_7064,N_1981,N_1164);
nor U7065 (N_7065,N_5529,N_3458);
nor U7066 (N_7066,N_2315,N_3196);
nand U7067 (N_7067,N_2616,N_2721);
or U7068 (N_7068,N_5531,N_3639);
nor U7069 (N_7069,N_5055,N_1838);
or U7070 (N_7070,N_3752,N_4619);
or U7071 (N_7071,N_1803,N_623);
or U7072 (N_7072,N_4016,N_206);
and U7073 (N_7073,N_3112,N_2862);
and U7074 (N_7074,N_1175,N_4127);
nand U7075 (N_7075,N_5432,N_5600);
nand U7076 (N_7076,N_1709,N_4076);
and U7077 (N_7077,N_407,N_3995);
and U7078 (N_7078,N_3312,N_5430);
and U7079 (N_7079,N_3136,N_3657);
nor U7080 (N_7080,N_3944,N_4719);
or U7081 (N_7081,N_5411,N_507);
or U7082 (N_7082,N_5356,N_5674);
nor U7083 (N_7083,N_1917,N_2217);
nand U7084 (N_7084,N_2194,N_704);
nand U7085 (N_7085,N_417,N_3942);
nor U7086 (N_7086,N_3572,N_4332);
or U7087 (N_7087,N_1105,N_3507);
and U7088 (N_7088,N_4658,N_1151);
and U7089 (N_7089,N_2902,N_5082);
or U7090 (N_7090,N_5134,N_5385);
and U7091 (N_7091,N_5987,N_3389);
or U7092 (N_7092,N_4516,N_678);
and U7093 (N_7093,N_1659,N_3874);
and U7094 (N_7094,N_220,N_4679);
and U7095 (N_7095,N_2075,N_1714);
nand U7096 (N_7096,N_4090,N_2192);
or U7097 (N_7097,N_1073,N_781);
nor U7098 (N_7098,N_4413,N_5010);
nor U7099 (N_7099,N_1514,N_1632);
nor U7100 (N_7100,N_1649,N_2364);
nor U7101 (N_7101,N_3313,N_1348);
nand U7102 (N_7102,N_2718,N_5598);
nor U7103 (N_7103,N_5652,N_1652);
xnor U7104 (N_7104,N_3133,N_5718);
or U7105 (N_7105,N_6239,N_5254);
and U7106 (N_7106,N_576,N_4167);
nor U7107 (N_7107,N_4930,N_2133);
and U7108 (N_7108,N_5398,N_5966);
or U7109 (N_7109,N_6054,N_3801);
or U7110 (N_7110,N_1422,N_3164);
nor U7111 (N_7111,N_833,N_4568);
and U7112 (N_7112,N_4718,N_1145);
nand U7113 (N_7113,N_125,N_4437);
and U7114 (N_7114,N_4318,N_828);
and U7115 (N_7115,N_5662,N_5294);
nor U7116 (N_7116,N_5107,N_2760);
nor U7117 (N_7117,N_5069,N_3603);
nor U7118 (N_7118,N_4729,N_672);
nand U7119 (N_7119,N_4403,N_4540);
xor U7120 (N_7120,N_1474,N_3526);
nor U7121 (N_7121,N_2983,N_5901);
nand U7122 (N_7122,N_4843,N_3863);
nand U7123 (N_7123,N_2119,N_4297);
nand U7124 (N_7124,N_1536,N_4246);
and U7125 (N_7125,N_6209,N_4649);
nor U7126 (N_7126,N_3487,N_2508);
nor U7127 (N_7127,N_5714,N_1684);
nor U7128 (N_7128,N_2796,N_3576);
xor U7129 (N_7129,N_4222,N_5418);
nand U7130 (N_7130,N_3825,N_274);
nand U7131 (N_7131,N_1233,N_3053);
and U7132 (N_7132,N_2612,N_4472);
or U7133 (N_7133,N_4248,N_1104);
or U7134 (N_7134,N_4876,N_5380);
nand U7135 (N_7135,N_4085,N_3726);
nor U7136 (N_7136,N_5917,N_1342);
nand U7137 (N_7137,N_3131,N_5062);
or U7138 (N_7138,N_3998,N_775);
and U7139 (N_7139,N_3510,N_5552);
nand U7140 (N_7140,N_2517,N_3017);
xor U7141 (N_7141,N_585,N_4478);
and U7142 (N_7142,N_3730,N_3026);
nor U7143 (N_7143,N_4975,N_5092);
or U7144 (N_7144,N_3815,N_4470);
or U7145 (N_7145,N_359,N_4352);
and U7146 (N_7146,N_5887,N_5409);
nor U7147 (N_7147,N_874,N_2030);
or U7148 (N_7148,N_2289,N_5158);
nor U7149 (N_7149,N_350,N_964);
and U7150 (N_7150,N_5763,N_3340);
nand U7151 (N_7151,N_4075,N_5339);
nor U7152 (N_7152,N_2482,N_6185);
nor U7153 (N_7153,N_4769,N_337);
nand U7154 (N_7154,N_1011,N_2531);
or U7155 (N_7155,N_2807,N_1229);
nor U7156 (N_7156,N_2166,N_2240);
and U7157 (N_7157,N_3343,N_3258);
nand U7158 (N_7158,N_4088,N_2737);
nor U7159 (N_7159,N_3460,N_5835);
nor U7160 (N_7160,N_1413,N_1480);
and U7161 (N_7161,N_2779,N_4043);
nor U7162 (N_7162,N_4144,N_267);
nand U7163 (N_7163,N_706,N_4380);
and U7164 (N_7164,N_3612,N_1420);
and U7165 (N_7165,N_5244,N_2609);
or U7166 (N_7166,N_3273,N_6034);
or U7167 (N_7167,N_4948,N_3846);
and U7168 (N_7168,N_5393,N_6013);
or U7169 (N_7169,N_4198,N_968);
nor U7170 (N_7170,N_2988,N_3991);
and U7171 (N_7171,N_3643,N_5841);
xor U7172 (N_7172,N_1762,N_5534);
or U7173 (N_7173,N_2909,N_1639);
or U7174 (N_7174,N_5262,N_285);
nor U7175 (N_7175,N_5309,N_3054);
and U7176 (N_7176,N_1729,N_3276);
xor U7177 (N_7177,N_4047,N_1017);
or U7178 (N_7178,N_5392,N_1726);
and U7179 (N_7179,N_3494,N_4343);
and U7180 (N_7180,N_3516,N_3345);
nor U7181 (N_7181,N_2632,N_2634);
and U7182 (N_7182,N_438,N_785);
xnor U7183 (N_7183,N_2987,N_4290);
nor U7184 (N_7184,N_4429,N_5728);
xor U7185 (N_7185,N_2545,N_5908);
nor U7186 (N_7186,N_1737,N_2227);
and U7187 (N_7187,N_885,N_1333);
or U7188 (N_7188,N_4956,N_6071);
nor U7189 (N_7189,N_4834,N_3377);
and U7190 (N_7190,N_4808,N_2962);
nor U7191 (N_7191,N_4917,N_4993);
and U7192 (N_7192,N_1509,N_5453);
and U7193 (N_7193,N_4737,N_5258);
and U7194 (N_7194,N_536,N_2449);
xor U7195 (N_7195,N_187,N_5802);
xnor U7196 (N_7196,N_5358,N_729);
xor U7197 (N_7197,N_4498,N_5988);
xor U7198 (N_7198,N_877,N_361);
and U7199 (N_7199,N_5572,N_5920);
nand U7200 (N_7200,N_3002,N_3182);
nor U7201 (N_7201,N_2293,N_4451);
or U7202 (N_7202,N_6084,N_5037);
xor U7203 (N_7203,N_4189,N_1040);
nor U7204 (N_7204,N_4936,N_5776);
and U7205 (N_7205,N_2597,N_243);
and U7206 (N_7206,N_1400,N_2181);
nand U7207 (N_7207,N_5355,N_2222);
nor U7208 (N_7208,N_4494,N_4019);
or U7209 (N_7209,N_4014,N_1615);
nand U7210 (N_7210,N_1279,N_2027);
or U7211 (N_7211,N_2381,N_916);
and U7212 (N_7212,N_6108,N_954);
nand U7213 (N_7213,N_4036,N_4465);
nor U7214 (N_7214,N_1756,N_4618);
nor U7215 (N_7215,N_2195,N_5911);
nor U7216 (N_7216,N_4570,N_2683);
nor U7217 (N_7217,N_2968,N_1120);
nand U7218 (N_7218,N_3610,N_4309);
or U7219 (N_7219,N_3904,N_2674);
and U7220 (N_7220,N_683,N_5830);
and U7221 (N_7221,N_3578,N_1392);
nand U7222 (N_7222,N_4584,N_1559);
or U7223 (N_7223,N_5808,N_5669);
xnor U7224 (N_7224,N_3365,N_2366);
or U7225 (N_7225,N_4554,N_4430);
nor U7226 (N_7226,N_75,N_5463);
nor U7227 (N_7227,N_4868,N_3383);
xnor U7228 (N_7228,N_5273,N_4230);
nor U7229 (N_7229,N_228,N_1039);
nor U7230 (N_7230,N_2984,N_2572);
or U7231 (N_7231,N_6067,N_3491);
and U7232 (N_7232,N_1707,N_2004);
and U7233 (N_7233,N_2076,N_2060);
or U7234 (N_7234,N_5540,N_1241);
and U7235 (N_7235,N_5354,N_5516);
nand U7236 (N_7236,N_1846,N_2414);
or U7237 (N_7237,N_3335,N_4696);
nand U7238 (N_7238,N_2996,N_2464);
nor U7239 (N_7239,N_179,N_2168);
nand U7240 (N_7240,N_2604,N_4951);
nand U7241 (N_7241,N_4964,N_4765);
nor U7242 (N_7242,N_2459,N_1992);
or U7243 (N_7243,N_3143,N_43);
nor U7244 (N_7244,N_794,N_1873);
nand U7245 (N_7245,N_5684,N_2080);
nand U7246 (N_7246,N_4921,N_1315);
xnor U7247 (N_7247,N_1721,N_3369);
and U7248 (N_7248,N_3154,N_1007);
and U7249 (N_7249,N_747,N_5160);
and U7250 (N_7250,N_2214,N_2602);
and U7251 (N_7251,N_1469,N_3067);
nand U7252 (N_7252,N_6078,N_4987);
xnor U7253 (N_7253,N_2308,N_6141);
nand U7254 (N_7254,N_5761,N_3940);
or U7255 (N_7255,N_4984,N_4329);
nor U7256 (N_7256,N_3128,N_4438);
xnor U7257 (N_7257,N_663,N_313);
and U7258 (N_7258,N_2305,N_2722);
nand U7259 (N_7259,N_5787,N_2417);
nor U7260 (N_7260,N_3262,N_1182);
or U7261 (N_7261,N_234,N_3333);
nor U7262 (N_7262,N_497,N_2820);
nor U7263 (N_7263,N_3822,N_1114);
or U7264 (N_7264,N_628,N_6040);
xnor U7265 (N_7265,N_1209,N_5677);
or U7266 (N_7266,N_3850,N_4530);
nand U7267 (N_7267,N_2529,N_4345);
or U7268 (N_7268,N_4242,N_4613);
and U7269 (N_7269,N_1355,N_5773);
nor U7270 (N_7270,N_2599,N_1606);
and U7271 (N_7271,N_4717,N_2472);
nor U7272 (N_7272,N_5096,N_3755);
or U7273 (N_7273,N_988,N_147);
or U7274 (N_7274,N_3886,N_1748);
or U7275 (N_7275,N_1388,N_6099);
and U7276 (N_7276,N_1512,N_962);
xnor U7277 (N_7277,N_3781,N_2568);
or U7278 (N_7278,N_4324,N_2465);
and U7279 (N_7279,N_1004,N_4988);
nor U7280 (N_7280,N_4286,N_4040);
nand U7281 (N_7281,N_2827,N_4145);
nand U7282 (N_7282,N_4362,N_5317);
nand U7283 (N_7283,N_4556,N_263);
or U7284 (N_7284,N_6147,N_2387);
nand U7285 (N_7285,N_1015,N_3888);
and U7286 (N_7286,N_4015,N_4648);
nor U7287 (N_7287,N_3031,N_914);
or U7288 (N_7288,N_1119,N_1437);
nand U7289 (N_7289,N_5502,N_72);
and U7290 (N_7290,N_5351,N_1111);
or U7291 (N_7291,N_994,N_140);
nor U7292 (N_7292,N_4654,N_5292);
and U7293 (N_7293,N_5607,N_1722);
xnor U7294 (N_7294,N_4153,N_4555);
nand U7295 (N_7295,N_2949,N_926);
and U7296 (N_7296,N_339,N_3973);
and U7297 (N_7297,N_5449,N_2713);
and U7298 (N_7298,N_1808,N_2183);
and U7299 (N_7299,N_956,N_5050);
or U7300 (N_7300,N_1088,N_3311);
nor U7301 (N_7301,N_5697,N_4046);
nand U7302 (N_7302,N_1882,N_19);
xor U7303 (N_7303,N_89,N_212);
and U7304 (N_7304,N_3282,N_2781);
or U7305 (N_7305,N_564,N_5031);
and U7306 (N_7306,N_464,N_4212);
or U7307 (N_7307,N_4937,N_6195);
and U7308 (N_7308,N_4273,N_1654);
xnor U7309 (N_7309,N_5375,N_2563);
nand U7310 (N_7310,N_1132,N_416);
or U7311 (N_7311,N_3257,N_5016);
nand U7312 (N_7312,N_2543,N_5496);
nand U7313 (N_7313,N_5706,N_5623);
or U7314 (N_7314,N_113,N_2622);
nand U7315 (N_7315,N_2813,N_333);
or U7316 (N_7316,N_130,N_400);
xor U7317 (N_7317,N_6228,N_5708);
xnor U7318 (N_7318,N_3239,N_3881);
nand U7319 (N_7319,N_3483,N_4084);
and U7320 (N_7320,N_2748,N_5225);
and U7321 (N_7321,N_510,N_3266);
and U7322 (N_7322,N_4289,N_1984);
nand U7323 (N_7323,N_2185,N_1881);
or U7324 (N_7324,N_5883,N_953);
or U7325 (N_7325,N_928,N_3906);
or U7326 (N_7326,N_4316,N_458);
or U7327 (N_7327,N_1533,N_3060);
nand U7328 (N_7328,N_2640,N_5046);
nor U7329 (N_7329,N_4199,N_1560);
xnor U7330 (N_7330,N_1200,N_4712);
and U7331 (N_7331,N_3955,N_1650);
nor U7332 (N_7332,N_5363,N_6123);
and U7333 (N_7333,N_4284,N_2853);
nor U7334 (N_7334,N_1385,N_1761);
nand U7335 (N_7335,N_3174,N_4259);
nand U7336 (N_7336,N_4802,N_5108);
nand U7337 (N_7337,N_1167,N_645);
or U7338 (N_7338,N_5344,N_56);
and U7339 (N_7339,N_2786,N_1631);
nand U7340 (N_7340,N_3844,N_1492);
or U7341 (N_7341,N_2516,N_1725);
nor U7342 (N_7342,N_5417,N_3422);
or U7343 (N_7343,N_3279,N_4726);
and U7344 (N_7344,N_4635,N_4721);
xnor U7345 (N_7345,N_2903,N_3283);
nand U7346 (N_7346,N_4059,N_2398);
nand U7347 (N_7347,N_2409,N_4042);
nor U7348 (N_7348,N_5460,N_487);
and U7349 (N_7349,N_204,N_210);
nand U7350 (N_7350,N_2310,N_4337);
nand U7351 (N_7351,N_1293,N_3334);
or U7352 (N_7352,N_1849,N_581);
and U7353 (N_7353,N_3408,N_1144);
and U7354 (N_7354,N_2405,N_5112);
and U7355 (N_7355,N_3948,N_1609);
xor U7356 (N_7356,N_992,N_1449);
nor U7357 (N_7357,N_1321,N_5284);
nand U7358 (N_7358,N_3065,N_5889);
or U7359 (N_7359,N_2826,N_208);
and U7360 (N_7360,N_95,N_5594);
and U7361 (N_7361,N_5660,N_1656);
nor U7362 (N_7362,N_707,N_5896);
and U7363 (N_7363,N_5526,N_5156);
or U7364 (N_7364,N_2379,N_1323);
and U7365 (N_7365,N_452,N_453);
nor U7366 (N_7366,N_6161,N_3743);
nor U7367 (N_7367,N_209,N_5940);
nand U7368 (N_7368,N_2675,N_5155);
nand U7369 (N_7369,N_973,N_2858);
nand U7370 (N_7370,N_2596,N_3317);
nor U7371 (N_7371,N_3204,N_5049);
and U7372 (N_7372,N_5132,N_358);
nand U7373 (N_7373,N_2190,N_1983);
nand U7374 (N_7374,N_2942,N_590);
nor U7375 (N_7375,N_5020,N_3900);
xor U7376 (N_7376,N_5422,N_1127);
or U7377 (N_7377,N_3412,N_3304);
nand U7378 (N_7378,N_2911,N_1895);
nand U7379 (N_7379,N_4123,N_3228);
nor U7380 (N_7380,N_3124,N_657);
nand U7381 (N_7381,N_2821,N_4268);
xnor U7382 (N_7382,N_3845,N_3597);
nand U7383 (N_7383,N_5,N_1307);
nor U7384 (N_7384,N_1822,N_2797);
and U7385 (N_7385,N_5843,N_4849);
nor U7386 (N_7386,N_1049,N_1286);
nor U7387 (N_7387,N_5912,N_3089);
or U7388 (N_7388,N_3127,N_5525);
xnor U7389 (N_7389,N_941,N_717);
and U7390 (N_7390,N_3363,N_1257);
and U7391 (N_7391,N_3977,N_4686);
or U7392 (N_7392,N_1697,N_5533);
nand U7393 (N_7393,N_3092,N_843);
or U7394 (N_7394,N_3269,N_1493);
nand U7395 (N_7395,N_5879,N_1951);
nand U7396 (N_7396,N_677,N_2555);
or U7397 (N_7397,N_4704,N_5440);
and U7398 (N_7398,N_4695,N_5946);
and U7399 (N_7399,N_5554,N_4385);
xnor U7400 (N_7400,N_959,N_3151);
nand U7401 (N_7401,N_3630,N_1122);
nor U7402 (N_7402,N_4645,N_4976);
nand U7403 (N_7403,N_377,N_2357);
nand U7404 (N_7404,N_3860,N_971);
nor U7405 (N_7405,N_5599,N_309);
or U7406 (N_7406,N_2750,N_1180);
and U7407 (N_7407,N_1188,N_5491);
nor U7408 (N_7408,N_4103,N_910);
or U7409 (N_7409,N_834,N_5519);
nor U7410 (N_7410,N_330,N_5984);
nand U7411 (N_7411,N_278,N_3949);
nand U7412 (N_7412,N_281,N_4955);
nor U7413 (N_7413,N_560,N_2138);
nand U7414 (N_7414,N_3352,N_4179);
xnor U7415 (N_7415,N_5303,N_5324);
or U7416 (N_7416,N_1414,N_1957);
and U7417 (N_7417,N_1202,N_1635);
nor U7418 (N_7418,N_2828,N_2736);
nor U7419 (N_7419,N_5005,N_723);
or U7420 (N_7420,N_1301,N_2694);
nand U7421 (N_7421,N_2436,N_6242);
nor U7422 (N_7422,N_4770,N_1173);
and U7423 (N_7423,N_2824,N_532);
nand U7424 (N_7424,N_524,N_991);
or U7425 (N_7425,N_3038,N_4919);
or U7426 (N_7426,N_955,N_817);
nand U7427 (N_7427,N_4793,N_4282);
nand U7428 (N_7428,N_4162,N_1636);
and U7429 (N_7429,N_1702,N_1837);
xnor U7430 (N_7430,N_1996,N_6052);
nand U7431 (N_7431,N_357,N_404);
or U7432 (N_7432,N_4024,N_1976);
or U7433 (N_7433,N_114,N_1856);
nor U7434 (N_7434,N_3049,N_3666);
and U7435 (N_7435,N_4685,N_5736);
nand U7436 (N_7436,N_4379,N_3985);
nor U7437 (N_7437,N_5494,N_297);
and U7438 (N_7438,N_1379,N_5105);
and U7439 (N_7439,N_3024,N_2882);
xor U7440 (N_7440,N_5338,N_4215);
xnor U7441 (N_7441,N_5359,N_1562);
or U7442 (N_7442,N_3265,N_4266);
or U7443 (N_7443,N_4700,N_6094);
or U7444 (N_7444,N_1809,N_2112);
and U7445 (N_7445,N_4787,N_5824);
nand U7446 (N_7446,N_177,N_1970);
nand U7447 (N_7447,N_733,N_1136);
nor U7448 (N_7448,N_1118,N_2577);
nor U7449 (N_7449,N_1967,N_1045);
or U7450 (N_7450,N_2512,N_906);
nor U7451 (N_7451,N_4166,N_2503);
nand U7452 (N_7452,N_3983,N_4009);
xnor U7453 (N_7453,N_448,N_1248);
or U7454 (N_7454,N_3898,N_2789);
xor U7455 (N_7455,N_863,N_2098);
nor U7456 (N_7456,N_2886,N_5998);
and U7457 (N_7457,N_2460,N_3199);
nor U7458 (N_7458,N_2163,N_5024);
or U7459 (N_7459,N_6204,N_2033);
xnor U7460 (N_7460,N_250,N_4452);
or U7461 (N_7461,N_3052,N_2541);
nand U7462 (N_7462,N_1847,N_4879);
or U7463 (N_7463,N_4641,N_2814);
and U7464 (N_7464,N_6132,N_866);
and U7465 (N_7465,N_6210,N_3650);
or U7466 (N_7466,N_441,N_4755);
nor U7467 (N_7467,N_2803,N_2352);
and U7468 (N_7468,N_1594,N_5099);
or U7469 (N_7469,N_5578,N_613);
xor U7470 (N_7470,N_5505,N_1870);
and U7471 (N_7471,N_4612,N_2540);
xor U7472 (N_7472,N_738,N_3088);
nand U7473 (N_7473,N_2457,N_1839);
and U7474 (N_7474,N_29,N_5538);
or U7475 (N_7475,N_5523,N_2410);
or U7476 (N_7476,N_2972,N_3872);
and U7477 (N_7477,N_4766,N_4599);
and U7478 (N_7478,N_5520,N_1728);
or U7479 (N_7479,N_3836,N_3294);
nor U7480 (N_7480,N_4453,N_1179);
nor U7481 (N_7481,N_3138,N_3789);
nand U7482 (N_7482,N_5894,N_639);
or U7483 (N_7483,N_5557,N_3281);
and U7484 (N_7484,N_5844,N_1907);
and U7485 (N_7485,N_5337,N_5298);
and U7486 (N_7486,N_3540,N_1253);
nand U7487 (N_7487,N_4622,N_4952);
and U7488 (N_7488,N_976,N_2919);
xnor U7489 (N_7489,N_4747,N_76);
or U7490 (N_7490,N_772,N_5001);
and U7491 (N_7491,N_2955,N_3571);
and U7492 (N_7492,N_1868,N_334);
nor U7493 (N_7493,N_518,N_2565);
nand U7494 (N_7494,N_4656,N_2209);
and U7495 (N_7495,N_2123,N_5482);
nor U7496 (N_7496,N_1804,N_3702);
nor U7497 (N_7497,N_3947,N_5095);
or U7498 (N_7498,N_908,N_6048);
nor U7499 (N_7499,N_782,N_5782);
xor U7500 (N_7500,N_2999,N_3816);
nor U7501 (N_7501,N_5964,N_3453);
nand U7502 (N_7502,N_2100,N_4475);
or U7503 (N_7503,N_4382,N_547);
xor U7504 (N_7504,N_5091,N_3148);
nand U7505 (N_7505,N_948,N_2874);
nand U7506 (N_7506,N_1935,N_5234);
or U7507 (N_7507,N_6036,N_4694);
and U7508 (N_7508,N_4436,N_3451);
nor U7509 (N_7509,N_2776,N_3862);
nor U7510 (N_7510,N_4319,N_3692);
nor U7511 (N_7511,N_3379,N_2510);
nor U7512 (N_7512,N_1896,N_2109);
nor U7513 (N_7513,N_1079,N_5676);
nor U7514 (N_7514,N_5293,N_2078);
nor U7515 (N_7515,N_831,N_2576);
nor U7516 (N_7516,N_6045,N_3509);
and U7517 (N_7517,N_2324,N_3769);
and U7518 (N_7518,N_2341,N_232);
or U7519 (N_7519,N_1550,N_2548);
and U7520 (N_7520,N_5232,N_2445);
nand U7521 (N_7521,N_2630,N_4908);
nor U7522 (N_7522,N_835,N_3183);
nor U7523 (N_7523,N_5322,N_2784);
and U7524 (N_7524,N_2322,N_4606);
and U7525 (N_7525,N_6223,N_1563);
nor U7526 (N_7526,N_786,N_2302);
xnor U7527 (N_7527,N_868,N_1356);
xnor U7528 (N_7528,N_3762,N_3683);
nand U7529 (N_7529,N_2313,N_4057);
nand U7530 (N_7530,N_1914,N_1274);
xnor U7531 (N_7531,N_4650,N_5436);
nand U7532 (N_7532,N_5224,N_750);
nor U7533 (N_7533,N_4999,N_3260);
and U7534 (N_7534,N_5289,N_3231);
nor U7535 (N_7535,N_4271,N_1658);
nand U7536 (N_7536,N_1593,N_921);
nand U7537 (N_7537,N_1198,N_4723);
or U7538 (N_7538,N_4073,N_1675);
xor U7539 (N_7539,N_2518,N_4672);
xor U7540 (N_7540,N_5240,N_2386);
and U7541 (N_7541,N_5038,N_5118);
nand U7542 (N_7542,N_4871,N_981);
nand U7543 (N_7543,N_2741,N_4195);
nand U7544 (N_7544,N_5026,N_4069);
nor U7545 (N_7545,N_3754,N_3651);
and U7546 (N_7546,N_503,N_5230);
and U7547 (N_7547,N_4082,N_1599);
or U7548 (N_7548,N_2923,N_5737);
xor U7549 (N_7549,N_1013,N_939);
nand U7550 (N_7550,N_3058,N_3882);
or U7551 (N_7551,N_5657,N_3873);
or U7552 (N_7552,N_553,N_4854);
or U7553 (N_7553,N_5614,N_214);
or U7554 (N_7554,N_5731,N_1667);
xor U7555 (N_7555,N_5606,N_3701);
nor U7556 (N_7556,N_1199,N_3965);
or U7557 (N_7557,N_4559,N_3216);
or U7558 (N_7558,N_3325,N_1451);
xnor U7559 (N_7559,N_4128,N_1565);
xnor U7560 (N_7560,N_5314,N_934);
nand U7561 (N_7561,N_4576,N_2619);
xor U7562 (N_7562,N_477,N_5408);
xor U7563 (N_7563,N_2520,N_4549);
and U7564 (N_7564,N_79,N_2200);
xnor U7565 (N_7565,N_3210,N_2763);
and U7566 (N_7566,N_6087,N_1484);
and U7567 (N_7567,N_4154,N_3524);
or U7568 (N_7568,N_2775,N_1025);
nor U7569 (N_7569,N_2961,N_1827);
nand U7570 (N_7570,N_1557,N_884);
nor U7571 (N_7571,N_5125,N_4149);
xor U7572 (N_7572,N_5093,N_2587);
and U7573 (N_7573,N_71,N_314);
nor U7574 (N_7574,N_6117,N_3938);
nor U7575 (N_7575,N_3638,N_3005);
nand U7576 (N_7576,N_1772,N_4223);
nand U7577 (N_7577,N_1160,N_2402);
xnor U7578 (N_7578,N_4346,N_2959);
or U7579 (N_7579,N_2608,N_801);
nand U7580 (N_7580,N_486,N_1436);
and U7581 (N_7581,N_251,N_4603);
xnor U7582 (N_7582,N_1125,N_1566);
nor U7583 (N_7583,N_1056,N_3799);
nand U7584 (N_7584,N_6219,N_608);
nor U7585 (N_7585,N_808,N_2618);
and U7586 (N_7586,N_1444,N_865);
nor U7587 (N_7587,N_4778,N_226);
xnor U7588 (N_7588,N_3247,N_1433);
or U7589 (N_7589,N_1706,N_4168);
nand U7590 (N_7590,N_3374,N_2973);
or U7591 (N_7591,N_198,N_5476);
and U7592 (N_7592,N_3566,N_1086);
or U7593 (N_7593,N_1292,N_1121);
or U7594 (N_7594,N_157,N_495);
and U7595 (N_7595,N_2927,N_4688);
nor U7596 (N_7596,N_51,N_3661);
and U7597 (N_7597,N_3214,N_1899);
nor U7598 (N_7598,N_4487,N_386);
or U7599 (N_7599,N_4200,N_6126);
or U7600 (N_7600,N_1753,N_3443);
xnor U7601 (N_7601,N_3520,N_3962);
and U7602 (N_7602,N_430,N_4564);
nand U7603 (N_7603,N_960,N_640);
nor U7604 (N_7604,N_5935,N_4476);
nor U7605 (N_7605,N_1699,N_3360);
and U7606 (N_7606,N_5434,N_3484);
nand U7607 (N_7607,N_2636,N_5199);
xor U7608 (N_7608,N_3842,N_1618);
nor U7609 (N_7609,N_1305,N_352);
nor U7610 (N_7610,N_3522,N_824);
and U7611 (N_7611,N_3226,N_4874);
nand U7612 (N_7612,N_6015,N_406);
or U7613 (N_7613,N_773,N_3388);
or U7614 (N_7614,N_4859,N_5486);
or U7615 (N_7615,N_1854,N_1387);
or U7616 (N_7616,N_3465,N_38);
xnor U7617 (N_7617,N_4962,N_3885);
or U7618 (N_7618,N_1810,N_5098);
and U7619 (N_7619,N_520,N_6202);
nand U7620 (N_7620,N_1551,N_2128);
or U7621 (N_7621,N_5165,N_4108);
and U7622 (N_7622,N_2480,N_53);
or U7623 (N_7623,N_5805,N_5475);
and U7624 (N_7624,N_897,N_2716);
or U7625 (N_7625,N_5506,N_2979);
nand U7626 (N_7626,N_4657,N_1817);
xnor U7627 (N_7627,N_3963,N_5173);
xnor U7628 (N_7628,N_5942,N_2426);
or U7629 (N_7629,N_4414,N_2533);
or U7630 (N_7630,N_4666,N_3315);
or U7631 (N_7631,N_300,N_1680);
and U7632 (N_7632,N_2869,N_449);
nor U7633 (N_7633,N_4277,N_3945);
nand U7634 (N_7634,N_3085,N_3222);
nand U7635 (N_7635,N_1470,N_3763);
nand U7636 (N_7636,N_428,N_1522);
or U7637 (N_7637,N_5323,N_857);
or U7638 (N_7638,N_673,N_5081);
nand U7639 (N_7639,N_5067,N_1024);
or U7640 (N_7640,N_549,N_1626);
or U7641 (N_7641,N_5947,N_2929);
nor U7642 (N_7642,N_491,N_3237);
and U7643 (N_7643,N_545,N_202);
nand U7644 (N_7644,N_2446,N_3331);
nor U7645 (N_7645,N_603,N_1438);
and U7646 (N_7646,N_48,N_1657);
and U7647 (N_7647,N_5671,N_4667);
nand U7648 (N_7648,N_106,N_2118);
nor U7649 (N_7649,N_5790,N_789);
nand U7650 (N_7650,N_5472,N_580);
nor U7651 (N_7651,N_3805,N_1455);
nand U7652 (N_7652,N_4086,N_6224);
or U7653 (N_7653,N_2575,N_979);
nand U7654 (N_7654,N_1975,N_1912);
or U7655 (N_7655,N_152,N_213);
nor U7656 (N_7656,N_4732,N_1059);
or U7657 (N_7657,N_5341,N_1821);
or U7658 (N_7658,N_6157,N_2443);
xor U7659 (N_7659,N_5646,N_4706);
xor U7660 (N_7660,N_832,N_3084);
or U7661 (N_7661,N_3814,N_896);
nor U7662 (N_7662,N_4781,N_1674);
xor U7663 (N_7663,N_2495,N_5511);
or U7664 (N_7664,N_6049,N_5910);
nand U7665 (N_7665,N_5711,N_5579);
and U7666 (N_7666,N_1236,N_748);
nand U7667 (N_7667,N_2285,N_4378);
and U7668 (N_7668,N_1378,N_6167);
xnor U7669 (N_7669,N_3828,N_5886);
nand U7670 (N_7670,N_3624,N_4186);
xnor U7671 (N_7671,N_3899,N_5175);
and U7672 (N_7672,N_100,N_1704);
nand U7673 (N_7673,N_1503,N_4226);
or U7674 (N_7674,N_5621,N_1341);
or U7675 (N_7675,N_69,N_1035);
nor U7676 (N_7676,N_4141,N_715);
or U7677 (N_7677,N_1244,N_3069);
nor U7678 (N_7678,N_172,N_1932);
or U7679 (N_7679,N_3353,N_6035);
nand U7680 (N_7680,N_426,N_3324);
nor U7681 (N_7681,N_4690,N_1197);
or U7682 (N_7682,N_2428,N_1217);
nand U7683 (N_7683,N_1377,N_4643);
or U7684 (N_7684,N_6146,N_6179);
nand U7685 (N_7685,N_1916,N_5466);
xor U7686 (N_7686,N_1439,N_5190);
or U7687 (N_7687,N_3493,N_1647);
nand U7688 (N_7688,N_4272,N_5859);
xor U7689 (N_7689,N_2733,N_6110);
nand U7690 (N_7690,N_556,N_5333);
nand U7691 (N_7691,N_742,N_1922);
and U7692 (N_7692,N_5870,N_5135);
and U7693 (N_7693,N_1883,N_746);
and U7694 (N_7694,N_4235,N_2534);
or U7695 (N_7695,N_2679,N_5639);
nand U7696 (N_7696,N_413,N_6227);
xor U7697 (N_7697,N_1300,N_2772);
and U7698 (N_7698,N_6234,N_4389);
nand U7699 (N_7699,N_4967,N_3142);
or U7700 (N_7700,N_3931,N_26);
nand U7701 (N_7701,N_1019,N_347);
nor U7702 (N_7702,N_4884,N_1616);
or U7703 (N_7703,N_4923,N_3362);
nor U7704 (N_7704,N_1165,N_360);
or U7705 (N_7705,N_5777,N_4509);
and U7706 (N_7706,N_4913,N_2625);
nand U7707 (N_7707,N_4571,N_4360);
nor U7708 (N_7708,N_983,N_4054);
or U7709 (N_7709,N_5403,N_3923);
or U7710 (N_7710,N_4017,N_1066);
and U7711 (N_7711,N_1242,N_3779);
nand U7712 (N_7712,N_1941,N_856);
nand U7713 (N_7713,N_5372,N_2105);
and U7714 (N_7714,N_5764,N_5858);
nor U7715 (N_7715,N_1776,N_4159);
or U7716 (N_7716,N_4731,N_627);
nand U7717 (N_7717,N_1044,N_1830);
nor U7718 (N_7718,N_1547,N_587);
or U7719 (N_7719,N_1998,N_3982);
nand U7720 (N_7720,N_5968,N_5980);
nand U7721 (N_7721,N_1691,N_4354);
nor U7722 (N_7722,N_17,N_1720);
nor U7723 (N_7723,N_5051,N_3600);
xnor U7724 (N_7724,N_2780,N_2110);
nor U7725 (N_7725,N_3682,N_2745);
xor U7726 (N_7726,N_3134,N_5437);
or U7727 (N_7727,N_2212,N_5792);
xor U7728 (N_7728,N_2173,N_4582);
nor U7729 (N_7729,N_2790,N_5571);
nor U7730 (N_7730,N_4983,N_2301);
xnor U7731 (N_7731,N_1893,N_3034);
nor U7732 (N_7732,N_2639,N_4736);
nor U7733 (N_7733,N_3457,N_6089);
xor U7734 (N_7734,N_2981,N_1973);
or U7735 (N_7735,N_2208,N_3922);
and U7736 (N_7736,N_2513,N_1365);
and U7737 (N_7737,N_1692,N_5617);
and U7738 (N_7738,N_1925,N_3837);
xnor U7739 (N_7739,N_4136,N_2709);
nand U7740 (N_7740,N_1075,N_3338);
and U7741 (N_7741,N_81,N_4524);
and U7742 (N_7742,N_1608,N_5670);
nand U7743 (N_7743,N_2031,N_4742);
nand U7744 (N_7744,N_5213,N_4035);
xor U7745 (N_7745,N_2808,N_800);
or U7746 (N_7746,N_4758,N_4944);
xnor U7747 (N_7747,N_6001,N_2251);
nand U7748 (N_7748,N_5556,N_6039);
and U7749 (N_7749,N_644,N_3568);
nor U7750 (N_7750,N_1479,N_3180);
nand U7751 (N_7751,N_4693,N_4106);
or U7752 (N_7752,N_3364,N_5732);
or U7753 (N_7753,N_5087,N_5694);
and U7754 (N_7754,N_3796,N_6010);
or U7755 (N_7755,N_5228,N_324);
or U7756 (N_7756,N_5659,N_961);
nand U7757 (N_7757,N_3158,N_2273);
or U7758 (N_7758,N_2970,N_3667);
xnor U7759 (N_7759,N_354,N_1872);
xor U7760 (N_7760,N_633,N_2477);
nor U7761 (N_7761,N_3217,N_3292);
and U7762 (N_7762,N_2933,N_3297);
or U7763 (N_7763,N_2490,N_1495);
or U7764 (N_7764,N_2852,N_133);
and U7765 (N_7765,N_2298,N_1431);
or U7766 (N_7766,N_4978,N_4663);
nor U7767 (N_7767,N_4339,N_385);
nor U7768 (N_7768,N_246,N_2139);
nor U7769 (N_7769,N_2254,N_3500);
and U7770 (N_7770,N_2461,N_3093);
nand U7771 (N_7771,N_2175,N_5854);
nand U7772 (N_7772,N_2353,N_4920);
or U7773 (N_7773,N_1574,N_4469);
and U7774 (N_7774,N_6162,N_2556);
and U7775 (N_7775,N_5006,N_3227);
nor U7776 (N_7776,N_345,N_986);
nand U7777 (N_7777,N_4409,N_5799);
and U7778 (N_7778,N_4558,N_606);
and U7779 (N_7779,N_5334,N_3117);
and U7780 (N_7780,N_4092,N_4895);
nor U7781 (N_7781,N_2479,N_2614);
nand U7782 (N_7782,N_411,N_1252);
nand U7783 (N_7783,N_3234,N_3200);
and U7784 (N_7784,N_1542,N_2611);
nor U7785 (N_7785,N_2610,N_4496);
xnor U7786 (N_7786,N_6092,N_4881);
nand U7787 (N_7787,N_3858,N_4701);
and U7788 (N_7788,N_3023,N_277);
and U7789 (N_7789,N_5569,N_5783);
or U7790 (N_7790,N_3225,N_1613);
or U7791 (N_7791,N_3404,N_974);
nand U7792 (N_7792,N_5266,N_5394);
and U7793 (N_7793,N_2463,N_2165);
nand U7794 (N_7794,N_795,N_1791);
nor U7795 (N_7795,N_15,N_3399);
nand U7796 (N_7796,N_4640,N_2336);
xor U7797 (N_7797,N_1026,N_3);
and U7798 (N_7798,N_3703,N_1000);
or U7799 (N_7799,N_5900,N_4206);
xnor U7800 (N_7800,N_3512,N_4121);
or U7801 (N_7801,N_6140,N_4308);
nor U7802 (N_7802,N_688,N_55);
and U7803 (N_7803,N_5332,N_3723);
nand U7804 (N_7804,N_2049,N_542);
nor U7805 (N_7805,N_5066,N_1603);
nor U7806 (N_7806,N_2904,N_1958);
or U7807 (N_7807,N_5140,N_3967);
xor U7808 (N_7808,N_4479,N_2667);
and U7809 (N_7809,N_10,N_614);
and U7810 (N_7810,N_1908,N_6077);
xnor U7811 (N_7811,N_1677,N_2867);
or U7812 (N_7812,N_4855,N_4431);
and U7813 (N_7813,N_6246,N_517);
or U7814 (N_7814,N_1371,N_790);
and U7815 (N_7815,N_3709,N_1174);
and U7816 (N_7816,N_2282,N_1641);
or U7817 (N_7817,N_1679,N_825);
nand U7818 (N_7818,N_2180,N_3175);
xor U7819 (N_7819,N_5353,N_743);
nand U7820 (N_7820,N_3532,N_3503);
nor U7821 (N_7821,N_4795,N_5919);
nor U7822 (N_7822,N_2532,N_635);
or U7823 (N_7823,N_5828,N_3867);
or U7824 (N_7824,N_5729,N_4756);
nor U7825 (N_7825,N_3957,N_5347);
nand U7826 (N_7826,N_2363,N_4233);
nand U7827 (N_7827,N_5054,N_3749);
nand U7828 (N_7828,N_5960,N_368);
and U7829 (N_7829,N_3795,N_6156);
nand U7830 (N_7830,N_5757,N_4807);
and U7831 (N_7831,N_3976,N_2437);
or U7832 (N_7832,N_4995,N_6112);
nor U7833 (N_7833,N_2687,N_4480);
nand U7834 (N_7834,N_3534,N_2442);
and U7835 (N_7835,N_5404,N_4563);
or U7836 (N_7836,N_5839,N_4142);
nand U7837 (N_7837,N_1835,N_5916);
nand U7838 (N_7838,N_3648,N_930);
nor U7839 (N_7839,N_6046,N_5586);
nand U7840 (N_7840,N_3474,N_1171);
or U7841 (N_7841,N_6008,N_4573);
and U7842 (N_7842,N_39,N_4320);
xnor U7843 (N_7843,N_949,N_2700);
xnor U7844 (N_7844,N_1447,N_1131);
and U7845 (N_7845,N_625,N_331);
and U7846 (N_7846,N_1999,N_820);
nor U7847 (N_7847,N_288,N_6166);
and U7848 (N_7848,N_85,N_5100);
or U7849 (N_7849,N_2203,N_1162);
or U7850 (N_7850,N_1361,N_4381);
nor U7851 (N_7851,N_1435,N_1226);
or U7852 (N_7852,N_2182,N_1681);
nand U7853 (N_7853,N_504,N_5631);
nand U7854 (N_7854,N_3187,N_2969);
and U7855 (N_7855,N_1621,N_450);
or U7856 (N_7856,N_2395,N_1227);
and U7857 (N_7857,N_1569,N_3933);
nand U7858 (N_7858,N_312,N_2785);
nor U7859 (N_7859,N_1094,N_3737);
nor U7860 (N_7860,N_4536,N_2102);
nor U7861 (N_7861,N_1270,N_2290);
or U7862 (N_7862,N_2805,N_592);
xnor U7863 (N_7863,N_4356,N_5312);
or U7864 (N_7864,N_4526,N_1446);
and U7865 (N_7865,N_1815,N_4291);
and U7866 (N_7866,N_2916,N_3157);
nor U7867 (N_7867,N_4862,N_127);
or U7868 (N_7868,N_3757,N_749);
nor U7869 (N_7869,N_2338,N_4066);
and U7870 (N_7870,N_5305,N_1773);
xnor U7871 (N_7871,N_809,N_158);
nor U7872 (N_7872,N_5028,N_3952);
or U7873 (N_7873,N_3654,N_5114);
and U7874 (N_7874,N_1031,N_1740);
nand U7875 (N_7875,N_3554,N_4158);
or U7876 (N_7876,N_5467,N_6063);
nand U7877 (N_7877,N_927,N_5391);
or U7878 (N_7878,N_6125,N_3656);
nor U7879 (N_7879,N_1237,N_2264);
nor U7880 (N_7880,N_5365,N_5963);
or U7881 (N_7881,N_3498,N_4508);
nand U7882 (N_7882,N_1936,N_5573);
nor U7883 (N_7883,N_4669,N_600);
nor U7884 (N_7884,N_5176,N_5837);
nor U7885 (N_7885,N_395,N_5197);
or U7886 (N_7886,N_5222,N_3788);
xor U7887 (N_7887,N_2450,N_1077);
or U7888 (N_7888,N_2526,N_3679);
nand U7889 (N_7889,N_3932,N_2323);
and U7890 (N_7890,N_1490,N_534);
and U7891 (N_7891,N_4493,N_2492);
nand U7892 (N_7892,N_1553,N_552);
nand U7893 (N_7893,N_1584,N_5907);
xnor U7894 (N_7894,N_6016,N_5008);
and U7895 (N_7895,N_4375,N_1051);
nor U7896 (N_7896,N_4761,N_2866);
and U7897 (N_7897,N_798,N_1834);
or U7898 (N_7898,N_2070,N_4147);
nor U7899 (N_7899,N_5831,N_2441);
and U7900 (N_7900,N_5397,N_3586);
nand U7901 (N_7901,N_2042,N_499);
or U7902 (N_7902,N_292,N_383);
nand U7903 (N_7903,N_5296,N_6003);
or U7904 (N_7904,N_1841,N_1003);
or U7905 (N_7905,N_2252,N_5562);
or U7906 (N_7906,N_764,N_879);
and U7907 (N_7907,N_2559,N_2551);
xnor U7908 (N_7908,N_1411,N_336);
nor U7909 (N_7909,N_5891,N_1546);
xnor U7910 (N_7910,N_6212,N_4133);
xor U7911 (N_7911,N_2053,N_5388);
xor U7912 (N_7912,N_2485,N_356);
xnor U7913 (N_7913,N_6178,N_1668);
and U7914 (N_7914,N_4202,N_685);
nand U7915 (N_7915,N_5285,N_2925);
and U7916 (N_7916,N_3675,N_1959);
and U7917 (N_7917,N_3587,N_1112);
or U7918 (N_7918,N_3580,N_4274);
nor U7919 (N_7919,N_618,N_3577);
and U7920 (N_7920,N_5975,N_5902);
xor U7921 (N_7921,N_1745,N_5048);
and U7922 (N_7922,N_423,N_73);
or U7923 (N_7923,N_2470,N_1768);
nand U7924 (N_7924,N_5961,N_4094);
nor U7925 (N_7925,N_5753,N_1710);
nand U7926 (N_7926,N_5876,N_3361);
xnor U7927 (N_7927,N_3549,N_1824);
and U7928 (N_7928,N_596,N_3588);
nor U7929 (N_7929,N_3386,N_1405);
nand U7930 (N_7930,N_1537,N_3746);
nand U7931 (N_7931,N_4989,N_2404);
xor U7932 (N_7932,N_1607,N_5921);
nand U7933 (N_7933,N_6096,N_1143);
nand U7934 (N_7934,N_1829,N_4405);
and U7935 (N_7935,N_3915,N_6082);
nand U7936 (N_7936,N_5760,N_3446);
or U7937 (N_7937,N_1076,N_1570);
nor U7938 (N_7938,N_4611,N_1644);
and U7939 (N_7939,N_3747,N_2274);
or U7940 (N_7940,N_1604,N_49);
nor U7941 (N_7941,N_112,N_5755);
nand U7942 (N_7942,N_1783,N_5846);
nor U7943 (N_7943,N_4125,N_2831);
xor U7944 (N_7944,N_3508,N_2283);
or U7945 (N_7945,N_2377,N_1813);
nand U7946 (N_7946,N_5373,N_4033);
xnor U7947 (N_7947,N_6237,N_4527);
nand U7948 (N_7948,N_3120,N_6029);
nand U7949 (N_7949,N_379,N_5171);
nand U7950 (N_7950,N_1653,N_3934);
nor U7951 (N_7951,N_6083,N_3623);
or U7952 (N_7952,N_2455,N_5813);
or U7953 (N_7953,N_1415,N_3984);
nor U7954 (N_7954,N_1166,N_99);
and U7955 (N_7955,N_1183,N_5288);
nand U7956 (N_7956,N_4018,N_2660);
or U7957 (N_7957,N_5553,N_420);
and U7958 (N_7958,N_5144,N_5874);
or U7959 (N_7959,N_607,N_642);
nor U7960 (N_7960,N_86,N_2937);
xnor U7961 (N_7961,N_6060,N_4518);
and U7962 (N_7962,N_2680,N_1376);
xnor U7963 (N_7963,N_5021,N_3935);
or U7964 (N_7964,N_5665,N_1851);
and U7965 (N_7965,N_3245,N_1892);
xnor U7966 (N_7966,N_4813,N_2052);
or U7967 (N_7967,N_4237,N_1712);
xor U7968 (N_7968,N_3527,N_1954);
nand U7969 (N_7969,N_6014,N_2552);
or U7970 (N_7970,N_5327,N_1423);
or U7971 (N_7971,N_6104,N_4050);
nor U7972 (N_7972,N_4961,N_2447);
nand U7973 (N_7973,N_1116,N_6037);
nand U7974 (N_7974,N_6199,N_5157);
xnor U7975 (N_7975,N_2334,N_4038);
nand U7976 (N_7976,N_1318,N_6155);
nor U7977 (N_7977,N_6190,N_3716);
xor U7978 (N_7978,N_1030,N_286);
or U7979 (N_7979,N_2879,N_1023);
nor U7980 (N_7980,N_2213,N_378);
nor U7981 (N_7981,N_6056,N_4664);
and U7982 (N_7982,N_2330,N_2871);
nand U7983 (N_7983,N_317,N_3941);
nor U7984 (N_7984,N_3477,N_4488);
nor U7985 (N_7985,N_2367,N_3240);
xnor U7986 (N_7986,N_3288,N_2661);
and U7987 (N_7987,N_1347,N_5075);
nand U7988 (N_7988,N_5348,N_5169);
nor U7989 (N_7989,N_5248,N_4471);
and U7990 (N_7990,N_696,N_2586);
nand U7991 (N_7991,N_5701,N_2939);
and U7992 (N_7992,N_5842,N_3165);
or U7993 (N_7993,N_1372,N_629);
nand U7994 (N_7994,N_3485,N_2569);
and U7995 (N_7995,N_4426,N_878);
and U7996 (N_7996,N_5080,N_4061);
nor U7997 (N_7997,N_5822,N_1651);
nand U7998 (N_7998,N_1412,N_4515);
nor U7999 (N_7999,N_1097,N_94);
nor U8000 (N_8000,N_2778,N_2816);
or U8001 (N_8001,N_2494,N_2232);
or U8002 (N_8002,N_3916,N_1222);
or U8003 (N_8003,N_1572,N_2311);
and U8004 (N_8004,N_6038,N_3149);
and U8005 (N_8005,N_2197,N_1801);
nor U8006 (N_8006,N_2320,N_1568);
or U8007 (N_8007,N_3426,N_2864);
nand U8008 (N_8008,N_5702,N_171);
nand U8009 (N_8009,N_3734,N_115);
nor U8010 (N_8010,N_2686,N_5013);
xor U8011 (N_8011,N_3946,N_1219);
or U8012 (N_8012,N_1592,N_3055);
xor U8013 (N_8013,N_4878,N_4981);
and U8014 (N_8014,N_4449,N_1988);
or U8015 (N_8015,N_6018,N_1338);
or U8016 (N_8016,N_4260,N_1945);
nor U8017 (N_8017,N_6043,N_4528);
xor U8018 (N_8018,N_5850,N_5147);
nor U8019 (N_8019,N_4604,N_2458);
and U8020 (N_8020,N_5555,N_1643);
and U8021 (N_8021,N_4708,N_5474);
or U8022 (N_8022,N_3804,N_1671);
and U8023 (N_8023,N_4832,N_2475);
and U8024 (N_8024,N_1532,N_3385);
nand U8025 (N_8025,N_4709,N_4789);
nand U8026 (N_8026,N_1192,N_2454);
or U8027 (N_8027,N_3756,N_4727);
or U8028 (N_8028,N_3823,N_5847);
or U8029 (N_8029,N_5950,N_1396);
or U8030 (N_8030,N_1235,N_2648);
nand U8031 (N_8031,N_5311,N_3068);
nand U8032 (N_8032,N_602,N_1476);
nand U8033 (N_8033,N_512,N_4156);
nor U8034 (N_8034,N_3992,N_3271);
and U8035 (N_8035,N_535,N_5439);
nor U8036 (N_8036,N_3785,N_1276);
nor U8037 (N_8037,N_2504,N_1100);
and U8038 (N_8038,N_4458,N_473);
or U8039 (N_8039,N_4589,N_1159);
nor U8040 (N_8040,N_3687,N_4245);
and U8041 (N_8041,N_3583,N_421);
nand U8042 (N_8042,N_2966,N_2239);
nand U8043 (N_8043,N_2230,N_1283);
or U8044 (N_8044,N_3563,N_5712);
xor U8045 (N_8045,N_2150,N_3859);
nor U8046 (N_8046,N_472,N_3080);
and U8047 (N_8047,N_1770,N_1383);
or U8048 (N_8048,N_1887,N_5029);
and U8049 (N_8049,N_5406,N_593);
nand U8050 (N_8050,N_1638,N_367);
xnor U8051 (N_8051,N_3691,N_2980);
nand U8052 (N_8052,N_3309,N_24);
nand U8053 (N_8053,N_1317,N_4714);
xor U8054 (N_8054,N_734,N_5478);
xnor U8055 (N_8055,N_3585,N_5986);
or U8056 (N_8056,N_257,N_3604);
and U8057 (N_8057,N_5283,N_4068);
nand U8058 (N_8058,N_5421,N_796);
and U8059 (N_8059,N_2081,N_5672);
xnor U8060 (N_8060,N_3808,N_2343);
nand U8061 (N_8061,N_873,N_3883);
nand U8062 (N_8062,N_103,N_269);
and U8063 (N_8063,N_2732,N_4151);
nor U8064 (N_8064,N_1234,N_414);
nand U8065 (N_8065,N_938,N_2201);
or U8066 (N_8066,N_2499,N_434);
or U8067 (N_8067,N_6148,N_1605);
nand U8068 (N_8068,N_3889,N_153);
and U8069 (N_8069,N_4130,N_5212);
or U8070 (N_8070,N_31,N_93);
or U8071 (N_8071,N_1780,N_2467);
or U8072 (N_8072,N_2012,N_2600);
nand U8073 (N_8073,N_777,N_2281);
xor U8074 (N_8074,N_5827,N_3741);
nor U8075 (N_8075,N_4434,N_4846);
nor U8076 (N_8076,N_5479,N_5518);
or U8077 (N_8077,N_6180,N_293);
xor U8078 (N_8078,N_3813,N_3427);
nand U8079 (N_8079,N_4454,N_6231);
nand U8080 (N_8080,N_4052,N_471);
and U8081 (N_8081,N_2677,N_810);
nand U8082 (N_8082,N_2845,N_1277);
or U8083 (N_8083,N_2900,N_5616);
and U8084 (N_8084,N_4926,N_900);
nor U8085 (N_8085,N_4011,N_4938);
xnor U8086 (N_8086,N_944,N_1441);
nor U8087 (N_8087,N_4368,N_5216);
nor U8088 (N_8088,N_3590,N_2219);
or U8089 (N_8089,N_5869,N_6186);
or U8090 (N_8090,N_3704,N_4390);
nand U8091 (N_8091,N_4782,N_4925);
and U8092 (N_8092,N_5680,N_4602);
xor U8093 (N_8093,N_2836,N_3248);
nand U8094 (N_8094,N_2218,N_289);
nand U8095 (N_8095,N_5888,N_4399);
or U8096 (N_8096,N_3447,N_5275);
or U8097 (N_8097,N_3033,N_2704);
nand U8098 (N_8098,N_363,N_1298);
nor U8099 (N_8099,N_4280,N_3513);
or U8100 (N_8100,N_102,N_20);
nor U8101 (N_8101,N_5378,N_594);
or U8102 (N_8102,N_3712,N_3628);
nor U8103 (N_8103,N_3596,N_5366);
nand U8104 (N_8104,N_435,N_1734);
nor U8105 (N_8105,N_3975,N_3896);
and U8106 (N_8106,N_5804,N_2172);
nor U8107 (N_8107,N_1155,N_2878);
and U8108 (N_8108,N_2215,N_2897);
and U8109 (N_8109,N_1792,N_5229);
and U8110 (N_8110,N_6095,N_804);
and U8111 (N_8111,N_5969,N_1259);
xnor U8112 (N_8112,N_5448,N_2216);
and U8113 (N_8113,N_3629,N_1501);
nand U8114 (N_8114,N_3396,N_3553);
or U8115 (N_8115,N_1359,N_3826);
nand U8116 (N_8116,N_2854,N_2585);
nor U8117 (N_8117,N_2840,N_730);
and U8118 (N_8118,N_58,N_5937);
nor U8119 (N_8119,N_2536,N_2114);
nand U8120 (N_8120,N_1092,N_2260);
and U8121 (N_8121,N_3444,N_2108);
nor U8122 (N_8122,N_5541,N_5301);
or U8123 (N_8123,N_4209,N_4295);
or U8124 (N_8124,N_5058,N_3717);
and U8125 (N_8125,N_2877,N_4079);
and U8126 (N_8126,N_4370,N_1021);
or U8127 (N_8127,N_1556,N_3495);
nor U8128 (N_8128,N_2635,N_6244);
and U8129 (N_8129,N_1696,N_2316);
nor U8130 (N_8130,N_1929,N_3707);
nand U8131 (N_8131,N_3278,N_3354);
xnor U8132 (N_8132,N_3831,N_3037);
xnor U8133 (N_8133,N_577,N_3832);
nand U8134 (N_8134,N_1802,N_3581);
or U8135 (N_8135,N_36,N_1373);
and U8136 (N_8136,N_931,N_4100);
or U8137 (N_8137,N_4486,N_70);
and U8138 (N_8138,N_3259,N_474);
or U8139 (N_8139,N_2863,N_2001);
and U8140 (N_8140,N_2142,N_905);
nand U8141 (N_8141,N_329,N_5634);
xnor U8142 (N_8142,N_506,N_6118);
nor U8143 (N_8143,N_3758,N_2452);
nor U8144 (N_8144,N_2982,N_2574);
nand U8145 (N_8145,N_2453,N_3218);
and U8146 (N_8146,N_2287,N_1068);
xnor U8147 (N_8147,N_3016,N_2122);
or U8148 (N_8148,N_5983,N_5414);
nor U8149 (N_8149,N_1786,N_1798);
nor U8150 (N_8150,N_4566,N_821);
nor U8151 (N_8151,N_4683,N_3448);
nor U8152 (N_8152,N_4392,N_118);
nor U8153 (N_8153,N_4972,N_2243);
nor U8154 (N_8154,N_2594,N_864);
xnor U8155 (N_8155,N_6245,N_2992);
and U8156 (N_8156,N_4557,N_4797);
nand U8157 (N_8157,N_2668,N_936);
nand U8158 (N_8158,N_2739,N_5768);
or U8159 (N_8159,N_2265,N_4835);
and U8160 (N_8160,N_4767,N_4285);
nand U8161 (N_8161,N_5678,N_4591);
nand U8162 (N_8162,N_5101,N_5259);
nand U8163 (N_8163,N_6249,N_2028);
nand U8164 (N_8164,N_2691,N_4253);
nand U8165 (N_8165,N_4958,N_4680);
or U8166 (N_8166,N_6106,N_4569);
and U8167 (N_8167,N_5036,N_5178);
nor U8168 (N_8168,N_3579,N_5390);
nor U8169 (N_8169,N_4957,N_5253);
or U8170 (N_8170,N_2,N_154);
and U8171 (N_8171,N_554,N_894);
and U8172 (N_8172,N_4689,N_3305);
or U8173 (N_8173,N_1894,N_5377);
or U8174 (N_8174,N_1749,N_4548);
or U8175 (N_8175,N_4512,N_3107);
nand U8176 (N_8176,N_872,N_6188);
or U8177 (N_8177,N_1461,N_1769);
nor U8178 (N_8178,N_2456,N_3481);
nand U8179 (N_8179,N_2418,N_3042);
nand U8180 (N_8180,N_2731,N_3014);
or U8181 (N_8181,N_4610,N_42);
or U8182 (N_8182,N_4590,N_1369);
and U8183 (N_8183,N_2684,N_3137);
nand U8184 (N_8184,N_1368,N_2064);
nor U8185 (N_8185,N_3192,N_6024);
xnor U8186 (N_8186,N_2890,N_2974);
or U8187 (N_8187,N_1694,N_3797);
or U8188 (N_8188,N_3162,N_1123);
nor U8189 (N_8189,N_5629,N_5130);
nor U8190 (N_8190,N_2844,N_2945);
and U8191 (N_8191,N_205,N_4803);
and U8192 (N_8192,N_2039,N_2751);
nor U8193 (N_8193,N_3966,N_1089);
or U8194 (N_8194,N_4325,N_3959);
nor U8195 (N_8195,N_1521,N_3812);
nor U8196 (N_8196,N_5930,N_1913);
nand U8197 (N_8197,N_126,N_3902);
nor U8198 (N_8198,N_4377,N_2328);
nor U8199 (N_8199,N_2151,N_6165);
nor U8200 (N_8200,N_4780,N_2747);
and U8201 (N_8201,N_4417,N_686);
nand U8202 (N_8202,N_3176,N_5587);
or U8203 (N_8203,N_6002,N_3536);
nand U8204 (N_8204,N_4858,N_1862);
and U8205 (N_8205,N_1850,N_4837);
or U8206 (N_8206,N_1067,N_2355);
or U8207 (N_8207,N_6101,N_3720);
or U8208 (N_8208,N_1176,N_2842);
nor U8209 (N_8209,N_1857,N_4652);
and U8210 (N_8210,N_753,N_396);
and U8211 (N_8211,N_2617,N_351);
nor U8212 (N_8212,N_5601,N_169);
nor U8213 (N_8213,N_6197,N_4074);
and U8214 (N_8214,N_185,N_2299);
nor U8215 (N_8215,N_5904,N_6090);
and U8216 (N_8216,N_5558,N_783);
nand U8217 (N_8217,N_1531,N_2650);
nand U8218 (N_8218,N_4675,N_818);
nand U8219 (N_8219,N_2509,N_5287);
or U8220 (N_8220,N_935,N_4210);
and U8221 (N_8221,N_1060,N_813);
and U8222 (N_8222,N_5451,N_5452);
or U8223 (N_8223,N_3019,N_1497);
nand U8224 (N_8224,N_5719,N_3185);
nor U8225 (N_8225,N_4080,N_2681);
or U8226 (N_8226,N_5471,N_3401);
nand U8227 (N_8227,N_4931,N_1676);
xor U8228 (N_8228,N_2633,N_5650);
and U8229 (N_8229,N_4070,N_4055);
and U8230 (N_8230,N_480,N_5204);
and U8231 (N_8231,N_3425,N_5971);
and U8232 (N_8232,N_4703,N_2342);
or U8233 (N_8233,N_4973,N_401);
nand U8234 (N_8234,N_6019,N_5566);
nor U8235 (N_8235,N_3064,N_1391);
or U8236 (N_8236,N_2131,N_3194);
xor U8237 (N_8237,N_229,N_1778);
or U8238 (N_8238,N_3431,N_942);
nand U8239 (N_8239,N_139,N_199);
nand U8240 (N_8240,N_2561,N_5085);
nand U8241 (N_8241,N_465,N_6193);
xnor U8242 (N_8242,N_4176,N_1993);
or U8243 (N_8243,N_658,N_5861);
xnor U8244 (N_8244,N_1588,N_145);
nand U8245 (N_8245,N_1496,N_2423);
and U8246 (N_8246,N_4757,N_5549);
and U8247 (N_8247,N_915,N_4840);
xor U8248 (N_8248,N_3669,N_1107);
xor U8249 (N_8249,N_5370,N_2558);
nand U8250 (N_8250,N_399,N_5649);
and U8251 (N_8251,N_4029,N_744);
nand U8252 (N_8252,N_2624,N_6160);
nor U8253 (N_8253,N_726,N_3930);
or U8254 (N_8254,N_4628,N_3877);
and U8255 (N_8255,N_2321,N_111);
xnor U8256 (N_8256,N_2220,N_1673);
nand U8257 (N_8257,N_2626,N_5754);
xnor U8258 (N_8258,N_5345,N_184);
nand U8259 (N_8259,N_6226,N_3555);
nand U8260 (N_8260,N_4447,N_1130);
and U8261 (N_8261,N_260,N_2478);
or U8262 (N_8262,N_4178,N_1683);
nand U8263 (N_8263,N_4614,N_47);
and U8264 (N_8264,N_4818,N_3901);
or U8265 (N_8265,N_219,N_5088);
nand U8266 (N_8266,N_2542,N_5416);
nor U8267 (N_8267,N_4000,N_1800);
nor U8268 (N_8268,N_3432,N_1478);
and U8269 (N_8269,N_5807,N_1265);
nor U8270 (N_8270,N_1807,N_392);
or U8271 (N_8271,N_4744,N_33);
xnor U8272 (N_8272,N_2880,N_3558);
or U8273 (N_8273,N_492,N_5079);
nand U8274 (N_8274,N_2671,N_5149);
xnor U8275 (N_8275,N_4404,N_3685);
or U8276 (N_8276,N_4810,N_303);
or U8277 (N_8277,N_1048,N_3827);
and U8278 (N_8278,N_5709,N_5086);
xnor U8279 (N_8279,N_2396,N_5462);
and U8280 (N_8280,N_2023,N_5595);
and U8281 (N_8281,N_741,N_2291);
or U8282 (N_8282,N_2250,N_3153);
nand U8283 (N_8283,N_2077,N_3751);
and U8284 (N_8284,N_1491,N_3342);
nand U8285 (N_8285,N_2538,N_3599);
nor U8286 (N_8286,N_3098,N_3349);
xor U8287 (N_8287,N_3251,N_1299);
nand U8288 (N_8288,N_1752,N_3641);
and U8289 (N_8289,N_403,N_3410);
nor U8290 (N_8290,N_913,N_5153);
nand U8291 (N_8291,N_3670,N_2276);
nand U8292 (N_8292,N_5882,N_1750);
or U8293 (N_8293,N_5508,N_1324);
xnor U8294 (N_8294,N_5438,N_2607);
nor U8295 (N_8295,N_4366,N_4353);
nor U8296 (N_8296,N_5039,N_762);
or U8297 (N_8297,N_886,N_3077);
or U8298 (N_8298,N_1327,N_4671);
or U8299 (N_8299,N_1254,N_2238);
and U8300 (N_8300,N_5306,N_3111);
nand U8301 (N_8301,N_1247,N_3519);
nand U8302 (N_8302,N_3433,N_5667);
nand U8303 (N_8303,N_4678,N_1462);
xor U8304 (N_8304,N_462,N_4456);
nor U8305 (N_8305,N_4574,N_2936);
nor U8306 (N_8306,N_1528,N_2724);
nand U8307 (N_8307,N_2067,N_1502);
or U8308 (N_8308,N_616,N_4030);
nor U8309 (N_8309,N_1567,N_4697);
xnor U8310 (N_8310,N_1687,N_1005);
xnor U8311 (N_8311,N_66,N_4809);
or U8312 (N_8312,N_5909,N_318);
nor U8313 (N_8313,N_4301,N_1640);
xor U8314 (N_8314,N_2971,N_6086);
nand U8315 (N_8315,N_2268,N_5078);
nor U8316 (N_8316,N_483,N_1477);
nor U8317 (N_8317,N_3523,N_966);
and U8318 (N_8318,N_822,N_5412);
or U8319 (N_8319,N_3285,N_5124);
and U8320 (N_8320,N_3195,N_4444);
nand U8321 (N_8321,N_1755,N_1458);
xnor U8322 (N_8322,N_170,N_5853);
nand U8323 (N_8323,N_2593,N_4466);
nor U8324 (N_8324,N_4699,N_1124);
and U8325 (N_8325,N_2876,N_3905);
xnor U8326 (N_8326,N_3171,N_4959);
or U8327 (N_8327,N_235,N_5589);
nor U8328 (N_8328,N_1203,N_4963);
and U8329 (N_8329,N_1345,N_1193);
or U8330 (N_8330,N_6057,N_1036);
nand U8331 (N_8331,N_4826,N_3631);
and U8332 (N_8332,N_2435,N_296);
or U8333 (N_8333,N_2669,N_543);
and U8334 (N_8334,N_1416,N_2907);
nor U8335 (N_8335,N_509,N_1897);
nand U8336 (N_8336,N_1308,N_3161);
and U8337 (N_8337,N_1353,N_3043);
and U8338 (N_8338,N_3249,N_2823);
nor U8339 (N_8339,N_3244,N_5849);
nand U8340 (N_8340,N_3463,N_4968);
and U8341 (N_8341,N_1934,N_5371);
or U8342 (N_8342,N_5316,N_711);
xor U8343 (N_8343,N_382,N_5331);
xor U8344 (N_8344,N_5207,N_5102);
nor U8345 (N_8345,N_3083,N_272);
and U8346 (N_8346,N_3406,N_6061);
nand U8347 (N_8347,N_4587,N_248);
nor U8348 (N_8348,N_2065,N_4034);
or U8349 (N_8349,N_3299,N_3492);
xor U8350 (N_8350,N_1498,N_5833);
and U8351 (N_8351,N_5788,N_4175);
and U8352 (N_8352,N_5565,N_2507);
xnor U8353 (N_8353,N_3775,N_3663);
nor U8354 (N_8354,N_2757,N_998);
or U8355 (N_8355,N_5605,N_1095);
nand U8356 (N_8356,N_2327,N_799);
and U8357 (N_8357,N_5191,N_4982);
and U8358 (N_8358,N_793,N_2473);
and U8359 (N_8359,N_3119,N_4684);
and U8360 (N_8360,N_3892,N_5336);
xnor U8361 (N_8361,N_5664,N_2583);
and U8362 (N_8362,N_3155,N_848);
nand U8363 (N_8363,N_2294,N_5868);
and U8364 (N_8364,N_2592,N_4373);
nand U8365 (N_8365,N_1320,N_2810);
or U8366 (N_8366,N_4240,N_611);
xor U8367 (N_8367,N_4021,N_1701);
nor U8368 (N_8368,N_2631,N_163);
xor U8369 (N_8369,N_384,N_3280);
or U8370 (N_8370,N_1724,N_1352);
xor U8371 (N_8371,N_5349,N_3435);
nand U8372 (N_8372,N_372,N_4457);
and U8373 (N_8373,N_2578,N_1771);
or U8374 (N_8374,N_3993,N_4888);
or U8375 (N_8375,N_3074,N_778);
nor U8376 (N_8376,N_5250,N_5043);
or U8377 (N_8377,N_4974,N_1858);
nand U8378 (N_8378,N_4027,N_4996);
nand U8379 (N_8379,N_5576,N_3169);
xor U8380 (N_8380,N_456,N_1296);
and U8381 (N_8381,N_2177,N_2657);
and U8382 (N_8382,N_2941,N_2726);
or U8383 (N_8383,N_1313,N_2339);
xor U8384 (N_8384,N_6097,N_88);
or U8385 (N_8385,N_1995,N_5721);
and U8386 (N_8386,N_3110,N_3489);
xor U8387 (N_8387,N_5803,N_2754);
nor U8388 (N_8388,N_2708,N_5369);
nor U8389 (N_8389,N_4143,N_97);
nor U8390 (N_8390,N_1831,N_5522);
nor U8391 (N_8391,N_4552,N_1879);
nand U8392 (N_8392,N_515,N_468);
and U8393 (N_8393,N_967,N_6059);
and U8394 (N_8394,N_4792,N_6088);
nor U8395 (N_8395,N_893,N_588);
or U8396 (N_8396,N_2059,N_514);
nor U8397 (N_8397,N_5163,N_5860);
nand U8398 (N_8398,N_3847,N_1220);
nor U8399 (N_8399,N_4966,N_2766);
nand U8400 (N_8400,N_4912,N_4112);
and U8401 (N_8401,N_221,N_1224);
nand U8402 (N_8402,N_2266,N_3284);
nor U8403 (N_8403,N_2229,N_5243);
and U8404 (N_8404,N_559,N_3156);
nand U8405 (N_8405,N_2091,N_2705);
nor U8406 (N_8406,N_4764,N_4129);
and U8407 (N_8407,N_2806,N_4728);
and U8408 (N_8408,N_4943,N_1297);
and U8409 (N_8409,N_1074,N_6203);
or U8410 (N_8410,N_2891,N_2147);
and U8411 (N_8411,N_4388,N_1735);
xnor U8412 (N_8412,N_2015,N_2306);
and U8413 (N_8413,N_5000,N_6139);
and U8414 (N_8414,N_1101,N_1205);
or U8415 (N_8415,N_2202,N_5551);
or U8416 (N_8416,N_3680,N_5848);
or U8417 (N_8417,N_571,N_4768);
nor U8418 (N_8418,N_4545,N_1002);
and U8419 (N_8419,N_985,N_3146);
xnor U8420 (N_8420,N_1310,N_8);
nor U8421 (N_8421,N_1404,N_2134);
or U8422 (N_8422,N_1280,N_3163);
nand U8423 (N_8423,N_3170,N_3633);
or U8424 (N_8424,N_4423,N_1963);
nor U8425 (N_8425,N_6026,N_1057);
nand U8426 (N_8426,N_1442,N_265);
xnor U8427 (N_8427,N_3145,N_5159);
xor U8428 (N_8428,N_875,N_190);
nor U8429 (N_8429,N_4491,N_2408);
nand U8430 (N_8430,N_1208,N_1459);
or U8431 (N_8431,N_3843,N_5580);
nor U8432 (N_8432,N_4300,N_3439);
nor U8433 (N_8433,N_3673,N_1991);
and U8434 (N_8434,N_1087,N_4597);
or U8435 (N_8435,N_2420,N_1946);
and U8436 (N_8436,N_3141,N_4104);
or U8437 (N_8437,N_298,N_5689);
and U8438 (N_8438,N_3012,N_279);
or U8439 (N_8439,N_3094,N_4481);
xor U8440 (N_8440,N_4081,N_4860);
nor U8441 (N_8441,N_2007,N_445);
nor U8442 (N_8442,N_3567,N_5170);
and U8443 (N_8443,N_523,N_4355);
or U8444 (N_8444,N_3891,N_1402);
xor U8445 (N_8445,N_4866,N_1288);
nor U8446 (N_8446,N_2017,N_2735);
and U8447 (N_8447,N_5994,N_4724);
or U8448 (N_8448,N_3848,N_5992);
and U8449 (N_8449,N_1294,N_3070);
nand U8450 (N_8450,N_1488,N_2462);
xnor U8451 (N_8451,N_4191,N_4990);
or U8452 (N_8452,N_4791,N_774);
nand U8453 (N_8453,N_5218,N_4998);
nand U8454 (N_8454,N_5581,N_3530);
nor U8455 (N_8455,N_3806,N_173);
nor U8456 (N_8456,N_3807,N_3890);
xor U8457 (N_8457,N_1685,N_2855);
nor U8458 (N_8458,N_3351,N_969);
nor U8459 (N_8459,N_5179,N_853);
or U8460 (N_8460,N_637,N_5138);
nand U8461 (N_8461,N_5687,N_1115);
or U8462 (N_8462,N_4830,N_6158);
or U8463 (N_8463,N_1997,N_150);
nor U8464 (N_8464,N_5700,N_3387);
nor U8465 (N_8465,N_3750,N_1070);
xor U8466 (N_8466,N_3479,N_5862);
or U8467 (N_8467,N_5150,N_4861);
nor U8468 (N_8468,N_5663,N_5172);
nand U8469 (N_8469,N_1468,N_46);
nand U8470 (N_8470,N_4134,N_5972);
or U8471 (N_8471,N_4267,N_6211);
nor U8472 (N_8472,N_4815,N_2424);
nor U8473 (N_8473,N_2714,N_1905);
nor U8474 (N_8474,N_2603,N_1494);
nor U8475 (N_8475,N_531,N_4227);
nand U8476 (N_8476,N_2164,N_572);
and U8477 (N_8477,N_4677,N_3371);
xnor U8478 (N_8478,N_1666,N_701);
nor U8479 (N_8479,N_5044,N_5183);
nor U8480 (N_8480,N_4172,N_494);
or U8481 (N_8481,N_5666,N_1287);
and U8482 (N_8482,N_2851,N_6079);
nor U8483 (N_8483,N_1148,N_1513);
nor U8484 (N_8484,N_2016,N_544);
and U8485 (N_8485,N_3693,N_141);
xnor U8486 (N_8486,N_604,N_4676);
nor U8487 (N_8487,N_671,N_3634);
nand U8488 (N_8488,N_5635,N_2522);
nand U8489 (N_8489,N_5192,N_1336);
nor U8490 (N_8490,N_408,N_5698);
nor U8491 (N_8491,N_2010,N_2579);
or U8492 (N_8492,N_3598,N_307);
nand U8493 (N_8493,N_4485,N_2822);
or U8494 (N_8494,N_5276,N_2159);
nand U8495 (N_8495,N_882,N_2116);
or U8496 (N_8496,N_1990,N_3233);
nand U8497 (N_8497,N_3322,N_5707);
or U8498 (N_8498,N_700,N_561);
and U8499 (N_8499,N_5018,N_1250);
or U8500 (N_8500,N_4255,N_5445);
and U8501 (N_8501,N_963,N_1330);
nand U8502 (N_8502,N_2135,N_461);
nor U8503 (N_8503,N_2271,N_3809);
nor U8504 (N_8504,N_6177,N_2228);
nand U8505 (N_8505,N_2697,N_2756);
nor U8506 (N_8506,N_4905,N_4567);
nor U8507 (N_8507,N_3742,N_3851);
nand U8508 (N_8508,N_5362,N_1987);
and U8509 (N_8509,N_4446,N_1877);
and U8510 (N_8510,N_1580,N_11);
nor U8511 (N_8511,N_5836,N_1601);
and U8512 (N_8512,N_4867,N_1747);
or U8513 (N_8513,N_4058,N_924);
nor U8514 (N_8514,N_5903,N_3358);
nor U8515 (N_8515,N_1463,N_2944);
or U8516 (N_8516,N_6196,N_1751);
nand U8517 (N_8517,N_641,N_193);
nor U8518 (N_8518,N_670,N_2652);
nand U8519 (N_8519,N_4138,N_5611);
xnor U8520 (N_8520,N_3496,N_4670);
and U8521 (N_8521,N_586,N_1705);
nor U8522 (N_8522,N_1263,N_1367);
or U8523 (N_8523,N_1239,N_1915);
xnor U8524 (N_8524,N_1972,N_5015);
nor U8525 (N_8525,N_4646,N_1113);
or U8526 (N_8526,N_4863,N_2412);
nand U8527 (N_8527,N_203,N_3126);
nor U8528 (N_8528,N_3803,N_344);
or U8529 (N_8529,N_2432,N_4759);
nand U8530 (N_8530,N_4519,N_4601);
and U8531 (N_8531,N_1508,N_4885);
or U8532 (N_8532,N_4062,N_2835);
or U8533 (N_8533,N_4896,N_4170);
nand U8534 (N_8534,N_1266,N_2666);
and U8535 (N_8535,N_1360,N_4182);
nor U8536 (N_8536,N_3391,N_3211);
and U8537 (N_8537,N_1366,N_1911);
or U8538 (N_8538,N_5636,N_6150);
nor U8539 (N_8539,N_912,N_5501);
nor U8540 (N_8540,N_2825,N_4607);
nand U8541 (N_8541,N_5072,N_615);
nor U8542 (N_8542,N_1306,N_3419);
nand U8543 (N_8543,N_626,N_2236);
nand U8544 (N_8544,N_3790,N_335);
xor U8545 (N_8545,N_698,N_4101);
xnor U8546 (N_8546,N_1243,N_3018);
nand U8547 (N_8547,N_5490,N_4720);
nor U8548 (N_8548,N_143,N_855);
or U8549 (N_8549,N_176,N_1424);
nand U8550 (N_8550,N_1950,N_5991);
nor U8551 (N_8551,N_4605,N_230);
or U8552 (N_8552,N_1394,N_2278);
nand U8553 (N_8553,N_1795,N_4950);
nor U8554 (N_8554,N_1781,N_3575);
and U8555 (N_8555,N_1825,N_929);
or U8556 (N_8556,N_3866,N_1050);
nor U8557 (N_8557,N_3970,N_1047);
xor U8558 (N_8558,N_4252,N_2069);
xor U8559 (N_8559,N_5999,N_68);
and U8560 (N_8560,N_6214,N_5625);
or U8561 (N_8561,N_2670,N_2524);
or U8562 (N_8562,N_4702,N_2573);
nand U8563 (N_8563,N_5189,N_584);
or U8564 (N_8564,N_2562,N_5982);
or U8565 (N_8565,N_3646,N_2801);
or U8566 (N_8566,N_898,N_5281);
nand U8567 (N_8567,N_725,N_5193);
xnor U8568 (N_8568,N_4415,N_1662);
or U8569 (N_8569,N_2160,N_4977);
or U8570 (N_8570,N_2768,N_2303);
and U8571 (N_8571,N_5747,N_5977);
or U8572 (N_8572,N_2137,N_2546);
nor U8573 (N_8573,N_1010,N_751);
nand U8574 (N_8574,N_759,N_1548);
and U8575 (N_8575,N_4784,N_4583);
nor U8576 (N_8576,N_6119,N_5944);
nand U8577 (N_8577,N_6153,N_6200);
and U8578 (N_8578,N_1150,N_2362);
xor U8579 (N_8579,N_3241,N_371);
and U8580 (N_8580,N_5932,N_2910);
or U8581 (N_8581,N_2892,N_5716);
or U8582 (N_8582,N_2967,N_3181);
and U8583 (N_8583,N_5608,N_3009);
nand U8584 (N_8584,N_5864,N_2994);
or U8585 (N_8585,N_2335,N_5544);
xor U8586 (N_8586,N_548,N_3129);
nor U8587 (N_8587,N_1630,N_4116);
or U8588 (N_8588,N_2729,N_3531);
or U8589 (N_8589,N_3430,N_780);
nand U8590 (N_8590,N_1375,N_3611);
and U8591 (N_8591,N_4551,N_3665);
nor U8592 (N_8592,N_4031,N_4735);
nand U8593 (N_8593,N_295,N_2505);
and U8594 (N_8594,N_1038,N_247);
nor U8595 (N_8595,N_5730,N_4004);
nor U8596 (N_8596,N_5433,N_4903);
or U8597 (N_8597,N_3653,N_1526);
or U8598 (N_8598,N_682,N_1290);
or U8599 (N_8599,N_5927,N_2259);
and U8600 (N_8600,N_3594,N_5820);
xnor U8601 (N_8601,N_1541,N_6074);
nand U8602 (N_8602,N_583,N_4707);
nor U8603 (N_8603,N_195,N_432);
and U8604 (N_8604,N_2712,N_6159);
nor U8605 (N_8605,N_3478,N_2468);
nand U8606 (N_8606,N_649,N_697);
nand U8607 (N_8607,N_4010,N_871);
or U8608 (N_8608,N_1736,N_1072);
nor U8609 (N_8609,N_1331,N_3705);
nand U8610 (N_8610,N_550,N_62);
nand U8611 (N_8611,N_4250,N_4596);
nand U8612 (N_8612,N_4902,N_2246);
nor U8613 (N_8613,N_4220,N_4196);
or U8614 (N_8614,N_5326,N_3025);
and U8615 (N_8615,N_5004,N_3911);
or U8616 (N_8616,N_4928,N_370);
nor U8617 (N_8617,N_4334,N_4448);
nand U8618 (N_8618,N_4261,N_2374);
or U8619 (N_8619,N_148,N_573);
xor U8620 (N_8620,N_5182,N_3090);
nand U8621 (N_8621,N_3560,N_3250);
nor U8622 (N_8622,N_1091,N_2549);
and U8623 (N_8623,N_1231,N_4831);
nor U8624 (N_8624,N_4137,N_181);
or U8625 (N_8625,N_2045,N_909);
nand U8626 (N_8626,N_3777,N_466);
nand U8627 (N_8627,N_5184,N_2225);
xor U8628 (N_8628,N_940,N_692);
or U8629 (N_8629,N_4421,N_4698);
nor U8630 (N_8630,N_1016,N_1275);
nand U8631 (N_8631,N_6233,N_1591);
nor U8632 (N_8632,N_6004,N_5117);
nor U8633 (N_8633,N_754,N_415);
xnor U8634 (N_8634,N_4091,N_880);
xnor U8635 (N_8635,N_2802,N_815);
or U8636 (N_8636,N_4525,N_952);
nand U8637 (N_8637,N_419,N_4753);
or U8638 (N_8638,N_993,N_135);
nor U8639 (N_8639,N_5597,N_2249);
or U8640 (N_8640,N_807,N_6064);
and U8641 (N_8641,N_4026,N_3887);
and U8642 (N_8642,N_2205,N_5032);
and U8643 (N_8643,N_3375,N_5832);
and U8644 (N_8644,N_1397,N_1018);
or U8645 (N_8645,N_5211,N_4314);
nor U8646 (N_8646,N_1408,N_1840);
or U8647 (N_8647,N_6120,N_256);
xnor U8648 (N_8648,N_1918,N_4225);
and U8649 (N_8649,N_4632,N_1295);
or U8650 (N_8650,N_2354,N_4039);
and U8651 (N_8651,N_4445,N_1819);
and U8652 (N_8652,N_2425,N_4344);
nand U8653 (N_8653,N_151,N_5704);
or U8654 (N_8654,N_5455,N_4315);
and U8655 (N_8655,N_3766,N_2187);
or U8656 (N_8656,N_104,N_5269);
or U8657 (N_8657,N_1517,N_1794);
nand U8658 (N_8658,N_1930,N_5726);
and U8659 (N_8659,N_722,N_850);
xor U8660 (N_8660,N_3729,N_977);
or U8661 (N_8661,N_4553,N_3421);
nand U8662 (N_8662,N_1577,N_4228);
nor U8663 (N_8663,N_2099,N_1978);
nor U8664 (N_8664,N_484,N_5821);
and U8665 (N_8665,N_1832,N_1523);
and U8666 (N_8666,N_3497,N_1719);
and U8667 (N_8667,N_792,N_3367);
or U8668 (N_8668,N_3394,N_3710);
and U8669 (N_8669,N_2272,N_2978);
nor U8670 (N_8670,N_2368,N_5381);
or U8671 (N_8671,N_5644,N_252);
or U8672 (N_8672,N_2849,N_2047);
nor U8673 (N_8673,N_268,N_3517);
or U8674 (N_8674,N_2783,N_137);
nor U8675 (N_8675,N_5195,N_3336);
nand U8676 (N_8676,N_4173,N_3937);
and U8677 (N_8677,N_1535,N_2237);
and U8678 (N_8678,N_4231,N_3461);
and U8679 (N_8679,N_1682,N_3645);
nand U8680 (N_8680,N_5727,N_1172);
nor U8681 (N_8681,N_1602,N_612);
xor U8682 (N_8682,N_2829,N_3263);
nand U8683 (N_8683,N_4954,N_6122);
nor U8684 (N_8684,N_4146,N_3318);
and U8685 (N_8685,N_109,N_1098);
nand U8686 (N_8686,N_932,N_1869);
and U8687 (N_8687,N_2125,N_3403);
or U8688 (N_8688,N_3528,N_950);
nand U8689 (N_8689,N_1816,N_2476);
nand U8690 (N_8690,N_4655,N_6154);
and U8691 (N_8691,N_2539,N_3081);
nand U8692 (N_8692,N_5282,N_2885);
nor U8693 (N_8693,N_620,N_1960);
or U8694 (N_8694,N_947,N_3943);
or U8695 (N_8695,N_5444,N_876);
and U8696 (N_8696,N_646,N_1081);
nor U8697 (N_8697,N_1848,N_3011);
and U8698 (N_8698,N_3254,N_451);
nand U8699 (N_8699,N_5515,N_5143);
nand U8700 (N_8700,N_3659,N_4321);
nand U8701 (N_8701,N_3722,N_4585);
nor U8702 (N_8702,N_4893,N_3438);
or U8703 (N_8703,N_1906,N_366);
nor U8704 (N_8704,N_2589,N_1885);
nand U8705 (N_8705,N_3470,N_5898);
or U8706 (N_8706,N_2394,N_5647);
or U8707 (N_8707,N_2715,N_718);
or U8708 (N_8708,N_3506,N_4269);
nor U8709 (N_8709,N_699,N_4386);
nand U8710 (N_8710,N_2170,N_3086);
nor U8711 (N_8711,N_6069,N_5785);
nor U8712 (N_8712,N_6247,N_4433);
xnor U8713 (N_8713,N_1207,N_2204);
nor U8714 (N_8714,N_911,N_5956);
or U8715 (N_8715,N_5318,N_5257);
nor U8716 (N_8716,N_3786,N_5290);
xor U8717 (N_8717,N_2743,N_2297);
or U8718 (N_8718,N_4262,N_3621);
nand U8719 (N_8719,N_2413,N_5683);
nor U8720 (N_8720,N_2223,N_3035);
and U8721 (N_8721,N_4037,N_4117);
and U8722 (N_8722,N_4148,N_5923);
or U8723 (N_8723,N_50,N_5814);
nor U8724 (N_8724,N_90,N_3514);
and U8725 (N_8725,N_732,N_1334);
nand U8726 (N_8726,N_3082,N_6225);
or U8727 (N_8727,N_1485,N_1384);
or U8728 (N_8728,N_3013,N_1739);
nand U8729 (N_8729,N_4864,N_3201);
and U8730 (N_8730,N_5738,N_3918);
nor U8731 (N_8731,N_1117,N_2692);
or U8732 (N_8732,N_224,N_1788);
nor U8733 (N_8733,N_4224,N_842);
xnor U8734 (N_8734,N_1700,N_5800);
xor U8735 (N_8735,N_1901,N_2930);
nand U8736 (N_8736,N_1796,N_5291);
nand U8737 (N_8737,N_5643,N_2245);
nand U8738 (N_8738,N_4122,N_5513);
nor U8739 (N_8739,N_3108,N_6243);
nor U8740 (N_8740,N_482,N_3420);
nor U8741 (N_8741,N_903,N_3876);
nor U8742 (N_8742,N_2013,N_4947);
nor U8743 (N_8743,N_373,N_5162);
nor U8744 (N_8744,N_1814,N_526);
nand U8745 (N_8745,N_2072,N_4847);
and U8746 (N_8746,N_2022,N_4636);
nand U8747 (N_8747,N_5778,N_6194);
or U8748 (N_8748,N_5535,N_5201);
nor U8749 (N_8749,N_194,N_6047);
nand U8750 (N_8750,N_2620,N_3328);
nor U8751 (N_8751,N_5368,N_388);
nand U8752 (N_8752,N_779,N_2392);
xor U8753 (N_8753,N_674,N_4828);
xnor U8754 (N_8754,N_4872,N_4687);
or U8755 (N_8755,N_4427,N_2615);
or U8756 (N_8756,N_3320,N_4213);
nand U8757 (N_8757,N_1573,N_1538);
and U8758 (N_8758,N_3625,N_2643);
nor U8759 (N_8759,N_123,N_619);
nand U8760 (N_8760,N_240,N_1695);
nor U8761 (N_8761,N_4734,N_1460);
or U8762 (N_8762,N_3356,N_3480);
and U8763 (N_8763,N_1471,N_5981);
and U8764 (N_8764,N_2292,N_2048);
xnor U8765 (N_8765,N_2319,N_2358);
or U8766 (N_8766,N_30,N_1096);
nand U8767 (N_8767,N_3960,N_4161);
nand U8768 (N_8768,N_1876,N_1448);
nand U8769 (N_8769,N_1128,N_1500);
nor U8770 (N_8770,N_5609,N_4335);
nand U8771 (N_8771,N_1425,N_5094);
nor U8772 (N_8772,N_1529,N_4779);
and U8773 (N_8773,N_5733,N_1169);
nand U8774 (N_8774,N_1027,N_3413);
or U8775 (N_8775,N_5995,N_4869);
or U8776 (N_8776,N_5141,N_3041);
or U8777 (N_8777,N_4933,N_1787);
nand U8778 (N_8778,N_91,N_2580);
nand U8779 (N_8779,N_3255,N_4561);
and U8780 (N_8780,N_2043,N_4441);
nor U8781 (N_8781,N_887,N_3212);
xnor U8782 (N_8782,N_6230,N_2773);
or U8783 (N_8783,N_2267,N_2998);
or U8784 (N_8784,N_4875,N_444);
xnor U8785 (N_8785,N_4391,N_5739);
and U8786 (N_8786,N_3647,N_1655);
nor U8787 (N_8787,N_4098,N_3618);
and U8788 (N_8788,N_4934,N_4072);
and U8789 (N_8789,N_3698,N_5321);
nand U8790 (N_8790,N_3028,N_1587);
nor U8791 (N_8791,N_5330,N_5514);
nand U8792 (N_8792,N_1504,N_1793);
nand U8793 (N_8793,N_2571,N_3059);
nor U8794 (N_8794,N_5003,N_3400);
or U8795 (N_8795,N_3839,N_6138);
or U8796 (N_8796,N_6072,N_1281);
and U8797 (N_8797,N_5604,N_1401);
and U8798 (N_8798,N_3854,N_1598);
or U8799 (N_8799,N_284,N_1058);
nand U8800 (N_8800,N_4418,N_34);
nand U8801 (N_8801,N_4630,N_5461);
nand U8802 (N_8802,N_2977,N_3246);
nand U8803 (N_8803,N_476,N_763);
xnor U8804 (N_8804,N_4806,N_5395);
nand U8805 (N_8805,N_5815,N_3209);
xor U8806 (N_8806,N_3542,N_3205);
nor U8807 (N_8807,N_4455,N_667);
nand U8808 (N_8808,N_5177,N_5407);
or U8809 (N_8809,N_791,N_3569);
nand U8810 (N_8810,N_5483,N_1475);
nor U8811 (N_8811,N_5632,N_3924);
and U8812 (N_8812,N_319,N_2601);
or U8813 (N_8813,N_1350,N_2755);
nor U8814 (N_8814,N_3897,N_5749);
nand U8815 (N_8815,N_5426,N_3895);
nor U8816 (N_8816,N_990,N_1034);
and U8817 (N_8817,N_1303,N_1962);
and U8818 (N_8818,N_3543,N_1304);
nand U8819 (N_8819,N_2235,N_4363);
and U8820 (N_8820,N_5577,N_3861);
and U8821 (N_8821,N_241,N_3096);
nand U8822 (N_8822,N_2144,N_1351);
and U8823 (N_8823,N_3840,N_5767);
and U8824 (N_8824,N_1754,N_4873);
nand U8825 (N_8825,N_4534,N_5023);
nand U8826 (N_8826,N_6208,N_215);
nand U8827 (N_8827,N_2440,N_3765);
nor U8828 (N_8828,N_242,N_570);
nor U8829 (N_8829,N_4932,N_5300);
xor U8830 (N_8830,N_5699,N_5203);
or U8831 (N_8831,N_1314,N_1759);
or U8832 (N_8832,N_3469,N_5521);
nor U8833 (N_8833,N_5713,N_6201);
and U8834 (N_8834,N_3853,N_2528);
nand U8835 (N_8835,N_2309,N_3551);
nand U8836 (N_8836,N_3376,N_6151);
nor U8837 (N_8837,N_182,N_1889);
nand U8838 (N_8838,N_1525,N_2938);
nor U8839 (N_8839,N_1805,N_3539);
nand U8840 (N_8840,N_2859,N_166);
and U8841 (N_8841,N_424,N_3591);
or U8842 (N_8842,N_3178,N_5464);
nor U8843 (N_8843,N_144,N_2537);
and U8844 (N_8844,N_4634,N_32);
or U8845 (N_8845,N_5261,N_3986);
nor U8846 (N_8846,N_5645,N_5675);
nand U8847 (N_8847,N_21,N_3405);
or U8848 (N_8848,N_3971,N_3350);
and U8849 (N_8849,N_823,N_2167);
or U8850 (N_8850,N_5235,N_3697);
xor U8851 (N_8851,N_6,N_5816);
and U8852 (N_8852,N_5022,N_3071);
or U8853 (N_8853,N_3582,N_3791);
and U8854 (N_8854,N_4135,N_3928);
and U8855 (N_8855,N_1942,N_5219);
or U8856 (N_8856,N_996,N_3718);
and U8857 (N_8857,N_283,N_136);
xor U8858 (N_8858,N_2082,N_3835);
nor U8859 (N_8859,N_4322,N_216);
or U8860 (N_8860,N_5806,N_752);
or U8861 (N_8861,N_3921,N_5915);
xnor U8862 (N_8862,N_2382,N_3696);
nand U8863 (N_8863,N_433,N_1139);
nand U8864 (N_8864,N_3989,N_3166);
and U8865 (N_8865,N_1890,N_1082);
or U8866 (N_8866,N_3914,N_5137);
nor U8867 (N_8867,N_5509,N_287);
nand U8868 (N_8868,N_2728,N_5934);
nor U8869 (N_8869,N_551,N_3784);
or U8870 (N_8870,N_1519,N_4980);
and U8871 (N_8871,N_3160,N_1965);
nor U8872 (N_8872,N_326,N_4504);
xor U8873 (N_8873,N_5014,N_5249);
nand U8874 (N_8874,N_4410,N_2057);
nor U8875 (N_8875,N_3652,N_485);
and U8876 (N_8876,N_5867,N_5429);
nor U8877 (N_8877,N_2304,N_4991);
xnor U8878 (N_8878,N_1552,N_4774);
and U8879 (N_8879,N_440,N_2068);
xnor U8880 (N_8880,N_4440,N_5237);
or U8881 (N_8881,N_2678,N_4814);
or U8882 (N_8882,N_2975,N_3099);
and U8883 (N_8883,N_4543,N_4105);
and U8884 (N_8884,N_4710,N_1417);
and U8885 (N_8885,N_4824,N_2146);
nand U8886 (N_8886,N_1715,N_3393);
nor U8887 (N_8887,N_2839,N_2868);
nor U8888 (N_8888,N_5893,N_5746);
nand U8889 (N_8889,N_4965,N_4099);
and U8890 (N_8890,N_1717,N_2875);
and U8891 (N_8891,N_5818,N_716);
nand U8892 (N_8892,N_647,N_757);
or U8893 (N_8893,N_4247,N_1741);
nor U8894 (N_8894,N_6105,N_4107);
nand U8895 (N_8895,N_5772,N_5613);
xnor U8896 (N_8896,N_1054,N_1633);
nand U8897 (N_8897,N_4804,N_310);
nor U8898 (N_8898,N_2188,N_2331);
or U8899 (N_8899,N_3719,N_9);
xor U8900 (N_8900,N_3958,N_4763);
nand U8901 (N_8901,N_1920,N_1223);
or U8902 (N_8902,N_138,N_1340);
and U8903 (N_8903,N_1693,N_578);
and U8904 (N_8904,N_4205,N_249);
or U8905 (N_8905,N_919,N_735);
xnor U8906 (N_8906,N_2369,N_2034);
and U8907 (N_8907,N_1126,N_5890);
nor U8908 (N_8908,N_5121,N_1527);
nand U8909 (N_8909,N_5536,N_1046);
nand U8910 (N_8910,N_1110,N_4109);
nand U8911 (N_8911,N_405,N_5402);
nand U8912 (N_8912,N_1921,N_5895);
nor U8913 (N_8913,N_4775,N_1228);
or U8914 (N_8914,N_16,N_4119);
nand U8915 (N_8915,N_1154,N_61);
nand U8916 (N_8916,N_6028,N_812);
nand U8917 (N_8917,N_2469,N_1109);
xor U8918 (N_8918,N_1670,N_2295);
nor U8919 (N_8919,N_4311,N_1319);
xnor U8920 (N_8920,N_3811,N_6051);
nor U8921 (N_8921,N_6130,N_1919);
nor U8922 (N_8922,N_6144,N_2411);
or U8923 (N_8923,N_2097,N_4063);
or U8924 (N_8924,N_328,N_119);
or U8925 (N_8925,N_4383,N_1482);
and U8926 (N_8926,N_2653,N_3436);
nor U8927 (N_8927,N_1866,N_4022);
xor U8928 (N_8928,N_3475,N_5823);
or U8929 (N_8929,N_5335,N_4165);
nor U8930 (N_8930,N_2740,N_2025);
or U8931 (N_8931,N_5620,N_1212);
and U8932 (N_8932,N_4171,N_2654);
nand U8933 (N_8933,N_6009,N_3997);
nor U8934 (N_8934,N_3672,N_2515);
and U8935 (N_8935,N_634,N_5357);
and U8936 (N_8936,N_566,N_601);
nand U8937 (N_8937,N_5568,N_6164);
nor U8938 (N_8938,N_2191,N_2818);
or U8939 (N_8939,N_2956,N_3671);
or U8940 (N_8940,N_1289,N_5119);
or U8941 (N_8941,N_14,N_4823);
and U8942 (N_8942,N_82,N_2934);
nand U8943 (N_8943,N_237,N_2415);
and U8944 (N_8944,N_881,N_1900);
or U8945 (N_8945,N_4428,N_327);
xnor U8946 (N_8946,N_2861,N_5459);
and U8947 (N_8947,N_3620,N_2914);
nor U8948 (N_8948,N_4424,N_5812);
nand U8949 (N_8949,N_5504,N_5974);
nand U8950 (N_8950,N_2770,N_5361);
nor U8951 (N_8951,N_180,N_3699);
nand U8952 (N_8952,N_3865,N_1309);
xor U8953 (N_8953,N_669,N_690);
or U8954 (N_8954,N_44,N_2360);
nor U8955 (N_8955,N_5724,N_1147);
xnor U8956 (N_8956,N_3939,N_2940);
or U8957 (N_8957,N_4093,N_923);
nand U8958 (N_8958,N_2905,N_1406);
nor U8959 (N_8959,N_4517,N_2535);
nand U8960 (N_8960,N_1029,N_3366);
and U8961 (N_8961,N_557,N_460);
nor U8962 (N_8962,N_656,N_92);
or U8963 (N_8963,N_1037,N_6011);
and U8964 (N_8964,N_2623,N_45);
nand U8965 (N_8965,N_5953,N_862);
xor U8966 (N_8966,N_4579,N_142);
nor U8967 (N_8967,N_5166,N_4020);
nor U8968 (N_8968,N_2018,N_5070);
and U8969 (N_8969,N_4820,N_1732);
nand U8970 (N_8970,N_1302,N_1910);
nor U8971 (N_8971,N_1716,N_1158);
nand U8972 (N_8972,N_186,N_2837);
and U8973 (N_8973,N_4401,N_3293);
nand U8974 (N_8974,N_3346,N_4715);
or U8975 (N_8975,N_2036,N_1646);
nand U8976 (N_8976,N_1354,N_4985);
and U8977 (N_8977,N_2130,N_5456);
or U8978 (N_8978,N_4600,N_107);
and U8979 (N_8979,N_2817,N_2588);
nand U8980 (N_8980,N_1362,N_5030);
nand U8981 (N_8981,N_3909,N_2141);
or U8982 (N_8982,N_4915,N_1106);
nor U8983 (N_8983,N_4776,N_4906);
nor U8984 (N_8984,N_2066,N_1466);
and U8985 (N_8985,N_178,N_728);
and U8986 (N_8986,N_2111,N_4181);
xnor U8987 (N_8987,N_1454,N_3738);
and U8988 (N_8988,N_1974,N_4986);
or U8989 (N_8989,N_3674,N_5619);
nand U8990 (N_8990,N_4942,N_1938);
or U8991 (N_8991,N_5979,N_3341);
and U8992 (N_8992,N_116,N_2040);
nand U8993 (N_8993,N_1624,N_5129);
or U8994 (N_8994,N_972,N_3256);
nand U8995 (N_8995,N_3286,N_183);
nand U8996 (N_8996,N_4357,N_3277);
or U8997 (N_8997,N_6121,N_3632);
or U8998 (N_8998,N_5210,N_3295);
xnor U8999 (N_8999,N_2378,N_6174);
xor U9000 (N_9000,N_2638,N_680);
or U9001 (N_9001,N_1486,N_4904);
nor U9002 (N_9002,N_4083,N_5035);
xor U9003 (N_9003,N_174,N_3676);
nor U9004 (N_9004,N_6007,N_4594);
nand U9005 (N_9005,N_997,N_4232);
or U9006 (N_9006,N_3760,N_1349);
nand U9007 (N_9007,N_393,N_5766);
xor U9008 (N_9008,N_6068,N_2954);
nor U9009 (N_9009,N_1855,N_4313);
nor U9010 (N_9010,N_1020,N_4922);
and U9011 (N_9011,N_5056,N_1099);
and U9012 (N_9012,N_5185,N_1871);
nor U9013 (N_9013,N_4644,N_1730);
or U9014 (N_9014,N_2856,N_1325);
xnor U9015 (N_9015,N_2161,N_3727);
nor U9016 (N_9016,N_5255,N_4625);
or U9017 (N_9017,N_4581,N_830);
or U9018 (N_9018,N_595,N_2002);
or U9019 (N_9019,N_5410,N_4044);
and U9020 (N_9020,N_1595,N_1985);
nor U9021 (N_9021,N_4351,N_5741);
nor U9022 (N_9022,N_6021,N_3793);
nor U9023 (N_9023,N_4541,N_568);
nand U9024 (N_9024,N_5819,N_1282);
and U9025 (N_9025,N_4140,N_2523);
and U9026 (N_9026,N_3972,N_1966);
and U9027 (N_9027,N_513,N_4095);
and U9028 (N_9028,N_6020,N_149);
or U9029 (N_9029,N_1904,N_5955);
nor U9030 (N_9030,N_5973,N_2734);
xor U9031 (N_9031,N_5654,N_5346);
xor U9032 (N_9032,N_1782,N_2800);
and U9033 (N_9033,N_3075,N_3437);
nor U9034 (N_9034,N_5367,N_4283);
nand U9035 (N_9035,N_5951,N_3454);
nor U9036 (N_9036,N_4416,N_271);
nor U9037 (N_9037,N_2471,N_5027);
or U9038 (N_9038,N_1170,N_22);
nor U9039 (N_9039,N_1137,N_4139);
xor U9040 (N_9040,N_3219,N_2095);
nor U9041 (N_9041,N_4890,N_2496);
nand U9042 (N_9042,N_4249,N_4505);
and U9043 (N_9043,N_2481,N_2145);
nand U9044 (N_9044,N_2730,N_2656);
xor U9045 (N_9045,N_481,N_1589);
nor U9046 (N_9046,N_3868,N_2037);
nand U9047 (N_9047,N_244,N_2280);
and U9048 (N_9048,N_622,N_2917);
or U9049 (N_9049,N_5167,N_2014);
or U9050 (N_9050,N_2101,N_6075);
xor U9051 (N_9051,N_2795,N_1581);
nor U9052 (N_9052,N_4406,N_1152);
xnor U9053 (N_9053,N_2024,N_3252);
nor U9054 (N_9054,N_2738,N_1909);
nand U9055 (N_9055,N_4349,N_5041);
and U9056 (N_9056,N_630,N_5263);
xor U9057 (N_9057,N_1540,N_3706);
nand U9058 (N_9058,N_3302,N_5524);
nor U9059 (N_9059,N_5517,N_852);
and U9060 (N_9060,N_5387,N_4805);
and U9061 (N_9061,N_4785,N_1927);
nor U9062 (N_9062,N_2438,N_5133);
xnor U9063 (N_9063,N_4887,N_5152);
or U9064 (N_9064,N_5174,N_2525);
nand U9065 (N_9065,N_84,N_1933);
nor U9066 (N_9066,N_2011,N_4160);
nor U9067 (N_9067,N_165,N_4842);
nor U9068 (N_9068,N_3573,N_3649);
nor U9069 (N_9069,N_5735,N_1711);
or U9070 (N_9070,N_4439,N_4811);
and U9071 (N_9071,N_4960,N_4064);
nor U9072 (N_9072,N_4633,N_4651);
and U9073 (N_9073,N_2932,N_4845);
and U9074 (N_9074,N_2020,N_3538);
nor U9075 (N_9075,N_4546,N_3471);
or U9076 (N_9076,N_1738,N_3097);
and U9077 (N_9077,N_539,N_2506);
nor U9078 (N_9078,N_259,N_4376);
nor U9079 (N_9079,N_5560,N_1969);
or U9080 (N_9080,N_4560,N_4258);
nand U9081 (N_9081,N_860,N_2270);
nand U9082 (N_9082,N_4490,N_740);
and U9083 (N_9083,N_3564,N_5270);
nor U9084 (N_9084,N_255,N_2511);
nor U9085 (N_9085,N_1505,N_4777);
nor U9086 (N_9086,N_270,N_844);
and U9087 (N_9087,N_4217,N_5774);
nand U9088 (N_9088,N_1291,N_2419);
nand U9089 (N_9089,N_3441,N_2351);
xnor U9090 (N_9090,N_4941,N_1823);
and U9091 (N_9091,N_538,N_3609);
or U9092 (N_9092,N_1464,N_5350);
nor U9093 (N_9093,N_1875,N_1554);
nor U9094 (N_9094,N_5447,N_5530);
nor U9095 (N_9095,N_4051,N_5633);
xor U9096 (N_9096,N_5574,N_2647);
nand U9097 (N_9097,N_1156,N_2258);
and U9098 (N_9098,N_3490,N_2198);
nor U9099 (N_9099,N_5532,N_4394);
nor U9100 (N_9100,N_3008,N_3994);
and U9101 (N_9101,N_5477,N_5415);
and U9102 (N_9102,N_1818,N_6080);
nor U9103 (N_9103,N_4013,N_4254);
and U9104 (N_9104,N_946,N_3188);
nor U9105 (N_9105,N_943,N_2263);
nand U9106 (N_9106,N_5885,N_1760);
nor U9107 (N_9107,N_1690,N_4891);
nand U9108 (N_9108,N_5786,N_1430);
and U9109 (N_9109,N_2032,N_3818);
nor U9110 (N_9110,N_3306,N_4799);
nand U9111 (N_9111,N_4407,N_3048);
or U9112 (N_9112,N_262,N_5488);
or U9113 (N_9113,N_282,N_4299);
nand U9114 (N_9114,N_3321,N_5077);
or U9115 (N_9115,N_5352,N_1326);
xnor U9116 (N_9116,N_5236,N_4738);
or U9117 (N_9117,N_4089,N_4894);
or U9118 (N_9118,N_2199,N_5797);
nand U9119 (N_9119,N_65,N_2157);
nor U9120 (N_9120,N_712,N_5007);
and U9121 (N_9121,N_902,N_2628);
nand U9122 (N_9122,N_346,N_5151);
xnor U9123 (N_9123,N_4393,N_1380);
and U9124 (N_9124,N_3894,N_6181);
nor U9125 (N_9125,N_2126,N_275);
or U9126 (N_9126,N_3619,N_1524);
and U9127 (N_9127,N_4889,N_63);
nor U9128 (N_9128,N_5186,N_4812);
nor U9129 (N_9129,N_2021,N_3123);
or U9130 (N_9130,N_2809,N_2794);
and U9131 (N_9131,N_4852,N_1269);
nand U9132 (N_9132,N_1764,N_1826);
or U9133 (N_9133,N_922,N_2514);
or U9134 (N_9134,N_387,N_591);
or U9135 (N_9135,N_1,N_2086);
and U9136 (N_9136,N_6216,N_4049);
nor U9137 (N_9137,N_5238,N_4193);
and U9138 (N_9138,N_4639,N_5962);
or U9139 (N_9139,N_5264,N_2129);
xor U9140 (N_9140,N_1129,N_5661);
and U9141 (N_9141,N_304,N_2530);
and U9142 (N_9142,N_5976,N_4949);
and U9143 (N_9143,N_3640,N_4586);
nor U9144 (N_9144,N_5274,N_4711);
nand U9145 (N_9145,N_803,N_239);
nand U9146 (N_9146,N_2347,N_5401);
or U9147 (N_9147,N_2269,N_2193);
or U9148 (N_9148,N_736,N_6134);
nor U9149 (N_9149,N_4411,N_2804);
nand U9150 (N_9150,N_2865,N_2771);
nand U9151 (N_9151,N_3664,N_5997);
or U9152 (N_9152,N_776,N_4495);
nand U9153 (N_9153,N_4623,N_2286);
and U9154 (N_9154,N_4111,N_2062);
xnor U9155 (N_9155,N_958,N_3953);
nor U9156 (N_9156,N_2793,N_4520);
or U9157 (N_9157,N_6152,N_3559);
nor U9158 (N_9158,N_1284,N_1429);
nor U9159 (N_9159,N_705,N_5936);
or U9160 (N_9160,N_1440,N_1285);
and U9161 (N_9161,N_5637,N_4746);
nand U9162 (N_9162,N_575,N_3147);
and U9163 (N_9163,N_5933,N_3397);
or U9164 (N_9164,N_2148,N_5206);
or U9165 (N_9165,N_679,N_5695);
or U9166 (N_9166,N_1251,N_2519);
nand U9167 (N_9167,N_4617,N_4608);
nand U9168 (N_9168,N_2707,N_5194);
nand U9169 (N_9169,N_2019,N_5278);
or U9170 (N_9170,N_4214,N_1065);
nor U9171 (N_9171,N_2706,N_1381);
or U9172 (N_9172,N_3150,N_122);
xor U9173 (N_9173,N_3787,N_2689);
and U9174 (N_9174,N_349,N_5145);
nor U9175 (N_9175,N_6093,N_121);
nand U9176 (N_9176,N_2991,N_4361);
nand U9177 (N_9177,N_5789,N_4851);
nand U9178 (N_9178,N_1390,N_2702);
xnor U9179 (N_9179,N_3533,N_3714);
and U9180 (N_9180,N_2672,N_320);
xnor U9181 (N_9181,N_37,N_3778);
nand U9182 (N_9182,N_4733,N_1940);
nand U9183 (N_9183,N_6113,N_5239);
and U9184 (N_9184,N_4501,N_1784);
nor U9185 (N_9185,N_3739,N_4844);
nand U9186 (N_9186,N_3202,N_3544);
or U9187 (N_9187,N_23,N_3593);
nor U9188 (N_9188,N_5762,N_167);
nand U9189 (N_9189,N_3100,N_3106);
and U9190 (N_9190,N_4953,N_1419);
and U9191 (N_9191,N_5925,N_1009);
and U9192 (N_9192,N_4492,N_4513);
xor U9193 (N_9193,N_4097,N_1539);
or U9194 (N_9194,N_2693,N_708);
and U9195 (N_9195,N_3511,N_1216);
or U9196 (N_9196,N_57,N_854);
nand U9197 (N_9197,N_3694,N_5382);
or U9198 (N_9198,N_5691,N_3290);
nor U9199 (N_9199,N_3114,N_2307);
and U9200 (N_9200,N_3776,N_6109);
and U9201 (N_9201,N_2120,N_676);
nor U9202 (N_9202,N_2058,N_5612);
and U9203 (N_9203,N_838,N_2349);
xor U9204 (N_9204,N_702,N_2003);
nand U9205 (N_9205,N_3030,N_380);
xnor U9206 (N_9206,N_3411,N_3677);
nor U9207 (N_9207,N_4762,N_6042);
nand U9208 (N_9208,N_1032,N_4994);
nand U9209 (N_9209,N_4152,N_2390);
nand U9210 (N_9210,N_1955,N_4474);
nand U9211 (N_9211,N_4857,N_5271);
nand U9212 (N_9212,N_2156,N_323);
nor U9213 (N_9213,N_261,N_5990);
nor U9214 (N_9214,N_6107,N_654);
or U9215 (N_9215,N_1516,N_1555);
or U9216 (N_9216,N_196,N_6128);
nor U9217 (N_9217,N_5122,N_661);
xor U9218 (N_9218,N_3355,N_3021);
nand U9219 (N_9219,N_2393,N_2486);
nor U9220 (N_9220,N_3173,N_77);
and U9221 (N_9221,N_1619,N_703);
or U9222 (N_9222,N_1852,N_1898);
nand U9223 (N_9223,N_4028,N_2946);
and U9224 (N_9224,N_253,N_6055);
and U9225 (N_9225,N_3468,N_500);
or U9226 (N_9226,N_4450,N_851);
or U9227 (N_9227,N_5497,N_4841);
nand U9228 (N_9228,N_2312,N_1578);
xnor U9229 (N_9229,N_4969,N_3561);
and U9230 (N_9230,N_5110,N_3230);
or U9231 (N_9231,N_3452,N_1206);
and U9232 (N_9232,N_847,N_1571);
nor U9233 (N_9233,N_227,N_5673);
xnor U9234 (N_9234,N_694,N_6142);
nor U9235 (N_9235,N_5881,N_3502);
nand U9236 (N_9236,N_2960,N_4800);
nand U9237 (N_9237,N_1611,N_2727);
and U9238 (N_9238,N_2870,N_5593);
and U9239 (N_9239,N_6213,N_4909);
xor U9240 (N_9240,N_1669,N_4500);
or U9241 (N_9241,N_1806,N_4326);
nand U9242 (N_9242,N_5209,N_4629);
or U9243 (N_9243,N_5120,N_5033);
xor U9244 (N_9244,N_5458,N_4238);
nor U9245 (N_9245,N_5002,N_5873);
nand U9246 (N_9246,N_582,N_3627);
or U9247 (N_9247,N_2711,N_3864);
xnor U9248 (N_9248,N_1612,N_3066);
and U9249 (N_9249,N_3545,N_508);
nand U9250 (N_9250,N_2762,N_4911);
nor U9251 (N_9251,N_3499,N_6221);
and U9252 (N_9252,N_5064,N_4786);
or U9253 (N_9253,N_5136,N_5089);
nand U9254 (N_9254,N_233,N_5242);
or U9255 (N_9255,N_1364,N_1888);
or U9256 (N_9256,N_2044,N_2695);
or U9257 (N_9257,N_4716,N_5794);
or U9258 (N_9258,N_4725,N_197);
or U9259 (N_9259,N_1939,N_4532);
nand U9260 (N_9260,N_1789,N_638);
nand U9261 (N_9261,N_3834,N_4341);
or U9262 (N_9262,N_3056,N_3272);
nand U9263 (N_9263,N_3841,N_3268);
nand U9264 (N_9264,N_4188,N_4562);
and U9265 (N_9265,N_849,N_1860);
or U9266 (N_9266,N_5958,N_3688);
nand U9267 (N_9267,N_2948,N_6183);
nor U9268 (N_9268,N_1774,N_6238);
nor U9269 (N_9269,N_2224,N_1204);
xnor U9270 (N_9270,N_925,N_4773);
or U9271 (N_9271,N_1196,N_1278);
nor U9272 (N_9272,N_5223,N_2950);
nand U9273 (N_9273,N_4395,N_1133);
and U9274 (N_9274,N_3029,N_2046);
or U9275 (N_9275,N_4239,N_4783);
xor U9276 (N_9276,N_1971,N_6111);
and U9277 (N_9277,N_3546,N_3525);
nand U9278 (N_9278,N_225,N_5585);
nand U9279 (N_9279,N_5127,N_1238);
nand U9280 (N_9280,N_597,N_5878);
or U9281 (N_9281,N_3167,N_1944);
nand U9282 (N_9282,N_892,N_2887);
nand U9283 (N_9283,N_811,N_1576);
nand U9284 (N_9284,N_5473,N_4865);
nor U9285 (N_9285,N_1843,N_4739);
nand U9286 (N_9286,N_3235,N_3152);
nor U9287 (N_9287,N_720,N_201);
xor U9288 (N_9288,N_4660,N_5769);
and U9289 (N_9289,N_867,N_3635);
and U9290 (N_9290,N_1410,N_2906);
xnor U9291 (N_9291,N_995,N_3462);
or U9292 (N_9292,N_3307,N_3907);
xnor U9293 (N_9293,N_5938,N_4216);
xnor U9294 (N_9294,N_1743,N_839);
and U9295 (N_9295,N_5780,N_5374);
nor U9296 (N_9296,N_758,N_5103);
nor U9297 (N_9297,N_390,N_156);
nand U9298 (N_9298,N_2009,N_5328);
nand U9299 (N_9299,N_3772,N_1785);
nor U9300 (N_9300,N_2211,N_3617);
xor U9301 (N_9301,N_579,N_1268);
nand U9302 (N_9302,N_3821,N_1610);
xor U9303 (N_9303,N_4819,N_4477);
and U9304 (N_9304,N_1214,N_533);
and U9305 (N_9305,N_6073,N_4722);
nand U9306 (N_9306,N_1733,N_2466);
xor U9307 (N_9307,N_895,N_5146);
or U9308 (N_9308,N_2915,N_5320);
nand U9309 (N_9309,N_5512,N_713);
nor U9310 (N_9310,N_1399,N_761);
nor U9311 (N_9311,N_5454,N_5503);
and U9312 (N_9312,N_3595,N_457);
and U9313 (N_9313,N_1625,N_5705);
and U9314 (N_9314,N_280,N_5781);
or U9315 (N_9315,N_2557,N_737);
xnor U9316 (N_9316,N_2262,N_162);
nor U9317 (N_9317,N_2000,N_5507);
nor U9318 (N_9318,N_1968,N_1481);
nor U9319 (N_9319,N_5965,N_2284);
nor U9320 (N_9320,N_5567,N_4821);
and U9321 (N_9321,N_2333,N_4263);
xor U9322 (N_9322,N_6032,N_3925);
nor U9323 (N_9323,N_2860,N_3416);
nor U9324 (N_9324,N_2314,N_4620);
nand U9325 (N_9325,N_5880,N_3296);
nand U9326 (N_9326,N_1357,N_2176);
or U9327 (N_9327,N_5267,N_1678);
or U9328 (N_9328,N_1506,N_1090);
and U9329 (N_9329,N_4588,N_745);
and U9330 (N_9330,N_5251,N_4918);
and U9331 (N_9331,N_1777,N_4665);
or U9332 (N_9332,N_5528,N_2383);
and U9333 (N_9333,N_1135,N_322);
or U9334 (N_9334,N_5618,N_5561);
and U9335 (N_9335,N_2746,N_5313);
nor U9336 (N_9336,N_1844,N_211);
or U9337 (N_9337,N_802,N_5742);
xor U9338 (N_9338,N_2376,N_3736);
xor U9339 (N_9339,N_290,N_1582);
nand U9340 (N_9340,N_3308,N_4833);
and U9341 (N_9341,N_52,N_4078);
nor U9342 (N_9342,N_1267,N_2701);
nand U9343 (N_9343,N_5775,N_6137);
and U9344 (N_9344,N_5202,N_4899);
nor U9345 (N_9345,N_2317,N_2898);
or U9346 (N_9346,N_6248,N_4897);
or U9347 (N_9347,N_1511,N_2325);
and U9348 (N_9348,N_1534,N_5442);
nor U9349 (N_9349,N_1140,N_338);
and U9350 (N_9350,N_299,N_4331);
nor U9351 (N_9351,N_2143,N_2056);
nand U9352 (N_9352,N_4916,N_5181);
and U9353 (N_9353,N_175,N_7);
or U9354 (N_9354,N_6091,N_2051);
nor U9355 (N_9355,N_1232,N_4177);
nand U9356 (N_9356,N_3920,N_1665);
or U9357 (N_9357,N_5825,N_1642);
and U9358 (N_9358,N_120,N_1102);
and U9359 (N_9359,N_3001,N_4945);
nand U9360 (N_9360,N_236,N_5343);
or U9361 (N_9361,N_3637,N_3903);
nor U9362 (N_9362,N_2234,N_5855);
and U9363 (N_9363,N_2241,N_826);
nand U9364 (N_9364,N_5148,N_2665);
xnor U9365 (N_9365,N_859,N_1836);
and U9366 (N_9366,N_3950,N_2957);
or U9367 (N_9367,N_1767,N_1891);
nor U9368 (N_9368,N_4880,N_5943);
and U9369 (N_9369,N_478,N_4333);
nor U9370 (N_9370,N_2399,N_5468);
nor U9371 (N_9371,N_3467,N_527);
and U9372 (N_9372,N_2127,N_4045);
nor U9373 (N_9373,N_2703,N_4510);
and U9374 (N_9374,N_3455,N_1157);
nor U9375 (N_9375,N_5591,N_2526);
xor U9376 (N_9376,N_89,N_4963);
and U9377 (N_9377,N_852,N_1903);
and U9378 (N_9378,N_5828,N_3305);
nand U9379 (N_9379,N_2393,N_502);
nor U9380 (N_9380,N_2790,N_3714);
or U9381 (N_9381,N_2237,N_4632);
or U9382 (N_9382,N_3157,N_2459);
nor U9383 (N_9383,N_6119,N_705);
or U9384 (N_9384,N_1021,N_729);
xnor U9385 (N_9385,N_1630,N_3183);
xnor U9386 (N_9386,N_719,N_31);
xor U9387 (N_9387,N_3073,N_2498);
nor U9388 (N_9388,N_2889,N_2217);
or U9389 (N_9389,N_5910,N_5419);
and U9390 (N_9390,N_52,N_24);
nand U9391 (N_9391,N_1978,N_147);
nand U9392 (N_9392,N_3686,N_1314);
nor U9393 (N_9393,N_3213,N_6134);
or U9394 (N_9394,N_6006,N_1660);
and U9395 (N_9395,N_882,N_2795);
nor U9396 (N_9396,N_3992,N_813);
or U9397 (N_9397,N_940,N_2563);
and U9398 (N_9398,N_6023,N_4218);
and U9399 (N_9399,N_5875,N_5360);
or U9400 (N_9400,N_6240,N_1151);
nor U9401 (N_9401,N_1729,N_4010);
or U9402 (N_9402,N_1654,N_4291);
nand U9403 (N_9403,N_4888,N_865);
nand U9404 (N_9404,N_3499,N_1156);
or U9405 (N_9405,N_2503,N_4033);
or U9406 (N_9406,N_3855,N_671);
nand U9407 (N_9407,N_2096,N_4120);
nand U9408 (N_9408,N_1046,N_5646);
nand U9409 (N_9409,N_988,N_5619);
and U9410 (N_9410,N_3656,N_3460);
nor U9411 (N_9411,N_5398,N_954);
or U9412 (N_9412,N_4492,N_4060);
or U9413 (N_9413,N_4553,N_4298);
nand U9414 (N_9414,N_140,N_1496);
nor U9415 (N_9415,N_3034,N_2302);
nand U9416 (N_9416,N_6042,N_3511);
or U9417 (N_9417,N_4886,N_4555);
nor U9418 (N_9418,N_5860,N_5208);
and U9419 (N_9419,N_3587,N_3548);
or U9420 (N_9420,N_884,N_423);
or U9421 (N_9421,N_1638,N_5745);
nor U9422 (N_9422,N_3307,N_880);
xnor U9423 (N_9423,N_709,N_838);
or U9424 (N_9424,N_2918,N_3610);
or U9425 (N_9425,N_5921,N_3726);
nand U9426 (N_9426,N_434,N_1242);
or U9427 (N_9427,N_2346,N_5251);
or U9428 (N_9428,N_3156,N_3660);
nand U9429 (N_9429,N_393,N_1988);
and U9430 (N_9430,N_784,N_1102);
or U9431 (N_9431,N_2004,N_3357);
or U9432 (N_9432,N_353,N_2168);
and U9433 (N_9433,N_1946,N_5124);
and U9434 (N_9434,N_3317,N_5397);
or U9435 (N_9435,N_2079,N_3614);
nor U9436 (N_9436,N_1887,N_3315);
and U9437 (N_9437,N_3333,N_5884);
nor U9438 (N_9438,N_4493,N_6139);
and U9439 (N_9439,N_1499,N_5719);
or U9440 (N_9440,N_3707,N_4955);
nand U9441 (N_9441,N_2830,N_4920);
xor U9442 (N_9442,N_3746,N_3172);
nor U9443 (N_9443,N_4703,N_4037);
xor U9444 (N_9444,N_3311,N_1370);
nor U9445 (N_9445,N_613,N_3900);
or U9446 (N_9446,N_820,N_4790);
nor U9447 (N_9447,N_2073,N_615);
or U9448 (N_9448,N_6142,N_5750);
nand U9449 (N_9449,N_3853,N_6220);
and U9450 (N_9450,N_5973,N_3109);
or U9451 (N_9451,N_2528,N_4872);
or U9452 (N_9452,N_1426,N_3832);
nand U9453 (N_9453,N_242,N_3435);
nand U9454 (N_9454,N_828,N_998);
or U9455 (N_9455,N_1964,N_3192);
or U9456 (N_9456,N_2257,N_1019);
nor U9457 (N_9457,N_536,N_1354);
or U9458 (N_9458,N_3091,N_2515);
nor U9459 (N_9459,N_5537,N_110);
and U9460 (N_9460,N_3481,N_6010);
nor U9461 (N_9461,N_1396,N_2088);
and U9462 (N_9462,N_2247,N_4560);
or U9463 (N_9463,N_5957,N_1235);
and U9464 (N_9464,N_1067,N_2509);
or U9465 (N_9465,N_1803,N_5103);
or U9466 (N_9466,N_4432,N_2311);
nor U9467 (N_9467,N_4929,N_5225);
nand U9468 (N_9468,N_3236,N_2391);
nor U9469 (N_9469,N_506,N_5121);
or U9470 (N_9470,N_296,N_6103);
and U9471 (N_9471,N_2399,N_2118);
nor U9472 (N_9472,N_1457,N_72);
and U9473 (N_9473,N_4965,N_1231);
nand U9474 (N_9474,N_202,N_1844);
nand U9475 (N_9475,N_406,N_683);
or U9476 (N_9476,N_3333,N_1828);
and U9477 (N_9477,N_1021,N_4345);
or U9478 (N_9478,N_2973,N_257);
nor U9479 (N_9479,N_97,N_35);
or U9480 (N_9480,N_361,N_5366);
and U9481 (N_9481,N_167,N_521);
or U9482 (N_9482,N_230,N_2844);
nor U9483 (N_9483,N_621,N_3173);
xor U9484 (N_9484,N_2376,N_6009);
nor U9485 (N_9485,N_3556,N_702);
nand U9486 (N_9486,N_4838,N_1416);
and U9487 (N_9487,N_5260,N_5427);
nand U9488 (N_9488,N_4331,N_4960);
xnor U9489 (N_9489,N_1068,N_5057);
or U9490 (N_9490,N_969,N_1769);
or U9491 (N_9491,N_2988,N_5173);
nand U9492 (N_9492,N_6218,N_5720);
nor U9493 (N_9493,N_3362,N_2784);
or U9494 (N_9494,N_2585,N_1124);
nand U9495 (N_9495,N_1937,N_436);
and U9496 (N_9496,N_1142,N_3352);
nand U9497 (N_9497,N_4062,N_5620);
xor U9498 (N_9498,N_4302,N_359);
xor U9499 (N_9499,N_4153,N_1406);
and U9500 (N_9500,N_3016,N_1916);
and U9501 (N_9501,N_2454,N_1225);
or U9502 (N_9502,N_5387,N_3460);
or U9503 (N_9503,N_6066,N_2850);
or U9504 (N_9504,N_3634,N_2230);
nand U9505 (N_9505,N_944,N_5845);
xor U9506 (N_9506,N_683,N_3408);
and U9507 (N_9507,N_4228,N_567);
and U9508 (N_9508,N_2131,N_2573);
nand U9509 (N_9509,N_5316,N_94);
and U9510 (N_9510,N_5477,N_3908);
nand U9511 (N_9511,N_32,N_3220);
or U9512 (N_9512,N_3760,N_435);
nand U9513 (N_9513,N_5392,N_4439);
or U9514 (N_9514,N_5446,N_5350);
or U9515 (N_9515,N_2722,N_6124);
and U9516 (N_9516,N_4776,N_337);
nor U9517 (N_9517,N_5699,N_2378);
nand U9518 (N_9518,N_5096,N_6174);
nor U9519 (N_9519,N_5376,N_1980);
nor U9520 (N_9520,N_1795,N_1020);
nor U9521 (N_9521,N_391,N_2224);
nand U9522 (N_9522,N_4712,N_5125);
and U9523 (N_9523,N_5650,N_3701);
nor U9524 (N_9524,N_5369,N_1323);
and U9525 (N_9525,N_5993,N_2437);
or U9526 (N_9526,N_1484,N_378);
nor U9527 (N_9527,N_173,N_2282);
nor U9528 (N_9528,N_6182,N_5119);
nand U9529 (N_9529,N_1565,N_3852);
or U9530 (N_9530,N_1672,N_23);
nor U9531 (N_9531,N_4307,N_3531);
and U9532 (N_9532,N_5775,N_5557);
nand U9533 (N_9533,N_509,N_81);
nor U9534 (N_9534,N_433,N_5520);
nor U9535 (N_9535,N_4182,N_3928);
and U9536 (N_9536,N_5196,N_5033);
nor U9537 (N_9537,N_77,N_1645);
nand U9538 (N_9538,N_1804,N_2577);
and U9539 (N_9539,N_6103,N_4652);
and U9540 (N_9540,N_5726,N_4287);
and U9541 (N_9541,N_5140,N_5493);
nand U9542 (N_9542,N_1182,N_324);
and U9543 (N_9543,N_4663,N_645);
or U9544 (N_9544,N_3538,N_3816);
and U9545 (N_9545,N_2384,N_5393);
or U9546 (N_9546,N_4100,N_3787);
and U9547 (N_9547,N_639,N_1158);
nand U9548 (N_9548,N_221,N_2765);
or U9549 (N_9549,N_817,N_5242);
nor U9550 (N_9550,N_4514,N_4513);
nor U9551 (N_9551,N_2589,N_1349);
xor U9552 (N_9552,N_4621,N_5770);
and U9553 (N_9553,N_867,N_2951);
and U9554 (N_9554,N_4048,N_4783);
or U9555 (N_9555,N_579,N_5680);
nor U9556 (N_9556,N_4915,N_3232);
and U9557 (N_9557,N_517,N_5212);
and U9558 (N_9558,N_1819,N_4405);
and U9559 (N_9559,N_2501,N_1921);
or U9560 (N_9560,N_5770,N_5579);
nand U9561 (N_9561,N_2646,N_246);
xnor U9562 (N_9562,N_3192,N_2628);
or U9563 (N_9563,N_6208,N_2031);
and U9564 (N_9564,N_1644,N_5115);
or U9565 (N_9565,N_5893,N_1285);
and U9566 (N_9566,N_1279,N_1091);
and U9567 (N_9567,N_2512,N_3750);
nand U9568 (N_9568,N_2839,N_4684);
or U9569 (N_9569,N_1030,N_3517);
nand U9570 (N_9570,N_1489,N_3957);
and U9571 (N_9571,N_2945,N_1576);
and U9572 (N_9572,N_3531,N_5760);
or U9573 (N_9573,N_2838,N_4670);
nor U9574 (N_9574,N_3729,N_3097);
nand U9575 (N_9575,N_5235,N_1150);
nor U9576 (N_9576,N_5109,N_3283);
or U9577 (N_9577,N_5030,N_3592);
nand U9578 (N_9578,N_5576,N_5149);
or U9579 (N_9579,N_1515,N_1029);
nand U9580 (N_9580,N_4206,N_4251);
nor U9581 (N_9581,N_2459,N_5667);
or U9582 (N_9582,N_4218,N_3631);
and U9583 (N_9583,N_594,N_1942);
or U9584 (N_9584,N_966,N_1271);
nor U9585 (N_9585,N_2707,N_3752);
nor U9586 (N_9586,N_2241,N_2303);
nand U9587 (N_9587,N_2974,N_3918);
xor U9588 (N_9588,N_4380,N_498);
nand U9589 (N_9589,N_4307,N_2081);
nand U9590 (N_9590,N_4969,N_5065);
nand U9591 (N_9591,N_5215,N_2122);
and U9592 (N_9592,N_444,N_3003);
and U9593 (N_9593,N_3270,N_6091);
and U9594 (N_9594,N_955,N_5381);
nand U9595 (N_9595,N_4739,N_2610);
or U9596 (N_9596,N_589,N_2147);
or U9597 (N_9597,N_4260,N_5012);
nor U9598 (N_9598,N_2747,N_4827);
and U9599 (N_9599,N_446,N_5229);
or U9600 (N_9600,N_5976,N_2986);
nor U9601 (N_9601,N_2991,N_3977);
and U9602 (N_9602,N_4025,N_747);
nor U9603 (N_9603,N_4758,N_1303);
xor U9604 (N_9604,N_818,N_3597);
nand U9605 (N_9605,N_6201,N_2775);
and U9606 (N_9606,N_3371,N_3072);
and U9607 (N_9607,N_942,N_2648);
nor U9608 (N_9608,N_6187,N_293);
or U9609 (N_9609,N_1015,N_1277);
xnor U9610 (N_9610,N_1454,N_5203);
nand U9611 (N_9611,N_1048,N_456);
nand U9612 (N_9612,N_2159,N_2789);
or U9613 (N_9613,N_128,N_585);
nor U9614 (N_9614,N_5032,N_5800);
or U9615 (N_9615,N_2480,N_97);
nor U9616 (N_9616,N_5511,N_4056);
xor U9617 (N_9617,N_238,N_4426);
nand U9618 (N_9618,N_5040,N_6161);
nor U9619 (N_9619,N_5302,N_581);
and U9620 (N_9620,N_3380,N_3748);
nor U9621 (N_9621,N_10,N_5313);
nand U9622 (N_9622,N_5925,N_5589);
nand U9623 (N_9623,N_4456,N_730);
nor U9624 (N_9624,N_3162,N_5665);
xnor U9625 (N_9625,N_3018,N_192);
or U9626 (N_9626,N_5827,N_955);
nor U9627 (N_9627,N_1225,N_4355);
nor U9628 (N_9628,N_5932,N_5858);
or U9629 (N_9629,N_4610,N_4561);
or U9630 (N_9630,N_5046,N_4977);
and U9631 (N_9631,N_1035,N_269);
nand U9632 (N_9632,N_2918,N_2678);
nand U9633 (N_9633,N_5246,N_1017);
nor U9634 (N_9634,N_5923,N_5875);
nand U9635 (N_9635,N_1322,N_2389);
or U9636 (N_9636,N_309,N_1248);
and U9637 (N_9637,N_735,N_4983);
and U9638 (N_9638,N_4416,N_5636);
or U9639 (N_9639,N_1931,N_5947);
or U9640 (N_9640,N_1062,N_2868);
nor U9641 (N_9641,N_4861,N_5832);
xor U9642 (N_9642,N_4175,N_5583);
and U9643 (N_9643,N_1712,N_936);
and U9644 (N_9644,N_1871,N_3921);
nand U9645 (N_9645,N_3517,N_6143);
and U9646 (N_9646,N_3275,N_5100);
nor U9647 (N_9647,N_4511,N_785);
xnor U9648 (N_9648,N_2751,N_5481);
nor U9649 (N_9649,N_5501,N_2221);
and U9650 (N_9650,N_1366,N_3573);
xor U9651 (N_9651,N_1250,N_5136);
nand U9652 (N_9652,N_4846,N_1541);
nand U9653 (N_9653,N_5458,N_1227);
and U9654 (N_9654,N_3426,N_3686);
and U9655 (N_9655,N_5215,N_1686);
nand U9656 (N_9656,N_5118,N_4250);
and U9657 (N_9657,N_5516,N_2911);
nor U9658 (N_9658,N_5642,N_3941);
nor U9659 (N_9659,N_4200,N_1067);
nor U9660 (N_9660,N_2768,N_548);
nor U9661 (N_9661,N_4078,N_2870);
and U9662 (N_9662,N_2320,N_5165);
nand U9663 (N_9663,N_1669,N_1688);
and U9664 (N_9664,N_1224,N_3508);
nor U9665 (N_9665,N_4069,N_646);
nand U9666 (N_9666,N_1260,N_4391);
and U9667 (N_9667,N_5086,N_428);
or U9668 (N_9668,N_5964,N_1198);
and U9669 (N_9669,N_4803,N_904);
and U9670 (N_9670,N_360,N_284);
nand U9671 (N_9671,N_616,N_5017);
and U9672 (N_9672,N_1728,N_2411);
or U9673 (N_9673,N_804,N_2264);
and U9674 (N_9674,N_5855,N_1690);
xor U9675 (N_9675,N_452,N_5694);
nand U9676 (N_9676,N_1565,N_1211);
or U9677 (N_9677,N_1931,N_5634);
nor U9678 (N_9678,N_4634,N_3720);
and U9679 (N_9679,N_3045,N_896);
xor U9680 (N_9680,N_5725,N_354);
nand U9681 (N_9681,N_5340,N_394);
and U9682 (N_9682,N_5270,N_4281);
and U9683 (N_9683,N_5679,N_2605);
and U9684 (N_9684,N_4935,N_278);
nor U9685 (N_9685,N_2712,N_5862);
xor U9686 (N_9686,N_2187,N_448);
and U9687 (N_9687,N_4902,N_3573);
nand U9688 (N_9688,N_1234,N_6163);
and U9689 (N_9689,N_4316,N_1145);
nand U9690 (N_9690,N_6185,N_1076);
xnor U9691 (N_9691,N_2562,N_5998);
and U9692 (N_9692,N_4638,N_3075);
and U9693 (N_9693,N_413,N_6235);
and U9694 (N_9694,N_64,N_5604);
xor U9695 (N_9695,N_3110,N_3540);
or U9696 (N_9696,N_2849,N_1384);
nand U9697 (N_9697,N_1467,N_4808);
and U9698 (N_9698,N_5254,N_1840);
nor U9699 (N_9699,N_6149,N_5886);
or U9700 (N_9700,N_6215,N_1389);
nor U9701 (N_9701,N_1669,N_4747);
nand U9702 (N_9702,N_3078,N_2747);
and U9703 (N_9703,N_2651,N_5607);
nand U9704 (N_9704,N_5113,N_3955);
or U9705 (N_9705,N_1257,N_6164);
xnor U9706 (N_9706,N_2868,N_5691);
and U9707 (N_9707,N_1566,N_1657);
nor U9708 (N_9708,N_5847,N_837);
nor U9709 (N_9709,N_2802,N_3229);
nor U9710 (N_9710,N_4355,N_4641);
and U9711 (N_9711,N_4887,N_4206);
or U9712 (N_9712,N_1003,N_177);
or U9713 (N_9713,N_2442,N_725);
and U9714 (N_9714,N_2606,N_5965);
xor U9715 (N_9715,N_1269,N_65);
xnor U9716 (N_9716,N_4150,N_4530);
or U9717 (N_9717,N_2125,N_5782);
nor U9718 (N_9718,N_5867,N_5250);
nor U9719 (N_9719,N_5520,N_4396);
or U9720 (N_9720,N_1976,N_6059);
xnor U9721 (N_9721,N_684,N_2692);
nor U9722 (N_9722,N_1039,N_5834);
nor U9723 (N_9723,N_5755,N_2882);
xor U9724 (N_9724,N_3582,N_6002);
xnor U9725 (N_9725,N_3892,N_3774);
or U9726 (N_9726,N_612,N_1022);
or U9727 (N_9727,N_1602,N_3260);
and U9728 (N_9728,N_6212,N_2170);
xor U9729 (N_9729,N_899,N_4532);
nand U9730 (N_9730,N_1009,N_117);
or U9731 (N_9731,N_1674,N_3333);
and U9732 (N_9732,N_6109,N_4597);
xor U9733 (N_9733,N_2035,N_2362);
and U9734 (N_9734,N_2891,N_757);
or U9735 (N_9735,N_4551,N_3798);
or U9736 (N_9736,N_4622,N_5092);
and U9737 (N_9737,N_8,N_971);
and U9738 (N_9738,N_2370,N_5001);
nor U9739 (N_9739,N_446,N_5443);
nor U9740 (N_9740,N_1956,N_4545);
nand U9741 (N_9741,N_2593,N_5219);
nor U9742 (N_9742,N_4529,N_6071);
or U9743 (N_9743,N_4158,N_5055);
nor U9744 (N_9744,N_3195,N_1548);
xor U9745 (N_9745,N_3376,N_3705);
and U9746 (N_9746,N_2088,N_4432);
or U9747 (N_9747,N_2652,N_1669);
nand U9748 (N_9748,N_2262,N_2011);
nand U9749 (N_9749,N_1201,N_5201);
nor U9750 (N_9750,N_2048,N_323);
and U9751 (N_9751,N_3769,N_2741);
nand U9752 (N_9752,N_976,N_1933);
or U9753 (N_9753,N_1613,N_651);
nand U9754 (N_9754,N_4127,N_4757);
xor U9755 (N_9755,N_4954,N_5795);
nand U9756 (N_9756,N_4509,N_4137);
xnor U9757 (N_9757,N_5871,N_2115);
and U9758 (N_9758,N_2306,N_1246);
xor U9759 (N_9759,N_4102,N_4394);
or U9760 (N_9760,N_4566,N_942);
nand U9761 (N_9761,N_1287,N_6214);
or U9762 (N_9762,N_207,N_833);
and U9763 (N_9763,N_2778,N_987);
xor U9764 (N_9764,N_5672,N_5014);
and U9765 (N_9765,N_3832,N_6191);
and U9766 (N_9766,N_3506,N_1300);
and U9767 (N_9767,N_1937,N_1940);
nand U9768 (N_9768,N_4256,N_838);
xnor U9769 (N_9769,N_1326,N_6166);
and U9770 (N_9770,N_3584,N_130);
nor U9771 (N_9771,N_766,N_3769);
or U9772 (N_9772,N_3231,N_974);
and U9773 (N_9773,N_3702,N_3115);
xor U9774 (N_9774,N_1743,N_1897);
nor U9775 (N_9775,N_6093,N_3673);
or U9776 (N_9776,N_4650,N_5586);
nand U9777 (N_9777,N_6154,N_3231);
xor U9778 (N_9778,N_4527,N_5988);
nor U9779 (N_9779,N_5247,N_1976);
or U9780 (N_9780,N_5758,N_1260);
nor U9781 (N_9781,N_4568,N_611);
nand U9782 (N_9782,N_3013,N_3845);
and U9783 (N_9783,N_3988,N_6225);
nand U9784 (N_9784,N_3635,N_1089);
and U9785 (N_9785,N_3741,N_3091);
nor U9786 (N_9786,N_5817,N_2995);
and U9787 (N_9787,N_4125,N_3587);
xnor U9788 (N_9788,N_6131,N_3605);
nor U9789 (N_9789,N_1894,N_2244);
or U9790 (N_9790,N_5874,N_622);
or U9791 (N_9791,N_2392,N_3398);
and U9792 (N_9792,N_5138,N_5780);
or U9793 (N_9793,N_171,N_5173);
nand U9794 (N_9794,N_5279,N_5388);
nand U9795 (N_9795,N_612,N_705);
or U9796 (N_9796,N_4525,N_2665);
xnor U9797 (N_9797,N_2856,N_3768);
and U9798 (N_9798,N_157,N_2388);
nand U9799 (N_9799,N_5891,N_5014);
and U9800 (N_9800,N_1789,N_978);
or U9801 (N_9801,N_4502,N_4863);
nor U9802 (N_9802,N_4079,N_2298);
and U9803 (N_9803,N_5245,N_2987);
nand U9804 (N_9804,N_3236,N_906);
nor U9805 (N_9805,N_4263,N_5640);
and U9806 (N_9806,N_1101,N_802);
and U9807 (N_9807,N_2610,N_3223);
xnor U9808 (N_9808,N_1072,N_2239);
nor U9809 (N_9809,N_4531,N_6041);
or U9810 (N_9810,N_5168,N_365);
or U9811 (N_9811,N_4519,N_4574);
and U9812 (N_9812,N_4801,N_5370);
nor U9813 (N_9813,N_626,N_188);
or U9814 (N_9814,N_3181,N_5007);
nor U9815 (N_9815,N_3389,N_512);
nand U9816 (N_9816,N_1078,N_5196);
nor U9817 (N_9817,N_4680,N_2406);
nor U9818 (N_9818,N_4142,N_3658);
or U9819 (N_9819,N_1789,N_1854);
or U9820 (N_9820,N_4381,N_6125);
or U9821 (N_9821,N_5919,N_3387);
and U9822 (N_9822,N_467,N_4552);
or U9823 (N_9823,N_446,N_5210);
nor U9824 (N_9824,N_50,N_928);
nand U9825 (N_9825,N_5933,N_6027);
nand U9826 (N_9826,N_2725,N_2046);
nor U9827 (N_9827,N_2890,N_4994);
xor U9828 (N_9828,N_4305,N_141);
xnor U9829 (N_9829,N_5606,N_3288);
and U9830 (N_9830,N_1409,N_2812);
or U9831 (N_9831,N_3909,N_4889);
nand U9832 (N_9832,N_5298,N_4883);
and U9833 (N_9833,N_137,N_2586);
or U9834 (N_9834,N_6232,N_3618);
nand U9835 (N_9835,N_454,N_3163);
xor U9836 (N_9836,N_2969,N_4534);
nor U9837 (N_9837,N_879,N_3909);
nor U9838 (N_9838,N_1704,N_4620);
nor U9839 (N_9839,N_4832,N_2640);
nand U9840 (N_9840,N_4824,N_5213);
nand U9841 (N_9841,N_5377,N_2261);
nor U9842 (N_9842,N_789,N_2812);
and U9843 (N_9843,N_5655,N_1889);
nor U9844 (N_9844,N_2643,N_3072);
nand U9845 (N_9845,N_5744,N_3338);
or U9846 (N_9846,N_208,N_3737);
and U9847 (N_9847,N_2867,N_1820);
nand U9848 (N_9848,N_625,N_5822);
xor U9849 (N_9849,N_4419,N_5818);
nand U9850 (N_9850,N_4174,N_1882);
nand U9851 (N_9851,N_2317,N_5484);
and U9852 (N_9852,N_1916,N_4729);
or U9853 (N_9853,N_4141,N_5202);
or U9854 (N_9854,N_5622,N_672);
and U9855 (N_9855,N_4753,N_3652);
nand U9856 (N_9856,N_3247,N_2025);
xor U9857 (N_9857,N_5196,N_2523);
nand U9858 (N_9858,N_3482,N_3380);
or U9859 (N_9859,N_5723,N_2381);
nand U9860 (N_9860,N_5975,N_311);
or U9861 (N_9861,N_2213,N_2629);
nor U9862 (N_9862,N_5338,N_4184);
and U9863 (N_9863,N_862,N_27);
nand U9864 (N_9864,N_4502,N_3859);
or U9865 (N_9865,N_4535,N_963);
nand U9866 (N_9866,N_5696,N_3181);
nor U9867 (N_9867,N_4541,N_6097);
and U9868 (N_9868,N_3267,N_667);
nand U9869 (N_9869,N_4105,N_2521);
and U9870 (N_9870,N_4976,N_2495);
nor U9871 (N_9871,N_6138,N_3208);
and U9872 (N_9872,N_6064,N_2185);
nor U9873 (N_9873,N_4422,N_649);
and U9874 (N_9874,N_2231,N_4348);
nand U9875 (N_9875,N_2602,N_4496);
or U9876 (N_9876,N_118,N_1449);
or U9877 (N_9877,N_1905,N_4448);
xor U9878 (N_9878,N_5465,N_3271);
xnor U9879 (N_9879,N_3446,N_3175);
nand U9880 (N_9880,N_691,N_319);
or U9881 (N_9881,N_4069,N_257);
xnor U9882 (N_9882,N_1022,N_6162);
or U9883 (N_9883,N_2465,N_523);
and U9884 (N_9884,N_2734,N_5740);
or U9885 (N_9885,N_5948,N_28);
or U9886 (N_9886,N_3339,N_2365);
nor U9887 (N_9887,N_1864,N_2384);
nor U9888 (N_9888,N_1787,N_1366);
nor U9889 (N_9889,N_1961,N_2286);
or U9890 (N_9890,N_2012,N_2323);
nor U9891 (N_9891,N_456,N_6146);
and U9892 (N_9892,N_1622,N_1888);
or U9893 (N_9893,N_3769,N_3875);
nor U9894 (N_9894,N_3719,N_133);
nand U9895 (N_9895,N_1766,N_1120);
nand U9896 (N_9896,N_939,N_1169);
xnor U9897 (N_9897,N_3997,N_1477);
nand U9898 (N_9898,N_3491,N_4492);
or U9899 (N_9899,N_4751,N_5246);
or U9900 (N_9900,N_3350,N_3713);
xor U9901 (N_9901,N_4092,N_1777);
nor U9902 (N_9902,N_617,N_5022);
nor U9903 (N_9903,N_5820,N_5339);
nand U9904 (N_9904,N_972,N_6147);
nor U9905 (N_9905,N_4946,N_4523);
nor U9906 (N_9906,N_4716,N_4158);
and U9907 (N_9907,N_4232,N_3590);
or U9908 (N_9908,N_2521,N_5328);
nand U9909 (N_9909,N_6248,N_5087);
or U9910 (N_9910,N_84,N_3814);
and U9911 (N_9911,N_5587,N_2696);
and U9912 (N_9912,N_4564,N_4415);
nor U9913 (N_9913,N_3399,N_4245);
and U9914 (N_9914,N_1590,N_4145);
and U9915 (N_9915,N_3575,N_425);
nor U9916 (N_9916,N_777,N_4159);
and U9917 (N_9917,N_1780,N_545);
or U9918 (N_9918,N_850,N_1162);
nor U9919 (N_9919,N_4452,N_6043);
or U9920 (N_9920,N_2272,N_185);
nor U9921 (N_9921,N_1805,N_2491);
or U9922 (N_9922,N_1304,N_1469);
nor U9923 (N_9923,N_2460,N_546);
nor U9924 (N_9924,N_1752,N_2160);
nor U9925 (N_9925,N_5762,N_1589);
and U9926 (N_9926,N_3626,N_3744);
or U9927 (N_9927,N_5192,N_2859);
or U9928 (N_9928,N_2697,N_170);
nand U9929 (N_9929,N_4666,N_4870);
nor U9930 (N_9930,N_807,N_713);
and U9931 (N_9931,N_3271,N_4379);
nor U9932 (N_9932,N_1455,N_5469);
nand U9933 (N_9933,N_5629,N_700);
nand U9934 (N_9934,N_2761,N_78);
nand U9935 (N_9935,N_1311,N_2892);
xor U9936 (N_9936,N_6019,N_357);
nor U9937 (N_9937,N_850,N_3800);
nand U9938 (N_9938,N_2249,N_5094);
nor U9939 (N_9939,N_3820,N_1364);
nor U9940 (N_9940,N_1542,N_2846);
nand U9941 (N_9941,N_6108,N_5987);
nand U9942 (N_9942,N_252,N_1271);
or U9943 (N_9943,N_517,N_4213);
nand U9944 (N_9944,N_4293,N_175);
xor U9945 (N_9945,N_3456,N_3798);
or U9946 (N_9946,N_1200,N_4770);
and U9947 (N_9947,N_5526,N_2504);
nand U9948 (N_9948,N_4692,N_2653);
and U9949 (N_9949,N_3099,N_2463);
or U9950 (N_9950,N_3469,N_67);
nand U9951 (N_9951,N_1738,N_1155);
nor U9952 (N_9952,N_1609,N_647);
and U9953 (N_9953,N_4186,N_2546);
and U9954 (N_9954,N_2280,N_5073);
or U9955 (N_9955,N_4302,N_6091);
nor U9956 (N_9956,N_1168,N_1915);
nand U9957 (N_9957,N_4941,N_4263);
and U9958 (N_9958,N_5199,N_138);
and U9959 (N_9959,N_3830,N_4662);
and U9960 (N_9960,N_5425,N_3173);
or U9961 (N_9961,N_2895,N_3765);
and U9962 (N_9962,N_3955,N_2168);
and U9963 (N_9963,N_3136,N_4418);
nor U9964 (N_9964,N_4947,N_2904);
or U9965 (N_9965,N_1806,N_4111);
or U9966 (N_9966,N_345,N_2879);
nor U9967 (N_9967,N_5785,N_4043);
and U9968 (N_9968,N_1896,N_5150);
nand U9969 (N_9969,N_1212,N_4301);
or U9970 (N_9970,N_5942,N_6021);
nor U9971 (N_9971,N_2314,N_5249);
or U9972 (N_9972,N_3871,N_1582);
xor U9973 (N_9973,N_868,N_2512);
nor U9974 (N_9974,N_2703,N_1925);
xor U9975 (N_9975,N_3780,N_231);
nand U9976 (N_9976,N_5180,N_4100);
or U9977 (N_9977,N_4808,N_5734);
nand U9978 (N_9978,N_3985,N_1953);
nand U9979 (N_9979,N_946,N_4504);
nand U9980 (N_9980,N_3871,N_4396);
xnor U9981 (N_9981,N_3029,N_2074);
or U9982 (N_9982,N_4718,N_1389);
xor U9983 (N_9983,N_256,N_1567);
or U9984 (N_9984,N_4873,N_2774);
nor U9985 (N_9985,N_961,N_2258);
nand U9986 (N_9986,N_3750,N_858);
nand U9987 (N_9987,N_4123,N_6244);
and U9988 (N_9988,N_46,N_3908);
xnor U9989 (N_9989,N_3621,N_3079);
nor U9990 (N_9990,N_1890,N_508);
and U9991 (N_9991,N_4741,N_6150);
nor U9992 (N_9992,N_4279,N_739);
or U9993 (N_9993,N_1855,N_1676);
nand U9994 (N_9994,N_3070,N_4327);
xor U9995 (N_9995,N_5101,N_3233);
or U9996 (N_9996,N_5206,N_3095);
or U9997 (N_9997,N_3259,N_5831);
and U9998 (N_9998,N_4944,N_5238);
or U9999 (N_9999,N_3788,N_4265);
or U10000 (N_10000,N_2667,N_3691);
and U10001 (N_10001,N_2092,N_2104);
or U10002 (N_10002,N_1215,N_5601);
nand U10003 (N_10003,N_5085,N_1381);
nand U10004 (N_10004,N_5813,N_1326);
nor U10005 (N_10005,N_137,N_1246);
nor U10006 (N_10006,N_5551,N_1322);
nor U10007 (N_10007,N_4279,N_4854);
nand U10008 (N_10008,N_330,N_1143);
nor U10009 (N_10009,N_4094,N_5787);
nand U10010 (N_10010,N_503,N_2529);
xor U10011 (N_10011,N_767,N_38);
nor U10012 (N_10012,N_1928,N_3186);
nor U10013 (N_10013,N_4790,N_155);
nor U10014 (N_10014,N_3182,N_614);
and U10015 (N_10015,N_4597,N_4173);
nand U10016 (N_10016,N_1816,N_4870);
xor U10017 (N_10017,N_163,N_2195);
or U10018 (N_10018,N_6031,N_4048);
or U10019 (N_10019,N_3573,N_4702);
nand U10020 (N_10020,N_2608,N_3633);
or U10021 (N_10021,N_2418,N_4434);
nor U10022 (N_10022,N_4748,N_165);
and U10023 (N_10023,N_2075,N_1206);
nor U10024 (N_10024,N_1111,N_1805);
and U10025 (N_10025,N_3345,N_5704);
nand U10026 (N_10026,N_800,N_664);
or U10027 (N_10027,N_1518,N_544);
and U10028 (N_10028,N_3395,N_673);
or U10029 (N_10029,N_2986,N_4172);
or U10030 (N_10030,N_4176,N_799);
nand U10031 (N_10031,N_2650,N_457);
or U10032 (N_10032,N_3489,N_5477);
xor U10033 (N_10033,N_4475,N_5255);
or U10034 (N_10034,N_5318,N_1364);
or U10035 (N_10035,N_575,N_6172);
nand U10036 (N_10036,N_5758,N_180);
nor U10037 (N_10037,N_238,N_5604);
or U10038 (N_10038,N_546,N_4380);
nor U10039 (N_10039,N_3827,N_4606);
nand U10040 (N_10040,N_1444,N_3864);
and U10041 (N_10041,N_117,N_2144);
nor U10042 (N_10042,N_3534,N_3283);
or U10043 (N_10043,N_2804,N_3120);
and U10044 (N_10044,N_3956,N_4446);
nor U10045 (N_10045,N_4462,N_4365);
xor U10046 (N_10046,N_52,N_984);
xnor U10047 (N_10047,N_5037,N_969);
nand U10048 (N_10048,N_2709,N_5025);
nand U10049 (N_10049,N_2243,N_5430);
nor U10050 (N_10050,N_2083,N_3340);
nand U10051 (N_10051,N_4161,N_925);
and U10052 (N_10052,N_3742,N_4710);
nand U10053 (N_10053,N_2659,N_354);
and U10054 (N_10054,N_5756,N_827);
or U10055 (N_10055,N_4336,N_3698);
and U10056 (N_10056,N_124,N_5103);
and U10057 (N_10057,N_579,N_5561);
nand U10058 (N_10058,N_3639,N_1118);
or U10059 (N_10059,N_2282,N_2917);
and U10060 (N_10060,N_4761,N_1532);
or U10061 (N_10061,N_5072,N_6244);
xnor U10062 (N_10062,N_2976,N_59);
and U10063 (N_10063,N_5789,N_5516);
nor U10064 (N_10064,N_5795,N_2118);
and U10065 (N_10065,N_1691,N_2384);
and U10066 (N_10066,N_4644,N_1449);
nor U10067 (N_10067,N_540,N_2401);
and U10068 (N_10068,N_2505,N_3776);
nor U10069 (N_10069,N_5003,N_5664);
xnor U10070 (N_10070,N_921,N_5870);
nand U10071 (N_10071,N_5295,N_3777);
nand U10072 (N_10072,N_1434,N_2600);
nor U10073 (N_10073,N_1861,N_2618);
and U10074 (N_10074,N_4993,N_460);
xor U10075 (N_10075,N_764,N_20);
nand U10076 (N_10076,N_3395,N_4166);
nor U10077 (N_10077,N_6133,N_553);
and U10078 (N_10078,N_3592,N_288);
nand U10079 (N_10079,N_4085,N_359);
and U10080 (N_10080,N_1046,N_1747);
nand U10081 (N_10081,N_824,N_1888);
nand U10082 (N_10082,N_5313,N_3462);
nor U10083 (N_10083,N_795,N_2753);
nand U10084 (N_10084,N_3918,N_3513);
nor U10085 (N_10085,N_4633,N_1850);
nand U10086 (N_10086,N_2754,N_1967);
nor U10087 (N_10087,N_122,N_5041);
xor U10088 (N_10088,N_2495,N_1268);
and U10089 (N_10089,N_3643,N_2040);
nand U10090 (N_10090,N_1443,N_2503);
nor U10091 (N_10091,N_6175,N_3530);
nand U10092 (N_10092,N_5564,N_2618);
or U10093 (N_10093,N_3137,N_6199);
nor U10094 (N_10094,N_1868,N_2071);
or U10095 (N_10095,N_2470,N_2460);
or U10096 (N_10096,N_1043,N_127);
nor U10097 (N_10097,N_5128,N_3893);
or U10098 (N_10098,N_5996,N_6005);
nand U10099 (N_10099,N_3160,N_1597);
nor U10100 (N_10100,N_2296,N_5729);
nand U10101 (N_10101,N_5190,N_2292);
or U10102 (N_10102,N_496,N_79);
nor U10103 (N_10103,N_6176,N_5786);
nor U10104 (N_10104,N_3863,N_3857);
nand U10105 (N_10105,N_945,N_2736);
and U10106 (N_10106,N_484,N_4337);
nand U10107 (N_10107,N_3981,N_2467);
or U10108 (N_10108,N_3929,N_3121);
or U10109 (N_10109,N_455,N_4739);
xor U10110 (N_10110,N_216,N_276);
nand U10111 (N_10111,N_3807,N_4225);
or U10112 (N_10112,N_636,N_2993);
and U10113 (N_10113,N_577,N_6237);
or U10114 (N_10114,N_4963,N_2468);
and U10115 (N_10115,N_1405,N_5609);
nor U10116 (N_10116,N_4414,N_5046);
and U10117 (N_10117,N_1213,N_2573);
nor U10118 (N_10118,N_1445,N_3573);
or U10119 (N_10119,N_5173,N_1853);
nor U10120 (N_10120,N_6085,N_4786);
and U10121 (N_10121,N_4189,N_4406);
and U10122 (N_10122,N_5364,N_3722);
nand U10123 (N_10123,N_239,N_4524);
xor U10124 (N_10124,N_1031,N_2165);
and U10125 (N_10125,N_4157,N_3136);
nor U10126 (N_10126,N_2005,N_2755);
or U10127 (N_10127,N_4651,N_2490);
and U10128 (N_10128,N_6143,N_1177);
and U10129 (N_10129,N_302,N_873);
and U10130 (N_10130,N_236,N_5429);
nor U10131 (N_10131,N_3501,N_3882);
or U10132 (N_10132,N_343,N_2507);
and U10133 (N_10133,N_2352,N_5305);
and U10134 (N_10134,N_6062,N_4949);
nand U10135 (N_10135,N_2233,N_665);
and U10136 (N_10136,N_5448,N_2936);
nand U10137 (N_10137,N_3530,N_4930);
and U10138 (N_10138,N_4979,N_2978);
or U10139 (N_10139,N_5151,N_3037);
nor U10140 (N_10140,N_2733,N_2539);
nor U10141 (N_10141,N_885,N_1096);
nand U10142 (N_10142,N_3824,N_1589);
nand U10143 (N_10143,N_847,N_534);
and U10144 (N_10144,N_1127,N_964);
and U10145 (N_10145,N_39,N_5025);
xor U10146 (N_10146,N_724,N_4759);
nor U10147 (N_10147,N_4496,N_4882);
or U10148 (N_10148,N_5054,N_1172);
nand U10149 (N_10149,N_2301,N_5933);
nor U10150 (N_10150,N_3310,N_3071);
xor U10151 (N_10151,N_1881,N_3178);
nand U10152 (N_10152,N_12,N_4324);
xor U10153 (N_10153,N_2132,N_4001);
nor U10154 (N_10154,N_2850,N_2252);
and U10155 (N_10155,N_585,N_2222);
or U10156 (N_10156,N_2209,N_1643);
nor U10157 (N_10157,N_4860,N_439);
and U10158 (N_10158,N_5087,N_4830);
or U10159 (N_10159,N_286,N_5412);
nand U10160 (N_10160,N_3330,N_4492);
nor U10161 (N_10161,N_4595,N_4436);
xor U10162 (N_10162,N_4171,N_2253);
or U10163 (N_10163,N_3058,N_5296);
and U10164 (N_10164,N_944,N_3446);
or U10165 (N_10165,N_3042,N_3444);
nor U10166 (N_10166,N_6204,N_844);
nand U10167 (N_10167,N_1923,N_1601);
and U10168 (N_10168,N_2284,N_2050);
nor U10169 (N_10169,N_6070,N_1950);
nor U10170 (N_10170,N_5665,N_5361);
xnor U10171 (N_10171,N_3528,N_5154);
xnor U10172 (N_10172,N_4500,N_2804);
nand U10173 (N_10173,N_1536,N_4970);
nor U10174 (N_10174,N_5548,N_1629);
nand U10175 (N_10175,N_1189,N_2003);
or U10176 (N_10176,N_1026,N_149);
nor U10177 (N_10177,N_1440,N_5262);
and U10178 (N_10178,N_2935,N_4701);
and U10179 (N_10179,N_4129,N_5745);
xor U10180 (N_10180,N_4830,N_1728);
or U10181 (N_10181,N_4908,N_3973);
nor U10182 (N_10182,N_5908,N_2822);
or U10183 (N_10183,N_4944,N_289);
and U10184 (N_10184,N_1842,N_857);
and U10185 (N_10185,N_3644,N_2619);
and U10186 (N_10186,N_4961,N_1191);
or U10187 (N_10187,N_1931,N_4646);
and U10188 (N_10188,N_334,N_2791);
and U10189 (N_10189,N_897,N_5591);
nor U10190 (N_10190,N_2769,N_2666);
xnor U10191 (N_10191,N_4111,N_2766);
or U10192 (N_10192,N_5342,N_1264);
and U10193 (N_10193,N_1922,N_3022);
nand U10194 (N_10194,N_2051,N_6207);
xor U10195 (N_10195,N_6182,N_1901);
or U10196 (N_10196,N_404,N_199);
nor U10197 (N_10197,N_3910,N_5383);
or U10198 (N_10198,N_1089,N_3864);
xor U10199 (N_10199,N_1575,N_3926);
nand U10200 (N_10200,N_3659,N_1206);
nand U10201 (N_10201,N_1699,N_5051);
xor U10202 (N_10202,N_6196,N_1763);
nor U10203 (N_10203,N_6129,N_1621);
or U10204 (N_10204,N_2525,N_4057);
or U10205 (N_10205,N_620,N_2616);
or U10206 (N_10206,N_4276,N_5318);
nor U10207 (N_10207,N_1712,N_1648);
and U10208 (N_10208,N_3865,N_6070);
nor U10209 (N_10209,N_1739,N_1115);
nand U10210 (N_10210,N_425,N_5746);
and U10211 (N_10211,N_68,N_3291);
or U10212 (N_10212,N_2059,N_1227);
or U10213 (N_10213,N_5832,N_3257);
and U10214 (N_10214,N_2173,N_2302);
nor U10215 (N_10215,N_1268,N_340);
nand U10216 (N_10216,N_5883,N_5890);
nand U10217 (N_10217,N_1097,N_4113);
nand U10218 (N_10218,N_822,N_982);
or U10219 (N_10219,N_4418,N_2491);
or U10220 (N_10220,N_1391,N_2599);
and U10221 (N_10221,N_655,N_2232);
or U10222 (N_10222,N_787,N_2982);
and U10223 (N_10223,N_2308,N_2701);
nand U10224 (N_10224,N_642,N_2574);
or U10225 (N_10225,N_4143,N_5324);
xor U10226 (N_10226,N_3379,N_2442);
nor U10227 (N_10227,N_1924,N_2517);
nor U10228 (N_10228,N_6062,N_2642);
nor U10229 (N_10229,N_4325,N_2183);
nand U10230 (N_10230,N_5627,N_6027);
and U10231 (N_10231,N_4459,N_3568);
xnor U10232 (N_10232,N_2147,N_470);
and U10233 (N_10233,N_4949,N_2513);
nor U10234 (N_10234,N_5498,N_3821);
or U10235 (N_10235,N_5301,N_5031);
nor U10236 (N_10236,N_4952,N_3302);
nand U10237 (N_10237,N_4089,N_3788);
or U10238 (N_10238,N_931,N_6131);
nand U10239 (N_10239,N_3845,N_3821);
and U10240 (N_10240,N_4451,N_2586);
and U10241 (N_10241,N_3656,N_876);
and U10242 (N_10242,N_4203,N_2464);
and U10243 (N_10243,N_1803,N_3926);
and U10244 (N_10244,N_540,N_5327);
nor U10245 (N_10245,N_5017,N_6210);
and U10246 (N_10246,N_4024,N_1744);
nand U10247 (N_10247,N_1183,N_970);
or U10248 (N_10248,N_4096,N_1342);
nor U10249 (N_10249,N_1537,N_4794);
nand U10250 (N_10250,N_269,N_3482);
or U10251 (N_10251,N_4024,N_3397);
nor U10252 (N_10252,N_822,N_4749);
and U10253 (N_10253,N_2884,N_2205);
xnor U10254 (N_10254,N_522,N_4942);
xor U10255 (N_10255,N_500,N_6027);
or U10256 (N_10256,N_5850,N_2751);
nand U10257 (N_10257,N_3075,N_219);
or U10258 (N_10258,N_88,N_2634);
nand U10259 (N_10259,N_1838,N_29);
or U10260 (N_10260,N_2690,N_4585);
nor U10261 (N_10261,N_4847,N_5636);
and U10262 (N_10262,N_4700,N_3879);
and U10263 (N_10263,N_5685,N_1750);
nand U10264 (N_10264,N_4104,N_3638);
nand U10265 (N_10265,N_411,N_6143);
nand U10266 (N_10266,N_5892,N_2829);
nand U10267 (N_10267,N_2919,N_700);
nor U10268 (N_10268,N_5907,N_3963);
xor U10269 (N_10269,N_5101,N_4185);
or U10270 (N_10270,N_352,N_1902);
and U10271 (N_10271,N_1599,N_1215);
nor U10272 (N_10272,N_6239,N_4935);
xor U10273 (N_10273,N_5784,N_695);
or U10274 (N_10274,N_4454,N_935);
nand U10275 (N_10275,N_1639,N_2950);
or U10276 (N_10276,N_1233,N_1610);
and U10277 (N_10277,N_5183,N_3074);
and U10278 (N_10278,N_1753,N_1567);
nor U10279 (N_10279,N_4396,N_1235);
or U10280 (N_10280,N_718,N_4553);
or U10281 (N_10281,N_3743,N_4464);
nand U10282 (N_10282,N_3398,N_5316);
nor U10283 (N_10283,N_962,N_4477);
or U10284 (N_10284,N_3144,N_5368);
nor U10285 (N_10285,N_825,N_5082);
nor U10286 (N_10286,N_407,N_3216);
nand U10287 (N_10287,N_4724,N_203);
or U10288 (N_10288,N_5810,N_647);
and U10289 (N_10289,N_1356,N_1228);
nand U10290 (N_10290,N_621,N_866);
nand U10291 (N_10291,N_3742,N_5465);
nor U10292 (N_10292,N_5449,N_39);
nor U10293 (N_10293,N_5639,N_4805);
and U10294 (N_10294,N_6123,N_2274);
and U10295 (N_10295,N_5307,N_1061);
or U10296 (N_10296,N_4745,N_634);
nor U10297 (N_10297,N_1700,N_3245);
nand U10298 (N_10298,N_3643,N_4833);
nand U10299 (N_10299,N_790,N_3596);
xor U10300 (N_10300,N_4150,N_1246);
or U10301 (N_10301,N_2989,N_230);
nor U10302 (N_10302,N_4351,N_3528);
or U10303 (N_10303,N_2942,N_3259);
and U10304 (N_10304,N_225,N_1995);
nor U10305 (N_10305,N_2115,N_2925);
nor U10306 (N_10306,N_595,N_596);
nand U10307 (N_10307,N_1385,N_3081);
nand U10308 (N_10308,N_3466,N_359);
nand U10309 (N_10309,N_868,N_702);
and U10310 (N_10310,N_2509,N_397);
nand U10311 (N_10311,N_1376,N_3691);
nand U10312 (N_10312,N_201,N_2753);
xnor U10313 (N_10313,N_3567,N_972);
and U10314 (N_10314,N_6235,N_4919);
nor U10315 (N_10315,N_5769,N_2027);
nand U10316 (N_10316,N_1366,N_1674);
nor U10317 (N_10317,N_8,N_2260);
or U10318 (N_10318,N_4156,N_2762);
xnor U10319 (N_10319,N_3339,N_275);
nor U10320 (N_10320,N_2752,N_5390);
or U10321 (N_10321,N_2,N_6123);
nand U10322 (N_10322,N_1049,N_1296);
nor U10323 (N_10323,N_2697,N_291);
or U10324 (N_10324,N_4026,N_95);
and U10325 (N_10325,N_5038,N_2847);
or U10326 (N_10326,N_338,N_3689);
nor U10327 (N_10327,N_2785,N_3055);
xor U10328 (N_10328,N_4922,N_5534);
or U10329 (N_10329,N_5410,N_1737);
xnor U10330 (N_10330,N_2542,N_2389);
xnor U10331 (N_10331,N_5655,N_5535);
nand U10332 (N_10332,N_4653,N_3546);
nand U10333 (N_10333,N_2022,N_1712);
or U10334 (N_10334,N_839,N_1048);
and U10335 (N_10335,N_5510,N_3182);
and U10336 (N_10336,N_1576,N_506);
and U10337 (N_10337,N_1110,N_5649);
and U10338 (N_10338,N_1873,N_4479);
or U10339 (N_10339,N_925,N_5152);
nor U10340 (N_10340,N_2303,N_196);
nor U10341 (N_10341,N_4494,N_3803);
nor U10342 (N_10342,N_2010,N_4185);
or U10343 (N_10343,N_4147,N_3302);
and U10344 (N_10344,N_795,N_148);
nand U10345 (N_10345,N_1303,N_1365);
or U10346 (N_10346,N_733,N_2439);
nor U10347 (N_10347,N_5567,N_5801);
xnor U10348 (N_10348,N_5645,N_3085);
xor U10349 (N_10349,N_549,N_1558);
or U10350 (N_10350,N_702,N_1098);
nand U10351 (N_10351,N_1928,N_1514);
nor U10352 (N_10352,N_1646,N_794);
or U10353 (N_10353,N_2389,N_3043);
or U10354 (N_10354,N_2724,N_1173);
nand U10355 (N_10355,N_4488,N_4142);
xnor U10356 (N_10356,N_5425,N_5502);
nor U10357 (N_10357,N_4159,N_1242);
nand U10358 (N_10358,N_883,N_2470);
nand U10359 (N_10359,N_961,N_6234);
nand U10360 (N_10360,N_1092,N_5537);
and U10361 (N_10361,N_4437,N_2199);
and U10362 (N_10362,N_4070,N_375);
nor U10363 (N_10363,N_2508,N_432);
nor U10364 (N_10364,N_5770,N_2248);
nor U10365 (N_10365,N_3636,N_3045);
nor U10366 (N_10366,N_3297,N_4760);
nand U10367 (N_10367,N_141,N_692);
xnor U10368 (N_10368,N_2193,N_4743);
and U10369 (N_10369,N_1377,N_3298);
nor U10370 (N_10370,N_2518,N_5256);
xnor U10371 (N_10371,N_674,N_3054);
nand U10372 (N_10372,N_3931,N_2882);
nand U10373 (N_10373,N_4044,N_413);
or U10374 (N_10374,N_1199,N_1220);
xor U10375 (N_10375,N_1420,N_481);
nand U10376 (N_10376,N_4935,N_4142);
nand U10377 (N_10377,N_3925,N_462);
nand U10378 (N_10378,N_626,N_2001);
and U10379 (N_10379,N_2707,N_1525);
and U10380 (N_10380,N_5155,N_4790);
nor U10381 (N_10381,N_5473,N_3459);
and U10382 (N_10382,N_451,N_4891);
or U10383 (N_10383,N_1755,N_3491);
nand U10384 (N_10384,N_712,N_5403);
nand U10385 (N_10385,N_6119,N_1926);
nand U10386 (N_10386,N_6019,N_5055);
nor U10387 (N_10387,N_6212,N_881);
nor U10388 (N_10388,N_5184,N_4707);
nand U10389 (N_10389,N_3549,N_1233);
and U10390 (N_10390,N_5344,N_5438);
nor U10391 (N_10391,N_1260,N_2972);
and U10392 (N_10392,N_5505,N_2184);
and U10393 (N_10393,N_1807,N_5841);
or U10394 (N_10394,N_5041,N_1201);
and U10395 (N_10395,N_2103,N_23);
nand U10396 (N_10396,N_1673,N_4283);
and U10397 (N_10397,N_3580,N_3569);
and U10398 (N_10398,N_5325,N_5218);
or U10399 (N_10399,N_3781,N_801);
nor U10400 (N_10400,N_5741,N_3865);
nand U10401 (N_10401,N_3699,N_600);
xnor U10402 (N_10402,N_938,N_544);
and U10403 (N_10403,N_1103,N_5400);
and U10404 (N_10404,N_1909,N_191);
nor U10405 (N_10405,N_2916,N_5064);
nand U10406 (N_10406,N_2909,N_2749);
nor U10407 (N_10407,N_2877,N_2315);
xor U10408 (N_10408,N_1377,N_4544);
or U10409 (N_10409,N_5955,N_3879);
or U10410 (N_10410,N_3729,N_325);
or U10411 (N_10411,N_5628,N_3459);
and U10412 (N_10412,N_5857,N_365);
nor U10413 (N_10413,N_4062,N_2013);
and U10414 (N_10414,N_5475,N_3781);
or U10415 (N_10415,N_3474,N_2195);
and U10416 (N_10416,N_2206,N_4897);
nor U10417 (N_10417,N_1373,N_3395);
nor U10418 (N_10418,N_1203,N_5214);
or U10419 (N_10419,N_2865,N_4473);
nor U10420 (N_10420,N_3873,N_2600);
nor U10421 (N_10421,N_1466,N_5308);
and U10422 (N_10422,N_476,N_5381);
nand U10423 (N_10423,N_4229,N_606);
or U10424 (N_10424,N_3388,N_1835);
nor U10425 (N_10425,N_591,N_2701);
nor U10426 (N_10426,N_364,N_2196);
and U10427 (N_10427,N_1031,N_4919);
xor U10428 (N_10428,N_2813,N_6134);
or U10429 (N_10429,N_1554,N_4007);
nor U10430 (N_10430,N_660,N_1438);
xnor U10431 (N_10431,N_1455,N_2486);
or U10432 (N_10432,N_5575,N_2965);
nand U10433 (N_10433,N_4250,N_3130);
nand U10434 (N_10434,N_766,N_5974);
nor U10435 (N_10435,N_4249,N_3073);
xor U10436 (N_10436,N_3406,N_1302);
nor U10437 (N_10437,N_1763,N_991);
and U10438 (N_10438,N_363,N_3613);
nor U10439 (N_10439,N_2030,N_3077);
nand U10440 (N_10440,N_425,N_2489);
nand U10441 (N_10441,N_5394,N_1561);
or U10442 (N_10442,N_360,N_2635);
or U10443 (N_10443,N_3419,N_4090);
nor U10444 (N_10444,N_2276,N_2310);
and U10445 (N_10445,N_1911,N_205);
nand U10446 (N_10446,N_4328,N_438);
nor U10447 (N_10447,N_1959,N_1956);
nor U10448 (N_10448,N_3157,N_2231);
or U10449 (N_10449,N_1560,N_3557);
and U10450 (N_10450,N_407,N_476);
xnor U10451 (N_10451,N_268,N_2894);
nor U10452 (N_10452,N_4194,N_1214);
and U10453 (N_10453,N_3375,N_4980);
nand U10454 (N_10454,N_4294,N_1166);
xnor U10455 (N_10455,N_2076,N_2826);
and U10456 (N_10456,N_6046,N_19);
nor U10457 (N_10457,N_4025,N_5374);
or U10458 (N_10458,N_779,N_5983);
and U10459 (N_10459,N_2707,N_5944);
and U10460 (N_10460,N_1747,N_5807);
and U10461 (N_10461,N_4641,N_232);
nand U10462 (N_10462,N_4586,N_3929);
nand U10463 (N_10463,N_2196,N_3885);
or U10464 (N_10464,N_6190,N_4213);
nand U10465 (N_10465,N_3417,N_4490);
nor U10466 (N_10466,N_6209,N_4652);
xnor U10467 (N_10467,N_569,N_3690);
nor U10468 (N_10468,N_6189,N_1398);
and U10469 (N_10469,N_1946,N_77);
or U10470 (N_10470,N_4540,N_5198);
and U10471 (N_10471,N_1048,N_6118);
or U10472 (N_10472,N_1878,N_3157);
and U10473 (N_10473,N_5171,N_1892);
nor U10474 (N_10474,N_487,N_2959);
xor U10475 (N_10475,N_146,N_371);
nor U10476 (N_10476,N_6008,N_941);
or U10477 (N_10477,N_5969,N_1122);
nand U10478 (N_10478,N_3975,N_4193);
nand U10479 (N_10479,N_4635,N_1311);
or U10480 (N_10480,N_1698,N_2610);
or U10481 (N_10481,N_2556,N_1532);
xnor U10482 (N_10482,N_1673,N_5714);
xnor U10483 (N_10483,N_118,N_3651);
and U10484 (N_10484,N_627,N_2684);
or U10485 (N_10485,N_4792,N_3391);
nand U10486 (N_10486,N_1363,N_5722);
or U10487 (N_10487,N_309,N_2277);
nand U10488 (N_10488,N_942,N_1640);
nor U10489 (N_10489,N_1631,N_6105);
nor U10490 (N_10490,N_4738,N_5943);
xnor U10491 (N_10491,N_3028,N_2661);
xor U10492 (N_10492,N_642,N_1773);
and U10493 (N_10493,N_5917,N_5679);
nand U10494 (N_10494,N_2008,N_5681);
nor U10495 (N_10495,N_2909,N_1061);
and U10496 (N_10496,N_2268,N_2974);
or U10497 (N_10497,N_2337,N_4856);
xor U10498 (N_10498,N_4129,N_1522);
nand U10499 (N_10499,N_4831,N_312);
nand U10500 (N_10500,N_585,N_1701);
xnor U10501 (N_10501,N_4140,N_2426);
and U10502 (N_10502,N_2392,N_776);
nand U10503 (N_10503,N_3999,N_1538);
or U10504 (N_10504,N_224,N_3698);
nand U10505 (N_10505,N_4401,N_5816);
and U10506 (N_10506,N_5479,N_4715);
nand U10507 (N_10507,N_660,N_3198);
or U10508 (N_10508,N_5961,N_5345);
or U10509 (N_10509,N_2464,N_1255);
nor U10510 (N_10510,N_4361,N_5506);
nor U10511 (N_10511,N_6132,N_5163);
nor U10512 (N_10512,N_6098,N_272);
nor U10513 (N_10513,N_5362,N_4958);
and U10514 (N_10514,N_5850,N_4866);
xnor U10515 (N_10515,N_150,N_2864);
and U10516 (N_10516,N_2311,N_4542);
xnor U10517 (N_10517,N_2934,N_161);
nand U10518 (N_10518,N_2673,N_5178);
xnor U10519 (N_10519,N_2396,N_561);
xor U10520 (N_10520,N_1343,N_5896);
or U10521 (N_10521,N_2982,N_2179);
and U10522 (N_10522,N_1252,N_175);
or U10523 (N_10523,N_3197,N_4847);
xnor U10524 (N_10524,N_2122,N_4754);
nand U10525 (N_10525,N_5623,N_2669);
nand U10526 (N_10526,N_5043,N_1456);
or U10527 (N_10527,N_4587,N_141);
or U10528 (N_10528,N_3814,N_6237);
nor U10529 (N_10529,N_3756,N_3003);
nor U10530 (N_10530,N_5934,N_2753);
and U10531 (N_10531,N_3051,N_2450);
or U10532 (N_10532,N_6237,N_380);
nand U10533 (N_10533,N_4304,N_2836);
nand U10534 (N_10534,N_2493,N_4868);
nor U10535 (N_10535,N_217,N_5755);
nor U10536 (N_10536,N_2614,N_1557);
or U10537 (N_10537,N_3469,N_3704);
or U10538 (N_10538,N_3688,N_49);
nor U10539 (N_10539,N_4281,N_3659);
nor U10540 (N_10540,N_4528,N_3298);
nor U10541 (N_10541,N_3124,N_5269);
or U10542 (N_10542,N_6065,N_1085);
and U10543 (N_10543,N_6111,N_4938);
or U10544 (N_10544,N_4299,N_519);
and U10545 (N_10545,N_1485,N_3536);
nand U10546 (N_10546,N_6249,N_380);
and U10547 (N_10547,N_4273,N_269);
or U10548 (N_10548,N_1029,N_3808);
nand U10549 (N_10549,N_2780,N_123);
and U10550 (N_10550,N_3214,N_579);
and U10551 (N_10551,N_5070,N_5564);
and U10552 (N_10552,N_668,N_28);
xnor U10553 (N_10553,N_2918,N_5352);
or U10554 (N_10554,N_1697,N_4428);
nor U10555 (N_10555,N_1004,N_1463);
or U10556 (N_10556,N_1561,N_5096);
nand U10557 (N_10557,N_1943,N_5969);
xnor U10558 (N_10558,N_1228,N_1067);
and U10559 (N_10559,N_2769,N_4394);
nor U10560 (N_10560,N_2414,N_5378);
nand U10561 (N_10561,N_6210,N_3258);
nand U10562 (N_10562,N_5427,N_2233);
and U10563 (N_10563,N_5195,N_5531);
and U10564 (N_10564,N_2795,N_2353);
nor U10565 (N_10565,N_6113,N_4761);
nor U10566 (N_10566,N_4254,N_5961);
and U10567 (N_10567,N_426,N_1872);
nor U10568 (N_10568,N_912,N_701);
nor U10569 (N_10569,N_2496,N_2668);
nor U10570 (N_10570,N_1493,N_2962);
or U10571 (N_10571,N_3139,N_1603);
nand U10572 (N_10572,N_2971,N_3772);
nand U10573 (N_10573,N_827,N_6044);
nand U10574 (N_10574,N_6059,N_4810);
and U10575 (N_10575,N_2779,N_1816);
nor U10576 (N_10576,N_4181,N_4377);
nand U10577 (N_10577,N_4016,N_2547);
or U10578 (N_10578,N_5245,N_5537);
nand U10579 (N_10579,N_1,N_496);
or U10580 (N_10580,N_4331,N_4272);
xnor U10581 (N_10581,N_5811,N_2809);
nand U10582 (N_10582,N_4165,N_4292);
and U10583 (N_10583,N_3264,N_3271);
xnor U10584 (N_10584,N_4467,N_5323);
nand U10585 (N_10585,N_5676,N_5680);
nand U10586 (N_10586,N_3828,N_4535);
and U10587 (N_10587,N_1077,N_3562);
and U10588 (N_10588,N_1282,N_1803);
and U10589 (N_10589,N_5248,N_4956);
nand U10590 (N_10590,N_4160,N_3921);
nand U10591 (N_10591,N_4763,N_5747);
nand U10592 (N_10592,N_5739,N_2408);
xor U10593 (N_10593,N_4519,N_1607);
xor U10594 (N_10594,N_5627,N_4944);
or U10595 (N_10595,N_1294,N_3705);
or U10596 (N_10596,N_2683,N_5355);
and U10597 (N_10597,N_1338,N_5178);
or U10598 (N_10598,N_1343,N_5482);
nand U10599 (N_10599,N_4599,N_4498);
nand U10600 (N_10600,N_872,N_3425);
nor U10601 (N_10601,N_2851,N_1722);
nand U10602 (N_10602,N_959,N_6125);
and U10603 (N_10603,N_470,N_3421);
and U10604 (N_10604,N_2432,N_3500);
nand U10605 (N_10605,N_2847,N_803);
nand U10606 (N_10606,N_5396,N_2238);
xor U10607 (N_10607,N_1449,N_3447);
nand U10608 (N_10608,N_4937,N_5812);
and U10609 (N_10609,N_3644,N_5451);
nor U10610 (N_10610,N_3686,N_2040);
nand U10611 (N_10611,N_2509,N_4413);
nor U10612 (N_10612,N_1322,N_4377);
nor U10613 (N_10613,N_5522,N_1566);
nand U10614 (N_10614,N_3938,N_3732);
nor U10615 (N_10615,N_3260,N_5662);
xnor U10616 (N_10616,N_6054,N_4743);
and U10617 (N_10617,N_3614,N_5652);
or U10618 (N_10618,N_1859,N_4588);
nor U10619 (N_10619,N_5609,N_3803);
nand U10620 (N_10620,N_990,N_1959);
and U10621 (N_10621,N_3804,N_3949);
xnor U10622 (N_10622,N_2511,N_2888);
nand U10623 (N_10623,N_1614,N_5363);
nand U10624 (N_10624,N_5716,N_1888);
or U10625 (N_10625,N_4115,N_3523);
and U10626 (N_10626,N_526,N_3634);
nor U10627 (N_10627,N_3435,N_1535);
or U10628 (N_10628,N_2849,N_3519);
or U10629 (N_10629,N_6100,N_2599);
and U10630 (N_10630,N_3739,N_599);
or U10631 (N_10631,N_2023,N_2359);
or U10632 (N_10632,N_388,N_153);
or U10633 (N_10633,N_1435,N_5871);
nand U10634 (N_10634,N_4938,N_3247);
or U10635 (N_10635,N_4590,N_3957);
and U10636 (N_10636,N_1137,N_4667);
and U10637 (N_10637,N_5315,N_54);
or U10638 (N_10638,N_4599,N_985);
or U10639 (N_10639,N_1602,N_2334);
nand U10640 (N_10640,N_4942,N_115);
xor U10641 (N_10641,N_5257,N_2425);
or U10642 (N_10642,N_1068,N_1180);
nor U10643 (N_10643,N_4127,N_3442);
nand U10644 (N_10644,N_1878,N_1874);
and U10645 (N_10645,N_5168,N_5614);
nand U10646 (N_10646,N_5489,N_4074);
nand U10647 (N_10647,N_2478,N_3138);
nor U10648 (N_10648,N_2744,N_132);
or U10649 (N_10649,N_3751,N_3322);
or U10650 (N_10650,N_5176,N_986);
and U10651 (N_10651,N_1342,N_1932);
xor U10652 (N_10652,N_2990,N_2549);
nor U10653 (N_10653,N_4398,N_1614);
or U10654 (N_10654,N_436,N_2828);
xnor U10655 (N_10655,N_534,N_769);
or U10656 (N_10656,N_4083,N_1938);
nand U10657 (N_10657,N_3077,N_1592);
nor U10658 (N_10658,N_3434,N_2179);
and U10659 (N_10659,N_1700,N_4505);
nand U10660 (N_10660,N_306,N_57);
nand U10661 (N_10661,N_5032,N_3775);
and U10662 (N_10662,N_1610,N_1950);
and U10663 (N_10663,N_2837,N_215);
and U10664 (N_10664,N_1305,N_3449);
nand U10665 (N_10665,N_1998,N_200);
and U10666 (N_10666,N_6235,N_5538);
xnor U10667 (N_10667,N_3427,N_5394);
nand U10668 (N_10668,N_4794,N_3684);
and U10669 (N_10669,N_4086,N_1132);
nand U10670 (N_10670,N_1087,N_5338);
nor U10671 (N_10671,N_668,N_3371);
or U10672 (N_10672,N_4451,N_4790);
or U10673 (N_10673,N_3464,N_1498);
xor U10674 (N_10674,N_3065,N_1210);
and U10675 (N_10675,N_5677,N_550);
and U10676 (N_10676,N_4571,N_2157);
and U10677 (N_10677,N_855,N_2684);
xnor U10678 (N_10678,N_2775,N_6077);
xnor U10679 (N_10679,N_3543,N_2422);
nor U10680 (N_10680,N_1334,N_573);
nor U10681 (N_10681,N_1076,N_5214);
or U10682 (N_10682,N_3387,N_2290);
xor U10683 (N_10683,N_3926,N_4686);
or U10684 (N_10684,N_749,N_4558);
nand U10685 (N_10685,N_2678,N_1850);
nor U10686 (N_10686,N_5106,N_2485);
nand U10687 (N_10687,N_5943,N_4582);
and U10688 (N_10688,N_4875,N_1974);
and U10689 (N_10689,N_1195,N_2994);
nand U10690 (N_10690,N_6009,N_5375);
nor U10691 (N_10691,N_4623,N_869);
or U10692 (N_10692,N_413,N_4916);
nand U10693 (N_10693,N_3098,N_3741);
xnor U10694 (N_10694,N_2702,N_939);
and U10695 (N_10695,N_2516,N_5107);
or U10696 (N_10696,N_3851,N_5558);
or U10697 (N_10697,N_5924,N_3898);
and U10698 (N_10698,N_395,N_1234);
nand U10699 (N_10699,N_3587,N_5288);
xor U10700 (N_10700,N_542,N_2342);
nor U10701 (N_10701,N_601,N_4725);
or U10702 (N_10702,N_4822,N_1231);
xor U10703 (N_10703,N_674,N_3502);
nor U10704 (N_10704,N_1669,N_499);
and U10705 (N_10705,N_5724,N_839);
nor U10706 (N_10706,N_242,N_3014);
nor U10707 (N_10707,N_378,N_3627);
or U10708 (N_10708,N_4921,N_913);
or U10709 (N_10709,N_209,N_1126);
nand U10710 (N_10710,N_3094,N_1795);
xnor U10711 (N_10711,N_2575,N_198);
nand U10712 (N_10712,N_1608,N_1859);
and U10713 (N_10713,N_3949,N_2476);
or U10714 (N_10714,N_3032,N_1998);
nor U10715 (N_10715,N_773,N_5443);
and U10716 (N_10716,N_3143,N_1650);
nor U10717 (N_10717,N_5084,N_5228);
or U10718 (N_10718,N_2355,N_1451);
nor U10719 (N_10719,N_5572,N_1778);
or U10720 (N_10720,N_439,N_2558);
nand U10721 (N_10721,N_249,N_2154);
nor U10722 (N_10722,N_1076,N_2812);
nand U10723 (N_10723,N_2594,N_2046);
or U10724 (N_10724,N_2899,N_2516);
or U10725 (N_10725,N_4226,N_2583);
nor U10726 (N_10726,N_5882,N_1486);
nand U10727 (N_10727,N_1230,N_62);
nand U10728 (N_10728,N_2542,N_933);
and U10729 (N_10729,N_5733,N_2448);
nand U10730 (N_10730,N_414,N_4935);
nand U10731 (N_10731,N_3674,N_4393);
xor U10732 (N_10732,N_5588,N_4527);
nor U10733 (N_10733,N_2488,N_2212);
nor U10734 (N_10734,N_1555,N_426);
xnor U10735 (N_10735,N_758,N_3991);
and U10736 (N_10736,N_1693,N_6111);
and U10737 (N_10737,N_622,N_4458);
nand U10738 (N_10738,N_5467,N_318);
and U10739 (N_10739,N_4844,N_4243);
and U10740 (N_10740,N_3870,N_2151);
nor U10741 (N_10741,N_4259,N_868);
and U10742 (N_10742,N_3136,N_648);
xnor U10743 (N_10743,N_665,N_4674);
nand U10744 (N_10744,N_5093,N_495);
xnor U10745 (N_10745,N_1805,N_1622);
or U10746 (N_10746,N_2815,N_328);
nand U10747 (N_10747,N_2030,N_674);
or U10748 (N_10748,N_962,N_2755);
or U10749 (N_10749,N_3804,N_1937);
nand U10750 (N_10750,N_4342,N_4507);
nand U10751 (N_10751,N_1706,N_3987);
and U10752 (N_10752,N_5080,N_4228);
nand U10753 (N_10753,N_948,N_47);
nand U10754 (N_10754,N_1525,N_2443);
or U10755 (N_10755,N_6034,N_1038);
nor U10756 (N_10756,N_4363,N_5563);
and U10757 (N_10757,N_2780,N_2868);
nand U10758 (N_10758,N_1383,N_1148);
or U10759 (N_10759,N_4916,N_1145);
or U10760 (N_10760,N_1074,N_5850);
nand U10761 (N_10761,N_1319,N_2423);
nor U10762 (N_10762,N_399,N_2013);
nor U10763 (N_10763,N_889,N_1696);
nor U10764 (N_10764,N_5824,N_5108);
nand U10765 (N_10765,N_3130,N_3228);
nor U10766 (N_10766,N_2620,N_5960);
and U10767 (N_10767,N_6129,N_4648);
and U10768 (N_10768,N_5752,N_89);
nor U10769 (N_10769,N_5910,N_1104);
and U10770 (N_10770,N_237,N_4975);
and U10771 (N_10771,N_4767,N_5990);
or U10772 (N_10772,N_5210,N_4221);
nand U10773 (N_10773,N_145,N_1184);
nand U10774 (N_10774,N_298,N_819);
nor U10775 (N_10775,N_5723,N_3925);
and U10776 (N_10776,N_843,N_2973);
nand U10777 (N_10777,N_4756,N_4213);
or U10778 (N_10778,N_740,N_926);
or U10779 (N_10779,N_3407,N_5055);
nand U10780 (N_10780,N_3878,N_256);
or U10781 (N_10781,N_5800,N_2113);
xnor U10782 (N_10782,N_4057,N_1825);
nor U10783 (N_10783,N_4995,N_4323);
xnor U10784 (N_10784,N_1007,N_1610);
nor U10785 (N_10785,N_1346,N_5811);
and U10786 (N_10786,N_1636,N_5114);
and U10787 (N_10787,N_2238,N_5246);
xor U10788 (N_10788,N_2451,N_5888);
and U10789 (N_10789,N_641,N_5111);
nand U10790 (N_10790,N_4426,N_5165);
nand U10791 (N_10791,N_5811,N_624);
nor U10792 (N_10792,N_4373,N_929);
nand U10793 (N_10793,N_4417,N_1719);
nand U10794 (N_10794,N_133,N_1669);
or U10795 (N_10795,N_557,N_3456);
xor U10796 (N_10796,N_6168,N_5568);
nand U10797 (N_10797,N_5875,N_2357);
or U10798 (N_10798,N_3088,N_5293);
nand U10799 (N_10799,N_407,N_2954);
nand U10800 (N_10800,N_2195,N_5233);
nor U10801 (N_10801,N_2395,N_3849);
or U10802 (N_10802,N_5786,N_534);
xor U10803 (N_10803,N_1039,N_2200);
or U10804 (N_10804,N_3387,N_5970);
nand U10805 (N_10805,N_4185,N_5726);
nor U10806 (N_10806,N_5455,N_4081);
and U10807 (N_10807,N_14,N_5090);
nor U10808 (N_10808,N_3054,N_3990);
or U10809 (N_10809,N_4478,N_6080);
and U10810 (N_10810,N_2776,N_693);
and U10811 (N_10811,N_2052,N_4414);
or U10812 (N_10812,N_1149,N_1066);
and U10813 (N_10813,N_1936,N_3398);
or U10814 (N_10814,N_5238,N_5985);
and U10815 (N_10815,N_81,N_1199);
and U10816 (N_10816,N_4697,N_1228);
nor U10817 (N_10817,N_5995,N_4774);
or U10818 (N_10818,N_3888,N_4441);
or U10819 (N_10819,N_6087,N_4706);
and U10820 (N_10820,N_5062,N_5043);
and U10821 (N_10821,N_4453,N_1302);
or U10822 (N_10822,N_1567,N_218);
nor U10823 (N_10823,N_5907,N_1377);
nor U10824 (N_10824,N_1933,N_2780);
nand U10825 (N_10825,N_2501,N_3130);
or U10826 (N_10826,N_3760,N_2057);
nand U10827 (N_10827,N_4291,N_1164);
nor U10828 (N_10828,N_3460,N_2136);
and U10829 (N_10829,N_5178,N_2140);
nand U10830 (N_10830,N_5056,N_1267);
or U10831 (N_10831,N_722,N_4637);
xor U10832 (N_10832,N_939,N_1016);
or U10833 (N_10833,N_4065,N_2658);
and U10834 (N_10834,N_75,N_5367);
xnor U10835 (N_10835,N_5090,N_1962);
xnor U10836 (N_10836,N_1263,N_3314);
or U10837 (N_10837,N_2307,N_2377);
or U10838 (N_10838,N_3702,N_1786);
or U10839 (N_10839,N_4414,N_5292);
xor U10840 (N_10840,N_1562,N_5479);
nor U10841 (N_10841,N_311,N_4527);
or U10842 (N_10842,N_5456,N_3688);
and U10843 (N_10843,N_2283,N_4625);
and U10844 (N_10844,N_798,N_1058);
nor U10845 (N_10845,N_3999,N_3000);
xnor U10846 (N_10846,N_4264,N_4309);
nor U10847 (N_10847,N_6079,N_2286);
nor U10848 (N_10848,N_1423,N_5678);
or U10849 (N_10849,N_1532,N_4721);
nor U10850 (N_10850,N_5530,N_3832);
or U10851 (N_10851,N_5814,N_4437);
nor U10852 (N_10852,N_6141,N_449);
nand U10853 (N_10853,N_3226,N_3838);
nor U10854 (N_10854,N_3080,N_5058);
and U10855 (N_10855,N_4629,N_3933);
or U10856 (N_10856,N_1025,N_4933);
xnor U10857 (N_10857,N_4241,N_4215);
nand U10858 (N_10858,N_2829,N_1837);
nor U10859 (N_10859,N_3701,N_4286);
nor U10860 (N_10860,N_1716,N_5817);
and U10861 (N_10861,N_4569,N_1595);
or U10862 (N_10862,N_5854,N_491);
nor U10863 (N_10863,N_896,N_4876);
nor U10864 (N_10864,N_3856,N_348);
nand U10865 (N_10865,N_4584,N_3073);
nand U10866 (N_10866,N_5246,N_4803);
nor U10867 (N_10867,N_3397,N_3089);
and U10868 (N_10868,N_5940,N_4818);
and U10869 (N_10869,N_2470,N_2190);
nor U10870 (N_10870,N_2979,N_5870);
and U10871 (N_10871,N_3105,N_5394);
or U10872 (N_10872,N_4200,N_3704);
nand U10873 (N_10873,N_5857,N_4910);
and U10874 (N_10874,N_3793,N_3318);
nor U10875 (N_10875,N_674,N_5038);
and U10876 (N_10876,N_5847,N_6114);
nand U10877 (N_10877,N_1353,N_4119);
or U10878 (N_10878,N_28,N_1308);
and U10879 (N_10879,N_2014,N_5371);
and U10880 (N_10880,N_3192,N_569);
nand U10881 (N_10881,N_6117,N_2598);
nand U10882 (N_10882,N_5365,N_3286);
or U10883 (N_10883,N_1833,N_2132);
nand U10884 (N_10884,N_465,N_2161);
nor U10885 (N_10885,N_1275,N_6216);
xor U10886 (N_10886,N_2858,N_1424);
or U10887 (N_10887,N_5742,N_5408);
nand U10888 (N_10888,N_1828,N_3128);
nor U10889 (N_10889,N_3239,N_5859);
nand U10890 (N_10890,N_3814,N_3369);
nand U10891 (N_10891,N_4647,N_2507);
nand U10892 (N_10892,N_1051,N_1034);
xor U10893 (N_10893,N_2161,N_5051);
or U10894 (N_10894,N_1485,N_3368);
nand U10895 (N_10895,N_4945,N_1354);
and U10896 (N_10896,N_1758,N_408);
xnor U10897 (N_10897,N_5281,N_4575);
nand U10898 (N_10898,N_800,N_456);
or U10899 (N_10899,N_3918,N_2955);
nor U10900 (N_10900,N_3397,N_894);
or U10901 (N_10901,N_2965,N_3009);
and U10902 (N_10902,N_3113,N_320);
nand U10903 (N_10903,N_1400,N_4658);
nor U10904 (N_10904,N_2368,N_821);
nand U10905 (N_10905,N_291,N_3619);
or U10906 (N_10906,N_4875,N_705);
xnor U10907 (N_10907,N_5078,N_1037);
and U10908 (N_10908,N_2673,N_2530);
and U10909 (N_10909,N_3456,N_591);
nand U10910 (N_10910,N_4049,N_3320);
nand U10911 (N_10911,N_3446,N_2063);
xor U10912 (N_10912,N_2775,N_4849);
or U10913 (N_10913,N_142,N_403);
xor U10914 (N_10914,N_3992,N_2334);
nor U10915 (N_10915,N_417,N_2721);
nor U10916 (N_10916,N_541,N_2710);
or U10917 (N_10917,N_5153,N_4626);
nor U10918 (N_10918,N_5145,N_1296);
or U10919 (N_10919,N_2880,N_3589);
and U10920 (N_10920,N_2388,N_1456);
nand U10921 (N_10921,N_3655,N_3359);
nand U10922 (N_10922,N_2792,N_5781);
nand U10923 (N_10923,N_1545,N_5031);
nor U10924 (N_10924,N_1678,N_1027);
xnor U10925 (N_10925,N_3267,N_2480);
or U10926 (N_10926,N_1718,N_2591);
and U10927 (N_10927,N_625,N_4939);
nand U10928 (N_10928,N_1113,N_1517);
nand U10929 (N_10929,N_3526,N_4391);
or U10930 (N_10930,N_6118,N_5834);
nand U10931 (N_10931,N_537,N_4295);
or U10932 (N_10932,N_3280,N_5539);
xor U10933 (N_10933,N_3012,N_5381);
and U10934 (N_10934,N_214,N_1540);
nand U10935 (N_10935,N_63,N_6203);
and U10936 (N_10936,N_5642,N_6056);
nor U10937 (N_10937,N_5008,N_3794);
or U10938 (N_10938,N_5840,N_1265);
nand U10939 (N_10939,N_3816,N_2534);
and U10940 (N_10940,N_5616,N_3466);
and U10941 (N_10941,N_109,N_5179);
nor U10942 (N_10942,N_2199,N_5456);
nand U10943 (N_10943,N_1544,N_1926);
xor U10944 (N_10944,N_2075,N_6017);
or U10945 (N_10945,N_1583,N_5665);
and U10946 (N_10946,N_1440,N_991);
or U10947 (N_10947,N_3866,N_1085);
xor U10948 (N_10948,N_2801,N_3362);
xnor U10949 (N_10949,N_1138,N_5781);
nor U10950 (N_10950,N_4939,N_1863);
and U10951 (N_10951,N_407,N_3660);
xor U10952 (N_10952,N_2113,N_6146);
xor U10953 (N_10953,N_1672,N_3539);
and U10954 (N_10954,N_4839,N_4808);
and U10955 (N_10955,N_4081,N_701);
and U10956 (N_10956,N_2406,N_3439);
xor U10957 (N_10957,N_4860,N_149);
xor U10958 (N_10958,N_2286,N_1898);
nor U10959 (N_10959,N_1945,N_2691);
nand U10960 (N_10960,N_4872,N_324);
or U10961 (N_10961,N_1096,N_836);
nor U10962 (N_10962,N_4799,N_2706);
or U10963 (N_10963,N_3155,N_5641);
and U10964 (N_10964,N_2979,N_3471);
and U10965 (N_10965,N_1859,N_4245);
nand U10966 (N_10966,N_2007,N_6090);
nand U10967 (N_10967,N_3687,N_6107);
nor U10968 (N_10968,N_4289,N_3938);
nor U10969 (N_10969,N_5073,N_6021);
or U10970 (N_10970,N_1344,N_2499);
and U10971 (N_10971,N_679,N_978);
and U10972 (N_10972,N_5586,N_459);
xnor U10973 (N_10973,N_5404,N_5238);
and U10974 (N_10974,N_3766,N_3715);
and U10975 (N_10975,N_5680,N_3236);
nand U10976 (N_10976,N_5434,N_3611);
xnor U10977 (N_10977,N_3409,N_3990);
nor U10978 (N_10978,N_3840,N_5877);
xor U10979 (N_10979,N_2265,N_5837);
or U10980 (N_10980,N_5633,N_421);
nand U10981 (N_10981,N_2380,N_1070);
nand U10982 (N_10982,N_4525,N_1236);
xor U10983 (N_10983,N_2181,N_3356);
nand U10984 (N_10984,N_592,N_4281);
and U10985 (N_10985,N_4892,N_2444);
and U10986 (N_10986,N_6023,N_2735);
nor U10987 (N_10987,N_395,N_4501);
nand U10988 (N_10988,N_840,N_2712);
nor U10989 (N_10989,N_2444,N_723);
nor U10990 (N_10990,N_5642,N_1710);
or U10991 (N_10991,N_5806,N_5069);
nand U10992 (N_10992,N_4409,N_2639);
and U10993 (N_10993,N_1847,N_5903);
or U10994 (N_10994,N_4205,N_1186);
and U10995 (N_10995,N_2803,N_783);
and U10996 (N_10996,N_5661,N_309);
nor U10997 (N_10997,N_3603,N_2852);
or U10998 (N_10998,N_5595,N_4338);
nor U10999 (N_10999,N_2750,N_231);
nand U11000 (N_11000,N_3817,N_5663);
or U11001 (N_11001,N_800,N_2260);
nor U11002 (N_11002,N_846,N_5125);
xnor U11003 (N_11003,N_4932,N_3487);
nor U11004 (N_11004,N_2697,N_3258);
and U11005 (N_11005,N_4162,N_5889);
nand U11006 (N_11006,N_3675,N_34);
nand U11007 (N_11007,N_3058,N_3847);
nor U11008 (N_11008,N_2446,N_723);
nand U11009 (N_11009,N_2978,N_4116);
nor U11010 (N_11010,N_1173,N_1968);
nand U11011 (N_11011,N_2738,N_2920);
nor U11012 (N_11012,N_4240,N_736);
and U11013 (N_11013,N_5947,N_2195);
and U11014 (N_11014,N_3190,N_4110);
nand U11015 (N_11015,N_2313,N_5272);
or U11016 (N_11016,N_4621,N_5762);
and U11017 (N_11017,N_1221,N_5625);
nand U11018 (N_11018,N_1106,N_5530);
nor U11019 (N_11019,N_1205,N_811);
or U11020 (N_11020,N_4281,N_5122);
nor U11021 (N_11021,N_755,N_4557);
nand U11022 (N_11022,N_5363,N_2135);
or U11023 (N_11023,N_1727,N_2236);
and U11024 (N_11024,N_2,N_2815);
or U11025 (N_11025,N_5876,N_4568);
and U11026 (N_11026,N_6025,N_906);
and U11027 (N_11027,N_6169,N_1155);
xor U11028 (N_11028,N_4539,N_2621);
nor U11029 (N_11029,N_2333,N_3061);
or U11030 (N_11030,N_1369,N_344);
xnor U11031 (N_11031,N_539,N_1500);
and U11032 (N_11032,N_3204,N_1166);
nand U11033 (N_11033,N_5594,N_3863);
or U11034 (N_11034,N_2669,N_673);
and U11035 (N_11035,N_2020,N_674);
or U11036 (N_11036,N_3642,N_2141);
and U11037 (N_11037,N_3018,N_3706);
nand U11038 (N_11038,N_941,N_2720);
and U11039 (N_11039,N_3990,N_1085);
and U11040 (N_11040,N_806,N_2724);
nor U11041 (N_11041,N_597,N_4325);
nand U11042 (N_11042,N_736,N_1452);
xor U11043 (N_11043,N_6067,N_2773);
nor U11044 (N_11044,N_5251,N_618);
and U11045 (N_11045,N_5222,N_1529);
or U11046 (N_11046,N_343,N_2720);
and U11047 (N_11047,N_5053,N_1883);
or U11048 (N_11048,N_399,N_4359);
xnor U11049 (N_11049,N_4467,N_6227);
or U11050 (N_11050,N_5718,N_3600);
xnor U11051 (N_11051,N_2518,N_4918);
or U11052 (N_11052,N_4488,N_4722);
xnor U11053 (N_11053,N_4753,N_1975);
or U11054 (N_11054,N_2783,N_3339);
nand U11055 (N_11055,N_529,N_1206);
nor U11056 (N_11056,N_1937,N_345);
and U11057 (N_11057,N_3892,N_6205);
or U11058 (N_11058,N_263,N_6011);
and U11059 (N_11059,N_2707,N_836);
nand U11060 (N_11060,N_2627,N_3752);
and U11061 (N_11061,N_1025,N_1909);
and U11062 (N_11062,N_1380,N_583);
or U11063 (N_11063,N_3669,N_3179);
or U11064 (N_11064,N_3104,N_5992);
and U11065 (N_11065,N_3527,N_30);
and U11066 (N_11066,N_361,N_1301);
and U11067 (N_11067,N_1140,N_4548);
nor U11068 (N_11068,N_4134,N_605);
and U11069 (N_11069,N_4996,N_2581);
nand U11070 (N_11070,N_1900,N_3736);
nor U11071 (N_11071,N_5993,N_814);
nor U11072 (N_11072,N_1175,N_646);
nand U11073 (N_11073,N_5910,N_480);
nand U11074 (N_11074,N_887,N_3425);
nor U11075 (N_11075,N_1034,N_658);
nand U11076 (N_11076,N_1602,N_2118);
or U11077 (N_11077,N_1208,N_2009);
and U11078 (N_11078,N_5205,N_21);
and U11079 (N_11079,N_1175,N_1954);
nor U11080 (N_11080,N_5787,N_4090);
and U11081 (N_11081,N_862,N_1336);
and U11082 (N_11082,N_2014,N_1400);
nor U11083 (N_11083,N_5747,N_4686);
or U11084 (N_11084,N_2668,N_4573);
or U11085 (N_11085,N_4097,N_3313);
nand U11086 (N_11086,N_4574,N_3104);
xnor U11087 (N_11087,N_284,N_3689);
nand U11088 (N_11088,N_6211,N_784);
nand U11089 (N_11089,N_645,N_3516);
or U11090 (N_11090,N_955,N_3815);
nor U11091 (N_11091,N_5005,N_2944);
and U11092 (N_11092,N_1017,N_2463);
nand U11093 (N_11093,N_3112,N_3339);
nor U11094 (N_11094,N_2143,N_3096);
and U11095 (N_11095,N_5280,N_502);
or U11096 (N_11096,N_1430,N_1777);
or U11097 (N_11097,N_4772,N_535);
xor U11098 (N_11098,N_2140,N_1);
nand U11099 (N_11099,N_409,N_157);
and U11100 (N_11100,N_1397,N_1517);
nand U11101 (N_11101,N_1470,N_4843);
nand U11102 (N_11102,N_2293,N_5968);
xnor U11103 (N_11103,N_1199,N_5131);
nand U11104 (N_11104,N_4146,N_2987);
nand U11105 (N_11105,N_629,N_3482);
nor U11106 (N_11106,N_2897,N_1544);
nor U11107 (N_11107,N_4204,N_4847);
xor U11108 (N_11108,N_2091,N_3613);
or U11109 (N_11109,N_5364,N_641);
and U11110 (N_11110,N_405,N_4015);
nand U11111 (N_11111,N_3508,N_3177);
nand U11112 (N_11112,N_4279,N_5993);
and U11113 (N_11113,N_4738,N_4381);
and U11114 (N_11114,N_5623,N_865);
nand U11115 (N_11115,N_13,N_1394);
or U11116 (N_11116,N_1631,N_4389);
and U11117 (N_11117,N_2993,N_5014);
nand U11118 (N_11118,N_3039,N_1318);
nor U11119 (N_11119,N_1392,N_4174);
xnor U11120 (N_11120,N_2110,N_1990);
nand U11121 (N_11121,N_1357,N_910);
nor U11122 (N_11122,N_2089,N_1805);
xnor U11123 (N_11123,N_5407,N_6171);
and U11124 (N_11124,N_3193,N_4255);
and U11125 (N_11125,N_598,N_275);
nand U11126 (N_11126,N_431,N_3089);
or U11127 (N_11127,N_2744,N_4687);
and U11128 (N_11128,N_468,N_3377);
nor U11129 (N_11129,N_2078,N_6245);
xor U11130 (N_11130,N_3383,N_1287);
nor U11131 (N_11131,N_4576,N_6008);
nand U11132 (N_11132,N_5281,N_840);
nor U11133 (N_11133,N_3435,N_4202);
and U11134 (N_11134,N_1021,N_5237);
and U11135 (N_11135,N_4483,N_1879);
xnor U11136 (N_11136,N_3804,N_2625);
xor U11137 (N_11137,N_3786,N_1789);
and U11138 (N_11138,N_1203,N_778);
and U11139 (N_11139,N_2804,N_5034);
and U11140 (N_11140,N_4060,N_1119);
and U11141 (N_11141,N_6003,N_2957);
nand U11142 (N_11142,N_4368,N_4131);
and U11143 (N_11143,N_3550,N_5644);
or U11144 (N_11144,N_1880,N_1736);
or U11145 (N_11145,N_4541,N_3925);
nand U11146 (N_11146,N_4208,N_6071);
nor U11147 (N_11147,N_5503,N_2101);
nor U11148 (N_11148,N_4703,N_3817);
or U11149 (N_11149,N_5577,N_2994);
and U11150 (N_11150,N_5766,N_943);
and U11151 (N_11151,N_3034,N_4224);
nor U11152 (N_11152,N_3480,N_97);
nand U11153 (N_11153,N_2603,N_2872);
and U11154 (N_11154,N_627,N_147);
nand U11155 (N_11155,N_1400,N_5413);
or U11156 (N_11156,N_5659,N_5564);
or U11157 (N_11157,N_110,N_2499);
or U11158 (N_11158,N_108,N_4188);
or U11159 (N_11159,N_5429,N_744);
nor U11160 (N_11160,N_5642,N_5719);
and U11161 (N_11161,N_4587,N_1070);
xnor U11162 (N_11162,N_478,N_5354);
nor U11163 (N_11163,N_4897,N_1356);
nor U11164 (N_11164,N_6011,N_126);
and U11165 (N_11165,N_4555,N_4807);
nand U11166 (N_11166,N_2179,N_5294);
nand U11167 (N_11167,N_53,N_4360);
or U11168 (N_11168,N_4654,N_3759);
and U11169 (N_11169,N_1183,N_1923);
nand U11170 (N_11170,N_1321,N_4854);
nand U11171 (N_11171,N_4995,N_3357);
nand U11172 (N_11172,N_5936,N_34);
nor U11173 (N_11173,N_5418,N_1335);
and U11174 (N_11174,N_5425,N_2444);
nor U11175 (N_11175,N_5831,N_1600);
nand U11176 (N_11176,N_3753,N_3414);
nor U11177 (N_11177,N_649,N_315);
nand U11178 (N_11178,N_3002,N_3844);
nor U11179 (N_11179,N_1717,N_3627);
nor U11180 (N_11180,N_3133,N_3274);
nor U11181 (N_11181,N_4048,N_5393);
or U11182 (N_11182,N_1930,N_1996);
and U11183 (N_11183,N_3604,N_1151);
and U11184 (N_11184,N_6193,N_1563);
nor U11185 (N_11185,N_2574,N_590);
nand U11186 (N_11186,N_5658,N_2609);
and U11187 (N_11187,N_4848,N_5446);
nand U11188 (N_11188,N_4117,N_3335);
xnor U11189 (N_11189,N_3723,N_3561);
and U11190 (N_11190,N_1065,N_6035);
or U11191 (N_11191,N_2608,N_4424);
or U11192 (N_11192,N_4437,N_2453);
or U11193 (N_11193,N_973,N_5598);
nand U11194 (N_11194,N_33,N_4555);
and U11195 (N_11195,N_753,N_2681);
nor U11196 (N_11196,N_5535,N_673);
nor U11197 (N_11197,N_805,N_1684);
nand U11198 (N_11198,N_3566,N_4428);
and U11199 (N_11199,N_2022,N_483);
or U11200 (N_11200,N_3070,N_4369);
nor U11201 (N_11201,N_2508,N_1741);
or U11202 (N_11202,N_3723,N_2488);
xor U11203 (N_11203,N_399,N_6017);
nand U11204 (N_11204,N_3755,N_1831);
or U11205 (N_11205,N_2145,N_18);
nor U11206 (N_11206,N_2315,N_3128);
xnor U11207 (N_11207,N_1402,N_4927);
nand U11208 (N_11208,N_922,N_5420);
and U11209 (N_11209,N_153,N_4892);
nor U11210 (N_11210,N_376,N_5984);
xnor U11211 (N_11211,N_3937,N_2310);
nand U11212 (N_11212,N_2744,N_2177);
or U11213 (N_11213,N_3280,N_4702);
or U11214 (N_11214,N_3431,N_97);
nor U11215 (N_11215,N_1846,N_14);
xnor U11216 (N_11216,N_3506,N_1564);
or U11217 (N_11217,N_2705,N_4170);
and U11218 (N_11218,N_3676,N_1123);
nor U11219 (N_11219,N_2357,N_235);
nor U11220 (N_11220,N_488,N_5830);
and U11221 (N_11221,N_3466,N_2637);
nand U11222 (N_11222,N_3515,N_3774);
nand U11223 (N_11223,N_2028,N_1857);
nor U11224 (N_11224,N_1813,N_462);
or U11225 (N_11225,N_5007,N_294);
or U11226 (N_11226,N_3406,N_1405);
and U11227 (N_11227,N_1546,N_662);
nor U11228 (N_11228,N_4040,N_292);
or U11229 (N_11229,N_5873,N_94);
or U11230 (N_11230,N_4006,N_1915);
nor U11231 (N_11231,N_1483,N_4089);
and U11232 (N_11232,N_2944,N_2025);
and U11233 (N_11233,N_4587,N_5730);
and U11234 (N_11234,N_5171,N_2172);
nor U11235 (N_11235,N_846,N_5101);
nand U11236 (N_11236,N_1946,N_3583);
nand U11237 (N_11237,N_221,N_6244);
nor U11238 (N_11238,N_845,N_1355);
or U11239 (N_11239,N_6019,N_2973);
xnor U11240 (N_11240,N_3060,N_3905);
or U11241 (N_11241,N_560,N_1106);
xor U11242 (N_11242,N_4101,N_2788);
or U11243 (N_11243,N_3632,N_725);
and U11244 (N_11244,N_5428,N_735);
xnor U11245 (N_11245,N_5679,N_363);
nand U11246 (N_11246,N_2752,N_5863);
and U11247 (N_11247,N_4889,N_1607);
and U11248 (N_11248,N_195,N_4164);
nor U11249 (N_11249,N_3650,N_5107);
and U11250 (N_11250,N_3032,N_2169);
xor U11251 (N_11251,N_62,N_5014);
or U11252 (N_11252,N_2199,N_952);
or U11253 (N_11253,N_6181,N_123);
nand U11254 (N_11254,N_4140,N_121);
xor U11255 (N_11255,N_3436,N_2193);
nand U11256 (N_11256,N_4166,N_1812);
and U11257 (N_11257,N_1209,N_252);
xnor U11258 (N_11258,N_79,N_6038);
nor U11259 (N_11259,N_2286,N_5044);
nor U11260 (N_11260,N_4867,N_5587);
and U11261 (N_11261,N_765,N_2333);
or U11262 (N_11262,N_2899,N_1197);
nor U11263 (N_11263,N_4427,N_2991);
or U11264 (N_11264,N_502,N_1545);
or U11265 (N_11265,N_487,N_257);
nor U11266 (N_11266,N_3521,N_997);
or U11267 (N_11267,N_1263,N_1986);
nor U11268 (N_11268,N_1746,N_1950);
nand U11269 (N_11269,N_131,N_1713);
nand U11270 (N_11270,N_1405,N_1851);
nor U11271 (N_11271,N_4326,N_4190);
and U11272 (N_11272,N_370,N_6133);
and U11273 (N_11273,N_5813,N_3869);
nor U11274 (N_11274,N_4416,N_372);
or U11275 (N_11275,N_3193,N_2753);
and U11276 (N_11276,N_4964,N_2669);
nand U11277 (N_11277,N_1391,N_5108);
nand U11278 (N_11278,N_1638,N_467);
nor U11279 (N_11279,N_5057,N_5502);
or U11280 (N_11280,N_370,N_372);
nor U11281 (N_11281,N_1152,N_222);
and U11282 (N_11282,N_963,N_5433);
and U11283 (N_11283,N_5158,N_762);
nand U11284 (N_11284,N_191,N_1707);
nor U11285 (N_11285,N_2601,N_1715);
and U11286 (N_11286,N_4330,N_3224);
nand U11287 (N_11287,N_3130,N_3123);
xor U11288 (N_11288,N_6032,N_4428);
and U11289 (N_11289,N_1943,N_504);
and U11290 (N_11290,N_2761,N_537);
nand U11291 (N_11291,N_4813,N_1589);
or U11292 (N_11292,N_384,N_5533);
nand U11293 (N_11293,N_1358,N_5840);
or U11294 (N_11294,N_4277,N_4921);
nor U11295 (N_11295,N_4935,N_5721);
nand U11296 (N_11296,N_112,N_4330);
nand U11297 (N_11297,N_1663,N_1167);
or U11298 (N_11298,N_127,N_2559);
nand U11299 (N_11299,N_1053,N_4454);
and U11300 (N_11300,N_988,N_5339);
or U11301 (N_11301,N_2887,N_5911);
xnor U11302 (N_11302,N_5242,N_4942);
and U11303 (N_11303,N_3180,N_5499);
nor U11304 (N_11304,N_1848,N_162);
or U11305 (N_11305,N_5690,N_4557);
nand U11306 (N_11306,N_5503,N_434);
and U11307 (N_11307,N_2161,N_4585);
xor U11308 (N_11308,N_4983,N_4475);
nand U11309 (N_11309,N_1249,N_1574);
nor U11310 (N_11310,N_4251,N_3838);
or U11311 (N_11311,N_1394,N_2228);
and U11312 (N_11312,N_2760,N_773);
and U11313 (N_11313,N_2453,N_4715);
or U11314 (N_11314,N_4066,N_1941);
nand U11315 (N_11315,N_6164,N_222);
or U11316 (N_11316,N_2245,N_658);
xnor U11317 (N_11317,N_5503,N_2224);
or U11318 (N_11318,N_3428,N_4796);
nor U11319 (N_11319,N_5013,N_536);
nand U11320 (N_11320,N_4398,N_3742);
and U11321 (N_11321,N_6035,N_5436);
or U11322 (N_11322,N_1923,N_1536);
and U11323 (N_11323,N_1158,N_510);
nand U11324 (N_11324,N_1091,N_235);
nand U11325 (N_11325,N_1561,N_752);
and U11326 (N_11326,N_4066,N_4882);
and U11327 (N_11327,N_6040,N_1369);
nand U11328 (N_11328,N_2721,N_881);
and U11329 (N_11329,N_5078,N_1951);
nand U11330 (N_11330,N_1243,N_4833);
xnor U11331 (N_11331,N_5769,N_876);
xnor U11332 (N_11332,N_942,N_4165);
or U11333 (N_11333,N_3450,N_6203);
or U11334 (N_11334,N_3884,N_2597);
and U11335 (N_11335,N_2785,N_2848);
nand U11336 (N_11336,N_3394,N_6212);
xnor U11337 (N_11337,N_3793,N_3973);
and U11338 (N_11338,N_1347,N_2852);
nand U11339 (N_11339,N_263,N_239);
xnor U11340 (N_11340,N_94,N_2602);
or U11341 (N_11341,N_3671,N_4857);
nor U11342 (N_11342,N_2789,N_1607);
nand U11343 (N_11343,N_4724,N_320);
or U11344 (N_11344,N_2096,N_1657);
and U11345 (N_11345,N_1437,N_4996);
nor U11346 (N_11346,N_3067,N_2954);
or U11347 (N_11347,N_3126,N_6161);
nor U11348 (N_11348,N_2493,N_4493);
xor U11349 (N_11349,N_2531,N_382);
or U11350 (N_11350,N_2836,N_2579);
and U11351 (N_11351,N_22,N_2612);
or U11352 (N_11352,N_4184,N_6152);
or U11353 (N_11353,N_5071,N_4942);
nor U11354 (N_11354,N_3775,N_3334);
nand U11355 (N_11355,N_4823,N_315);
nand U11356 (N_11356,N_576,N_5714);
nand U11357 (N_11357,N_59,N_1860);
nand U11358 (N_11358,N_4321,N_3327);
nor U11359 (N_11359,N_5305,N_951);
or U11360 (N_11360,N_3953,N_1824);
xor U11361 (N_11361,N_1752,N_2491);
and U11362 (N_11362,N_5618,N_4898);
nand U11363 (N_11363,N_66,N_4488);
and U11364 (N_11364,N_1170,N_1545);
or U11365 (N_11365,N_520,N_1950);
or U11366 (N_11366,N_910,N_4567);
nor U11367 (N_11367,N_3767,N_2018);
xnor U11368 (N_11368,N_423,N_60);
xor U11369 (N_11369,N_1831,N_601);
nand U11370 (N_11370,N_2631,N_4123);
nand U11371 (N_11371,N_6235,N_633);
and U11372 (N_11372,N_4479,N_5972);
nor U11373 (N_11373,N_1618,N_1504);
and U11374 (N_11374,N_2117,N_6185);
or U11375 (N_11375,N_2657,N_1342);
or U11376 (N_11376,N_4222,N_3015);
and U11377 (N_11377,N_5460,N_311);
nor U11378 (N_11378,N_2824,N_6194);
nand U11379 (N_11379,N_5776,N_5942);
or U11380 (N_11380,N_5330,N_1537);
nor U11381 (N_11381,N_4707,N_3525);
or U11382 (N_11382,N_62,N_2388);
xor U11383 (N_11383,N_760,N_3814);
nand U11384 (N_11384,N_5348,N_1402);
nand U11385 (N_11385,N_6170,N_4453);
nor U11386 (N_11386,N_4065,N_438);
and U11387 (N_11387,N_2299,N_5678);
or U11388 (N_11388,N_4273,N_4668);
or U11389 (N_11389,N_5302,N_1546);
and U11390 (N_11390,N_919,N_976);
or U11391 (N_11391,N_3354,N_4549);
nor U11392 (N_11392,N_3715,N_5119);
or U11393 (N_11393,N_4710,N_5064);
nor U11394 (N_11394,N_1137,N_5483);
nor U11395 (N_11395,N_5754,N_1168);
nand U11396 (N_11396,N_3432,N_4313);
or U11397 (N_11397,N_5264,N_2460);
nand U11398 (N_11398,N_2625,N_3083);
or U11399 (N_11399,N_230,N_3839);
and U11400 (N_11400,N_4686,N_4642);
or U11401 (N_11401,N_3205,N_328);
nand U11402 (N_11402,N_3586,N_3344);
xnor U11403 (N_11403,N_915,N_5178);
and U11404 (N_11404,N_4145,N_3321);
nand U11405 (N_11405,N_1539,N_3490);
and U11406 (N_11406,N_5564,N_5646);
or U11407 (N_11407,N_2153,N_2105);
nand U11408 (N_11408,N_973,N_3517);
and U11409 (N_11409,N_3454,N_1844);
nor U11410 (N_11410,N_4783,N_3656);
and U11411 (N_11411,N_2205,N_5164);
or U11412 (N_11412,N_1615,N_2953);
or U11413 (N_11413,N_5107,N_891);
xor U11414 (N_11414,N_4812,N_2467);
or U11415 (N_11415,N_2157,N_6069);
nand U11416 (N_11416,N_2268,N_5819);
nand U11417 (N_11417,N_4893,N_1041);
xnor U11418 (N_11418,N_5148,N_2692);
and U11419 (N_11419,N_2209,N_1343);
nor U11420 (N_11420,N_973,N_1099);
and U11421 (N_11421,N_2408,N_5755);
xor U11422 (N_11422,N_2823,N_4387);
nand U11423 (N_11423,N_1853,N_222);
nand U11424 (N_11424,N_4717,N_3434);
nor U11425 (N_11425,N_5194,N_5288);
nand U11426 (N_11426,N_1983,N_3417);
nor U11427 (N_11427,N_5389,N_3831);
nor U11428 (N_11428,N_4906,N_3890);
xnor U11429 (N_11429,N_743,N_2025);
nand U11430 (N_11430,N_4899,N_590);
and U11431 (N_11431,N_3889,N_1311);
xor U11432 (N_11432,N_4018,N_462);
and U11433 (N_11433,N_4087,N_1903);
nand U11434 (N_11434,N_2570,N_5295);
nor U11435 (N_11435,N_6000,N_5790);
and U11436 (N_11436,N_4428,N_3733);
and U11437 (N_11437,N_3365,N_3823);
and U11438 (N_11438,N_1199,N_1567);
nand U11439 (N_11439,N_4070,N_981);
or U11440 (N_11440,N_1432,N_4248);
nand U11441 (N_11441,N_4833,N_4598);
and U11442 (N_11442,N_3393,N_2849);
xor U11443 (N_11443,N_4462,N_4973);
nand U11444 (N_11444,N_5406,N_5223);
nand U11445 (N_11445,N_5648,N_1427);
xor U11446 (N_11446,N_6141,N_4014);
nand U11447 (N_11447,N_1193,N_3410);
or U11448 (N_11448,N_5095,N_739);
or U11449 (N_11449,N_2512,N_1312);
xnor U11450 (N_11450,N_4195,N_4450);
or U11451 (N_11451,N_912,N_4677);
and U11452 (N_11452,N_3103,N_497);
and U11453 (N_11453,N_3379,N_6005);
nand U11454 (N_11454,N_4759,N_4431);
or U11455 (N_11455,N_3577,N_6111);
nand U11456 (N_11456,N_5870,N_1111);
nor U11457 (N_11457,N_2777,N_2737);
or U11458 (N_11458,N_733,N_4985);
xnor U11459 (N_11459,N_238,N_4396);
nand U11460 (N_11460,N_4030,N_1937);
and U11461 (N_11461,N_2291,N_5499);
nand U11462 (N_11462,N_3190,N_2384);
nor U11463 (N_11463,N_3511,N_176);
nor U11464 (N_11464,N_1680,N_2137);
nor U11465 (N_11465,N_2333,N_220);
nor U11466 (N_11466,N_1115,N_5847);
and U11467 (N_11467,N_3229,N_4059);
nor U11468 (N_11468,N_3793,N_1945);
nor U11469 (N_11469,N_378,N_1357);
or U11470 (N_11470,N_5448,N_6055);
xor U11471 (N_11471,N_2032,N_5086);
or U11472 (N_11472,N_5337,N_5995);
and U11473 (N_11473,N_3737,N_3813);
nor U11474 (N_11474,N_2990,N_1414);
nor U11475 (N_11475,N_2726,N_2662);
xnor U11476 (N_11476,N_850,N_4991);
nor U11477 (N_11477,N_1907,N_3396);
nor U11478 (N_11478,N_4346,N_5786);
or U11479 (N_11479,N_2163,N_2291);
nand U11480 (N_11480,N_2248,N_5648);
and U11481 (N_11481,N_4263,N_261);
and U11482 (N_11482,N_2235,N_763);
nor U11483 (N_11483,N_5375,N_1527);
nand U11484 (N_11484,N_4021,N_5042);
nand U11485 (N_11485,N_5851,N_4710);
or U11486 (N_11486,N_5319,N_5093);
or U11487 (N_11487,N_2929,N_5277);
or U11488 (N_11488,N_5557,N_5194);
and U11489 (N_11489,N_4064,N_4553);
nor U11490 (N_11490,N_1317,N_3660);
and U11491 (N_11491,N_3914,N_1835);
nor U11492 (N_11492,N_2611,N_326);
and U11493 (N_11493,N_5514,N_5221);
and U11494 (N_11494,N_2527,N_1021);
nand U11495 (N_11495,N_6119,N_2424);
or U11496 (N_11496,N_404,N_1300);
nand U11497 (N_11497,N_6125,N_5654);
or U11498 (N_11498,N_4783,N_4460);
and U11499 (N_11499,N_3187,N_932);
and U11500 (N_11500,N_5838,N_5237);
or U11501 (N_11501,N_149,N_3398);
nand U11502 (N_11502,N_2637,N_2913);
or U11503 (N_11503,N_848,N_4904);
nor U11504 (N_11504,N_3686,N_4528);
nand U11505 (N_11505,N_5352,N_2873);
or U11506 (N_11506,N_466,N_4563);
or U11507 (N_11507,N_2469,N_160);
and U11508 (N_11508,N_4845,N_583);
or U11509 (N_11509,N_4770,N_5032);
nor U11510 (N_11510,N_3700,N_737);
nor U11511 (N_11511,N_6182,N_4546);
or U11512 (N_11512,N_356,N_2961);
or U11513 (N_11513,N_3796,N_1196);
or U11514 (N_11514,N_1749,N_4401);
nor U11515 (N_11515,N_57,N_3537);
nor U11516 (N_11516,N_5545,N_6165);
nor U11517 (N_11517,N_4952,N_4590);
nor U11518 (N_11518,N_4071,N_2045);
nand U11519 (N_11519,N_1227,N_3356);
or U11520 (N_11520,N_5105,N_3850);
nor U11521 (N_11521,N_3482,N_3438);
nand U11522 (N_11522,N_5449,N_1204);
nand U11523 (N_11523,N_2554,N_5867);
and U11524 (N_11524,N_768,N_5469);
or U11525 (N_11525,N_4852,N_2283);
and U11526 (N_11526,N_6227,N_81);
nor U11527 (N_11527,N_3777,N_4962);
nor U11528 (N_11528,N_5531,N_5213);
nor U11529 (N_11529,N_3112,N_4847);
nand U11530 (N_11530,N_5402,N_4803);
nand U11531 (N_11531,N_2646,N_4249);
nand U11532 (N_11532,N_1971,N_878);
nor U11533 (N_11533,N_693,N_2964);
nand U11534 (N_11534,N_5670,N_1080);
and U11535 (N_11535,N_1176,N_4874);
nand U11536 (N_11536,N_1502,N_6061);
nand U11537 (N_11537,N_1374,N_960);
and U11538 (N_11538,N_4148,N_5755);
nor U11539 (N_11539,N_2986,N_613);
nor U11540 (N_11540,N_4269,N_3044);
nand U11541 (N_11541,N_3194,N_1926);
nor U11542 (N_11542,N_5180,N_361);
xnor U11543 (N_11543,N_5987,N_3918);
and U11544 (N_11544,N_5072,N_5958);
and U11545 (N_11545,N_5948,N_2137);
nand U11546 (N_11546,N_2830,N_2769);
and U11547 (N_11547,N_5979,N_1117);
and U11548 (N_11548,N_724,N_5606);
nand U11549 (N_11549,N_3880,N_1601);
or U11550 (N_11550,N_217,N_1443);
and U11551 (N_11551,N_5516,N_1689);
nor U11552 (N_11552,N_2945,N_5365);
nand U11553 (N_11553,N_4875,N_5785);
nor U11554 (N_11554,N_1625,N_688);
nand U11555 (N_11555,N_985,N_6133);
nor U11556 (N_11556,N_2907,N_4725);
nor U11557 (N_11557,N_2330,N_6107);
and U11558 (N_11558,N_2263,N_2440);
nor U11559 (N_11559,N_5419,N_4361);
and U11560 (N_11560,N_2397,N_95);
or U11561 (N_11561,N_1673,N_5145);
nand U11562 (N_11562,N_6204,N_3690);
or U11563 (N_11563,N_6120,N_4671);
nand U11564 (N_11564,N_130,N_1428);
nor U11565 (N_11565,N_5007,N_4466);
or U11566 (N_11566,N_3118,N_4378);
nand U11567 (N_11567,N_2225,N_165);
and U11568 (N_11568,N_4746,N_5670);
and U11569 (N_11569,N_5661,N_3186);
nor U11570 (N_11570,N_159,N_5830);
and U11571 (N_11571,N_3365,N_5550);
nand U11572 (N_11572,N_148,N_2155);
nor U11573 (N_11573,N_2487,N_2608);
and U11574 (N_11574,N_4313,N_1764);
nand U11575 (N_11575,N_353,N_1418);
nor U11576 (N_11576,N_3879,N_5357);
nand U11577 (N_11577,N_5943,N_4609);
and U11578 (N_11578,N_129,N_5305);
nor U11579 (N_11579,N_3282,N_1663);
and U11580 (N_11580,N_3929,N_5924);
and U11581 (N_11581,N_421,N_3256);
or U11582 (N_11582,N_2093,N_324);
nor U11583 (N_11583,N_4912,N_44);
and U11584 (N_11584,N_3986,N_5993);
or U11585 (N_11585,N_523,N_2358);
and U11586 (N_11586,N_3009,N_2350);
nand U11587 (N_11587,N_937,N_749);
or U11588 (N_11588,N_890,N_958);
and U11589 (N_11589,N_4501,N_1813);
or U11590 (N_11590,N_1501,N_3787);
nor U11591 (N_11591,N_1635,N_5133);
nor U11592 (N_11592,N_3351,N_4072);
nor U11593 (N_11593,N_494,N_1610);
or U11594 (N_11594,N_5829,N_1766);
or U11595 (N_11595,N_2314,N_4479);
nor U11596 (N_11596,N_1985,N_3674);
nand U11597 (N_11597,N_5752,N_2184);
nor U11598 (N_11598,N_6131,N_232);
or U11599 (N_11599,N_543,N_3247);
and U11600 (N_11600,N_682,N_3231);
nor U11601 (N_11601,N_5610,N_3485);
and U11602 (N_11602,N_4588,N_4623);
or U11603 (N_11603,N_5765,N_3855);
nand U11604 (N_11604,N_5955,N_2983);
nand U11605 (N_11605,N_1238,N_1078);
nand U11606 (N_11606,N_5117,N_391);
or U11607 (N_11607,N_2081,N_3955);
and U11608 (N_11608,N_4736,N_2567);
or U11609 (N_11609,N_1680,N_2195);
nor U11610 (N_11610,N_5123,N_3992);
xor U11611 (N_11611,N_3947,N_3288);
nand U11612 (N_11612,N_1662,N_3098);
xnor U11613 (N_11613,N_3486,N_1945);
nand U11614 (N_11614,N_1949,N_406);
nor U11615 (N_11615,N_4913,N_6232);
or U11616 (N_11616,N_5632,N_2832);
xor U11617 (N_11617,N_6072,N_1686);
nor U11618 (N_11618,N_2460,N_5702);
nand U11619 (N_11619,N_3372,N_2557);
or U11620 (N_11620,N_2509,N_3556);
and U11621 (N_11621,N_5562,N_473);
nand U11622 (N_11622,N_827,N_5363);
and U11623 (N_11623,N_4825,N_2665);
nand U11624 (N_11624,N_2380,N_5060);
nor U11625 (N_11625,N_5587,N_217);
nand U11626 (N_11626,N_2532,N_1313);
nor U11627 (N_11627,N_806,N_4601);
and U11628 (N_11628,N_4619,N_2236);
nor U11629 (N_11629,N_1743,N_338);
nand U11630 (N_11630,N_4420,N_6049);
or U11631 (N_11631,N_4895,N_885);
or U11632 (N_11632,N_2214,N_2019);
xnor U11633 (N_11633,N_5800,N_2472);
or U11634 (N_11634,N_5789,N_5937);
nand U11635 (N_11635,N_6065,N_5326);
nand U11636 (N_11636,N_1370,N_1657);
and U11637 (N_11637,N_204,N_6181);
or U11638 (N_11638,N_3005,N_5516);
nand U11639 (N_11639,N_5665,N_4111);
xor U11640 (N_11640,N_5452,N_1161);
or U11641 (N_11641,N_2773,N_1769);
and U11642 (N_11642,N_2867,N_4782);
nand U11643 (N_11643,N_3208,N_3334);
or U11644 (N_11644,N_3813,N_2139);
nand U11645 (N_11645,N_5769,N_917);
and U11646 (N_11646,N_5530,N_4504);
or U11647 (N_11647,N_2246,N_1620);
nand U11648 (N_11648,N_2532,N_6196);
and U11649 (N_11649,N_4892,N_1900);
xor U11650 (N_11650,N_4016,N_2957);
nand U11651 (N_11651,N_4751,N_4504);
or U11652 (N_11652,N_1584,N_6152);
xor U11653 (N_11653,N_1599,N_2243);
and U11654 (N_11654,N_5145,N_167);
or U11655 (N_11655,N_4502,N_3396);
or U11656 (N_11656,N_4436,N_6158);
nor U11657 (N_11657,N_4095,N_5327);
and U11658 (N_11658,N_1417,N_1563);
nand U11659 (N_11659,N_1098,N_1596);
nor U11660 (N_11660,N_4570,N_5369);
nor U11661 (N_11661,N_38,N_3236);
and U11662 (N_11662,N_2401,N_3746);
nor U11663 (N_11663,N_4403,N_2266);
nor U11664 (N_11664,N_2896,N_3295);
nand U11665 (N_11665,N_5408,N_297);
nand U11666 (N_11666,N_4002,N_4923);
nor U11667 (N_11667,N_2617,N_705);
nor U11668 (N_11668,N_3614,N_2012);
nand U11669 (N_11669,N_5990,N_4687);
and U11670 (N_11670,N_5110,N_2817);
nor U11671 (N_11671,N_621,N_3206);
nor U11672 (N_11672,N_2413,N_4743);
or U11673 (N_11673,N_1874,N_690);
or U11674 (N_11674,N_4580,N_2987);
and U11675 (N_11675,N_5107,N_2362);
nand U11676 (N_11676,N_405,N_2571);
nand U11677 (N_11677,N_597,N_1953);
or U11678 (N_11678,N_5458,N_2733);
and U11679 (N_11679,N_5060,N_3524);
or U11680 (N_11680,N_4230,N_1106);
nor U11681 (N_11681,N_3753,N_2398);
and U11682 (N_11682,N_177,N_4305);
xnor U11683 (N_11683,N_1380,N_4182);
nor U11684 (N_11684,N_4027,N_2630);
nand U11685 (N_11685,N_1617,N_1714);
nor U11686 (N_11686,N_987,N_900);
and U11687 (N_11687,N_3320,N_3721);
or U11688 (N_11688,N_4186,N_184);
nand U11689 (N_11689,N_3534,N_2938);
nand U11690 (N_11690,N_2474,N_33);
and U11691 (N_11691,N_858,N_6237);
and U11692 (N_11692,N_1781,N_1160);
and U11693 (N_11693,N_1536,N_5069);
xnor U11694 (N_11694,N_3942,N_3002);
and U11695 (N_11695,N_3993,N_4082);
and U11696 (N_11696,N_1479,N_1487);
nor U11697 (N_11697,N_3469,N_1414);
and U11698 (N_11698,N_6085,N_5608);
or U11699 (N_11699,N_3913,N_1599);
or U11700 (N_11700,N_417,N_5007);
nor U11701 (N_11701,N_1447,N_2131);
nor U11702 (N_11702,N_1576,N_1850);
and U11703 (N_11703,N_6099,N_6167);
nor U11704 (N_11704,N_405,N_3963);
or U11705 (N_11705,N_2711,N_264);
nor U11706 (N_11706,N_1919,N_3322);
nand U11707 (N_11707,N_655,N_4632);
nand U11708 (N_11708,N_4594,N_5255);
xor U11709 (N_11709,N_1037,N_3998);
or U11710 (N_11710,N_1680,N_5906);
xnor U11711 (N_11711,N_5062,N_4125);
or U11712 (N_11712,N_529,N_1528);
nor U11713 (N_11713,N_2143,N_649);
and U11714 (N_11714,N_4178,N_1417);
or U11715 (N_11715,N_1057,N_6193);
and U11716 (N_11716,N_176,N_1340);
and U11717 (N_11717,N_4987,N_3979);
or U11718 (N_11718,N_929,N_1247);
xnor U11719 (N_11719,N_1120,N_990);
or U11720 (N_11720,N_497,N_4672);
and U11721 (N_11721,N_2230,N_1269);
and U11722 (N_11722,N_3445,N_2877);
xor U11723 (N_11723,N_5021,N_1619);
xor U11724 (N_11724,N_653,N_1466);
nand U11725 (N_11725,N_5999,N_760);
and U11726 (N_11726,N_5806,N_3281);
and U11727 (N_11727,N_5718,N_611);
and U11728 (N_11728,N_4363,N_1347);
or U11729 (N_11729,N_4113,N_2086);
nand U11730 (N_11730,N_6008,N_821);
nor U11731 (N_11731,N_5490,N_1757);
or U11732 (N_11732,N_3431,N_1314);
or U11733 (N_11733,N_4503,N_524);
nor U11734 (N_11734,N_5828,N_622);
nor U11735 (N_11735,N_4560,N_4725);
or U11736 (N_11736,N_5314,N_4425);
xor U11737 (N_11737,N_2361,N_3152);
nand U11738 (N_11738,N_4959,N_3965);
nand U11739 (N_11739,N_1452,N_4368);
and U11740 (N_11740,N_2017,N_2487);
nand U11741 (N_11741,N_4813,N_3031);
nand U11742 (N_11742,N_1518,N_341);
or U11743 (N_11743,N_1129,N_3202);
nand U11744 (N_11744,N_10,N_1497);
and U11745 (N_11745,N_2463,N_3634);
and U11746 (N_11746,N_444,N_420);
and U11747 (N_11747,N_5844,N_1632);
or U11748 (N_11748,N_338,N_1562);
nand U11749 (N_11749,N_361,N_3580);
nor U11750 (N_11750,N_1700,N_4897);
nor U11751 (N_11751,N_1061,N_5689);
nor U11752 (N_11752,N_861,N_1339);
nand U11753 (N_11753,N_4391,N_221);
or U11754 (N_11754,N_745,N_2479);
or U11755 (N_11755,N_5212,N_6138);
nor U11756 (N_11756,N_528,N_3161);
nand U11757 (N_11757,N_972,N_5408);
and U11758 (N_11758,N_6106,N_3736);
and U11759 (N_11759,N_452,N_2657);
nor U11760 (N_11760,N_3371,N_6057);
nor U11761 (N_11761,N_5339,N_3638);
nand U11762 (N_11762,N_423,N_5813);
nand U11763 (N_11763,N_3116,N_1299);
nand U11764 (N_11764,N_919,N_4242);
nand U11765 (N_11765,N_4229,N_267);
or U11766 (N_11766,N_1598,N_4625);
nand U11767 (N_11767,N_2414,N_398);
or U11768 (N_11768,N_1156,N_1678);
or U11769 (N_11769,N_1847,N_1193);
or U11770 (N_11770,N_2316,N_3135);
and U11771 (N_11771,N_705,N_5216);
or U11772 (N_11772,N_2414,N_4330);
nor U11773 (N_11773,N_5331,N_5682);
nand U11774 (N_11774,N_4156,N_3219);
nor U11775 (N_11775,N_4548,N_2080);
and U11776 (N_11776,N_1156,N_5915);
nand U11777 (N_11777,N_2787,N_5153);
nor U11778 (N_11778,N_1617,N_2038);
xnor U11779 (N_11779,N_5231,N_3028);
nand U11780 (N_11780,N_6229,N_6133);
nand U11781 (N_11781,N_434,N_4441);
and U11782 (N_11782,N_579,N_4916);
and U11783 (N_11783,N_3275,N_5474);
nor U11784 (N_11784,N_238,N_5899);
and U11785 (N_11785,N_6088,N_5859);
and U11786 (N_11786,N_2710,N_2669);
xor U11787 (N_11787,N_43,N_4107);
and U11788 (N_11788,N_1491,N_1222);
or U11789 (N_11789,N_106,N_2946);
nor U11790 (N_11790,N_3510,N_3047);
or U11791 (N_11791,N_3786,N_482);
and U11792 (N_11792,N_5325,N_1267);
or U11793 (N_11793,N_4901,N_5445);
or U11794 (N_11794,N_3306,N_1273);
and U11795 (N_11795,N_4416,N_683);
and U11796 (N_11796,N_5454,N_252);
nand U11797 (N_11797,N_4929,N_3975);
nand U11798 (N_11798,N_6117,N_4473);
nor U11799 (N_11799,N_3675,N_5575);
or U11800 (N_11800,N_2981,N_2756);
nand U11801 (N_11801,N_2478,N_4272);
or U11802 (N_11802,N_670,N_5331);
nand U11803 (N_11803,N_3731,N_4646);
or U11804 (N_11804,N_3097,N_5408);
or U11805 (N_11805,N_1596,N_1035);
xnor U11806 (N_11806,N_3626,N_3014);
nand U11807 (N_11807,N_4404,N_2386);
or U11808 (N_11808,N_541,N_5229);
nand U11809 (N_11809,N_353,N_4377);
or U11810 (N_11810,N_2487,N_1372);
or U11811 (N_11811,N_4583,N_2653);
or U11812 (N_11812,N_3110,N_4440);
xor U11813 (N_11813,N_2481,N_5182);
or U11814 (N_11814,N_1388,N_4253);
and U11815 (N_11815,N_3559,N_6067);
nor U11816 (N_11816,N_6105,N_5584);
xor U11817 (N_11817,N_5424,N_503);
or U11818 (N_11818,N_3716,N_2504);
or U11819 (N_11819,N_322,N_4183);
or U11820 (N_11820,N_43,N_6127);
or U11821 (N_11821,N_3956,N_1803);
or U11822 (N_11822,N_4509,N_5067);
and U11823 (N_11823,N_6058,N_1662);
and U11824 (N_11824,N_717,N_1766);
nand U11825 (N_11825,N_2185,N_4643);
or U11826 (N_11826,N_2467,N_2885);
and U11827 (N_11827,N_361,N_3702);
nor U11828 (N_11828,N_3808,N_6005);
or U11829 (N_11829,N_4487,N_2974);
nor U11830 (N_11830,N_5324,N_123);
or U11831 (N_11831,N_4027,N_2373);
or U11832 (N_11832,N_973,N_4893);
nor U11833 (N_11833,N_5019,N_150);
nor U11834 (N_11834,N_655,N_2428);
or U11835 (N_11835,N_434,N_3313);
nor U11836 (N_11836,N_3952,N_2545);
nand U11837 (N_11837,N_3950,N_4008);
nand U11838 (N_11838,N_1490,N_2664);
xor U11839 (N_11839,N_2824,N_1856);
or U11840 (N_11840,N_4106,N_921);
nand U11841 (N_11841,N_3143,N_5244);
nor U11842 (N_11842,N_3688,N_4536);
xnor U11843 (N_11843,N_4431,N_3654);
and U11844 (N_11844,N_770,N_4493);
nand U11845 (N_11845,N_1857,N_5688);
nand U11846 (N_11846,N_384,N_84);
or U11847 (N_11847,N_5987,N_160);
or U11848 (N_11848,N_4196,N_2255);
xor U11849 (N_11849,N_4514,N_3359);
nor U11850 (N_11850,N_4632,N_5161);
nor U11851 (N_11851,N_2728,N_765);
xnor U11852 (N_11852,N_1607,N_3294);
nand U11853 (N_11853,N_3900,N_1558);
or U11854 (N_11854,N_4973,N_2943);
nand U11855 (N_11855,N_2843,N_5533);
nand U11856 (N_11856,N_2800,N_1479);
or U11857 (N_11857,N_289,N_5356);
or U11858 (N_11858,N_4784,N_6248);
and U11859 (N_11859,N_4518,N_4792);
nor U11860 (N_11860,N_937,N_93);
and U11861 (N_11861,N_577,N_2178);
or U11862 (N_11862,N_3342,N_2845);
and U11863 (N_11863,N_4313,N_4977);
xnor U11864 (N_11864,N_1857,N_6203);
nor U11865 (N_11865,N_2633,N_5634);
nand U11866 (N_11866,N_4537,N_1904);
nor U11867 (N_11867,N_2069,N_3750);
nor U11868 (N_11868,N_5194,N_3478);
nand U11869 (N_11869,N_793,N_2657);
nand U11870 (N_11870,N_3170,N_1782);
or U11871 (N_11871,N_134,N_5471);
or U11872 (N_11872,N_3504,N_103);
or U11873 (N_11873,N_3226,N_654);
nor U11874 (N_11874,N_1755,N_874);
or U11875 (N_11875,N_1721,N_6030);
xor U11876 (N_11876,N_395,N_5377);
nor U11877 (N_11877,N_5479,N_5027);
or U11878 (N_11878,N_5709,N_5194);
and U11879 (N_11879,N_5845,N_3735);
or U11880 (N_11880,N_6158,N_3736);
nor U11881 (N_11881,N_2004,N_4819);
xnor U11882 (N_11882,N_1480,N_4289);
and U11883 (N_11883,N_3759,N_5786);
and U11884 (N_11884,N_5530,N_3687);
nand U11885 (N_11885,N_5287,N_381);
xnor U11886 (N_11886,N_3285,N_1544);
nor U11887 (N_11887,N_4269,N_5791);
nand U11888 (N_11888,N_1541,N_5000);
nand U11889 (N_11889,N_1678,N_1949);
and U11890 (N_11890,N_1211,N_1173);
nand U11891 (N_11891,N_2933,N_468);
or U11892 (N_11892,N_3531,N_3262);
nand U11893 (N_11893,N_4569,N_1154);
nand U11894 (N_11894,N_1409,N_5843);
and U11895 (N_11895,N_1702,N_2236);
or U11896 (N_11896,N_1985,N_3017);
xor U11897 (N_11897,N_1727,N_700);
nand U11898 (N_11898,N_1913,N_186);
nor U11899 (N_11899,N_3671,N_707);
nor U11900 (N_11900,N_4907,N_5486);
and U11901 (N_11901,N_5766,N_5892);
nand U11902 (N_11902,N_1354,N_3483);
or U11903 (N_11903,N_982,N_5879);
nor U11904 (N_11904,N_1994,N_2900);
nor U11905 (N_11905,N_4804,N_4246);
nor U11906 (N_11906,N_5207,N_4153);
or U11907 (N_11907,N_5158,N_4415);
nand U11908 (N_11908,N_991,N_1148);
or U11909 (N_11909,N_969,N_2281);
or U11910 (N_11910,N_6230,N_108);
and U11911 (N_11911,N_2186,N_2051);
or U11912 (N_11912,N_1852,N_4921);
nor U11913 (N_11913,N_1071,N_1717);
or U11914 (N_11914,N_4842,N_3766);
nand U11915 (N_11915,N_436,N_6146);
nor U11916 (N_11916,N_2869,N_1253);
or U11917 (N_11917,N_895,N_4271);
and U11918 (N_11918,N_6204,N_3053);
or U11919 (N_11919,N_971,N_5791);
nand U11920 (N_11920,N_3058,N_144);
and U11921 (N_11921,N_4661,N_4742);
nor U11922 (N_11922,N_4536,N_1765);
nand U11923 (N_11923,N_3054,N_346);
xor U11924 (N_11924,N_438,N_3401);
or U11925 (N_11925,N_1510,N_5734);
nand U11926 (N_11926,N_2193,N_1769);
nor U11927 (N_11927,N_5060,N_6166);
or U11928 (N_11928,N_5665,N_4857);
or U11929 (N_11929,N_3414,N_708);
and U11930 (N_11930,N_5245,N_1275);
nand U11931 (N_11931,N_3625,N_5289);
xnor U11932 (N_11932,N_6109,N_1838);
or U11933 (N_11933,N_2405,N_2234);
nor U11934 (N_11934,N_4259,N_216);
nor U11935 (N_11935,N_4494,N_417);
nor U11936 (N_11936,N_4977,N_386);
nor U11937 (N_11937,N_884,N_871);
nor U11938 (N_11938,N_720,N_2357);
or U11939 (N_11939,N_5507,N_2423);
nand U11940 (N_11940,N_4980,N_988);
nand U11941 (N_11941,N_4136,N_2127);
nand U11942 (N_11942,N_4849,N_3695);
and U11943 (N_11943,N_2552,N_421);
and U11944 (N_11944,N_5212,N_1953);
nor U11945 (N_11945,N_262,N_2405);
or U11946 (N_11946,N_2766,N_2468);
and U11947 (N_11947,N_5878,N_5971);
and U11948 (N_11948,N_3058,N_4059);
and U11949 (N_11949,N_4450,N_5427);
nor U11950 (N_11950,N_3432,N_5896);
or U11951 (N_11951,N_2183,N_4017);
or U11952 (N_11952,N_4952,N_3399);
nand U11953 (N_11953,N_5442,N_6168);
or U11954 (N_11954,N_4845,N_2181);
nor U11955 (N_11955,N_1840,N_958);
or U11956 (N_11956,N_4820,N_1652);
or U11957 (N_11957,N_1161,N_4940);
or U11958 (N_11958,N_5107,N_6221);
and U11959 (N_11959,N_1947,N_5802);
nand U11960 (N_11960,N_5075,N_3765);
or U11961 (N_11961,N_4499,N_4021);
and U11962 (N_11962,N_1482,N_2167);
xor U11963 (N_11963,N_2625,N_1477);
and U11964 (N_11964,N_1580,N_180);
and U11965 (N_11965,N_802,N_2080);
nor U11966 (N_11966,N_3729,N_231);
and U11967 (N_11967,N_2070,N_5610);
or U11968 (N_11968,N_3823,N_5865);
or U11969 (N_11969,N_2300,N_3701);
nor U11970 (N_11970,N_1137,N_2979);
and U11971 (N_11971,N_623,N_310);
xor U11972 (N_11972,N_3655,N_1918);
or U11973 (N_11973,N_3373,N_4230);
nand U11974 (N_11974,N_2588,N_3769);
nor U11975 (N_11975,N_3066,N_1618);
nor U11976 (N_11976,N_371,N_6148);
or U11977 (N_11977,N_1629,N_4049);
nor U11978 (N_11978,N_1202,N_3274);
or U11979 (N_11979,N_4644,N_803);
nor U11980 (N_11980,N_4615,N_3100);
or U11981 (N_11981,N_3707,N_4894);
and U11982 (N_11982,N_196,N_3451);
or U11983 (N_11983,N_528,N_4329);
and U11984 (N_11984,N_5244,N_4377);
or U11985 (N_11985,N_3941,N_3501);
nor U11986 (N_11986,N_3732,N_2011);
nand U11987 (N_11987,N_5342,N_3584);
nand U11988 (N_11988,N_633,N_5574);
xor U11989 (N_11989,N_2778,N_2558);
nor U11990 (N_11990,N_3106,N_4020);
nor U11991 (N_11991,N_4997,N_3988);
or U11992 (N_11992,N_284,N_3634);
nand U11993 (N_11993,N_5939,N_2403);
or U11994 (N_11994,N_1043,N_5847);
and U11995 (N_11995,N_1133,N_1224);
nor U11996 (N_11996,N_1954,N_1900);
xor U11997 (N_11997,N_3918,N_2086);
nor U11998 (N_11998,N_285,N_3645);
nor U11999 (N_11999,N_1041,N_1568);
xnor U12000 (N_12000,N_2083,N_6103);
or U12001 (N_12001,N_969,N_4650);
xnor U12002 (N_12002,N_5489,N_3098);
nand U12003 (N_12003,N_6156,N_2499);
nor U12004 (N_12004,N_1982,N_864);
and U12005 (N_12005,N_2302,N_399);
or U12006 (N_12006,N_278,N_2190);
nor U12007 (N_12007,N_1593,N_3839);
or U12008 (N_12008,N_4987,N_3892);
nand U12009 (N_12009,N_2198,N_4407);
and U12010 (N_12010,N_1704,N_4316);
nand U12011 (N_12011,N_946,N_3427);
and U12012 (N_12012,N_3732,N_1169);
or U12013 (N_12013,N_6130,N_1773);
or U12014 (N_12014,N_4870,N_3758);
and U12015 (N_12015,N_1440,N_3851);
nor U12016 (N_12016,N_1795,N_2137);
nor U12017 (N_12017,N_5677,N_2453);
and U12018 (N_12018,N_2790,N_2363);
and U12019 (N_12019,N_3618,N_1250);
or U12020 (N_12020,N_301,N_6214);
nand U12021 (N_12021,N_4195,N_1506);
nand U12022 (N_12022,N_3259,N_5355);
or U12023 (N_12023,N_5528,N_2276);
nor U12024 (N_12024,N_5972,N_3198);
nand U12025 (N_12025,N_4706,N_2690);
xor U12026 (N_12026,N_3082,N_762);
nand U12027 (N_12027,N_4831,N_4393);
xnor U12028 (N_12028,N_495,N_6162);
nand U12029 (N_12029,N_1034,N_3688);
nor U12030 (N_12030,N_5302,N_5576);
and U12031 (N_12031,N_1406,N_6107);
or U12032 (N_12032,N_3911,N_5370);
nor U12033 (N_12033,N_2062,N_508);
nor U12034 (N_12034,N_1877,N_4317);
or U12035 (N_12035,N_4593,N_82);
nand U12036 (N_12036,N_568,N_2498);
or U12037 (N_12037,N_2340,N_5231);
nor U12038 (N_12038,N_4506,N_5626);
nor U12039 (N_12039,N_4827,N_3661);
and U12040 (N_12040,N_5586,N_857);
and U12041 (N_12041,N_4509,N_4546);
and U12042 (N_12042,N_2641,N_5825);
and U12043 (N_12043,N_5928,N_4193);
nand U12044 (N_12044,N_3447,N_2825);
nand U12045 (N_12045,N_828,N_464);
or U12046 (N_12046,N_1554,N_1062);
or U12047 (N_12047,N_4618,N_5116);
and U12048 (N_12048,N_4531,N_6134);
nand U12049 (N_12049,N_1050,N_4141);
nor U12050 (N_12050,N_2933,N_563);
or U12051 (N_12051,N_2581,N_536);
nand U12052 (N_12052,N_3649,N_3355);
nor U12053 (N_12053,N_874,N_1112);
or U12054 (N_12054,N_1313,N_920);
and U12055 (N_12055,N_5465,N_5855);
nor U12056 (N_12056,N_2788,N_2648);
nand U12057 (N_12057,N_2659,N_2239);
or U12058 (N_12058,N_3844,N_3933);
nand U12059 (N_12059,N_2145,N_781);
nand U12060 (N_12060,N_4597,N_3278);
and U12061 (N_12061,N_4054,N_6192);
and U12062 (N_12062,N_3109,N_6146);
and U12063 (N_12063,N_3570,N_3689);
or U12064 (N_12064,N_4566,N_2368);
and U12065 (N_12065,N_3527,N_4289);
or U12066 (N_12066,N_2164,N_2525);
or U12067 (N_12067,N_5828,N_5438);
and U12068 (N_12068,N_6124,N_5215);
xor U12069 (N_12069,N_3492,N_2853);
nand U12070 (N_12070,N_3018,N_5364);
or U12071 (N_12071,N_1096,N_5786);
nor U12072 (N_12072,N_5108,N_6107);
nor U12073 (N_12073,N_4375,N_4494);
and U12074 (N_12074,N_4945,N_4149);
and U12075 (N_12075,N_6215,N_772);
xnor U12076 (N_12076,N_5127,N_4065);
and U12077 (N_12077,N_326,N_4212);
xor U12078 (N_12078,N_2464,N_3201);
and U12079 (N_12079,N_2758,N_3731);
or U12080 (N_12080,N_873,N_4846);
nor U12081 (N_12081,N_4971,N_4107);
nor U12082 (N_12082,N_3368,N_2365);
nor U12083 (N_12083,N_2771,N_4908);
or U12084 (N_12084,N_5038,N_3394);
or U12085 (N_12085,N_4347,N_2830);
nor U12086 (N_12086,N_4764,N_177);
nand U12087 (N_12087,N_1363,N_3544);
nand U12088 (N_12088,N_3614,N_1744);
or U12089 (N_12089,N_5842,N_6099);
and U12090 (N_12090,N_6172,N_2865);
and U12091 (N_12091,N_5314,N_4163);
nor U12092 (N_12092,N_2786,N_4013);
and U12093 (N_12093,N_4436,N_6248);
or U12094 (N_12094,N_492,N_1265);
nor U12095 (N_12095,N_3313,N_3566);
nor U12096 (N_12096,N_3855,N_4148);
and U12097 (N_12097,N_251,N_4567);
or U12098 (N_12098,N_6032,N_1081);
xor U12099 (N_12099,N_5523,N_492);
and U12100 (N_12100,N_2809,N_5625);
or U12101 (N_12101,N_4639,N_725);
nor U12102 (N_12102,N_1879,N_5251);
nand U12103 (N_12103,N_4896,N_5882);
nor U12104 (N_12104,N_4217,N_4663);
nand U12105 (N_12105,N_1785,N_167);
nand U12106 (N_12106,N_2555,N_2994);
or U12107 (N_12107,N_3714,N_4595);
or U12108 (N_12108,N_1746,N_3745);
nor U12109 (N_12109,N_4836,N_6223);
and U12110 (N_12110,N_2364,N_5212);
xnor U12111 (N_12111,N_83,N_2795);
nor U12112 (N_12112,N_956,N_1461);
and U12113 (N_12113,N_682,N_5931);
or U12114 (N_12114,N_2800,N_392);
xor U12115 (N_12115,N_4814,N_5152);
and U12116 (N_12116,N_4070,N_1398);
and U12117 (N_12117,N_4881,N_4873);
nor U12118 (N_12118,N_4730,N_5795);
nor U12119 (N_12119,N_2531,N_2360);
or U12120 (N_12120,N_1187,N_347);
nor U12121 (N_12121,N_2263,N_4767);
xor U12122 (N_12122,N_1126,N_2890);
and U12123 (N_12123,N_4529,N_258);
xor U12124 (N_12124,N_5290,N_2325);
and U12125 (N_12125,N_5138,N_2576);
nor U12126 (N_12126,N_1742,N_4841);
nor U12127 (N_12127,N_2189,N_1009);
and U12128 (N_12128,N_422,N_2577);
or U12129 (N_12129,N_5489,N_357);
and U12130 (N_12130,N_873,N_5095);
nand U12131 (N_12131,N_5300,N_5267);
xor U12132 (N_12132,N_3355,N_2055);
or U12133 (N_12133,N_1862,N_5448);
or U12134 (N_12134,N_3741,N_3530);
nand U12135 (N_12135,N_4125,N_5539);
or U12136 (N_12136,N_87,N_4535);
nor U12137 (N_12137,N_4208,N_4165);
xnor U12138 (N_12138,N_4183,N_3472);
or U12139 (N_12139,N_4668,N_5377);
or U12140 (N_12140,N_3300,N_4414);
or U12141 (N_12141,N_46,N_2830);
xnor U12142 (N_12142,N_862,N_2323);
and U12143 (N_12143,N_580,N_5418);
nor U12144 (N_12144,N_1298,N_1970);
or U12145 (N_12145,N_5763,N_5066);
nor U12146 (N_12146,N_575,N_2047);
xnor U12147 (N_12147,N_3166,N_19);
and U12148 (N_12148,N_5278,N_5804);
and U12149 (N_12149,N_2382,N_2219);
nand U12150 (N_12150,N_5053,N_2446);
or U12151 (N_12151,N_3156,N_1394);
xnor U12152 (N_12152,N_2881,N_2901);
nor U12153 (N_12153,N_5604,N_4249);
or U12154 (N_12154,N_3530,N_3726);
xor U12155 (N_12155,N_846,N_3871);
xnor U12156 (N_12156,N_3182,N_4350);
nand U12157 (N_12157,N_1458,N_6153);
or U12158 (N_12158,N_355,N_2042);
nor U12159 (N_12159,N_3537,N_116);
nor U12160 (N_12160,N_1801,N_5278);
or U12161 (N_12161,N_5185,N_4519);
nand U12162 (N_12162,N_3667,N_1888);
nor U12163 (N_12163,N_4279,N_3351);
nor U12164 (N_12164,N_4056,N_3289);
or U12165 (N_12165,N_5647,N_4502);
nor U12166 (N_12166,N_2402,N_4139);
or U12167 (N_12167,N_3242,N_4842);
nand U12168 (N_12168,N_1676,N_727);
and U12169 (N_12169,N_3695,N_1565);
nand U12170 (N_12170,N_5248,N_2372);
or U12171 (N_12171,N_5058,N_3382);
nand U12172 (N_12172,N_4160,N_809);
nor U12173 (N_12173,N_3423,N_1475);
and U12174 (N_12174,N_4154,N_2971);
and U12175 (N_12175,N_923,N_1052);
xnor U12176 (N_12176,N_2478,N_1010);
and U12177 (N_12177,N_4493,N_5521);
nor U12178 (N_12178,N_4585,N_4441);
and U12179 (N_12179,N_1445,N_133);
nand U12180 (N_12180,N_790,N_5220);
and U12181 (N_12181,N_4352,N_3635);
nor U12182 (N_12182,N_1848,N_1041);
nor U12183 (N_12183,N_2435,N_5069);
nor U12184 (N_12184,N_3835,N_629);
nor U12185 (N_12185,N_635,N_6116);
xor U12186 (N_12186,N_522,N_2367);
nand U12187 (N_12187,N_2720,N_3841);
and U12188 (N_12188,N_4115,N_1083);
or U12189 (N_12189,N_3560,N_5541);
and U12190 (N_12190,N_4056,N_2239);
nand U12191 (N_12191,N_496,N_3165);
nand U12192 (N_12192,N_5667,N_2209);
or U12193 (N_12193,N_2402,N_3987);
nand U12194 (N_12194,N_599,N_2706);
nand U12195 (N_12195,N_1586,N_62);
nor U12196 (N_12196,N_4522,N_4958);
or U12197 (N_12197,N_5162,N_1137);
or U12198 (N_12198,N_5930,N_1779);
nand U12199 (N_12199,N_4867,N_2261);
or U12200 (N_12200,N_5037,N_1797);
and U12201 (N_12201,N_6225,N_3170);
nand U12202 (N_12202,N_584,N_838);
nor U12203 (N_12203,N_4226,N_4921);
or U12204 (N_12204,N_3307,N_2366);
and U12205 (N_12205,N_2795,N_3116);
nor U12206 (N_12206,N_3209,N_2913);
nor U12207 (N_12207,N_4926,N_4703);
nand U12208 (N_12208,N_280,N_2406);
and U12209 (N_12209,N_4858,N_2295);
nand U12210 (N_12210,N_4832,N_5736);
nor U12211 (N_12211,N_993,N_5215);
xnor U12212 (N_12212,N_649,N_476);
and U12213 (N_12213,N_4335,N_3306);
nor U12214 (N_12214,N_5148,N_2433);
or U12215 (N_12215,N_3970,N_1937);
and U12216 (N_12216,N_5290,N_1391);
and U12217 (N_12217,N_1816,N_1110);
nand U12218 (N_12218,N_4446,N_5098);
and U12219 (N_12219,N_4066,N_5252);
or U12220 (N_12220,N_1963,N_3733);
nand U12221 (N_12221,N_409,N_5946);
nor U12222 (N_12222,N_4124,N_5205);
nand U12223 (N_12223,N_2804,N_1298);
nor U12224 (N_12224,N_5553,N_2729);
nand U12225 (N_12225,N_6096,N_2674);
nor U12226 (N_12226,N_4653,N_2372);
nor U12227 (N_12227,N_5770,N_648);
nor U12228 (N_12228,N_1940,N_4020);
or U12229 (N_12229,N_2603,N_1162);
or U12230 (N_12230,N_2368,N_4426);
and U12231 (N_12231,N_165,N_5473);
nor U12232 (N_12232,N_1223,N_5177);
nor U12233 (N_12233,N_3333,N_5923);
xor U12234 (N_12234,N_5400,N_5514);
and U12235 (N_12235,N_1094,N_2799);
nor U12236 (N_12236,N_1957,N_2884);
or U12237 (N_12237,N_4496,N_2458);
nand U12238 (N_12238,N_2882,N_172);
nand U12239 (N_12239,N_415,N_1324);
nand U12240 (N_12240,N_567,N_1498);
nand U12241 (N_12241,N_1269,N_3304);
nor U12242 (N_12242,N_611,N_1247);
xnor U12243 (N_12243,N_1521,N_3951);
or U12244 (N_12244,N_608,N_3969);
nor U12245 (N_12245,N_4570,N_1070);
or U12246 (N_12246,N_2571,N_2405);
and U12247 (N_12247,N_1260,N_392);
nand U12248 (N_12248,N_4851,N_69);
and U12249 (N_12249,N_894,N_4391);
and U12250 (N_12250,N_3940,N_1097);
and U12251 (N_12251,N_310,N_5652);
nand U12252 (N_12252,N_1486,N_3594);
xnor U12253 (N_12253,N_5792,N_6083);
xnor U12254 (N_12254,N_2827,N_5135);
or U12255 (N_12255,N_2485,N_5686);
or U12256 (N_12256,N_4336,N_1298);
and U12257 (N_12257,N_2351,N_4805);
nor U12258 (N_12258,N_3010,N_5897);
xnor U12259 (N_12259,N_5879,N_1018);
and U12260 (N_12260,N_1626,N_4988);
nand U12261 (N_12261,N_531,N_3436);
nor U12262 (N_12262,N_4581,N_1458);
or U12263 (N_12263,N_5733,N_3454);
nand U12264 (N_12264,N_3265,N_3376);
or U12265 (N_12265,N_231,N_3368);
nor U12266 (N_12266,N_318,N_5375);
or U12267 (N_12267,N_2380,N_370);
and U12268 (N_12268,N_2917,N_2361);
and U12269 (N_12269,N_1173,N_427);
nor U12270 (N_12270,N_3281,N_5973);
nand U12271 (N_12271,N_1132,N_3230);
nand U12272 (N_12272,N_1373,N_2431);
and U12273 (N_12273,N_139,N_2462);
and U12274 (N_12274,N_4407,N_3422);
nor U12275 (N_12275,N_3251,N_3479);
or U12276 (N_12276,N_2090,N_3804);
xnor U12277 (N_12277,N_2791,N_2030);
xor U12278 (N_12278,N_4872,N_4691);
and U12279 (N_12279,N_3989,N_5702);
or U12280 (N_12280,N_848,N_4825);
nand U12281 (N_12281,N_1132,N_1059);
and U12282 (N_12282,N_2425,N_2869);
nand U12283 (N_12283,N_6050,N_1432);
and U12284 (N_12284,N_426,N_5554);
and U12285 (N_12285,N_558,N_2866);
nor U12286 (N_12286,N_912,N_4347);
and U12287 (N_12287,N_606,N_1422);
or U12288 (N_12288,N_6050,N_2059);
and U12289 (N_12289,N_4051,N_3697);
nand U12290 (N_12290,N_2288,N_4721);
nor U12291 (N_12291,N_3339,N_4860);
or U12292 (N_12292,N_1047,N_5973);
and U12293 (N_12293,N_3634,N_145);
or U12294 (N_12294,N_5602,N_2305);
nand U12295 (N_12295,N_318,N_2509);
and U12296 (N_12296,N_2974,N_5003);
nand U12297 (N_12297,N_904,N_4313);
xnor U12298 (N_12298,N_3670,N_3286);
or U12299 (N_12299,N_5968,N_1140);
or U12300 (N_12300,N_2854,N_3865);
nand U12301 (N_12301,N_3071,N_3900);
or U12302 (N_12302,N_1981,N_3911);
or U12303 (N_12303,N_4973,N_2097);
or U12304 (N_12304,N_1095,N_4156);
nand U12305 (N_12305,N_1603,N_3355);
and U12306 (N_12306,N_1324,N_4191);
and U12307 (N_12307,N_3936,N_2185);
nor U12308 (N_12308,N_5218,N_5740);
nor U12309 (N_12309,N_5632,N_843);
or U12310 (N_12310,N_4115,N_4399);
and U12311 (N_12311,N_2103,N_2691);
and U12312 (N_12312,N_2603,N_2117);
and U12313 (N_12313,N_3756,N_2855);
nor U12314 (N_12314,N_1503,N_1948);
or U12315 (N_12315,N_522,N_4680);
and U12316 (N_12316,N_2270,N_1996);
or U12317 (N_12317,N_46,N_1577);
and U12318 (N_12318,N_2149,N_4949);
and U12319 (N_12319,N_3864,N_6122);
and U12320 (N_12320,N_3917,N_419);
and U12321 (N_12321,N_379,N_4862);
nand U12322 (N_12322,N_5188,N_1446);
xnor U12323 (N_12323,N_4418,N_1160);
or U12324 (N_12324,N_154,N_1574);
or U12325 (N_12325,N_337,N_5840);
nor U12326 (N_12326,N_522,N_2460);
nor U12327 (N_12327,N_1337,N_2854);
nor U12328 (N_12328,N_5155,N_3995);
nand U12329 (N_12329,N_4242,N_4375);
and U12330 (N_12330,N_3559,N_2513);
nor U12331 (N_12331,N_1609,N_5207);
or U12332 (N_12332,N_2590,N_705);
or U12333 (N_12333,N_3458,N_3269);
or U12334 (N_12334,N_3365,N_4725);
or U12335 (N_12335,N_5651,N_1910);
and U12336 (N_12336,N_1204,N_4060);
and U12337 (N_12337,N_4322,N_4060);
nor U12338 (N_12338,N_1704,N_4722);
nor U12339 (N_12339,N_4886,N_2768);
xnor U12340 (N_12340,N_6071,N_6168);
nand U12341 (N_12341,N_1134,N_334);
xnor U12342 (N_12342,N_1213,N_4413);
nand U12343 (N_12343,N_481,N_4747);
and U12344 (N_12344,N_5843,N_5102);
nand U12345 (N_12345,N_3928,N_6068);
or U12346 (N_12346,N_6141,N_5109);
nand U12347 (N_12347,N_1465,N_3928);
and U12348 (N_12348,N_5819,N_410);
or U12349 (N_12349,N_5120,N_5151);
nand U12350 (N_12350,N_4329,N_1551);
nand U12351 (N_12351,N_5546,N_3789);
and U12352 (N_12352,N_5152,N_3326);
xor U12353 (N_12353,N_790,N_2095);
nand U12354 (N_12354,N_1399,N_2256);
or U12355 (N_12355,N_4379,N_2830);
or U12356 (N_12356,N_1737,N_233);
nand U12357 (N_12357,N_1438,N_353);
and U12358 (N_12358,N_5339,N_4793);
and U12359 (N_12359,N_2965,N_3292);
or U12360 (N_12360,N_1542,N_4994);
or U12361 (N_12361,N_2536,N_5887);
nand U12362 (N_12362,N_2960,N_1350);
and U12363 (N_12363,N_2504,N_4376);
and U12364 (N_12364,N_5410,N_4685);
or U12365 (N_12365,N_2552,N_3552);
xor U12366 (N_12366,N_206,N_1813);
or U12367 (N_12367,N_5914,N_5869);
nand U12368 (N_12368,N_3063,N_4301);
nand U12369 (N_12369,N_585,N_5177);
nor U12370 (N_12370,N_291,N_3853);
nor U12371 (N_12371,N_6209,N_3133);
and U12372 (N_12372,N_4434,N_217);
nand U12373 (N_12373,N_3173,N_1383);
or U12374 (N_12374,N_3043,N_3141);
nand U12375 (N_12375,N_5555,N_419);
xor U12376 (N_12376,N_2747,N_6028);
and U12377 (N_12377,N_1554,N_4796);
or U12378 (N_12378,N_2849,N_2748);
and U12379 (N_12379,N_2847,N_5047);
nor U12380 (N_12380,N_3978,N_5924);
nand U12381 (N_12381,N_4946,N_4404);
nor U12382 (N_12382,N_5660,N_314);
and U12383 (N_12383,N_5142,N_2103);
nor U12384 (N_12384,N_317,N_2885);
and U12385 (N_12385,N_2457,N_643);
nor U12386 (N_12386,N_4497,N_5558);
or U12387 (N_12387,N_4582,N_3117);
xor U12388 (N_12388,N_1881,N_6045);
and U12389 (N_12389,N_5293,N_5157);
or U12390 (N_12390,N_6099,N_3740);
and U12391 (N_12391,N_3753,N_5230);
and U12392 (N_12392,N_1316,N_2435);
or U12393 (N_12393,N_2640,N_1635);
nand U12394 (N_12394,N_2351,N_2150);
or U12395 (N_12395,N_5057,N_2499);
and U12396 (N_12396,N_894,N_776);
and U12397 (N_12397,N_2998,N_1786);
or U12398 (N_12398,N_3965,N_1462);
nand U12399 (N_12399,N_6151,N_2008);
xor U12400 (N_12400,N_751,N_3025);
nor U12401 (N_12401,N_3115,N_1543);
xor U12402 (N_12402,N_1260,N_3205);
nor U12403 (N_12403,N_3816,N_2220);
nor U12404 (N_12404,N_5987,N_5669);
and U12405 (N_12405,N_3541,N_3056);
nor U12406 (N_12406,N_830,N_1998);
or U12407 (N_12407,N_2794,N_1026);
and U12408 (N_12408,N_1038,N_5307);
or U12409 (N_12409,N_769,N_1856);
nor U12410 (N_12410,N_5860,N_2127);
and U12411 (N_12411,N_1612,N_6028);
and U12412 (N_12412,N_2923,N_5633);
nor U12413 (N_12413,N_3150,N_4549);
and U12414 (N_12414,N_3523,N_1259);
nor U12415 (N_12415,N_3475,N_4135);
xnor U12416 (N_12416,N_5084,N_1328);
and U12417 (N_12417,N_5278,N_1195);
nor U12418 (N_12418,N_340,N_6067);
xnor U12419 (N_12419,N_1551,N_2968);
or U12420 (N_12420,N_1471,N_384);
or U12421 (N_12421,N_4310,N_844);
and U12422 (N_12422,N_54,N_1979);
and U12423 (N_12423,N_4042,N_2816);
nand U12424 (N_12424,N_6042,N_6163);
or U12425 (N_12425,N_2022,N_2427);
nor U12426 (N_12426,N_322,N_1562);
or U12427 (N_12427,N_1994,N_2791);
nand U12428 (N_12428,N_944,N_3493);
and U12429 (N_12429,N_1630,N_3429);
or U12430 (N_12430,N_4472,N_4169);
or U12431 (N_12431,N_5268,N_1675);
and U12432 (N_12432,N_1337,N_3842);
and U12433 (N_12433,N_5501,N_686);
or U12434 (N_12434,N_1375,N_1827);
nand U12435 (N_12435,N_2826,N_3007);
or U12436 (N_12436,N_5324,N_5454);
nor U12437 (N_12437,N_6112,N_1992);
nand U12438 (N_12438,N_3071,N_1509);
and U12439 (N_12439,N_3122,N_3912);
nor U12440 (N_12440,N_179,N_6067);
or U12441 (N_12441,N_5395,N_708);
nand U12442 (N_12442,N_4234,N_1002);
and U12443 (N_12443,N_4257,N_3322);
nand U12444 (N_12444,N_3455,N_6246);
and U12445 (N_12445,N_488,N_4107);
and U12446 (N_12446,N_814,N_633);
nor U12447 (N_12447,N_1677,N_5884);
xnor U12448 (N_12448,N_4080,N_4059);
nand U12449 (N_12449,N_5911,N_2353);
and U12450 (N_12450,N_5483,N_5623);
and U12451 (N_12451,N_4068,N_5352);
and U12452 (N_12452,N_5163,N_1511);
or U12453 (N_12453,N_4548,N_965);
or U12454 (N_12454,N_2943,N_4031);
nor U12455 (N_12455,N_2766,N_5367);
and U12456 (N_12456,N_380,N_4498);
nand U12457 (N_12457,N_1480,N_764);
nand U12458 (N_12458,N_2157,N_2756);
nor U12459 (N_12459,N_1824,N_391);
and U12460 (N_12460,N_2280,N_1337);
nor U12461 (N_12461,N_1126,N_5131);
and U12462 (N_12462,N_3261,N_5368);
nand U12463 (N_12463,N_5702,N_4240);
or U12464 (N_12464,N_49,N_5848);
and U12465 (N_12465,N_4732,N_1719);
nor U12466 (N_12466,N_5343,N_1250);
nor U12467 (N_12467,N_5719,N_3652);
nand U12468 (N_12468,N_3352,N_820);
xnor U12469 (N_12469,N_4795,N_2676);
nor U12470 (N_12470,N_3114,N_164);
and U12471 (N_12471,N_4243,N_3241);
and U12472 (N_12472,N_1880,N_5752);
and U12473 (N_12473,N_4730,N_5455);
xnor U12474 (N_12474,N_2750,N_1696);
and U12475 (N_12475,N_3946,N_4167);
nor U12476 (N_12476,N_3805,N_2926);
nand U12477 (N_12477,N_2189,N_5448);
xor U12478 (N_12478,N_3335,N_5705);
nand U12479 (N_12479,N_1218,N_2362);
nor U12480 (N_12480,N_6071,N_658);
xor U12481 (N_12481,N_5091,N_1996);
nand U12482 (N_12482,N_4077,N_1108);
or U12483 (N_12483,N_2425,N_416);
xnor U12484 (N_12484,N_5362,N_6027);
and U12485 (N_12485,N_5182,N_4959);
and U12486 (N_12486,N_3699,N_6136);
nor U12487 (N_12487,N_2690,N_4659);
or U12488 (N_12488,N_5874,N_3491);
nor U12489 (N_12489,N_178,N_560);
nor U12490 (N_12490,N_4557,N_5533);
or U12491 (N_12491,N_5014,N_806);
and U12492 (N_12492,N_4826,N_4987);
nor U12493 (N_12493,N_5703,N_1674);
xor U12494 (N_12494,N_2446,N_5910);
nand U12495 (N_12495,N_6072,N_2658);
or U12496 (N_12496,N_3501,N_1960);
nor U12497 (N_12497,N_1232,N_1865);
xnor U12498 (N_12498,N_3603,N_4015);
nor U12499 (N_12499,N_6002,N_4824);
nor U12500 (N_12500,N_10990,N_8171);
nand U12501 (N_12501,N_10126,N_10996);
nor U12502 (N_12502,N_9863,N_8563);
or U12503 (N_12503,N_11698,N_8744);
nand U12504 (N_12504,N_10856,N_11130);
nor U12505 (N_12505,N_7856,N_6972);
or U12506 (N_12506,N_8980,N_8658);
and U12507 (N_12507,N_7616,N_9909);
or U12508 (N_12508,N_6405,N_6445);
and U12509 (N_12509,N_12407,N_8641);
and U12510 (N_12510,N_12147,N_6279);
or U12511 (N_12511,N_9423,N_6710);
or U12512 (N_12512,N_12481,N_7171);
nor U12513 (N_12513,N_8079,N_9810);
nand U12514 (N_12514,N_11544,N_11811);
nand U12515 (N_12515,N_10736,N_7658);
nor U12516 (N_12516,N_11630,N_8804);
and U12517 (N_12517,N_8342,N_8584);
xnor U12518 (N_12518,N_9195,N_9029);
nand U12519 (N_12519,N_10848,N_9739);
or U12520 (N_12520,N_7520,N_10163);
or U12521 (N_12521,N_9603,N_9101);
nor U12522 (N_12522,N_12001,N_9702);
and U12523 (N_12523,N_10506,N_12156);
and U12524 (N_12524,N_11383,N_7688);
nand U12525 (N_12525,N_12495,N_8047);
xnor U12526 (N_12526,N_10059,N_11503);
nand U12527 (N_12527,N_10751,N_7791);
nor U12528 (N_12528,N_7403,N_11739);
or U12529 (N_12529,N_11604,N_8531);
nand U12530 (N_12530,N_10263,N_10554);
nor U12531 (N_12531,N_8059,N_11056);
or U12532 (N_12532,N_12297,N_10620);
nand U12533 (N_12533,N_9849,N_6630);
nand U12534 (N_12534,N_10282,N_7001);
or U12535 (N_12535,N_10179,N_11438);
xor U12536 (N_12536,N_11559,N_9271);
nand U12537 (N_12537,N_9819,N_7752);
or U12538 (N_12538,N_7093,N_7214);
nand U12539 (N_12539,N_10431,N_12019);
or U12540 (N_12540,N_8739,N_10063);
nor U12541 (N_12541,N_7301,N_10693);
and U12542 (N_12542,N_9738,N_7138);
xnor U12543 (N_12543,N_8397,N_11568);
or U12544 (N_12544,N_7430,N_6595);
nand U12545 (N_12545,N_8711,N_9696);
or U12546 (N_12546,N_11081,N_9770);
nor U12547 (N_12547,N_8912,N_10820);
nand U12548 (N_12548,N_12225,N_7822);
and U12549 (N_12549,N_9677,N_6996);
nand U12550 (N_12550,N_11267,N_6690);
or U12551 (N_12551,N_8615,N_9232);
or U12552 (N_12552,N_10151,N_11395);
nor U12553 (N_12553,N_11289,N_9994);
nand U12554 (N_12554,N_10199,N_11737);
nand U12555 (N_12555,N_6418,N_9530);
xnor U12556 (N_12556,N_7627,N_9543);
xor U12557 (N_12557,N_9735,N_9208);
or U12558 (N_12558,N_10955,N_6439);
and U12559 (N_12559,N_10393,N_8892);
nor U12560 (N_12560,N_11144,N_6505);
and U12561 (N_12561,N_10572,N_6417);
or U12562 (N_12562,N_7153,N_12293);
or U12563 (N_12563,N_6513,N_10476);
nand U12564 (N_12564,N_9560,N_8273);
and U12565 (N_12565,N_7998,N_11935);
nand U12566 (N_12566,N_11152,N_10907);
nor U12567 (N_12567,N_9321,N_12275);
or U12568 (N_12568,N_8411,N_10709);
nand U12569 (N_12569,N_6744,N_9577);
nor U12570 (N_12570,N_12318,N_7186);
and U12571 (N_12571,N_6788,N_9507);
nand U12572 (N_12572,N_9796,N_11984);
nand U12573 (N_12573,N_7061,N_7131);
or U12574 (N_12574,N_9668,N_8412);
and U12575 (N_12575,N_6306,N_11147);
and U12576 (N_12576,N_11259,N_8599);
nand U12577 (N_12577,N_6498,N_7742);
and U12578 (N_12578,N_12434,N_10436);
nor U12579 (N_12579,N_6725,N_8959);
nand U12580 (N_12580,N_11354,N_11591);
or U12581 (N_12581,N_11932,N_9744);
and U12582 (N_12582,N_7374,N_8286);
and U12583 (N_12583,N_8021,N_10912);
nand U12584 (N_12584,N_11906,N_11250);
nor U12585 (N_12585,N_11046,N_12155);
or U12586 (N_12586,N_9072,N_9965);
or U12587 (N_12587,N_12020,N_11852);
xnor U12588 (N_12588,N_6886,N_11367);
and U12589 (N_12589,N_11966,N_7031);
or U12590 (N_12590,N_11150,N_9771);
nor U12591 (N_12591,N_10133,N_9108);
and U12592 (N_12592,N_10192,N_6460);
nand U12593 (N_12593,N_11765,N_11990);
nand U12594 (N_12594,N_8318,N_7431);
nor U12595 (N_12595,N_9769,N_7866);
xnor U12596 (N_12596,N_6922,N_9049);
nand U12597 (N_12597,N_12014,N_10272);
xnor U12598 (N_12598,N_12497,N_9383);
nor U12599 (N_12599,N_11177,N_7708);
and U12600 (N_12600,N_8924,N_9716);
and U12601 (N_12601,N_11457,N_9631);
nand U12602 (N_12602,N_10313,N_9526);
or U12603 (N_12603,N_9276,N_9432);
nor U12604 (N_12604,N_12024,N_7059);
nor U12605 (N_12605,N_11458,N_10827);
or U12606 (N_12606,N_8201,N_11263);
or U12607 (N_12607,N_10985,N_7718);
xor U12608 (N_12608,N_7490,N_9806);
nand U12609 (N_12609,N_6815,N_9193);
and U12610 (N_12610,N_11404,N_11044);
and U12611 (N_12611,N_9439,N_8652);
nor U12612 (N_12612,N_7286,N_11114);
and U12613 (N_12613,N_8815,N_8438);
nand U12614 (N_12614,N_9681,N_6539);
nand U12615 (N_12615,N_11134,N_10354);
or U12616 (N_12616,N_11532,N_8379);
nor U12617 (N_12617,N_11403,N_6586);
nand U12618 (N_12618,N_8339,N_8713);
nand U12619 (N_12619,N_11620,N_9902);
and U12620 (N_12620,N_10857,N_8962);
nor U12621 (N_12621,N_7462,N_7048);
nand U12622 (N_12622,N_10363,N_9873);
nor U12623 (N_12623,N_6607,N_8170);
nand U12624 (N_12624,N_7152,N_8164);
and U12625 (N_12625,N_7532,N_9467);
nand U12626 (N_12626,N_11857,N_9643);
nor U12627 (N_12627,N_10988,N_10102);
and U12628 (N_12628,N_6311,N_11304);
nor U12629 (N_12629,N_7834,N_7289);
nor U12630 (N_12630,N_7287,N_6394);
nand U12631 (N_12631,N_11531,N_7255);
nand U12632 (N_12632,N_10097,N_7134);
nand U12633 (N_12633,N_7422,N_7934);
or U12634 (N_12634,N_9199,N_6546);
or U12635 (N_12635,N_7121,N_8583);
nand U12636 (N_12636,N_8348,N_6759);
nand U12637 (N_12637,N_12267,N_8462);
nor U12638 (N_12638,N_9002,N_6923);
or U12639 (N_12639,N_11116,N_7961);
and U12640 (N_12640,N_9135,N_6383);
or U12641 (N_12641,N_6957,N_11791);
xnor U12642 (N_12642,N_7720,N_10697);
or U12643 (N_12643,N_6365,N_7836);
nand U12644 (N_12644,N_11092,N_11062);
nand U12645 (N_12645,N_11702,N_9688);
nand U12646 (N_12646,N_8272,N_10608);
or U12647 (N_12647,N_12272,N_9273);
and U12648 (N_12648,N_8754,N_7022);
nor U12649 (N_12649,N_11355,N_12454);
nor U12650 (N_12650,N_9297,N_12447);
xnor U12651 (N_12651,N_8520,N_8146);
nand U12652 (N_12652,N_10305,N_7544);
and U12653 (N_12653,N_10541,N_9646);
or U12654 (N_12654,N_8690,N_11157);
nor U12655 (N_12655,N_10831,N_8724);
nor U12656 (N_12656,N_6628,N_11901);
nor U12657 (N_12657,N_11802,N_10713);
nand U12658 (N_12658,N_7936,N_10438);
or U12659 (N_12659,N_8865,N_8137);
nand U12660 (N_12660,N_8507,N_11965);
nand U12661 (N_12661,N_11836,N_12443);
nand U12662 (N_12662,N_6415,N_10062);
nand U12663 (N_12663,N_11710,N_8904);
or U12664 (N_12664,N_7772,N_11431);
nor U12665 (N_12665,N_9761,N_8909);
or U12666 (N_12666,N_6600,N_11330);
and U12667 (N_12667,N_8642,N_9309);
nor U12668 (N_12668,N_12484,N_11807);
and U12669 (N_12669,N_8194,N_11659);
or U12670 (N_12670,N_7256,N_12159);
xor U12671 (N_12671,N_8922,N_9246);
nand U12672 (N_12672,N_6359,N_7614);
nand U12673 (N_12673,N_7940,N_6562);
nor U12674 (N_12674,N_10471,N_10411);
nor U12675 (N_12675,N_9568,N_10316);
nand U12676 (N_12676,N_6254,N_10984);
or U12677 (N_12677,N_11337,N_10729);
nand U12678 (N_12678,N_9822,N_10833);
nand U12679 (N_12679,N_11970,N_7865);
nand U12680 (N_12680,N_12106,N_10362);
or U12681 (N_12681,N_9351,N_11838);
nand U12682 (N_12682,N_11401,N_11317);
or U12683 (N_12683,N_6728,N_6327);
nand U12684 (N_12684,N_9093,N_10081);
and U12685 (N_12685,N_8993,N_8045);
xor U12686 (N_12686,N_6693,N_11641);
nand U12687 (N_12687,N_11927,N_7113);
nand U12688 (N_12688,N_7232,N_11615);
and U12689 (N_12689,N_7514,N_12065);
nor U12690 (N_12690,N_12033,N_6494);
nor U12691 (N_12691,N_10061,N_9686);
nand U12692 (N_12692,N_9957,N_8384);
or U12693 (N_12693,N_8099,N_9892);
nor U12694 (N_12694,N_8787,N_11947);
nor U12695 (N_12695,N_9375,N_11366);
nand U12696 (N_12696,N_7862,N_7041);
and U12697 (N_12697,N_11724,N_12448);
and U12698 (N_12698,N_8293,N_12455);
nor U12699 (N_12699,N_7917,N_6763);
nand U12700 (N_12700,N_8064,N_11002);
or U12701 (N_12701,N_8179,N_11775);
nand U12702 (N_12702,N_6873,N_11786);
and U12703 (N_12703,N_7308,N_12498);
nand U12704 (N_12704,N_12486,N_9165);
nor U12705 (N_12705,N_6372,N_11118);
or U12706 (N_12706,N_7326,N_7864);
and U12707 (N_12707,N_10499,N_6518);
nor U12708 (N_12708,N_7460,N_8317);
and U12709 (N_12709,N_9240,N_9176);
nor U12710 (N_12710,N_7533,N_12394);
and U12711 (N_12711,N_8032,N_9364);
nand U12712 (N_12712,N_6751,N_7410);
and U12713 (N_12713,N_10773,N_6574);
and U12714 (N_12714,N_7058,N_8082);
nor U12715 (N_12715,N_9112,N_11041);
xnor U12716 (N_12716,N_7154,N_12286);
nand U12717 (N_12717,N_11439,N_8351);
nand U12718 (N_12718,N_10705,N_9807);
nand U12719 (N_12719,N_8155,N_9975);
nor U12720 (N_12720,N_7637,N_11509);
or U12721 (N_12721,N_8609,N_11708);
or U12722 (N_12722,N_10546,N_7174);
and U12723 (N_12723,N_7105,N_10986);
nand U12724 (N_12724,N_7238,N_12485);
and U12725 (N_12725,N_11562,N_8631);
nor U12726 (N_12726,N_11393,N_8848);
nand U12727 (N_12727,N_7758,N_6268);
or U12728 (N_12728,N_12128,N_10403);
xor U12729 (N_12729,N_12456,N_10226);
nor U12730 (N_12730,N_8634,N_7439);
nand U12731 (N_12731,N_10973,N_11050);
nand U12732 (N_12732,N_8648,N_12276);
nand U12733 (N_12733,N_12058,N_9050);
nand U12734 (N_12734,N_7505,N_11280);
and U12735 (N_12735,N_8928,N_11960);
or U12736 (N_12736,N_10526,N_7398);
xnor U12737 (N_12737,N_8366,N_8673);
nand U12738 (N_12738,N_9591,N_7359);
or U12739 (N_12739,N_8537,N_8797);
nor U12740 (N_12740,N_11587,N_7903);
and U12741 (N_12741,N_9928,N_8855);
and U12742 (N_12742,N_10543,N_10629);
and U12743 (N_12743,N_10614,N_6508);
nor U12744 (N_12744,N_8221,N_8259);
or U12745 (N_12745,N_6576,N_7361);
xor U12746 (N_12746,N_9486,N_8292);
xnor U12747 (N_12747,N_11226,N_6904);
nand U12748 (N_12748,N_7555,N_11803);
nand U12749 (N_12749,N_8911,N_12314);
nand U12750 (N_12750,N_7399,N_8251);
or U12751 (N_12751,N_11879,N_6387);
or U12752 (N_12752,N_6784,N_6726);
nor U12753 (N_12753,N_11779,N_12414);
nand U12754 (N_12754,N_11262,N_10035);
nand U12755 (N_12755,N_10392,N_8432);
nor U12756 (N_12756,N_8112,N_7055);
nand U12757 (N_12757,N_7319,N_9977);
or U12758 (N_12758,N_7795,N_11109);
or U12759 (N_12759,N_11703,N_11281);
nand U12760 (N_12760,N_10410,N_10220);
nor U12761 (N_12761,N_9508,N_12183);
nand U12762 (N_12762,N_9647,N_8161);
and U12763 (N_12763,N_8310,N_6499);
xor U12764 (N_12764,N_11482,N_11411);
xor U12765 (N_12765,N_12209,N_7633);
nand U12766 (N_12766,N_12228,N_9934);
nor U12767 (N_12767,N_7989,N_7139);
nand U12768 (N_12768,N_9649,N_12442);
nor U12769 (N_12769,N_11969,N_6644);
or U12770 (N_12770,N_7007,N_8502);
and U12771 (N_12771,N_10974,N_7250);
and U12772 (N_12772,N_9830,N_12433);
nor U12773 (N_12773,N_8316,N_7878);
and U12774 (N_12774,N_7142,N_10415);
nor U12775 (N_12775,N_11751,N_11917);
or U12776 (N_12776,N_8486,N_12358);
xnor U12777 (N_12777,N_10329,N_10348);
and U12778 (N_12778,N_7788,N_6698);
or U12779 (N_12779,N_6421,N_6457);
nor U12780 (N_12780,N_8886,N_6376);
nand U12781 (N_12781,N_9398,N_10374);
and U12782 (N_12782,N_7911,N_8223);
or U12783 (N_12783,N_7479,N_9684);
or U12784 (N_12784,N_11821,N_6472);
nor U12785 (N_12785,N_9039,N_9987);
or U12786 (N_12786,N_6567,N_11972);
and U12787 (N_12787,N_8174,N_7782);
and U12788 (N_12788,N_6834,N_10383);
or U12789 (N_12789,N_9085,N_7798);
and U12790 (N_12790,N_11223,N_7670);
and U12791 (N_12791,N_11916,N_11264);
or U12792 (N_12792,N_11706,N_8610);
nand U12793 (N_12793,N_8710,N_7833);
or U12794 (N_12794,N_11047,N_9671);
or U12795 (N_12795,N_9694,N_8481);
and U12796 (N_12796,N_10452,N_8190);
or U12797 (N_12797,N_10710,N_9918);
nor U12798 (N_12798,N_8463,N_10609);
or U12799 (N_12799,N_9227,N_7295);
nor U12800 (N_12800,N_11139,N_9588);
and U12801 (N_12801,N_11851,N_8620);
xor U12802 (N_12802,N_9125,N_9053);
nand U12803 (N_12803,N_9318,N_11859);
and U12804 (N_12804,N_11074,N_9664);
nand U12805 (N_12805,N_10594,N_11808);
nor U12806 (N_12806,N_11774,N_7129);
or U12807 (N_12807,N_12409,N_9118);
nand U12808 (N_12808,N_10665,N_12406);
or U12809 (N_12809,N_8514,N_10838);
and U12810 (N_12810,N_12154,N_8452);
and U12811 (N_12811,N_10702,N_9510);
or U12812 (N_12812,N_11886,N_10749);
or U12813 (N_12813,N_6920,N_11876);
nand U12814 (N_12814,N_10889,N_9481);
nor U12815 (N_12815,N_8343,N_8844);
nor U12816 (N_12816,N_11484,N_7068);
and U12817 (N_12817,N_6310,N_6645);
nand U12818 (N_12818,N_6691,N_11396);
or U12819 (N_12819,N_6816,N_10006);
xor U12820 (N_12820,N_7133,N_6428);
nor U12821 (N_12821,N_11212,N_6536);
and U12822 (N_12822,N_8624,N_9949);
or U12823 (N_12823,N_9211,N_8162);
nor U12824 (N_12824,N_11974,N_11605);
nand U12825 (N_12825,N_6866,N_8943);
nor U12826 (N_12826,N_11685,N_10574);
and U12827 (N_12827,N_10615,N_11288);
nand U12828 (N_12828,N_10727,N_7169);
or U12829 (N_12829,N_8607,N_10291);
nor U12830 (N_12830,N_10205,N_7426);
xnor U12831 (N_12831,N_7081,N_8381);
xor U12832 (N_12832,N_11809,N_6900);
nand U12833 (N_12833,N_10145,N_10724);
and U12834 (N_12834,N_11406,N_7993);
xor U12835 (N_12835,N_6269,N_12417);
or U12836 (N_12836,N_6578,N_7922);
and U12837 (N_12837,N_8346,N_10701);
or U12838 (N_12838,N_9847,N_10079);
and U12839 (N_12839,N_6288,N_9636);
xor U12840 (N_12840,N_7707,N_6361);
and U12841 (N_12841,N_8908,N_8800);
nor U12842 (N_12842,N_11442,N_10409);
nand U12843 (N_12843,N_11909,N_8947);
nor U12844 (N_12844,N_6799,N_9615);
nor U12845 (N_12845,N_9275,N_9008);
nand U12846 (N_12846,N_7760,N_12064);
nand U12847 (N_12847,N_9590,N_9673);
xor U12848 (N_12848,N_9220,N_9434);
or U12849 (N_12849,N_6363,N_11185);
or U12850 (N_12850,N_6629,N_10553);
xnor U12851 (N_12851,N_9492,N_11186);
nand U12852 (N_12852,N_7952,N_9366);
nand U12853 (N_12853,N_9194,N_7107);
nor U12854 (N_12854,N_10349,N_11162);
nand U12855 (N_12855,N_10739,N_10008);
and U12856 (N_12856,N_9479,N_6274);
and U12857 (N_12857,N_10288,N_6503);
nand U12858 (N_12858,N_8277,N_7740);
nor U12859 (N_12859,N_7728,N_7956);
or U12860 (N_12860,N_8906,N_6750);
or U12861 (N_12861,N_9904,N_6429);
or U12862 (N_12862,N_7318,N_6414);
nor U12863 (N_12863,N_10290,N_6331);
nor U12864 (N_12864,N_10661,N_9997);
or U12865 (N_12865,N_7665,N_7787);
xor U12866 (N_12866,N_8399,N_7401);
nand U12867 (N_12867,N_9840,N_11324);
nor U12868 (N_12868,N_6885,N_11371);
and U12869 (N_12869,N_10723,N_11426);
nor U12870 (N_12870,N_10603,N_7043);
and U12871 (N_12871,N_7870,N_11976);
and U12872 (N_12872,N_11837,N_6646);
nand U12873 (N_12873,N_9400,N_11741);
nor U12874 (N_12874,N_7100,N_8418);
xnor U12875 (N_12875,N_8020,N_7280);
nor U12876 (N_12876,N_11433,N_11329);
nor U12877 (N_12877,N_10832,N_7316);
or U12878 (N_12878,N_9571,N_7645);
nor U12879 (N_12879,N_6842,N_9466);
or U12880 (N_12880,N_9421,N_6863);
or U12881 (N_12881,N_11883,N_12346);
or U12882 (N_12882,N_9198,N_10576);
nor U12883 (N_12883,N_11720,N_6860);
and U12884 (N_12884,N_6982,N_8600);
and U12885 (N_12885,N_11609,N_10561);
and U12886 (N_12886,N_12298,N_9523);
or U12887 (N_12887,N_6822,N_9473);
and U12888 (N_12888,N_10235,N_11543);
or U12889 (N_12889,N_7756,N_6263);
xnor U12890 (N_12890,N_11508,N_8499);
or U12891 (N_12891,N_10125,N_8357);
nor U12892 (N_12892,N_7766,N_11348);
or U12893 (N_12893,N_12076,N_11138);
or U12894 (N_12894,N_7775,N_10886);
and U12895 (N_12895,N_7643,N_8106);
nand U12896 (N_12896,N_10419,N_9009);
or U12897 (N_12897,N_11266,N_7392);
or U12898 (N_12898,N_8382,N_8720);
and U12899 (N_12899,N_8842,N_6389);
xor U12900 (N_12900,N_11670,N_10873);
nand U12901 (N_12901,N_8781,N_8365);
nand U12902 (N_12902,N_7114,N_9151);
or U12903 (N_12903,N_10200,N_6851);
or U12904 (N_12904,N_8846,N_7698);
nand U12905 (N_12905,N_7717,N_8860);
nand U12906 (N_12906,N_10007,N_11474);
and U12907 (N_12907,N_6401,N_10478);
or U12908 (N_12908,N_10157,N_9940);
and U12909 (N_12909,N_8245,N_11296);
nor U12910 (N_12910,N_8903,N_11583);
nand U12911 (N_12911,N_6287,N_8374);
xnor U12912 (N_12912,N_7842,N_12196);
nand U12913 (N_12913,N_8241,N_11633);
and U12914 (N_12914,N_12244,N_9147);
nand U12915 (N_12915,N_7877,N_10483);
nor U12916 (N_12916,N_11364,N_8453);
nor U12917 (N_12917,N_12334,N_8459);
xnor U12918 (N_12918,N_11608,N_9252);
and U12919 (N_12919,N_8042,N_9846);
or U12920 (N_12920,N_11010,N_10598);
nand U12921 (N_12921,N_6326,N_8466);
or U12922 (N_12922,N_7881,N_11196);
and U12923 (N_12923,N_7542,N_7466);
and U12924 (N_12924,N_9119,N_12206);
nand U12925 (N_12925,N_8519,N_8256);
nand U12926 (N_12926,N_10915,N_7144);
nor U12927 (N_12927,N_7828,N_8538);
nand U12928 (N_12928,N_10654,N_8629);
and U12929 (N_12929,N_7680,N_11582);
nand U12930 (N_12930,N_6350,N_8338);
and U12931 (N_12931,N_12083,N_10071);
nand U12932 (N_12932,N_10947,N_12371);
nand U12933 (N_12933,N_8252,N_9470);
nand U12934 (N_12934,N_10028,N_11475);
nor U12935 (N_12935,N_12023,N_8033);
xnor U12936 (N_12936,N_6837,N_6843);
nand U12937 (N_12937,N_11008,N_11497);
xor U12938 (N_12938,N_6380,N_9561);
and U12939 (N_12939,N_6798,N_9784);
and U12940 (N_12940,N_12323,N_7654);
nand U12941 (N_12941,N_10261,N_8644);
nor U12942 (N_12942,N_8883,N_11199);
nor U12943 (N_12943,N_8113,N_8523);
nor U12944 (N_12944,N_11174,N_10798);
nand U12945 (N_12945,N_12171,N_8024);
nor U12946 (N_12946,N_8508,N_10711);
or U12947 (N_12947,N_10088,N_11505);
or U12948 (N_12948,N_9123,N_7411);
nor U12949 (N_12949,N_10646,N_10787);
xnor U12950 (N_12950,N_7071,N_6531);
nor U12951 (N_12951,N_9650,N_10781);
or U12952 (N_12952,N_9237,N_11561);
nand U12953 (N_12953,N_7005,N_9792);
or U12954 (N_12954,N_7729,N_10861);
nor U12955 (N_12955,N_10496,N_12333);
xor U12956 (N_12956,N_11217,N_11360);
and U12957 (N_12957,N_9841,N_7497);
or U12958 (N_12958,N_10124,N_11104);
xnor U12959 (N_12959,N_11934,N_8732);
nor U12960 (N_12960,N_12243,N_11486);
nor U12961 (N_12961,N_7003,N_11129);
xnor U12962 (N_12962,N_8166,N_11764);
or U12963 (N_12963,N_7328,N_11241);
nand U12964 (N_12964,N_6519,N_10236);
xor U12965 (N_12965,N_7586,N_10258);
and U12966 (N_12966,N_9828,N_6696);
nor U12967 (N_12967,N_8701,N_9419);
and U12968 (N_12968,N_8810,N_7716);
and U12969 (N_12969,N_9299,N_11137);
or U12970 (N_12970,N_8666,N_8013);
and U12971 (N_12971,N_10304,N_6487);
nand U12972 (N_12972,N_11992,N_10753);
nand U12973 (N_12973,N_8345,N_8173);
or U12974 (N_12974,N_8262,N_10965);
and U12975 (N_12975,N_7919,N_9245);
nand U12976 (N_12976,N_7813,N_8497);
and U12977 (N_12977,N_8283,N_8671);
nor U12978 (N_12978,N_10152,N_11000);
nor U12979 (N_12979,N_6330,N_8645);
and U12980 (N_12980,N_9864,N_11629);
and U12981 (N_12981,N_9669,N_11014);
or U12982 (N_12982,N_11142,N_12254);
and U12983 (N_12983,N_8260,N_7996);
and U12984 (N_12984,N_7216,N_9184);
and U12985 (N_12985,N_12292,N_9778);
and U12986 (N_12986,N_11790,N_8555);
or U12987 (N_12987,N_9926,N_10641);
nand U12988 (N_12988,N_11613,N_7969);
xnor U12989 (N_12989,N_9930,N_6903);
or U12990 (N_12990,N_9882,N_7346);
or U12991 (N_12991,N_12086,N_8882);
nor U12992 (N_12992,N_11908,N_8258);
and U12993 (N_12993,N_7179,N_11090);
xor U12994 (N_12994,N_9109,N_7743);
and U12995 (N_12995,N_6818,N_8821);
or U12996 (N_12996,N_7168,N_8480);
nor U12997 (N_12997,N_8455,N_8132);
nor U12998 (N_12998,N_11812,N_9156);
nor U12999 (N_12999,N_6345,N_8680);
nor U13000 (N_13000,N_6754,N_8937);
xnor U13001 (N_13001,N_8731,N_9293);
and U13002 (N_13002,N_10037,N_12252);
nand U13003 (N_13003,N_7202,N_7569);
nor U13004 (N_13004,N_9884,N_8498);
and U13005 (N_13005,N_8877,N_8605);
or U13006 (N_13006,N_6611,N_10726);
and U13007 (N_13007,N_8057,N_9566);
or U13008 (N_13008,N_9972,N_9316);
xor U13009 (N_13009,N_10001,N_8515);
nor U13010 (N_13010,N_9935,N_8898);
nor U13011 (N_13011,N_9953,N_8248);
and U13012 (N_13012,N_7019,N_11953);
or U13013 (N_13013,N_7858,N_10811);
xnor U13014 (N_13014,N_8108,N_11548);
and U13015 (N_13015,N_8953,N_7733);
or U13016 (N_13016,N_12170,N_7899);
or U13017 (N_13017,N_11871,N_9027);
or U13018 (N_13018,N_9903,N_11516);
and U13019 (N_13019,N_7607,N_11664);
and U13020 (N_13020,N_6955,N_11788);
nor U13021 (N_13021,N_9833,N_7260);
and U13022 (N_13022,N_11378,N_10539);
and U13023 (N_13023,N_10042,N_9497);
or U13024 (N_13024,N_10164,N_11878);
xnor U13025 (N_13025,N_9665,N_12162);
nand U13026 (N_13026,N_10273,N_11444);
or U13027 (N_13027,N_11578,N_7500);
nor U13028 (N_13028,N_11762,N_10252);
xnor U13029 (N_13029,N_7176,N_6991);
nand U13030 (N_13030,N_6681,N_7002);
and U13031 (N_13031,N_8159,N_10479);
and U13032 (N_13032,N_7939,N_6560);
nand U13033 (N_13033,N_8424,N_12088);
nand U13034 (N_13034,N_10065,N_8373);
xor U13035 (N_13035,N_6817,N_8429);
nand U13036 (N_13036,N_7692,N_8279);
nand U13037 (N_13037,N_8368,N_7262);
and U13038 (N_13038,N_8232,N_12097);
nand U13039 (N_13039,N_9178,N_8142);
nor U13040 (N_13040,N_12153,N_12130);
and U13041 (N_13041,N_6366,N_11690);
nand U13042 (N_13042,N_7781,N_7850);
and U13043 (N_13043,N_6705,N_11776);
nand U13044 (N_13044,N_9687,N_7838);
or U13045 (N_13045,N_8550,N_9868);
or U13046 (N_13046,N_9393,N_6902);
nand U13047 (N_13047,N_9901,N_10552);
nand U13048 (N_13048,N_6719,N_9848);
xnor U13049 (N_13049,N_10107,N_7641);
nor U13050 (N_13050,N_7324,N_10473);
or U13051 (N_13051,N_10160,N_8447);
and U13052 (N_13052,N_8760,N_11445);
or U13053 (N_13053,N_6608,N_11911);
and U13054 (N_13054,N_11825,N_6775);
and U13055 (N_13055,N_10768,N_6992);
or U13056 (N_13056,N_6720,N_10025);
nor U13057 (N_13057,N_12466,N_11640);
nor U13058 (N_13058,N_7572,N_7618);
nand U13059 (N_13059,N_9092,N_11409);
nand U13060 (N_13060,N_7471,N_9655);
nand U13061 (N_13061,N_10900,N_7651);
nor U13062 (N_13062,N_6599,N_8031);
and U13063 (N_13063,N_11958,N_8404);
xnor U13064 (N_13064,N_7282,N_8733);
nor U13065 (N_13065,N_9116,N_9757);
nand U13066 (N_13066,N_11725,N_10266);
or U13067 (N_13067,N_9790,N_9785);
or U13068 (N_13068,N_8125,N_6684);
nor U13069 (N_13069,N_10231,N_11530);
nand U13070 (N_13070,N_6284,N_11435);
nor U13071 (N_13071,N_12480,N_11463);
and U13072 (N_13072,N_7266,N_8006);
or U13073 (N_13073,N_11131,N_7137);
and U13074 (N_13074,N_7684,N_10021);
xnor U13075 (N_13075,N_10780,N_8309);
or U13076 (N_13076,N_12013,N_7487);
and U13077 (N_13077,N_7036,N_8849);
xnor U13078 (N_13078,N_6970,N_6565);
nand U13079 (N_13079,N_7052,N_11255);
and U13080 (N_13080,N_6556,N_10956);
nand U13081 (N_13081,N_9457,N_9795);
or U13082 (N_13082,N_11987,N_11660);
nand U13083 (N_13083,N_6448,N_10346);
or U13084 (N_13084,N_11286,N_8764);
nand U13085 (N_13085,N_7985,N_12059);
and U13086 (N_13086,N_11227,N_7650);
nand U13087 (N_13087,N_8741,N_12304);
or U13088 (N_13088,N_10099,N_8696);
nand U13089 (N_13089,N_10995,N_10423);
and U13090 (N_13090,N_9059,N_12268);
nand U13091 (N_13091,N_8702,N_11884);
and U13092 (N_13092,N_7060,N_10825);
nor U13093 (N_13093,N_8311,N_6480);
or U13094 (N_13094,N_8192,N_7944);
or U13095 (N_13095,N_11233,N_7872);
nand U13096 (N_13096,N_6432,N_8363);
or U13097 (N_13097,N_9756,N_10408);
and U13098 (N_13098,N_11332,N_10627);
and U13099 (N_13099,N_10905,N_11350);
and U13100 (N_13100,N_10529,N_9355);
nor U13101 (N_13101,N_6849,N_9545);
or U13102 (N_13102,N_11727,N_10041);
nor U13103 (N_13103,N_7943,N_8813);
or U13104 (N_13104,N_9783,N_7777);
nor U13105 (N_13105,N_9985,N_8917);
nand U13106 (N_13106,N_9323,N_8971);
xor U13107 (N_13107,N_7368,N_6589);
nor U13108 (N_13108,N_6631,N_10639);
nor U13109 (N_13109,N_8655,N_10384);
xor U13110 (N_13110,N_7299,N_11318);
nor U13111 (N_13111,N_12198,N_9462);
nor U13112 (N_13112,N_10105,N_12440);
nand U13113 (N_13113,N_9660,N_6358);
nor U13114 (N_13114,N_8851,N_7964);
xnor U13115 (N_13115,N_8703,N_7596);
nor U13116 (N_13116,N_12190,N_11555);
nor U13117 (N_13117,N_10254,N_7078);
and U13118 (N_13118,N_10318,N_11918);
and U13119 (N_13119,N_11473,N_8532);
nand U13120 (N_13120,N_10610,N_10013);
and U13121 (N_13121,N_7547,N_11540);
nor U13122 (N_13122,N_8988,N_8934);
and U13123 (N_13123,N_10275,N_6341);
or U13124 (N_13124,N_11524,N_11059);
nor U13125 (N_13125,N_12220,N_7937);
or U13126 (N_13126,N_10480,N_6946);
nor U13127 (N_13127,N_12216,N_6597);
nand U13128 (N_13128,N_10844,N_11537);
xor U13129 (N_13129,N_12120,N_11526);
and U13130 (N_13130,N_8875,N_9324);
nand U13131 (N_13131,N_12353,N_6470);
xor U13132 (N_13132,N_8561,N_7843);
and U13133 (N_13133,N_10066,N_10286);
or U13134 (N_13134,N_8199,N_6639);
nor U13135 (N_13135,N_7181,N_10161);
nand U13136 (N_13136,N_6626,N_6406);
nor U13137 (N_13137,N_12459,N_9551);
nor U13138 (N_13138,N_9249,N_9070);
or U13139 (N_13139,N_10270,N_10528);
nand U13140 (N_13140,N_9521,N_9877);
and U13141 (N_13141,N_11325,N_10330);
and U13142 (N_13142,N_7653,N_9140);
nor U13143 (N_13143,N_9041,N_12307);
nor U13144 (N_13144,N_11520,N_6606);
nand U13145 (N_13145,N_6791,N_7432);
and U13146 (N_13146,N_7784,N_11754);
nor U13147 (N_13147,N_11224,N_11347);
nor U13148 (N_13148,N_11761,N_9939);
and U13149 (N_13149,N_7674,N_10014);
nor U13150 (N_13150,N_11701,N_11870);
nor U13151 (N_13151,N_7463,N_10433);
nor U13152 (N_13152,N_9448,N_9071);
or U13153 (N_13153,N_11327,N_11341);
or U13154 (N_13154,N_8434,N_10223);
nor U13155 (N_13155,N_11869,N_8972);
nand U13156 (N_13156,N_7565,N_7499);
nor U13157 (N_13157,N_9047,N_7744);
and U13158 (N_13158,N_9110,N_10010);
nor U13159 (N_13159,N_12336,N_9493);
nand U13160 (N_13160,N_8557,N_10043);
xnor U13161 (N_13161,N_9415,N_6315);
or U13162 (N_13162,N_11523,N_9013);
or U13163 (N_13163,N_11417,N_11057);
nor U13164 (N_13164,N_10015,N_7384);
and U13165 (N_13165,N_9883,N_8872);
and U13166 (N_13166,N_9727,N_11500);
nor U13167 (N_13167,N_6980,N_9074);
and U13168 (N_13168,N_6884,N_7933);
nor U13169 (N_13169,N_8471,N_9161);
and U13170 (N_13170,N_7507,N_10551);
or U13171 (N_13171,N_10502,N_12269);
and U13172 (N_13172,N_12361,N_7579);
nor U13173 (N_13173,N_10123,N_9399);
or U13174 (N_13174,N_8868,N_8921);
nor U13175 (N_13175,N_8541,N_6260);
xnor U13176 (N_13176,N_10847,N_11920);
or U13177 (N_13177,N_6422,N_6368);
nor U13178 (N_13178,N_11416,N_10355);
xnor U13179 (N_13179,N_8358,N_8472);
and U13180 (N_13180,N_8437,N_9689);
and U13181 (N_13181,N_11564,N_8896);
nand U13182 (N_13182,N_8678,N_6846);
nand U13183 (N_13183,N_6969,N_10867);
nand U13184 (N_13184,N_11556,N_6475);
or U13185 (N_13185,N_11939,N_9710);
nand U13186 (N_13186,N_7304,N_11861);
nand U13187 (N_13187,N_9608,N_10943);
xnor U13188 (N_13188,N_7464,N_12152);
or U13189 (N_13189,N_11673,N_10334);
nor U13190 (N_13190,N_11070,N_10795);
nor U13191 (N_13191,N_9150,N_6879);
nand U13192 (N_13192,N_12113,N_8504);
xor U13193 (N_13193,N_7011,N_11307);
nand U13194 (N_13194,N_9980,N_7599);
and U13195 (N_13195,N_12302,N_7621);
and U13196 (N_13196,N_10851,N_10398);
or U13197 (N_13197,N_11955,N_6727);
nand U13198 (N_13198,N_9426,N_12000);
nor U13199 (N_13199,N_7894,N_10052);
nor U13200 (N_13200,N_12347,N_7534);
xor U13201 (N_13201,N_6400,N_9254);
or U13202 (N_13202,N_8588,N_10583);
nor U13203 (N_13203,N_7610,N_11801);
and U13204 (N_13204,N_10169,N_10842);
and U13205 (N_13205,N_11735,N_8041);
and U13206 (N_13206,N_11632,N_7723);
nand U13207 (N_13207,N_10703,N_7379);
nor U13208 (N_13208,N_11335,N_7636);
or U13209 (N_13209,N_10993,N_9304);
and U13210 (N_13210,N_11195,N_7185);
and U13211 (N_13211,N_10439,N_12303);
xnor U13212 (N_13212,N_7159,N_8585);
nor U13213 (N_13213,N_7274,N_7868);
nor U13214 (N_13214,N_8964,N_11156);
xor U13215 (N_13215,N_10754,N_12110);
xor U13216 (N_13216,N_8439,N_10714);
xnor U13217 (N_13217,N_11030,N_8567);
nand U13218 (N_13218,N_10904,N_11924);
nand U13219 (N_13219,N_12261,N_10684);
nor U13220 (N_13220,N_11694,N_9044);
nand U13221 (N_13221,N_10835,N_11033);
or U13222 (N_13222,N_8274,N_9765);
and U13223 (N_13223,N_11681,N_7315);
or U13224 (N_13224,N_10396,N_9191);
nor U13225 (N_13225,N_12041,N_12009);
nor U13226 (N_13226,N_8177,N_11203);
and U13227 (N_13227,N_12393,N_12316);
and U13228 (N_13228,N_6571,N_9392);
or U13229 (N_13229,N_11345,N_8743);
nand U13230 (N_13230,N_10232,N_6979);
nor U13231 (N_13231,N_12437,N_7590);
or U13232 (N_13232,N_9742,N_7415);
and U13233 (N_13233,N_6514,N_9292);
nand U13234 (N_13234,N_11191,N_9159);
nor U13235 (N_13235,N_9347,N_8839);
nor U13236 (N_13236,N_10799,N_12164);
nand U13237 (N_13237,N_11421,N_9812);
and U13238 (N_13238,N_9431,N_9674);
or U13239 (N_13239,N_7521,N_7300);
or U13240 (N_13240,N_8748,N_8712);
and U13241 (N_13241,N_9988,N_7909);
and U13242 (N_13242,N_6408,N_8361);
nand U13243 (N_13243,N_8869,N_9896);
and U13244 (N_13244,N_11243,N_12080);
xor U13245 (N_13245,N_6984,N_10488);
nor U13246 (N_13246,N_10340,N_9968);
nor U13247 (N_13247,N_9925,N_6512);
nand U13248 (N_13248,N_10147,N_8398);
nand U13249 (N_13249,N_9691,N_7908);
nor U13250 (N_13250,N_6634,N_11847);
and U13251 (N_13251,N_10936,N_12223);
nand U13252 (N_13252,N_7130,N_6520);
nand U13253 (N_13253,N_11132,N_10575);
and U13254 (N_13254,N_8352,N_8775);
and U13255 (N_13255,N_11988,N_6975);
xnor U13256 (N_13256,N_11446,N_8792);
and U13257 (N_13257,N_8406,N_7251);
and U13258 (N_13258,N_6594,N_8355);
and U13259 (N_13259,N_8985,N_7504);
or U13260 (N_13260,N_9797,N_10663);
nand U13261 (N_13261,N_12034,N_8951);
nor U13262 (N_13262,N_6785,N_11252);
or U13263 (N_13263,N_9381,N_11784);
or U13264 (N_13264,N_6664,N_9499);
nand U13265 (N_13265,N_12322,N_9335);
nand U13266 (N_13266,N_12401,N_10017);
nor U13267 (N_13267,N_8327,N_12410);
and U13268 (N_13268,N_12197,N_10301);
nor U13269 (N_13269,N_8289,N_7686);
or U13270 (N_13270,N_8965,N_6702);
and U13271 (N_13271,N_7570,N_12335);
xor U13272 (N_13272,N_10883,N_10345);
nor U13273 (N_13273,N_8154,N_9946);
or U13274 (N_13274,N_7450,N_10852);
and U13275 (N_13275,N_11058,N_12042);
and U13276 (N_13276,N_9310,N_6458);
and U13277 (N_13277,N_9064,N_9820);
or U13278 (N_13278,N_12161,N_6931);
nor U13279 (N_13279,N_11709,N_10573);
nor U13280 (N_13280,N_12217,N_11951);
and U13281 (N_13281,N_7049,N_12062);
nand U13282 (N_13282,N_11359,N_7404);
or U13283 (N_13283,N_7248,N_7024);
nand U13284 (N_13284,N_11082,N_7904);
and U13285 (N_13285,N_7199,N_12032);
nand U13286 (N_13286,N_10294,N_9175);
nor U13287 (N_13287,N_8598,N_10173);
and U13288 (N_13288,N_9951,N_7975);
nor U13289 (N_13289,N_9277,N_7406);
nor U13290 (N_13290,N_8889,N_9937);
xnor U13291 (N_13291,N_11225,N_9487);
nand U13292 (N_13292,N_7642,N_10373);
nand U13293 (N_13293,N_8827,N_10899);
nand U13294 (N_13294,N_7496,N_11235);
and U13295 (N_13295,N_7965,N_10375);
or U13296 (N_13296,N_7895,N_10868);
or U13297 (N_13297,N_7683,N_8749);
xor U13298 (N_13298,N_8253,N_9122);
and U13299 (N_13299,N_11914,N_7254);
nor U13300 (N_13300,N_8204,N_12326);
nand U13301 (N_13301,N_10140,N_6493);
xor U13302 (N_13302,N_10819,N_8983);
nand U13303 (N_13303,N_8410,N_6896);
nor U13304 (N_13304,N_9565,N_8026);
or U13305 (N_13305,N_11522,N_10527);
nand U13306 (N_13306,N_7959,N_10796);
nand U13307 (N_13307,N_7901,N_9805);
xor U13308 (N_13308,N_7212,N_7597);
and U13309 (N_13309,N_7855,N_10117);
or U13310 (N_13310,N_12079,N_12037);
nor U13311 (N_13311,N_12351,N_8281);
nand U13312 (N_13312,N_7609,N_6764);
nor U13313 (N_13313,N_7341,N_10870);
or U13314 (N_13314,N_6362,N_11101);
xor U13315 (N_13315,N_10946,N_6558);
xnor U13316 (N_13316,N_7844,N_8955);
or U13317 (N_13317,N_11771,N_12226);
nor U13318 (N_13318,N_11303,N_9158);
and U13319 (N_13319,N_7620,N_12202);
nor U13320 (N_13320,N_7818,N_6515);
and U13321 (N_13321,N_9260,N_9929);
and U13322 (N_13322,N_6393,N_9168);
xnor U13323 (N_13323,N_10808,N_12416);
nand U13324 (N_13324,N_9725,N_8981);
and U13325 (N_13325,N_10158,N_11674);
nor U13326 (N_13326,N_8156,N_7851);
and U13327 (N_13327,N_7164,N_11386);
nand U13328 (N_13328,N_8239,N_9042);
nand U13329 (N_13329,N_10850,N_10067);
nand U13330 (N_13330,N_10777,N_8043);
nor U13331 (N_13331,N_9891,N_9418);
nand U13332 (N_13332,N_8202,N_6911);
nor U13333 (N_13333,N_9266,N_9549);
or U13334 (N_13334,N_10662,N_11460);
xor U13335 (N_13335,N_11625,N_8656);
nor U13336 (N_13336,N_6324,N_10756);
or U13337 (N_13337,N_9853,N_11513);
nor U13338 (N_13338,N_9976,N_9023);
and U13339 (N_13339,N_11815,N_10156);
nor U13340 (N_13340,N_7079,N_9201);
nor U13341 (N_13341,N_6486,N_9413);
xnor U13342 (N_13342,N_11677,N_6827);
xnor U13343 (N_13343,N_11249,N_7433);
nor U13344 (N_13344,N_12066,N_11297);
or U13345 (N_13345,N_6459,N_8544);
or U13346 (N_13346,N_9169,N_7082);
nor U13347 (N_13347,N_8606,N_6716);
or U13348 (N_13348,N_8707,N_7025);
nand U13349 (N_13349,N_6907,N_10350);
xnor U13350 (N_13350,N_8275,N_11389);
and U13351 (N_13351,N_12004,N_9888);
nand U13352 (N_13352,N_9908,N_12366);
or U13353 (N_13353,N_9422,N_11919);
xor U13354 (N_13354,N_9215,N_8197);
nor U13355 (N_13355,N_7296,N_9038);
xor U13356 (N_13356,N_7412,N_12005);
and U13357 (N_13357,N_9713,N_9417);
or U13358 (N_13358,N_6772,N_6786);
and U13359 (N_13359,N_11584,N_6479);
nor U13360 (N_13360,N_9190,N_8752);
and U13361 (N_13361,N_10296,N_6688);
and U13362 (N_13362,N_8751,N_8115);
xnor U13363 (N_13363,N_10494,N_11361);
and U13364 (N_13364,N_11061,N_11183);
xor U13365 (N_13365,N_12174,N_9405);
nand U13366 (N_13366,N_9982,N_9464);
nor U13367 (N_13367,N_9210,N_7611);
nor U13368 (N_13368,N_10888,N_11107);
xnor U13369 (N_13369,N_10743,N_6768);
xnor U13370 (N_13370,N_10660,N_9931);
or U13371 (N_13371,N_10456,N_8581);
nand U13372 (N_13372,N_6841,N_7381);
nor U13373 (N_13373,N_11610,N_7126);
or U13374 (N_13374,N_7830,N_8556);
or U13375 (N_13375,N_11387,N_9866);
and U13376 (N_13376,N_6767,N_10580);
and U13377 (N_13377,N_9350,N_7949);
nand U13378 (N_13378,N_6875,N_6836);
nor U13379 (N_13379,N_7132,N_7783);
and U13380 (N_13380,N_10916,N_6667);
or U13381 (N_13381,N_9519,N_10534);
nor U13382 (N_13382,N_8861,N_10651);
xnor U13383 (N_13383,N_7298,N_10972);
nand U13384 (N_13384,N_7032,N_8149);
nand U13385 (N_13385,N_9712,N_6820);
nand U13386 (N_13386,N_10137,N_11099);
or U13387 (N_13387,N_7584,N_7884);
xor U13388 (N_13388,N_7157,N_11163);
and U13389 (N_13389,N_9453,N_9145);
nand U13390 (N_13390,N_8769,N_12463);
or U13391 (N_13391,N_7382,N_7149);
and U13392 (N_13392,N_12476,N_7035);
and U13393 (N_13393,N_10806,N_7924);
nor U13394 (N_13394,N_11818,N_12308);
nand U13395 (N_13395,N_7339,N_6641);
xor U13396 (N_13396,N_10209,N_12477);
or U13397 (N_13397,N_10036,N_12148);
nor U13398 (N_13398,N_7028,N_11476);
nand U13399 (N_13399,N_11936,N_9754);
or U13400 (N_13400,N_6461,N_9700);
or U13401 (N_13401,N_12232,N_11766);
and U13402 (N_13402,N_10864,N_9307);
and U13403 (N_13403,N_8958,N_9117);
nor U13404 (N_13404,N_8185,N_11394);
and U13405 (N_13405,N_10253,N_8096);
or U13406 (N_13406,N_11427,N_9576);
xnor U13407 (N_13407,N_9632,N_7320);
xor U13408 (N_13408,N_11423,N_10032);
nand U13409 (N_13409,N_9204,N_6588);
nor U13410 (N_13410,N_9328,N_8360);
nand U13411 (N_13411,N_7691,N_12006);
or U13412 (N_13412,N_7593,N_12390);
nor U13413 (N_13413,N_11684,N_11106);
and U13414 (N_13414,N_8559,N_7713);
or U13415 (N_13415,N_9638,N_6659);
xnor U13416 (N_13416,N_10255,N_12342);
and U13417 (N_13417,N_8271,N_9026);
nand U13418 (N_13418,N_11995,N_9675);
or U13419 (N_13419,N_12141,N_11299);
nor U13420 (N_13420,N_12363,N_10866);
or U13421 (N_13421,N_10394,N_9751);
nand U13422 (N_13422,N_7468,N_10095);
nor U13423 (N_13423,N_11778,N_12093);
nand U13424 (N_13424,N_6715,N_7962);
and U13425 (N_13425,N_6328,N_10481);
xor U13426 (N_13426,N_10172,N_11542);
nor U13427 (N_13427,N_7806,N_9075);
nor U13428 (N_13428,N_8878,N_6289);
or U13429 (N_13429,N_9045,N_7682);
nand U13430 (N_13430,N_6582,N_11023);
nor U13431 (N_13431,N_6348,N_8102);
or U13432 (N_13432,N_9578,N_9917);
and U13433 (N_13433,N_8029,N_9787);
nor U13434 (N_13434,N_7796,N_12189);
or U13435 (N_13435,N_10664,N_10607);
or U13436 (N_13436,N_12491,N_7696);
or U13437 (N_13437,N_7522,N_11577);
or U13438 (N_13438,N_10038,N_12280);
or U13439 (N_13439,N_6555,N_9274);
nand U13440 (N_13440,N_11648,N_6983);
nor U13441 (N_13441,N_12386,N_10680);
nand U13442 (N_13442,N_6521,N_6371);
nand U13443 (N_13443,N_12085,N_7103);
nor U13444 (N_13444,N_7017,N_6674);
or U13445 (N_13445,N_11078,N_6853);
nand U13446 (N_13446,N_10619,N_8334);
and U13447 (N_13447,N_8140,N_10118);
nand U13448 (N_13448,N_12438,N_8094);
nand U13449 (N_13449,N_11110,N_6283);
nor U13450 (N_13450,N_12378,N_6794);
nor U13451 (N_13451,N_9253,N_10814);
xnor U13452 (N_13452,N_7209,N_9295);
nor U13453 (N_13453,N_9056,N_9016);
xor U13454 (N_13454,N_11650,N_11067);
nand U13455 (N_13455,N_8297,N_8717);
or U13456 (N_13456,N_9973,N_11260);
xnor U13457 (N_13457,N_10696,N_7014);
or U13458 (N_13458,N_11451,N_9741);
and U13459 (N_13459,N_7735,N_10446);
nor U13460 (N_13460,N_10901,N_10060);
nor U13461 (N_13461,N_8061,N_10468);
nand U13462 (N_13462,N_10241,N_7340);
or U13463 (N_13463,N_9802,N_9410);
nand U13464 (N_13464,N_10428,N_8664);
or U13465 (N_13465,N_8038,N_8880);
or U13466 (N_13466,N_8843,N_6909);
and U13467 (N_13467,N_10689,N_10853);
and U13468 (N_13468,N_10911,N_9958);
and U13469 (N_13469,N_8580,N_12213);
nand U13470 (N_13470,N_11704,N_12214);
nor U13471 (N_13471,N_8784,N_7671);
xnor U13472 (N_13472,N_9241,N_10859);
nand U13473 (N_13473,N_9437,N_8377);
nor U13474 (N_13474,N_7918,N_11713);
nand U13475 (N_13475,N_9676,N_7396);
xnor U13476 (N_13476,N_8736,N_7145);
and U13477 (N_13477,N_7263,N_7902);
or U13478 (N_13478,N_8394,N_6420);
or U13479 (N_13479,N_8484,N_7594);
and U13480 (N_13480,N_8897,N_10367);
and U13481 (N_13481,N_8997,N_6739);
nor U13482 (N_13482,N_7362,N_11276);
nor U13483 (N_13483,N_6755,N_11004);
nor U13484 (N_13484,N_10260,N_11964);
xor U13485 (N_13485,N_9443,N_11980);
nor U13486 (N_13486,N_10632,N_6489);
nor U13487 (N_13487,N_9278,N_9225);
nand U13488 (N_13488,N_7929,N_8451);
xor U13489 (N_13489,N_8931,N_10950);
and U13490 (N_13490,N_11331,N_10818);
nand U13491 (N_13491,N_6872,N_9504);
nor U13492 (N_13492,N_12300,N_11519);
nor U13493 (N_13493,N_10103,N_7541);
nand U13494 (N_13494,N_10498,N_9535);
or U13495 (N_13495,N_7757,N_10735);
nand U13496 (N_13496,N_7170,N_12483);
xnor U13497 (N_13497,N_7625,N_9629);
and U13498 (N_13498,N_6985,N_12029);
xor U13499 (N_13499,N_10422,N_10992);
nor U13500 (N_13500,N_10489,N_10718);
nor U13501 (N_13501,N_11792,N_12051);
or U13502 (N_13502,N_8246,N_11257);
or U13503 (N_13503,N_11084,N_10389);
nand U13504 (N_13504,N_6723,N_8415);
nand U13505 (N_13505,N_7070,N_8564);
nand U13506 (N_13506,N_12327,N_10823);
xor U13507 (N_13507,N_6712,N_7355);
and U13508 (N_13508,N_7726,N_7515);
and U13509 (N_13509,N_11944,N_10982);
and U13510 (N_13510,N_6890,N_7963);
or U13511 (N_13511,N_9436,N_7160);
xor U13512 (N_13512,N_11733,N_8729);
nor U13513 (N_13513,N_8649,N_8326);
nand U13514 (N_13514,N_7023,N_8063);
or U13515 (N_13515,N_11298,N_9514);
or U13516 (N_13516,N_7067,N_8995);
nor U13517 (N_13517,N_10605,N_6427);
or U13518 (N_13518,N_6509,N_9587);
nor U13519 (N_13519,N_11855,N_7099);
or U13520 (N_13520,N_7336,N_6309);
nor U13521 (N_13521,N_8160,N_8948);
nor U13522 (N_13522,N_10863,N_12201);
and U13523 (N_13523,N_10759,N_7863);
or U13524 (N_13524,N_9124,N_7372);
and U13525 (N_13525,N_11595,N_6648);
and U13526 (N_13526,N_7920,N_8811);
and U13527 (N_13527,N_7012,N_9912);
and U13528 (N_13528,N_11265,N_10734);
nor U13529 (N_13529,N_8684,N_9839);
nor U13530 (N_13530,N_10217,N_9518);
and U13531 (N_13531,N_9991,N_6473);
nor U13532 (N_13532,N_8667,N_9438);
nand U13533 (N_13533,N_8208,N_8230);
or U13534 (N_13534,N_7879,N_11981);
nor U13535 (N_13535,N_8089,N_9711);
nand U13536 (N_13536,N_10585,N_7290);
nor U13537 (N_13537,N_10182,N_12082);
and U13538 (N_13538,N_10371,N_11202);
nor U13539 (N_13539,N_12233,N_9993);
nor U13540 (N_13540,N_12073,N_8441);
and U13541 (N_13541,N_9998,N_8536);
nand U13542 (N_13542,N_9300,N_8134);
or U13543 (N_13543,N_12398,N_11305);
nor U13544 (N_13544,N_7269,N_11830);
and U13545 (N_13545,N_9661,N_8774);
nand U13546 (N_13546,N_8467,N_8653);
nor U13547 (N_13547,N_12090,N_11658);
xor U13548 (N_13548,N_7600,N_7281);
or U13549 (N_13549,N_7664,N_9944);
nand U13550 (N_13550,N_10323,N_11336);
nand U13551 (N_13551,N_6782,N_11923);
nand U13552 (N_13552,N_9808,N_9031);
xnor U13553 (N_13553,N_9517,N_10746);
and U13554 (N_13554,N_6941,N_7178);
nor U13555 (N_13555,N_12096,N_7391);
nor U13556 (N_13556,N_6803,N_12224);
or U13557 (N_13557,N_8028,N_12138);
nand U13558 (N_13558,N_6738,N_11273);
nand U13559 (N_13559,N_7536,N_11636);
or U13560 (N_13560,N_8054,N_8854);
and U13561 (N_13561,N_10508,N_6411);
nor U13562 (N_13562,N_11546,N_7045);
or U13563 (N_13563,N_10779,N_9800);
xnor U13564 (N_13564,N_9870,N_9403);
and U13565 (N_13565,N_6444,N_12238);
and U13566 (N_13566,N_9995,N_8400);
and U13567 (N_13567,N_6416,N_11245);
or U13568 (N_13568,N_6867,N_9825);
nor U13569 (N_13569,N_9472,N_10618);
and U13570 (N_13570,N_8009,N_7297);
or U13571 (N_13571,N_11888,N_6699);
nand U13572 (N_13572,N_8954,N_6824);
nor U13573 (N_13573,N_7427,N_11817);
xnor U13574 (N_13574,N_10854,N_11714);
nand U13575 (N_13575,N_10119,N_8530);
nand U13576 (N_13576,N_7366,N_7095);
or U13577 (N_13577,N_10178,N_8905);
and U13578 (N_13578,N_7414,N_8049);
nand U13579 (N_13579,N_9662,N_7897);
and U13580 (N_13580,N_9622,N_6355);
nand U13581 (N_13581,N_9585,N_10484);
nor U13582 (N_13582,N_12157,N_7293);
or U13583 (N_13583,N_11091,N_12295);
and U13584 (N_13584,N_8970,N_8577);
nor U13585 (N_13585,N_10047,N_8758);
or U13586 (N_13586,N_9384,N_9984);
and U13587 (N_13587,N_12234,N_10213);
and U13588 (N_13588,N_11581,N_8535);
nor U13589 (N_13589,N_10557,N_8294);
and U13590 (N_13590,N_6367,N_11160);
xnor U13591 (N_13591,N_10128,N_9693);
nor U13592 (N_13592,N_9533,N_10645);
and U13593 (N_13593,N_8996,N_8055);
nand U13594 (N_13594,N_9722,N_10593);
or U13595 (N_13595,N_6452,N_10400);
nor U13596 (N_13596,N_11621,N_9572);
or U13597 (N_13597,N_9163,N_6692);
or U13598 (N_13598,N_11124,N_12039);
nand U13599 (N_13599,N_8093,N_12175);
and U13600 (N_13600,N_7349,N_7913);
or U13601 (N_13601,N_8986,N_11994);
xor U13602 (N_13602,N_9921,N_10490);
nor U13603 (N_13603,N_10344,N_7503);
nand U13604 (N_13604,N_9610,N_11579);
and U13605 (N_13605,N_8974,N_7930);
or U13606 (N_13606,N_6552,N_11495);
and U13607 (N_13607,N_6769,N_11487);
nand U13608 (N_13608,N_9942,N_8367);
nor U13609 (N_13609,N_9658,N_11275);
and U13610 (N_13610,N_7428,N_6928);
nand U13611 (N_13611,N_12050,N_11365);
nand U13612 (N_13612,N_8386,N_7242);
nand U13613 (N_13613,N_6986,N_10144);
xor U13614 (N_13614,N_11738,N_12166);
or U13615 (N_13615,N_9724,N_6482);
or U13616 (N_13616,N_9948,N_7829);
xnor U13617 (N_13617,N_12101,N_8939);
nor U13618 (N_13618,N_12100,N_9875);
and U13619 (N_13619,N_8172,N_9442);
or U13620 (N_13620,N_9594,N_11462);
nand U13621 (N_13621,N_10299,N_8693);
nand U13622 (N_13622,N_8639,N_10846);
xor U13623 (N_13623,N_7568,N_10892);
or U13624 (N_13624,N_8935,N_8572);
nor U13625 (N_13625,N_6625,N_10679);
nand U13626 (N_13626,N_10026,N_10948);
nand U13627 (N_13627,N_11370,N_6812);
nor U13628 (N_13628,N_6926,N_9256);
and U13629 (N_13629,N_7193,N_11678);
and U13630 (N_13630,N_9051,N_8828);
nor U13631 (N_13631,N_8184,N_7375);
or U13632 (N_13632,N_6757,N_11277);
nor U13633 (N_13633,N_10688,N_11949);
nand U13634 (N_13634,N_9267,N_11731);
or U13635 (N_13635,N_11220,N_10447);
or U13636 (N_13636,N_9171,N_11029);
or U13637 (N_13637,N_8888,N_8436);
and U13638 (N_13638,N_7845,N_6500);
xor U13639 (N_13639,N_6713,N_6953);
or U13640 (N_13640,N_7526,N_11381);
xnor U13641 (N_13641,N_7089,N_7792);
nor U13642 (N_13642,N_10782,N_6998);
nor U13643 (N_13643,N_11149,N_9843);
nor U13644 (N_13644,N_11912,N_8923);
nand U13645 (N_13645,N_7360,N_10979);
nor U13646 (N_13646,N_9389,N_10121);
or U13647 (N_13647,N_12127,N_8786);
nor U13648 (N_13648,N_11491,N_7397);
nor U13649 (N_13649,N_9762,N_9488);
nand U13650 (N_13650,N_9983,N_7472);
nor U13651 (N_13651,N_8856,N_11415);
and U13652 (N_13652,N_11108,N_7861);
nand U13653 (N_13653,N_9301,N_8209);
nand U13654 (N_13654,N_8335,N_9387);
and U13655 (N_13655,N_7669,N_11853);
or U13656 (N_13656,N_9390,N_7088);
and U13657 (N_13657,N_7817,N_11098);
nand U13658 (N_13658,N_7091,N_7292);
nand U13659 (N_13659,N_6838,N_9911);
nor U13660 (N_13660,N_12435,N_12137);
nand U13661 (N_13661,N_7976,N_6658);
nand U13662 (N_13662,N_10658,N_11862);
nor U13663 (N_13663,N_7672,N_7309);
nor U13664 (N_13664,N_8548,N_11639);
and U13665 (N_13665,N_12099,N_9454);
nor U13666 (N_13666,N_7552,N_6862);
nor U13667 (N_13667,N_7502,N_12026);
nor U13668 (N_13668,N_6881,N_7278);
and U13669 (N_13669,N_12215,N_12192);
or U13670 (N_13670,N_10171,N_6878);
xnor U13671 (N_13671,N_11742,N_8565);
and U13672 (N_13672,N_10155,N_12126);
or U13673 (N_13673,N_8925,N_8200);
nor U13674 (N_13674,N_10612,N_9542);
or U13675 (N_13675,N_9200,N_6995);
nand U13676 (N_13676,N_8396,N_11665);
nand U13677 (N_13677,N_12103,N_7173);
or U13678 (N_13678,N_7945,N_7098);
or U13679 (N_13679,N_8823,N_9789);
nor U13680 (N_13680,N_8638,N_11933);
or U13681 (N_13681,N_7732,N_7333);
nor U13682 (N_13682,N_8973,N_10757);
nor U13683 (N_13683,N_8044,N_7567);
and U13684 (N_13684,N_7648,N_8611);
nand U13685 (N_13685,N_11020,N_10306);
nand U13686 (N_13686,N_6603,N_11795);
nor U13687 (N_13687,N_12241,N_12475);
nand U13688 (N_13688,N_7230,N_11055);
nand U13689 (N_13689,N_10211,N_9874);
nand U13690 (N_13690,N_8697,N_12178);
nand U13691 (N_13691,N_7823,N_8183);
or U13692 (N_13692,N_7871,N_8375);
xnor U13693 (N_13693,N_10638,N_10533);
and U13694 (N_13694,N_8261,N_10890);
xnor U13695 (N_13695,N_8718,N_12204);
and U13696 (N_13696,N_7710,N_10699);
nand U13697 (N_13697,N_9595,N_8558);
nor U13698 (N_13698,N_6964,N_9376);
or U13699 (N_13699,N_11236,N_7612);
or U13700 (N_13700,N_10969,N_7204);
nand U13701 (N_13701,N_8562,N_11750);
nor U13702 (N_13702,N_11063,N_10525);
nand U13703 (N_13703,N_6252,N_7013);
nand U13704 (N_13704,N_11586,N_8070);
nor U13705 (N_13705,N_7461,N_11719);
nor U13706 (N_13706,N_6290,N_8282);
xnor U13707 (N_13707,N_8136,N_12102);
nor U13708 (N_13708,N_8950,N_6404);
or U13709 (N_13709,N_11301,N_7465);
and U13710 (N_13710,N_6548,N_7722);
xor U13711 (N_13711,N_8234,N_7562);
nor U13712 (N_13712,N_8837,N_7000);
and U13713 (N_13713,N_6749,N_10005);
nand U13714 (N_13714,N_10387,N_12262);
and U13715 (N_13715,N_8918,N_10999);
and U13716 (N_13716,N_11626,N_7429);
nor U13717 (N_13717,N_7029,N_7220);
nand U13718 (N_13718,N_11021,N_11283);
and U13719 (N_13719,N_8314,N_9793);
and U13720 (N_13720,N_10504,N_6868);
nand U13721 (N_13721,N_9914,N_11828);
or U13722 (N_13722,N_10039,N_6906);
and U13723 (N_13723,N_9601,N_12359);
nor U13724 (N_13724,N_11991,N_8211);
nor U13725 (N_13725,N_7218,N_10836);
nand U13726 (N_13726,N_12273,N_7473);
and U13727 (N_13727,N_6338,N_8505);
and U13728 (N_13728,N_9062,N_6901);
nor U13729 (N_13729,N_7501,N_8428);
nand U13730 (N_13730,N_6774,N_8617);
or U13731 (N_13731,N_6364,N_11900);
nor U13732 (N_13732,N_6258,N_6929);
nand U13733 (N_13733,N_10210,N_11278);
nor U13734 (N_13734,N_7687,N_8669);
nand U13735 (N_13735,N_10563,N_11313);
xnor U13736 (N_13736,N_10197,N_10695);
xor U13737 (N_13737,N_12279,N_8679);
nand U13738 (N_13738,N_8586,N_12246);
nor U13739 (N_13739,N_10971,N_7891);
or U13740 (N_13740,N_12015,N_10377);
nor U13741 (N_13741,N_9100,N_9231);
xor U13742 (N_13742,N_9144,N_11036);
nor U13743 (N_13743,N_8907,N_6510);
and U13744 (N_13744,N_7285,N_8187);
and U13745 (N_13745,N_12288,N_10094);
nor U13746 (N_13746,N_12402,N_10463);
nor U13747 (N_13747,N_11077,N_10687);
nor U13748 (N_13748,N_11209,N_11194);
nor U13749 (N_13749,N_10370,N_10510);
nand U13750 (N_13750,N_7474,N_8517);
nor U13751 (N_13751,N_11026,N_11390);
nand U13752 (N_13752,N_9547,N_11576);
nor U13753 (N_13753,N_7524,N_12256);
or U13754 (N_13754,N_9032,N_12482);
or U13755 (N_13755,N_11810,N_9342);
xnor U13756 (N_13756,N_11311,N_8737);
or U13757 (N_13757,N_10317,N_7984);
and U13758 (N_13758,N_7420,N_12160);
nor U13759 (N_13759,N_7679,N_10945);
nand U13760 (N_13760,N_11011,N_10758);
nor U13761 (N_13761,N_10240,N_11590);
nand U13762 (N_13762,N_9799,N_11206);
and U13763 (N_13763,N_7476,N_10769);
nor U13764 (N_13764,N_9001,N_8304);
or U13765 (N_13765,N_10523,N_8312);
and U13766 (N_13766,N_10589,N_11344);
nand U13767 (N_13767,N_10045,N_12423);
nand U13768 (N_13768,N_7739,N_11240);
or U13769 (N_13769,N_8771,N_11716);
nand U13770 (N_13770,N_8465,N_12352);
nand U13771 (N_13771,N_8165,N_8302);
nand U13772 (N_13772,N_6802,N_10653);
nand U13773 (N_13773,N_7598,N_7265);
nand U13774 (N_13774,N_10430,N_6870);
or U13775 (N_13775,N_7771,N_11699);
nor U13776 (N_13776,N_8135,N_10783);
and U13777 (N_13777,N_7892,N_10636);
xnor U13778 (N_13778,N_7745,N_6381);
or U13779 (N_13779,N_10944,N_6547);
nand U13780 (N_13780,N_12488,N_10807);
nor U13781 (N_13781,N_7955,N_8086);
nor U13782 (N_13782,N_6797,N_8578);
or U13783 (N_13783,N_11319,N_8300);
nand U13784 (N_13784,N_7180,N_11529);
nand U13785 (N_13785,N_8469,N_8349);
xor U13786 (N_13786,N_7378,N_11261);
nand U13787 (N_13787,N_6334,N_12257);
nor U13788 (N_13788,N_8547,N_11045);
nand U13789 (N_13789,N_9747,N_7311);
or U13790 (N_13790,N_11145,N_9251);
or U13791 (N_13791,N_7141,N_9552);
xor U13792 (N_13792,N_7416,N_6930);
and U13793 (N_13793,N_7451,N_10830);
or U13794 (N_13794,N_6590,N_7363);
or U13795 (N_13795,N_9311,N_7516);
nand U13796 (N_13796,N_6806,N_6356);
and U13797 (N_13797,N_8107,N_6619);
and U13798 (N_13798,N_11789,N_8306);
nor U13799 (N_13799,N_8735,N_9801);
nand U13800 (N_13800,N_11326,N_10595);
or U13801 (N_13801,N_11290,N_10940);
nand U13802 (N_13802,N_10535,N_9257);
and U13803 (N_13803,N_8372,N_6966);
nand U13804 (N_13804,N_6905,N_8687);
or U13805 (N_13805,N_9501,N_7923);
xnor U13806 (N_13806,N_7258,N_9567);
nand U13807 (N_13807,N_8092,N_8890);
nand U13808 (N_13808,N_6977,N_11657);
nor U13809 (N_13809,N_12211,N_10148);
nor U13810 (N_13810,N_12116,N_10800);
or U13811 (N_13811,N_8590,N_11753);
nand U13812 (N_13812,N_8824,N_8280);
and U13813 (N_13813,N_8413,N_11024);
nand U13814 (N_13814,N_9599,N_9030);
or U13815 (N_13815,N_6469,N_9794);
and U13816 (N_13816,N_8217,N_7854);
xnor U13817 (N_13817,N_7021,N_12425);
or U13818 (N_13818,N_12397,N_10776);
or U13819 (N_13819,N_11176,N_11661);
nor U13820 (N_13820,N_9089,N_11333);
xnor U13821 (N_13821,N_6402,N_10635);
xnor U13822 (N_13822,N_11414,N_10801);
nor U13823 (N_13823,N_11697,N_6952);
nand U13824 (N_13824,N_11087,N_7640);
nand U13825 (N_13825,N_8944,N_12131);
xor U13826 (N_13826,N_11618,N_7213);
and U13827 (N_13827,N_12021,N_6549);
or U13828 (N_13828,N_10271,N_11899);
nand U13829 (N_13829,N_10186,N_7456);
or U13830 (N_13830,N_10449,N_10437);
nor U13831 (N_13831,N_8133,N_7106);
nand U13832 (N_13832,N_7436,N_8331);
nor U13833 (N_13833,N_7753,N_7531);
xnor U13834 (N_13834,N_9932,N_7896);
nor U13835 (N_13835,N_9531,N_9349);
and U13836 (N_13836,N_7231,N_12077);
or U13837 (N_13837,N_8853,N_6273);
nand U13838 (N_13838,N_7268,N_6828);
or U13839 (N_13839,N_6543,N_10712);
or U13840 (N_13840,N_9766,N_6478);
nand U13841 (N_13841,N_6999,N_8371);
nand U13842 (N_13842,N_8885,N_11717);
and U13843 (N_13843,N_11379,N_11957);
and U13844 (N_13844,N_6942,N_6501);
nand U13845 (N_13845,N_7549,N_10300);
or U13846 (N_13846,N_9854,N_6678);
and U13847 (N_13847,N_7811,N_11001);
and U13848 (N_13848,N_11589,N_10656);
xor U13849 (N_13849,N_7846,N_7454);
or U13850 (N_13850,N_8138,N_7135);
or U13851 (N_13851,N_9731,N_11747);
nand U13852 (N_13852,N_8460,N_11816);
and U13853 (N_13853,N_11407,N_8695);
nor U13854 (N_13854,N_8738,N_11285);
or U13855 (N_13855,N_8229,N_7442);
xor U13856 (N_13856,N_11892,N_10096);
xor U13857 (N_13857,N_10070,N_11115);
nor U13858 (N_13858,N_6733,N_7763);
or U13859 (N_13859,N_9017,N_8464);
xnor U13860 (N_13860,N_8337,N_12227);
nor U13861 (N_13861,N_12283,N_6671);
nand U13862 (N_13862,N_11873,N_8444);
nand U13863 (N_13863,N_7697,N_9391);
nand U13864 (N_13864,N_8266,N_10333);
nor U13865 (N_13865,N_6789,N_9441);
nor U13866 (N_13866,N_10218,N_9320);
nand U13867 (N_13867,N_9040,N_9068);
and U13868 (N_13868,N_9209,N_10668);
nand U13869 (N_13869,N_6384,N_8832);
nor U13870 (N_13870,N_8150,N_11525);
nand U13871 (N_13871,N_9569,N_9597);
or U13872 (N_13872,N_6871,N_9476);
nor U13873 (N_13873,N_7201,N_6581);
or U13874 (N_13874,N_7369,N_10002);
and U13875 (N_13875,N_9491,N_7629);
and U13876 (N_13876,N_8244,N_8570);
or U13877 (N_13877,N_8573,N_7721);
xor U13878 (N_13878,N_6497,N_9319);
nor U13879 (N_13879,N_8403,N_7898);
nor U13880 (N_13880,N_7244,N_8494);
and U13881 (N_13881,N_6618,N_10244);
and U13882 (N_13882,N_7364,N_8966);
xnor U13883 (N_13883,N_11569,N_9527);
or U13884 (N_13884,N_10766,N_8062);
xor U13885 (N_13885,N_7385,N_9938);
nand U13886 (N_13886,N_12360,N_11248);
and U13887 (N_13887,N_11284,N_11518);
or U13888 (N_13888,N_8100,N_10624);
nand U13889 (N_13889,N_9139,N_11872);
and U13890 (N_13890,N_9337,N_11175);
or U13891 (N_13891,N_6948,N_11122);
nor U13892 (N_13892,N_11155,N_10056);
xor U13893 (N_13893,N_10569,N_9707);
nor U13894 (N_13894,N_11172,N_10429);
and U13895 (N_13895,N_7405,N_8691);
nand U13896 (N_13896,N_6354,N_8370);
and U13897 (N_13897,N_6305,N_6307);
nor U13898 (N_13898,N_10308,N_8957);
nor U13899 (N_13899,N_10809,N_6981);
nor U13900 (N_13900,N_8067,N_11231);
or U13901 (N_13901,N_10089,N_6272);
xnor U13902 (N_13902,N_6504,N_6557);
nand U13903 (N_13903,N_10778,N_10894);
nor U13904 (N_13904,N_9234,N_7768);
and U13905 (N_13905,N_8780,N_10465);
nand U13906 (N_13906,N_7950,N_9550);
and U13907 (N_13907,N_7970,N_6829);
and U13908 (N_13908,N_11963,N_11545);
nand U13909 (N_13909,N_10074,N_9698);
xor U13910 (N_13910,N_6989,N_7774);
nand U13911 (N_13911,N_10150,N_12415);
nand U13912 (N_13912,N_6541,N_8007);
nor U13913 (N_13913,N_12460,N_8812);
nand U13914 (N_13914,N_7327,N_12242);
nor U13915 (N_13915,N_6431,N_7034);
and U13916 (N_13916,N_12496,N_11638);
or U13917 (N_13917,N_12462,N_9913);
nand U13918 (N_13918,N_7972,N_8915);
nor U13919 (N_13919,N_10637,N_11470);
and U13920 (N_13920,N_9378,N_8819);
nor U13921 (N_13921,N_11071,N_8017);
or U13922 (N_13922,N_8817,N_7306);
xor U13923 (N_13923,N_7417,N_11154);
nor U13924 (N_13924,N_8785,N_8225);
nand U13925 (N_13925,N_6773,N_10675);
and U13926 (N_13926,N_9440,N_8960);
nand U13927 (N_13927,N_9107,N_6976);
and U13928 (N_13928,N_9554,N_7207);
nand U13929 (N_13929,N_10442,N_7117);
xor U13930 (N_13930,N_8433,N_6282);
and U13931 (N_13931,N_8867,N_11374);
nor U13932 (N_13932,N_8236,N_9264);
and U13933 (N_13933,N_9563,N_10180);
nand U13934 (N_13934,N_9087,N_10112);
nor U13935 (N_13935,N_9152,N_10927);
nor U13936 (N_13936,N_8299,N_6250);
and U13937 (N_13937,N_11654,N_7979);
nor U13938 (N_13938,N_7663,N_10193);
and U13939 (N_13939,N_11466,N_7358);
nor U13940 (N_13940,N_11968,N_6529);
or U13941 (N_13941,N_9346,N_12349);
nor U13942 (N_13942,N_11854,N_11696);
xnor U13943 (N_13943,N_6437,N_7800);
nor U13944 (N_13944,N_8350,N_8445);
xor U13945 (N_13945,N_8270,N_8157);
and U13946 (N_13946,N_10616,N_8409);
and U13947 (N_13947,N_9652,N_12199);
nor U13948 (N_13948,N_11352,N_10339);
xor U13949 (N_13949,N_9704,N_10303);
or U13950 (N_13950,N_11405,N_8402);
or U13951 (N_13951,N_7042,N_9218);
or U13952 (N_13952,N_7272,N_8956);
and U13953 (N_13953,N_7506,N_6443);
nand U13954 (N_13954,N_10432,N_9734);
nand U13955 (N_13955,N_8163,N_7110);
and U13956 (N_13956,N_9046,N_7564);
nand U13957 (N_13957,N_10351,N_12167);
nor U13958 (N_13958,N_7388,N_9173);
and U13959 (N_13959,N_12061,N_7084);
nor U13960 (N_13960,N_7347,N_6516);
nor U13961 (N_13961,N_7958,N_8829);
nor U13962 (N_13962,N_8167,N_6714);
and U13963 (N_13963,N_7478,N_9459);
and U13964 (N_13964,N_9174,N_11682);
xor U13965 (N_13965,N_12208,N_8233);
nand U13966 (N_13966,N_9834,N_10785);
and U13967 (N_13967,N_11796,N_10730);
or U13968 (N_13968,N_10692,N_10243);
and U13969 (N_13969,N_6292,N_10069);
nor U13970 (N_13970,N_7981,N_9012);
or U13971 (N_13971,N_10212,N_9927);
and U13972 (N_13972,N_8876,N_10268);
nor U13973 (N_13973,N_11839,N_10184);
or U13974 (N_13974,N_7094,N_7737);
xnor U13975 (N_13975,N_10544,N_11856);
nor U13976 (N_13976,N_9451,N_6876);
nor U13977 (N_13977,N_6848,N_11440);
or U13978 (N_13978,N_9471,N_6596);
and U13979 (N_13979,N_8431,N_7946);
nor U13980 (N_13980,N_8715,N_7407);
nand U13981 (N_13981,N_8496,N_11601);
and U13982 (N_13982,N_6329,N_11506);
nor U13983 (N_13983,N_11328,N_6891);
and U13984 (N_13984,N_11646,N_8461);
nor U13985 (N_13985,N_10633,N_9654);
nor U13986 (N_13986,N_11820,N_8685);
nor U13987 (N_13987,N_9605,N_10845);
nand U13988 (N_13988,N_11866,N_11651);
and U13989 (N_13989,N_6915,N_7797);
and U13990 (N_13990,N_6485,N_7151);
nor U13991 (N_13991,N_12251,N_8625);
and U13992 (N_13992,N_7667,N_11306);
or U13993 (N_13993,N_7793,N_8243);
and U13994 (N_13994,N_11881,N_6819);
and U13995 (N_13995,N_12144,N_9740);
nand U13996 (N_13996,N_7563,N_11493);
xnor U13997 (N_13997,N_8852,N_12107);
nor U13998 (N_13998,N_12028,N_7329);
nor U13999 (N_13999,N_6783,N_6642);
and U14000 (N_14000,N_11551,N_10804);
nand U14001 (N_14001,N_11962,N_8111);
and U14002 (N_14002,N_10440,N_9084);
nand U14003 (N_14003,N_10204,N_10493);
nand U14004 (N_14004,N_6944,N_11715);
xnor U14005 (N_14005,N_7291,N_7646);
nor U14006 (N_14006,N_8324,N_8740);
nor U14007 (N_14007,N_10168,N_7194);
nand U14008 (N_14008,N_7967,N_11950);
and U14009 (N_14009,N_11891,N_9247);
and U14010 (N_14010,N_9261,N_9052);
nor U14011 (N_14011,N_9095,N_7761);
and U14012 (N_14012,N_8633,N_9111);
nor U14013 (N_14013,N_12413,N_8203);
and U14014 (N_14014,N_10707,N_11842);
or U14015 (N_14015,N_9755,N_7027);
or U14016 (N_14016,N_7253,N_10515);
nor U14017 (N_14017,N_8932,N_6927);
or U14018 (N_14018,N_12194,N_10450);
nor U14019 (N_14019,N_9791,N_9186);
xnor U14020 (N_14020,N_9196,N_9475);
or U14021 (N_14021,N_8238,N_7175);
nor U14022 (N_14022,N_10098,N_8074);
nor U14023 (N_14023,N_12452,N_7968);
or U14024 (N_14024,N_8643,N_7469);
nor U14025 (N_14025,N_10592,N_7233);
and U14026 (N_14026,N_9268,N_11655);
nand U14027 (N_14027,N_6554,N_11229);
or U14028 (N_14028,N_10765,N_11783);
and U14029 (N_14029,N_6887,N_7750);
nor U14030 (N_14030,N_9573,N_11244);
nand U14031 (N_14031,N_7810,N_8489);
nand U14032 (N_14032,N_10876,N_11999);
nor U14033 (N_14033,N_9425,N_11834);
or U14034 (N_14034,N_9936,N_10762);
and U14035 (N_14035,N_11885,N_8487);
nand U14036 (N_14036,N_6623,N_10048);
xnor U14037 (N_14037,N_11937,N_11009);
nand U14038 (N_14038,N_10514,N_6924);
xnor U14039 (N_14039,N_10091,N_12313);
nor U14040 (N_14040,N_9149,N_8158);
nand U14041 (N_14041,N_9685,N_10382);
and U14042 (N_14042,N_10492,N_7849);
and U14043 (N_14043,N_11017,N_11449);
xnor U14044 (N_14044,N_8088,N_11903);
xnor U14045 (N_14045,N_6580,N_9018);
nand U14046 (N_14046,N_8757,N_6793);
xor U14047 (N_14047,N_8940,N_11752);
or U14048 (N_14048,N_7992,N_7853);
or U14049 (N_14049,N_12306,N_9943);
nor U14050 (N_14050,N_8307,N_11874);
and U14051 (N_14051,N_11418,N_7445);
nor U14052 (N_14052,N_11571,N_7455);
nand U14053 (N_14053,N_11841,N_7546);
nand U14054 (N_14054,N_7649,N_11349);
nand U14055 (N_14055,N_11339,N_10196);
nor U14056 (N_14056,N_11362,N_11572);
xor U14057 (N_14057,N_9106,N_12108);
or U14058 (N_14058,N_9798,N_11282);
nand U14059 (N_14059,N_9468,N_6932);
nand U14060 (N_14060,N_8704,N_9990);
nand U14061 (N_14061,N_11088,N_11246);
nor U14062 (N_14062,N_11049,N_11182);
nand U14063 (N_14063,N_10219,N_10975);
and U14064 (N_14064,N_8627,N_8000);
or U14065 (N_14065,N_10755,N_12114);
and U14066 (N_14066,N_7997,N_11718);
or U14067 (N_14067,N_8576,N_11606);
and U14068 (N_14068,N_7695,N_12419);
nand U14069 (N_14069,N_11600,N_6680);
or U14070 (N_14070,N_11675,N_6490);
nor U14071 (N_14071,N_8347,N_11054);
or U14072 (N_14072,N_10343,N_9950);
nand U14073 (N_14073,N_8706,N_11356);
or U14074 (N_14074,N_10791,N_7978);
nand U14075 (N_14075,N_7540,N_10467);
and U14076 (N_14076,N_8881,N_7140);
and U14077 (N_14077,N_10314,N_12151);
nand U14078 (N_14078,N_9659,N_11269);
nand U14079 (N_14079,N_7789,N_6398);
or U14080 (N_14080,N_10376,N_8773);
nor U14081 (N_14081,N_7712,N_7491);
nand U14082 (N_14082,N_8568,N_11617);
or U14083 (N_14083,N_8593,N_10311);
xnor U14084 (N_14084,N_9556,N_10222);
and U14085 (N_14085,N_8369,N_8240);
nor U14086 (N_14086,N_10678,N_8900);
and U14087 (N_14087,N_11797,N_8816);
nand U14088 (N_14088,N_8768,N_8414);
and U14089 (N_14089,N_12087,N_8295);
or U14090 (N_14090,N_11726,N_6277);
and U14091 (N_14091,N_10895,N_9511);
or U14092 (N_14092,N_10378,N_6647);
or U14093 (N_14093,N_8831,N_6913);
nor U14094 (N_14094,N_8650,N_9945);
and U14095 (N_14095,N_12098,N_11100);
nand U14096 (N_14096,N_7097,N_12230);
or U14097 (N_14097,N_9617,N_6278);
nand U14098 (N_14098,N_10335,N_10875);
and U14099 (N_14099,N_9296,N_10874);
or U14100 (N_14100,N_11959,N_11612);
and U14101 (N_14101,N_11940,N_7883);
or U14102 (N_14102,N_9579,N_7816);
nor U14103 (N_14103,N_10519,N_9498);
nand U14104 (N_14104,N_9726,N_9330);
nand U14105 (N_14105,N_8858,N_10183);
nand U14106 (N_14106,N_6391,N_9287);
nand U14107 (N_14107,N_10691,N_7108);
nor U14108 (N_14108,N_8692,N_11121);
or U14109 (N_14109,N_6323,N_6700);
nor U14110 (N_14110,N_8035,N_10530);
and U14111 (N_14111,N_7009,N_8265);
and U14112 (N_14112,N_11270,N_8320);
and U14113 (N_14113,N_10970,N_9331);
nor U14114 (N_14114,N_8016,N_6392);
nor U14115 (N_14115,N_11671,N_9133);
xor U14116 (N_14116,N_11996,N_9974);
and U14117 (N_14117,N_9243,N_10797);
and U14118 (N_14118,N_8677,N_8212);
or U14119 (N_14119,N_8490,N_6568);
nand U14120 (N_14120,N_9014,N_10324);
nand U14121 (N_14121,N_6477,N_8777);
or U14122 (N_14122,N_7332,N_11173);
nor U14123 (N_14123,N_11997,N_10309);
or U14124 (N_14124,N_12468,N_7196);
or U14125 (N_14125,N_9226,N_7734);
or U14126 (N_14126,N_9358,N_8721);
nor U14127 (N_14127,N_12075,N_7730);
xnor U14128 (N_14128,N_7820,N_8722);
nor U14129 (N_14129,N_11902,N_6551);
nand U14130 (N_14130,N_10328,N_6663);
or U14131 (N_14131,N_8168,N_11758);
and U14132 (N_14132,N_7755,N_8296);
nor U14133 (N_14133,N_11712,N_8574);
nor U14134 (N_14134,N_7148,N_11669);
or U14135 (N_14135,N_11623,N_7839);
nor U14136 (N_14136,N_8727,N_9340);
or U14137 (N_14137,N_9456,N_11166);
or U14138 (N_14138,N_6517,N_6732);
and U14139 (N_14139,N_9416,N_6833);
or U14140 (N_14140,N_7668,N_9270);
nor U14141 (N_14141,N_9876,N_10738);
or U14142 (N_14142,N_6669,N_6262);
xor U14143 (N_14143,N_6430,N_7063);
nand U14144 (N_14144,N_7837,N_8791);
or U14145 (N_14145,N_6779,N_11499);
xnor U14146 (N_14146,N_8539,N_11494);
nor U14147 (N_14147,N_9447,N_9115);
nand U14148 (N_14148,N_12450,N_9207);
or U14149 (N_14149,N_11253,N_6917);
nor U14150 (N_14150,N_8604,N_9509);
nand U14151 (N_14151,N_7069,N_12176);
nand U14152 (N_14152,N_9205,N_7150);
or U14153 (N_14153,N_10278,N_7006);
nor U14154 (N_14154,N_7246,N_7786);
nor U14155 (N_14155,N_9865,N_10122);
or U14156 (N_14156,N_6522,N_11086);
or U14157 (N_14157,N_10040,N_10100);
xnor U14158 (N_14158,N_12207,N_9750);
nand U14159 (N_14159,N_8389,N_11565);
nand U14160 (N_14160,N_9525,N_8969);
nand U14161 (N_14161,N_7725,N_9782);
xnor U14162 (N_14162,N_8926,N_12036);
xnor U14163 (N_14163,N_8614,N_10198);
nor U14164 (N_14164,N_8616,N_7601);
or U14165 (N_14165,N_6811,N_11450);
nor U14166 (N_14166,N_7457,N_10698);
and U14167 (N_14167,N_11003,N_7685);
or U14168 (N_14168,N_7259,N_7805);
and U14169 (N_14169,N_11558,N_9143);
nand U14170 (N_14170,N_11622,N_11197);
and U14171 (N_14171,N_12328,N_11119);
and U14172 (N_14172,N_7631,N_6908);
nand U14173 (N_14173,N_11954,N_11805);
nor U14174 (N_14174,N_11823,N_11849);
xnor U14175 (N_14175,N_8826,N_12184);
nand U14176 (N_14176,N_11425,N_6471);
nor U14177 (N_14177,N_7119,N_9363);
nand U14178 (N_14178,N_6636,N_9584);
and U14179 (N_14179,N_6672,N_7056);
xor U14180 (N_14180,N_10880,N_6921);
nand U14181 (N_14181,N_6620,N_8023);
or U14182 (N_14182,N_6753,N_6741);
xor U14183 (N_14183,N_7203,N_10722);
nor U14184 (N_14184,N_11397,N_8114);
xnor U14185 (N_14185,N_12053,N_6476);
nand U14186 (N_14186,N_7741,N_11867);
and U14187 (N_14187,N_6943,N_8255);
nor U14188 (N_14188,N_7085,N_9621);
xnor U14189 (N_14189,N_12432,N_10621);
nand U14190 (N_14190,N_12278,N_9979);
nor U14191 (N_14191,N_6792,N_9298);
or U14192 (N_14192,N_11436,N_11471);
nor U14193 (N_14193,N_8651,N_6934);
nor U14194 (N_14194,N_9368,N_9695);
and U14195 (N_14195,N_6317,N_9719);
or U14196 (N_14196,N_12119,N_8303);
or U14197 (N_14197,N_9313,N_10630);
nand U14198 (N_14198,N_9826,N_9553);
or U14199 (N_14199,N_6261,N_8213);
nor U14200 (N_14200,N_8332,N_6638);
or U14201 (N_14201,N_7660,N_8385);
or U14202 (N_14202,N_9614,N_10878);
nand U14203 (N_14203,N_8040,N_6990);
or U14204 (N_14204,N_8264,N_8354);
and U14205 (N_14205,N_8503,N_7192);
nor U14206 (N_14206,N_9382,N_9730);
nor U14207 (N_14207,N_9113,N_9449);
xor U14208 (N_14208,N_8513,N_10655);
nand U14209 (N_14209,N_12245,N_6910);
and U14210 (N_14210,N_8533,N_9396);
nand U14211 (N_14211,N_8492,N_6285);
and U14212 (N_14212,N_7066,N_12057);
nor U14213 (N_14213,N_8298,N_10677);
or U14214 (N_14214,N_10033,N_11373);
nor U14215 (N_14215,N_6737,N_8267);
nand U14216 (N_14216,N_9367,N_8601);
and U14217 (N_14217,N_7764,N_12399);
xnor U14218 (N_14218,N_11448,N_8902);
xnor U14219 (N_14219,N_8910,N_10685);
or U14220 (N_14220,N_9986,N_8942);
nand U14221 (N_14221,N_11746,N_12312);
nor U14222 (N_14222,N_11833,N_9103);
xnor U14223 (N_14223,N_6770,N_11644);
and U14224 (N_14224,N_6396,N_10149);
and U14225 (N_14225,N_9203,N_9005);
nor U14226 (N_14226,N_6462,N_8362);
nand U14227 (N_14227,N_6545,N_6835);
xnor U14228 (N_14228,N_8128,N_11420);
or U14229 (N_14229,N_10932,N_11748);
or U14230 (N_14230,N_9564,N_12115);
or U14231 (N_14231,N_6614,N_9714);
nor U14232 (N_14232,N_10897,N_8308);
or U14233 (N_14233,N_12345,N_8073);
nand U14234 (N_14234,N_7662,N_8765);
or U14235 (N_14235,N_7334,N_9513);
nand U14236 (N_14236,N_8037,N_9607);
nor U14237 (N_14237,N_7847,N_11377);
nand U14238 (N_14238,N_7435,N_10937);
xnor U14239 (N_14239,N_10626,N_11705);
or U14240 (N_14240,N_11693,N_7551);
xnor U14241 (N_14241,N_9344,N_7731);
nor U14242 (N_14242,N_10659,N_12453);
nor U14243 (N_14243,N_10540,N_6780);
and U14244 (N_14244,N_11006,N_10657);
nand U14245 (N_14245,N_8198,N_6602);
or U14246 (N_14246,N_9920,N_6481);
nor U14247 (N_14247,N_10427,N_10215);
nor U14248 (N_14248,N_8793,N_10050);
nand U14249 (N_14249,N_10087,N_9906);
or U14250 (N_14250,N_11794,N_6865);
xnor U14251 (N_14251,N_10027,N_10464);
nor U14252 (N_14252,N_7706,N_7941);
nor U14253 (N_14253,N_8686,N_6276);
and U14254 (N_14254,N_12465,N_7595);
nand U14255 (N_14255,N_6748,N_6736);
nand U14256 (N_14256,N_12263,N_8579);
nand U14257 (N_14257,N_10954,N_6937);
nor U14258 (N_14258,N_11592,N_8440);
nand U14259 (N_14259,N_7889,N_6321);
nor U14260 (N_14260,N_11459,N_12350);
nand U14261 (N_14261,N_11358,N_8391);
or U14262 (N_14262,N_8571,N_6796);
or U14263 (N_14263,N_7916,N_10930);
nor U14264 (N_14264,N_8833,N_9736);
nor U14265 (N_14265,N_6810,N_8753);
or U14266 (N_14266,N_6852,N_11588);
xor U14267 (N_14267,N_9433,N_9967);
nand U14268 (N_14268,N_6271,N_11627);
and U14269 (N_14269,N_12478,N_7807);
xnor U14270 (N_14270,N_9458,N_7785);
xor U14271 (N_14271,N_11095,N_9132);
xnor U14272 (N_14272,N_10555,N_9890);
and U14273 (N_14273,N_11315,N_9540);
nand U14274 (N_14274,N_10077,N_12449);
nand U14275 (N_14275,N_7523,N_8745);
or U14276 (N_14276,N_8901,N_11193);
nand U14277 (N_14277,N_8478,N_9809);
or U14278 (N_14278,N_6967,N_9202);
and U14279 (N_14279,N_12095,N_9737);
and U14280 (N_14280,N_6813,N_7815);
nor U14281 (N_14281,N_8919,N_11165);
nand U14282 (N_14282,N_9851,N_12458);
nand U14283 (N_14283,N_6525,N_6752);
nor U14284 (N_14284,N_7146,N_10673);
nand U14285 (N_14285,N_9079,N_10834);
nand U14286 (N_14286,N_6655,N_10877);
nand U14287 (N_14287,N_8050,N_11353);
nor U14288 (N_14288,N_11048,N_7635);
or U14289 (N_14289,N_9602,N_7801);
nand U14290 (N_14290,N_8668,N_9505);
nand U14291 (N_14291,N_6787,N_7576);
nand U14292 (N_14292,N_7482,N_12337);
and U14293 (N_14293,N_11692,N_9096);
and U14294 (N_14294,N_12055,N_12430);
and U14295 (N_14295,N_10669,N_8807);
nor U14296 (N_14296,N_9128,N_10957);
nor U14297 (N_14297,N_6740,N_10500);
nor U14298 (N_14298,N_9137,N_11978);
and U14299 (N_14299,N_12368,N_7229);
or U14300 (N_14300,N_10865,N_11585);
or U14301 (N_14301,N_11607,N_7747);
and U14302 (N_14302,N_9142,N_9429);
or U14303 (N_14303,N_7156,N_8945);
nand U14304 (N_14304,N_8426,N_11016);
or U14305 (N_14305,N_6729,N_7128);
nor U14306 (N_14306,N_6605,N_9315);
or U14307 (N_14307,N_9073,N_10542);
and U14308 (N_14308,N_7104,N_6593);
nand U14309 (N_14309,N_12457,N_9217);
or U14310 (N_14310,N_12441,N_11570);
xor U14311 (N_14311,N_12025,N_11800);
and U14312 (N_14312,N_12018,N_8124);
and U14313 (N_14313,N_12377,N_12205);
nand U14314 (N_14314,N_8608,N_12250);
or U14315 (N_14315,N_6301,N_11400);
and U14316 (N_14316,N_10251,N_11863);
and U14317 (N_14317,N_12229,N_11875);
and U14318 (N_14318,N_9394,N_11504);
nand U14319 (N_14319,N_8215,N_7880);
nor U14320 (N_14320,N_7073,N_8022);
and U14321 (N_14321,N_7814,N_9482);
nor U14322 (N_14322,N_10331,N_6374);
nand U14323 (N_14323,N_8803,N_11596);
xor U14324 (N_14324,N_7912,N_12219);
and U14325 (N_14325,N_10565,N_9850);
xnor U14326 (N_14326,N_11392,N_11549);
or U14327 (N_14327,N_12035,N_6683);
xor U14328 (N_14328,N_8994,N_11140);
nand U14329 (N_14329,N_8709,N_11538);
nand U14330 (N_14330,N_6897,N_8699);
nand U14331 (N_14331,N_10803,N_9090);
and U14332 (N_14332,N_12181,N_6534);
nand U14333 (N_14333,N_12180,N_11777);
or U14334 (N_14334,N_10676,N_6721);
xnor U14335 (N_14335,N_8961,N_6654);
xnor U14336 (N_14336,N_9033,N_11691);
nand U14337 (N_14337,N_6776,N_11769);
nor U14338 (N_14338,N_11428,N_11515);
nor U14339 (N_14339,N_12179,N_9279);
nor U14340 (N_14340,N_10581,N_8894);
and U14341 (N_14341,N_10591,N_7453);
nor U14342 (N_14342,N_8425,N_10216);
or U14343 (N_14343,N_11464,N_12105);
xnor U14344 (N_14344,N_6677,N_7387);
or U14345 (N_14345,N_11271,N_9512);
nor U14346 (N_14346,N_8841,N_12139);
nand U14347 (N_14347,N_10564,N_8500);
or U14348 (N_14348,N_10185,N_9155);
nand U14349 (N_14349,N_10959,N_6805);
nand U14350 (N_14350,N_11169,N_7365);
and U14351 (N_14351,N_11188,N_8936);
or U14352 (N_14352,N_10745,N_7313);
and U14353 (N_14353,N_9541,N_11268);
nand U14354 (N_14354,N_9626,N_7489);
nand U14355 (N_14355,N_12320,N_7350);
or U14356 (N_14356,N_8814,N_7371);
nor U14357 (N_14357,N_12274,N_11032);
nand U14358 (N_14358,N_7288,N_7249);
nor U14359 (N_14359,N_8560,N_10262);
nor U14360 (N_14360,N_10963,N_8529);
nor U14361 (N_14361,N_12310,N_9359);
xnor U14362 (N_14362,N_11780,N_6299);
nand U14363 (N_14363,N_12472,N_9385);
nor U14364 (N_14364,N_8801,N_9954);
nand U14365 (N_14365,N_8139,N_11228);
or U14366 (N_14366,N_8145,N_8495);
nand U14367 (N_14367,N_8288,N_6960);
nor U14368 (N_14368,N_11323,N_11772);
nor U14369 (N_14369,N_11025,N_8417);
xor U14370 (N_14370,N_6899,N_7799);
or U14371 (N_14371,N_6949,N_10239);
and U14372 (N_14372,N_7188,N_6563);
nand U14373 (N_14373,N_9083,N_10951);
nor U14374 (N_14374,N_9562,N_6466);
and U14375 (N_14375,N_8982,N_8967);
nor U14376 (N_14376,N_8796,N_10453);
nor U14377 (N_14377,N_12003,N_9923);
nand U14378 (N_14378,N_7557,N_6892);
nor U14379 (N_14379,N_7400,N_12294);
nand U14380 (N_14380,N_8895,N_8072);
nand U14381 (N_14381,N_10012,N_12403);
nand U14382 (N_14382,N_6293,N_10159);
nor U14383 (N_14383,N_6709,N_10080);
or U14384 (N_14384,N_10229,N_9500);
nor U14385 (N_14385,N_10812,N_10898);
or U14386 (N_14386,N_8845,N_8862);
or U14387 (N_14387,N_11687,N_7525);
or U14388 (N_14388,N_9465,N_11614);
or U14389 (N_14389,N_11334,N_12427);
or U14390 (N_14390,N_9097,N_6343);
nand U14391 (N_14391,N_7986,N_6449);
and U14392 (N_14392,N_6346,N_7125);
nor U14393 (N_14393,N_11079,N_6657);
and U14394 (N_14394,N_11672,N_11946);
nand U14395 (N_14395,N_10083,N_7101);
and U14396 (N_14396,N_9055,N_12091);
nand U14397 (N_14397,N_6963,N_10558);
or U14398 (N_14398,N_11141,N_7380);
xor U14399 (N_14399,N_9538,N_11128);
and U14400 (N_14400,N_11256,N_7240);
and U14401 (N_14401,N_11689,N_8750);
or U14402 (N_14402,N_7644,N_9081);
or U14403 (N_14403,N_6809,N_7724);
or U14404 (N_14404,N_8542,N_9604);
xor U14405 (N_14405,N_10760,N_6689);
and U14406 (N_14406,N_6579,N_6651);
nor U14407 (N_14407,N_11922,N_10414);
and U14408 (N_14408,N_11340,N_10885);
nand U14409 (N_14409,N_8938,N_10924);
nor U14410 (N_14410,N_6436,N_10794);
and U14411 (N_14411,N_12030,N_9238);
nor U14412 (N_14412,N_9345,N_7147);
xnor U14413 (N_14413,N_8491,N_6496);
nand U14414 (N_14414,N_10366,N_6604);
nor U14415 (N_14415,N_6312,N_10588);
nor U14416 (N_14416,N_9616,N_8836);
nor U14417 (N_14417,N_7458,N_8130);
or U14418 (N_14418,N_10742,N_7619);
and U14419 (N_14419,N_11480,N_6339);
nand U14420 (N_14420,N_12404,N_8646);
or U14421 (N_14421,N_8196,N_12143);
nor U14422 (N_14422,N_12078,N_9536);
or U14423 (N_14423,N_9126,N_11097);
nor U14424 (N_14424,N_8630,N_12473);
nor U14425 (N_14425,N_9764,N_10399);
nand U14426 (N_14426,N_10320,N_10085);
nor U14427 (N_14427,N_11051,N_11563);
nand U14428 (N_14428,N_11804,N_6468);
xnor U14429 (N_14429,N_8688,N_12074);
nand U14430 (N_14430,N_7112,N_12129);
nand U14431 (N_14431,N_9057,N_12348);
or U14432 (N_14432,N_11782,N_12133);
nand U14433 (N_14433,N_9388,N_11380);
xor U14434 (N_14434,N_11443,N_8597);
nand U14435 (N_14435,N_7527,N_8186);
nand U14436 (N_14436,N_10004,N_8526);
and U14437 (N_14437,N_7344,N_9753);
nand U14438 (N_14438,N_9402,N_8511);
nor U14439 (N_14439,N_11930,N_10606);
nor U14440 (N_14440,N_12499,N_11294);
nand U14441 (N_14441,N_7932,N_7517);
nand U14442 (N_14442,N_7841,N_11083);
and U14443 (N_14443,N_7325,N_9678);
xnor U14444 (N_14444,N_7323,N_6665);
or U14445 (N_14445,N_9586,N_11517);
nor U14446 (N_14446,N_8952,N_6997);
and U14447 (N_14447,N_12109,N_10849);
xnor U14448 (N_14448,N_8420,N_10631);
and U14449 (N_14449,N_11251,N_9672);
nand U14450 (N_14450,N_6613,N_8485);
and U14451 (N_14451,N_7198,N_8387);
and U14452 (N_14452,N_9408,N_12258);
and U14453 (N_14453,N_9348,N_8018);
and U14454 (N_14454,N_12282,N_7190);
nor U14455 (N_14455,N_6378,N_12047);
nor U14456 (N_14456,N_7342,N_6523);
xnor U14457 (N_14457,N_10532,N_7875);
nor U14458 (N_14458,N_10840,N_10920);
xor U14459 (N_14459,N_7790,N_11550);
xor U14460 (N_14460,N_12054,N_12370);
or U14461 (N_14461,N_9015,N_11295);
or U14462 (N_14462,N_8206,N_12060);
nand U14463 (N_14463,N_11921,N_9183);
nand U14464 (N_14464,N_11942,N_9922);
nand U14465 (N_14465,N_12264,N_8913);
nor U14466 (N_14466,N_11184,N_9259);
nor U14467 (N_14467,N_8874,N_11072);
and U14468 (N_14468,N_9170,N_11840);
and U14469 (N_14469,N_12068,N_6535);
xnor U14470 (N_14470,N_8596,N_6530);
or U14471 (N_14471,N_9281,N_9966);
nor U14472 (N_14472,N_12287,N_12329);
nand U14473 (N_14473,N_9907,N_10737);
or U14474 (N_14474,N_8788,N_6971);
nand U14475 (N_14475,N_10142,N_12056);
nor U14476 (N_14476,N_11745,N_10520);
and U14477 (N_14477,N_8443,N_6936);
and U14478 (N_14478,N_11575,N_12493);
or U14479 (N_14479,N_9153,N_8501);
nand U14480 (N_14480,N_11454,N_6397);
and U14481 (N_14481,N_7545,N_10454);
or U14482 (N_14482,N_10611,N_12382);
or U14483 (N_14483,N_6708,N_6412);
nand U14484 (N_14484,N_7446,N_7977);
or U14485 (N_14485,N_11831,N_11158);
and U14486 (N_14486,N_9302,N_9035);
nand U14487 (N_14487,N_8632,N_7483);
nor U14488 (N_14488,N_11200,N_6650);
xor U14489 (N_14489,N_9286,N_8330);
and U14490 (N_14490,N_8522,N_8482);
nand U14491 (N_14491,N_7907,N_12356);
nor U14492 (N_14492,N_8488,N_9338);
nand U14493 (N_14493,N_9130,N_6675);
nor U14494 (N_14494,N_8822,N_8319);
nor U14495 (N_14495,N_9146,N_9099);
xnor U14496 (N_14496,N_11181,N_7077);
or U14497 (N_14497,N_9138,N_11363);
and U14498 (N_14498,N_8628,N_9611);
nand U14499 (N_14499,N_6492,N_9222);
nand U14500 (N_14500,N_9592,N_11408);
nand U14501 (N_14501,N_10837,N_7016);
nor U14502 (N_14502,N_11662,N_10933);
or U14503 (N_14503,N_10505,N_9326);
and U14504 (N_14504,N_7245,N_10412);
or U14505 (N_14505,N_9339,N_6939);
and U14506 (N_14506,N_10764,N_11287);
and U14507 (N_14507,N_10228,N_7310);
nand U14508 (N_14508,N_12188,N_9154);
xor U14509 (N_14509,N_12031,N_7356);
nor U14510 (N_14510,N_6379,N_6434);
xnor U14511 (N_14511,N_6612,N_8778);
and U14512 (N_14512,N_7928,N_11910);
or U14513 (N_14513,N_10202,N_11743);
nand U14514 (N_14514,N_6893,N_10828);
and U14515 (N_14515,N_10964,N_11481);
or U14516 (N_14516,N_12421,N_11593);
nand U14517 (N_14517,N_9373,N_10365);
or U14518 (N_14518,N_6253,N_12420);
and U14519 (N_14519,N_10841,N_7040);
and U14520 (N_14520,N_10358,N_7257);
nor U14521 (N_14521,N_7699,N_11642);
xor U14522 (N_14522,N_10072,N_11759);
xor U14523 (N_14523,N_12017,N_10556);
or U14524 (N_14524,N_10640,N_8873);
or U14525 (N_14525,N_9322,N_10497);
or U14526 (N_14526,N_10443,N_9478);
and U14527 (N_14527,N_9022,N_12374);
nand U14528 (N_14528,N_10076,N_6386);
or U14529 (N_14529,N_6673,N_7602);
xor U14530 (N_14530,N_9989,N_11514);
nand U14531 (N_14531,N_11028,N_10919);
nor U14532 (N_14532,N_10643,N_10790);
nor U14533 (N_14533,N_10976,N_8660);
and U14534 (N_14534,N_9651,N_6895);
nand U14535 (N_14535,N_7498,N_12343);
and U14536 (N_14536,N_7444,N_9414);
nand U14537 (N_14537,N_10826,N_9024);
and U14538 (N_14538,N_10987,N_11734);
or U14539 (N_14539,N_10191,N_8675);
or U14540 (N_14540,N_7386,N_11143);
nand U14541 (N_14541,N_9430,N_10744);
nand U14542 (N_14542,N_9570,N_11534);
xnor U14543 (N_14543,N_10700,N_9855);
and U14544 (N_14544,N_12094,N_9612);
and U14545 (N_14545,N_10201,N_11343);
and U14546 (N_14546,N_11093,N_7893);
and U14547 (N_14547,N_10022,N_8759);
xor U14548 (N_14548,N_6325,N_10503);
and U14549 (N_14549,N_11219,N_7277);
or U14550 (N_14550,N_11254,N_9758);
nand U14551 (N_14551,N_6255,N_8046);
and U14552 (N_14552,N_11897,N_11085);
xor U14553 (N_14553,N_9859,N_8148);
nand U14554 (N_14554,N_11103,N_6265);
and U14555 (N_14555,N_10524,N_9411);
nand U14556 (N_14556,N_6847,N_7748);
nand U14557 (N_14557,N_8726,N_10092);
nand U14558 (N_14558,N_10817,N_11167);
and U14559 (N_14559,N_7440,N_10287);
nor U14560 (N_14560,N_12395,N_11080);
or U14561 (N_14561,N_10582,N_7452);
nor U14562 (N_14562,N_11151,N_11035);
nor U14563 (N_14563,N_10003,N_8224);
nor U14564 (N_14564,N_10136,N_12376);
xnor U14565 (N_14565,N_9377,N_11749);
nand U14566 (N_14566,N_12372,N_8621);
nand U14567 (N_14567,N_7004,N_8336);
nand U14568 (N_14568,N_8659,N_9856);
xnor U14569 (N_14569,N_11925,N_12168);
or U14570 (N_14570,N_6874,N_10441);
and U14571 (N_14571,N_11422,N_12118);
and U14572 (N_14572,N_12200,N_12290);
xnor U14573 (N_14573,N_10336,N_7638);
and U14574 (N_14574,N_9897,N_8329);
nor U14575 (N_14575,N_7558,N_6781);
or U14576 (N_14576,N_6370,N_8144);
nor U14577 (N_14577,N_9362,N_8449);
xnor U14578 (N_14578,N_9832,N_9811);
or U14579 (N_14579,N_12387,N_8014);
nor U14580 (N_14580,N_12408,N_6801);
nand U14581 (N_14581,N_8012,N_11843);
or U14582 (N_14582,N_7155,N_6403);
nand U14583 (N_14583,N_8587,N_10379);
xor U14584 (N_14584,N_6766,N_11793);
nand U14585 (N_14585,N_7661,N_12461);
or U14586 (N_14586,N_11806,N_6742);
nor U14587 (N_14587,N_6898,N_7303);
nor U14588 (N_14588,N_10939,N_7681);
or U14589 (N_14589,N_8268,N_11864);
nand U14590 (N_14590,N_10968,N_11034);
or U14591 (N_14591,N_7111,N_9803);
nor U14592 (N_14592,N_11490,N_10250);
nand U14593 (N_14593,N_10642,N_8975);
or U14594 (N_14594,N_6537,N_6974);
nor U14595 (N_14595,N_7927,N_6532);
nor U14596 (N_14596,N_7840,N_7702);
and U14597 (N_14597,N_10910,N_7395);
and U14598 (N_14598,N_10538,N_10560);
nand U14599 (N_14599,N_7224,N_9420);
and U14600 (N_14600,N_7812,N_11787);
and U14601 (N_14601,N_6303,N_8662);
and U14602 (N_14602,N_9867,N_7065);
or U14603 (N_14603,N_11890,N_10586);
or U14604 (N_14604,N_8976,N_7656);
nand U14605 (N_14605,N_7434,N_11915);
and U14606 (N_14606,N_9706,N_10326);
or U14607 (N_14607,N_10997,N_9474);
nand U14608 (N_14608,N_10928,N_7819);
nor U14609 (N_14609,N_10321,N_9164);
xnor U14610 (N_14610,N_11272,N_7182);
or U14611 (N_14611,N_9701,N_6701);
nor U14612 (N_14612,N_7109,N_9058);
or U14613 (N_14613,N_11928,N_12011);
or U14614 (N_14614,N_9899,N_9996);
or U14615 (N_14615,N_9881,N_7488);
and U14616 (N_14616,N_12439,N_6407);
or U14617 (N_14617,N_9162,N_7994);
nand U14618 (N_14618,N_12186,N_12007);
or U14619 (N_14619,N_11441,N_7348);
nand U14620 (N_14620,N_11512,N_10189);
or U14621 (N_14621,N_10023,N_8087);
and U14622 (N_14622,N_9094,N_9294);
or U14623 (N_14623,N_10991,N_7759);
nor U14624 (N_14624,N_9623,N_8095);
and U14625 (N_14625,N_8870,N_12112);
or U14626 (N_14626,N_9709,N_11889);
nor U14627 (N_14627,N_12424,N_9528);
and U14628 (N_14628,N_6919,N_9104);
nor U14629 (N_14629,N_11567,N_8929);
nand U14630 (N_14630,N_6319,N_7438);
or U14631 (N_14631,N_6336,N_6446);
or U14632 (N_14632,N_10302,N_6342);
nand U14633 (N_14633,N_8376,N_10203);
and U14634 (N_14634,N_9697,N_8592);
and U14635 (N_14635,N_6959,N_9469);
and U14636 (N_14636,N_9558,N_10906);
nor U14637 (N_14637,N_10921,N_10115);
or U14638 (N_14638,N_10064,N_6635);
or U14639 (N_14639,N_7513,N_8676);
nand U14640 (N_14640,N_6839,N_11597);
or U14641 (N_14641,N_10981,N_9098);
nand U14642 (N_14642,N_8034,N_8393);
nand U14643 (N_14643,N_10051,N_8683);
xnor U14644 (N_14644,N_10451,N_7548);
nand U14645 (N_14645,N_6617,N_6912);
nand U14646 (N_14646,N_6304,N_8665);
nand U14647 (N_14647,N_12317,N_10721);
and U14648 (N_14648,N_10325,N_10571);
nor U14649 (N_14649,N_7530,N_9772);
and U14650 (N_14650,N_7235,N_7767);
nor U14651 (N_14651,N_10683,N_11904);
and U14652 (N_14652,N_10625,N_9515);
nand U14653 (N_14653,N_9192,N_8989);
or U14654 (N_14654,N_8189,N_7580);
xnor U14655 (N_14655,N_10143,N_8011);
and U14656 (N_14656,N_7423,N_11159);
and U14657 (N_14657,N_10120,N_10545);
nand U14658 (N_14658,N_9019,N_9386);
nand U14659 (N_14659,N_11430,N_8091);
or U14660 (N_14660,N_10725,N_10516);
xor U14661 (N_14661,N_8483,N_6440);
or U14662 (N_14662,N_9177,N_6425);
and U14663 (N_14663,N_9580,N_8820);
and U14664 (N_14664,N_6706,N_6264);
nand U14665 (N_14665,N_8575,N_8476);
and U14666 (N_14666,N_7677,N_10390);
and U14667 (N_14667,N_9748,N_7353);
xnor U14668 (N_14668,N_11755,N_10511);
or U14669 (N_14669,N_10327,N_10650);
nand U14670 (N_14670,N_9078,N_9034);
and U14671 (N_14671,N_11975,N_8122);
nor U14672 (N_14672,N_11039,N_10110);
or U14673 (N_14673,N_10177,N_9224);
or U14674 (N_14674,N_6333,N_12092);
nand U14675 (N_14675,N_8705,N_8278);
and U14676 (N_14676,N_10485,N_11384);
and U14677 (N_14677,N_7529,N_8510);
or U14678 (N_14678,N_10269,N_11447);
nor U14679 (N_14679,N_10341,N_12444);
nand U14680 (N_14680,N_10078,N_10285);
nor U14681 (N_14681,N_8176,N_9559);
or U14682 (N_14682,N_10686,N_7183);
and U14683 (N_14683,N_8056,N_7208);
nor U14684 (N_14684,N_12089,N_8528);
nand U14685 (N_14685,N_6377,N_10224);
and U14686 (N_14686,N_6637,N_11429);
nand U14687 (N_14687,N_10871,N_6954);
and U14688 (N_14688,N_10165,N_8626);
nor U14689 (N_14689,N_10416,N_12446);
nand U14690 (N_14690,N_11201,N_10562);
and U14691 (N_14691,N_11215,N_9353);
nor U14692 (N_14692,N_7925,N_9905);
nor U14693 (N_14693,N_8353,N_10283);
and U14694 (N_14694,N_12422,N_7184);
xnor U14695 (N_14695,N_6375,N_8005);
or U14696 (N_14696,N_10462,N_6854);
or U14697 (N_14697,N_7634,N_7980);
nor U14698 (N_14698,N_10862,N_8847);
xnor U14699 (N_14699,N_6409,N_6438);
nor U14700 (N_14700,N_11178,N_9648);
nor U14701 (N_14701,N_6540,N_9639);
and U14702 (N_14702,N_7779,N_10405);
or U14703 (N_14703,N_11127,N_12259);
and U14704 (N_14704,N_9941,N_7852);
nor U14705 (N_14705,N_12373,N_12388);
nand U14706 (N_14706,N_9842,N_8636);
nand U14707 (N_14707,N_8048,N_11198);
and U14708 (N_14708,N_11580,N_6524);
nand U14709 (N_14709,N_9557,N_11102);
nand U14710 (N_14710,N_11767,N_12365);
nand U14711 (N_14711,N_10597,N_6666);
or U14712 (N_14712,N_7191,N_7165);
and U14713 (N_14713,N_6550,N_11037);
or U14714 (N_14714,N_10961,N_7352);
nand U14715 (N_14715,N_7437,N_8249);
nor U14716 (N_14716,N_12277,N_7247);
nor U14717 (N_14717,N_11238,N_9657);
or U14718 (N_14718,N_6447,N_10221);
xnor U14719 (N_14719,N_9705,N_8566);
xor U14720 (N_14720,N_9365,N_7583);
nand U14721 (N_14721,N_11552,N_6382);
and U14722 (N_14722,N_8647,N_10466);
nor U14723 (N_14723,N_10839,N_6747);
nand U14724 (N_14724,N_6495,N_12412);
or U14725 (N_14725,N_9280,N_7827);
nand U14726 (N_14726,N_7973,N_9609);
or U14727 (N_14727,N_9088,N_7064);
or U14728 (N_14728,N_6399,N_7831);
and U14729 (N_14729,N_9952,N_7511);
nand U14730 (N_14730,N_9212,N_11667);
and U14731 (N_14731,N_12195,N_7217);
and U14732 (N_14732,N_12340,N_12354);
xor U14733 (N_14733,N_8949,N_9004);
nor U14734 (N_14734,N_11663,N_11369);
and U14735 (N_14735,N_8322,N_9760);
nor U14736 (N_14736,N_7738,N_8871);
xnor U14737 (N_14737,N_12291,N_8118);
nand U14738 (N_14738,N_7337,N_11375);
nor U14739 (N_14739,N_10267,N_11952);
nand U14740 (N_14740,N_6686,N_7886);
nand U14741 (N_14741,N_9818,N_9895);
nor U14742 (N_14742,N_7769,N_8341);
and U14743 (N_14743,N_10601,N_8287);
or U14744 (N_14744,N_12381,N_8008);
nand U14745 (N_14745,N_11986,N_7228);
nor U14746 (N_14746,N_8182,N_11239);
or U14747 (N_14747,N_10644,N_10279);
nor U14748 (N_14748,N_8090,N_6587);
nand U14749 (N_14749,N_10075,N_12231);
xor U14750 (N_14750,N_8946,N_11896);
and U14751 (N_14751,N_10470,N_11312);
or U14752 (N_14752,N_10284,N_7694);
nand U14753 (N_14753,N_8419,N_10670);
or U14754 (N_14754,N_6335,N_9077);
nor U14755 (N_14755,N_12008,N_11711);
nor U14756 (N_14756,N_8301,N_11012);
nand U14757 (N_14757,N_10455,N_11507);
nor U14758 (N_14758,N_11982,N_6561);
nand U14759 (N_14759,N_6592,N_11314);
nor U14760 (N_14760,N_8479,N_8077);
or U14761 (N_14761,N_8635,N_12362);
and U14762 (N_14762,N_7589,N_9157);
nand U14763 (N_14763,N_6318,N_9869);
or U14764 (N_14764,N_8475,N_9250);
and U14765 (N_14765,N_9774,N_11602);
or U14766 (N_14766,N_11485,N_11649);
and U14767 (N_14767,N_7885,N_8105);
nand U14768 (N_14768,N_10672,N_8546);
nor U14769 (N_14769,N_6724,N_7302);
nor U14770 (N_14770,N_10353,N_6320);
xor U14771 (N_14771,N_8719,N_7470);
or U14772 (N_14772,N_7338,N_11424);
and U14773 (N_14773,N_8291,N_8790);
and U14774 (N_14774,N_12299,N_10337);
or U14775 (N_14775,N_9969,N_9037);
nand U14776 (N_14776,N_12492,N_7205);
nand U14777 (N_14777,N_7116,N_9814);
nand U14778 (N_14778,N_8525,N_7773);
and U14779 (N_14779,N_6474,N_6679);
nand U14780 (N_14780,N_9354,N_7413);
and U14781 (N_14781,N_10190,N_10952);
nand U14782 (N_14782,N_10578,N_10127);
nand U14783 (N_14783,N_12210,N_9288);
or U14784 (N_14784,N_11945,N_7754);
nor U14785 (N_14785,N_10926,N_9642);
and U14786 (N_14786,N_10486,N_9827);
nand U14787 (N_14787,N_7666,N_9007);
nand U14788 (N_14788,N_9961,N_6656);
or U14789 (N_14789,N_10602,N_10116);
xnor U14790 (N_14790,N_8941,N_6585);
or U14791 (N_14791,N_10084,N_9325);
nand U14792 (N_14792,N_9619,N_6883);
or U14793 (N_14793,N_12237,N_11432);
nand U14794 (N_14794,N_11557,N_11382);
and U14795 (N_14795,N_10548,N_10360);
or U14796 (N_14796,N_7441,N_10821);
and U14797 (N_14797,N_11728,N_9428);
or U14798 (N_14798,N_8612,N_11478);
nor U14799 (N_14799,N_8654,N_10141);
or U14800 (N_14800,N_9844,N_9401);
and U14801 (N_14801,N_6566,N_7033);
and U14802 (N_14802,N_7632,N_12142);
and U14803 (N_14803,N_9043,N_10129);
and U14804 (N_14804,N_7389,N_8766);
or U14805 (N_14805,N_6256,N_12002);
nor U14806 (N_14806,N_8364,N_7177);
nor U14807 (N_14807,N_10113,N_9924);
nor U14808 (N_14808,N_6633,N_11893);
xnor U14809 (N_14809,N_8254,N_8619);
or U14810 (N_14810,N_9506,N_9333);
or U14811 (N_14811,N_9248,N_6947);
or U14812 (N_14812,N_11291,N_7143);
or U14813 (N_14813,N_11218,N_9236);
nor U14814 (N_14814,N_10893,N_8027);
and U14815 (N_14815,N_11216,N_7226);
or U14816 (N_14816,N_11898,N_7447);
and U14817 (N_14817,N_8747,N_6450);
or U14818 (N_14818,N_9670,N_7475);
and U14819 (N_14819,N_10747,N_6369);
and U14820 (N_14820,N_6825,N_9189);
nand U14821 (N_14821,N_9114,N_7122);
nor U14822 (N_14822,N_6280,N_9185);
xnor U14823 (N_14823,N_10767,N_7273);
nand U14824 (N_14824,N_9371,N_12111);
nor U14825 (N_14825,N_7550,N_7038);
nor U14826 (N_14826,N_10153,N_10208);
or U14827 (N_14827,N_10600,N_8730);
or U14828 (N_14828,N_6888,N_9862);
nand U14829 (N_14829,N_9999,N_7241);
and U14830 (N_14830,N_9915,N_9290);
and U14831 (N_14831,N_12247,N_11242);
nand U14832 (N_14832,N_6559,N_11346);
or U14833 (N_14833,N_6859,N_7948);
or U14834 (N_14834,N_8226,N_11763);
xor U14835 (N_14835,N_11189,N_7582);
and U14836 (N_14836,N_8237,N_11813);
nor U14837 (N_14837,N_8477,N_7693);
nand U14838 (N_14838,N_6300,N_7409);
and U14839 (N_14839,N_9776,N_11868);
xor U14840 (N_14840,N_9718,N_10748);
nand U14841 (N_14841,N_9683,N_11013);
and U14842 (N_14842,N_10247,N_6978);
nor U14843 (N_14843,N_6653,N_6542);
nor U14844 (N_14844,N_11533,N_8081);
or U14845 (N_14845,N_9773,N_6640);
nand U14846 (N_14846,N_7556,N_6958);
and U14847 (N_14847,N_6703,N_9025);
nand U14848 (N_14848,N_8151,N_8175);
or U14849 (N_14849,N_8992,N_8789);
or U14850 (N_14850,N_10264,N_9606);
nand U14851 (N_14851,N_9780,N_7275);
and U14852 (N_14852,N_10879,N_10536);
nand U14853 (N_14853,N_10843,N_9312);
nand U14854 (N_14854,N_8085,N_12255);
nand U14855 (N_14855,N_7322,N_10474);
and U14856 (N_14856,N_7080,N_10902);
and U14857 (N_14857,N_8126,N_7971);
and U14858 (N_14858,N_10934,N_7553);
or U14859 (N_14859,N_9356,N_12436);
and U14860 (N_14860,N_8930,N_8117);
or U14861 (N_14861,N_8674,N_10872);
nor U14862 (N_14862,N_12187,N_8899);
nand U14863 (N_14863,N_12027,N_11316);
nor U14864 (N_14864,N_11566,N_7345);
or U14865 (N_14865,N_8104,N_7508);
nor U14866 (N_14866,N_12392,N_6257);
and U14867 (N_14867,N_10230,N_7351);
and U14868 (N_14868,N_10101,N_6583);
and U14869 (N_14869,N_7905,N_9919);
or U14870 (N_14870,N_10319,N_8383);
xor U14871 (N_14871,N_6643,N_9635);
or U14872 (N_14872,N_7770,N_6456);
nor U14873 (N_14873,N_7615,N_9060);
and U14874 (N_14874,N_7485,N_11413);
xor U14875 (N_14875,N_10170,N_10537);
nand U14876 (N_14876,N_8207,N_10207);
and U14877 (N_14877,N_12321,N_7252);
nor U14878 (N_14878,N_8359,N_8121);
nor U14879 (N_14879,N_9263,N_9933);
or U14880 (N_14880,N_10381,N_9282);
nor U14881 (N_14881,N_7210,N_9824);
or U14882 (N_14882,N_7906,N_11826);
xor U14883 (N_14883,N_11686,N_11829);
and U14884 (N_14884,N_12355,N_6538);
and U14885 (N_14885,N_8131,N_7046);
and U14886 (N_14886,N_7857,N_9021);
nand U14887 (N_14887,N_6845,N_8802);
and U14888 (N_14888,N_6344,N_11338);
nor U14889 (N_14889,N_10941,N_12270);
nand U14890 (N_14890,N_6777,N_7577);
xnor U14891 (N_14891,N_8830,N_8805);
nor U14892 (N_14892,N_7957,N_10566);
or U14893 (N_14893,N_9831,N_9065);
nor U14894 (N_14894,N_8734,N_9269);
nand U14895 (N_14895,N_8030,N_7776);
nor U14896 (N_14896,N_10407,N_12380);
nor U14897 (N_14897,N_8622,N_10587);
and U14898 (N_14898,N_8218,N_6352);
nor U14899 (N_14899,N_11208,N_10922);
and U14900 (N_14900,N_11053,N_11961);
xnor U14901 (N_14901,N_7575,N_8884);
and U14902 (N_14902,N_9960,N_9679);
and U14903 (N_14903,N_12471,N_11170);
or U14904 (N_14904,N_9484,N_11094);
or U14905 (N_14905,N_7086,N_10046);
nor U14906 (N_14906,N_11560,N_7592);
nand U14907 (N_14907,N_7678,N_12052);
and U14908 (N_14908,N_7543,N_8698);
nand U14909 (N_14909,N_10347,N_6765);
nand U14910 (N_14910,N_11453,N_9618);
nor U14911 (N_14911,N_6889,N_10860);
nor U14912 (N_14912,N_8723,N_8051);
nor U14913 (N_14913,N_12146,N_8066);
nand U14914 (N_14914,N_8214,N_8435);
or U14915 (N_14915,N_8762,N_9858);
and U14916 (N_14916,N_9845,N_12040);
nor U14917 (N_14917,N_10418,N_12235);
and U14918 (N_14918,N_6291,N_12212);
and U14919 (N_14919,N_7714,N_11391);
nand U14920 (N_14920,N_11237,N_7124);
and U14921 (N_14921,N_12411,N_11730);
nand U14922 (N_14922,N_7581,N_11385);
and U14923 (N_14923,N_8978,N_7751);
or U14924 (N_14924,N_9490,N_11168);
and U14925 (N_14925,N_11040,N_7803);
and U14926 (N_14926,N_6441,N_11865);
nand U14927 (N_14927,N_9291,N_6423);
and U14928 (N_14928,N_8039,N_10274);
nor U14929 (N_14929,N_6731,N_12364);
nand U14930 (N_14930,N_11985,N_11824);
nand U14931 (N_14931,N_7335,N_6695);
and U14932 (N_14932,N_7047,N_6601);
or U14933 (N_14933,N_11845,N_7215);
nand U14934 (N_14934,N_10720,N_6821);
or U14935 (N_14935,N_11768,N_9412);
nand U14936 (N_14936,N_6553,N_12185);
or U14937 (N_14937,N_11342,N_10068);
nor U14938 (N_14938,N_6266,N_8442);
xnor U14939 (N_14939,N_7983,N_11695);
and U14940 (N_14940,N_9460,N_8933);
nor U14941 (N_14941,N_12044,N_8835);
nand U14942 (N_14942,N_8180,N_10245);
and U14943 (N_14943,N_6298,N_8454);
nor U14944 (N_14944,N_9745,N_7162);
or U14945 (N_14945,N_9837,N_9067);
or U14946 (N_14946,N_6627,N_10356);
and U14947 (N_14947,N_8119,N_9838);
nand U14948 (N_14948,N_7623,N_10967);
nand U14949 (N_14949,N_7118,N_8468);
xnor U14950 (N_14950,N_7270,N_7835);
and U14951 (N_14951,N_7484,N_10073);
and U14952 (N_14952,N_6313,N_10482);
xor U14953 (N_14953,N_10256,N_10475);
or U14954 (N_14954,N_10057,N_11547);
nand U14955 (N_14955,N_9255,N_7158);
or U14956 (N_14956,N_12311,N_6616);
nand U14957 (N_14957,N_6831,N_10372);
nor U14958 (N_14958,N_6808,N_9496);
and U14959 (N_14959,N_11535,N_10131);
nor U14960 (N_14960,N_8991,N_8591);
or U14961 (N_14961,N_10617,N_7566);
xor U14962 (N_14962,N_12289,N_9063);
and U14963 (N_14963,N_6267,N_9180);
and U14964 (N_14964,N_10512,N_11634);
or U14965 (N_14965,N_10829,N_7383);
and U14966 (N_14966,N_12071,N_9857);
or U14967 (N_14967,N_12203,N_6682);
or U14968 (N_14968,N_10518,N_10477);
and U14969 (N_14969,N_12330,N_7486);
nor U14970 (N_14970,N_11760,N_10788);
nand U14971 (N_14971,N_10741,N_10388);
nand U14972 (N_14972,N_7587,N_7343);
or U14973 (N_14973,N_9963,N_11180);
xor U14974 (N_14974,N_10855,N_7539);
nand U14975 (N_14975,N_11065,N_8222);
and U14976 (N_14976,N_9813,N_7394);
and U14977 (N_14977,N_10034,N_11019);
or U14978 (N_14978,N_7859,N_12049);
nand U14979 (N_14979,N_10577,N_6572);
nor U14980 (N_14980,N_11136,N_11376);
xor U14981 (N_14981,N_7459,N_7120);
nand U14982 (N_14982,N_10238,N_12193);
xnor U14983 (N_14983,N_7538,N_7848);
or U14984 (N_14984,N_7655,N_7942);
or U14985 (N_14985,N_11164,N_8235);
nor U14986 (N_14986,N_12467,N_7222);
nand U14987 (N_14987,N_9775,N_7200);
nor U14988 (N_14988,N_8825,N_6761);
nand U14989 (N_14989,N_11320,N_6858);
nand U14990 (N_14990,N_10487,N_9182);
or U14991 (N_14991,N_7026,N_9916);
nand U14992 (N_14992,N_10858,N_7935);
and U14993 (N_14993,N_8407,N_7115);
nor U14994 (N_14994,N_7510,N_12239);
nand U14995 (N_14995,N_10445,N_11527);
nor U14996 (N_14996,N_8421,N_10425);
nand U14997 (N_14997,N_10980,N_7900);
nor U14998 (N_14998,N_7628,N_11835);
nor U14999 (N_14999,N_6385,N_12221);
nand U15000 (N_15000,N_7573,N_6938);
or U15001 (N_15001,N_7276,N_9489);
nor U15002 (N_15002,N_10977,N_9852);
xor U15003 (N_15003,N_12012,N_11205);
nor U15004 (N_15004,N_12121,N_8755);
and U15005 (N_15005,N_7072,N_7560);
or U15006 (N_15006,N_7987,N_6722);
or U15007 (N_15007,N_6771,N_7243);
or U15008 (N_15008,N_9733,N_12309);
or U15009 (N_15009,N_6956,N_11190);
nand U15010 (N_15010,N_10918,N_9188);
nor U15011 (N_15011,N_6807,N_10652);
nor U15012 (N_15012,N_8227,N_11492);
xor U15013 (N_15013,N_9495,N_8004);
or U15014 (N_15014,N_7999,N_9329);
xor U15015 (N_15015,N_6442,N_6707);
nor U15016 (N_15016,N_9244,N_12067);
xnor U15017 (N_15017,N_9233,N_11300);
nor U15018 (N_15018,N_7630,N_11279);
and U15019 (N_15019,N_10289,N_7167);
nor U15020 (N_15020,N_7537,N_11653);
nor U15021 (N_15021,N_8927,N_10248);
nand U15022 (N_15022,N_6584,N_10380);
and U15023 (N_15023,N_9682,N_8799);
or U15024 (N_15024,N_8776,N_6622);
nand U15025 (N_15025,N_9020,N_10130);
or U15026 (N_15026,N_9637,N_11781);
nand U15027 (N_15027,N_7279,N_9872);
or U15028 (N_15028,N_8543,N_6668);
and U15029 (N_15029,N_11998,N_10792);
nor U15030 (N_15030,N_9160,N_10114);
nand U15031 (N_15031,N_6826,N_7197);
and U15032 (N_15032,N_10246,N_12281);
and U15033 (N_15033,N_7690,N_7921);
nor U15034 (N_15034,N_10771,N_9265);
xor U15035 (N_15035,N_8408,N_8076);
nor U15036 (N_15036,N_7357,N_11770);
nand U15037 (N_15037,N_7402,N_6270);
nor U15038 (N_15038,N_9127,N_8552);
nand U15039 (N_15039,N_10966,N_10297);
and U15040 (N_15040,N_10016,N_9076);
nand U15041 (N_15041,N_9341,N_11042);
or U15042 (N_15042,N_8458,N_7715);
and U15043 (N_15043,N_10166,N_12385);
nor U15044 (N_15044,N_11539,N_11483);
nor U15045 (N_15045,N_9166,N_9666);
or U15046 (N_15046,N_12357,N_9221);
or U15047 (N_15047,N_8521,N_6988);
and U15048 (N_15048,N_11887,N_10740);
and U15049 (N_15049,N_9435,N_11860);
nand U15050 (N_15050,N_9768,N_7990);
and U15051 (N_15051,N_11721,N_8524);
or U15052 (N_15052,N_7887,N_10111);
and U15053 (N_15053,N_7264,N_11973);
and U15054 (N_15054,N_8623,N_7931);
nor U15055 (N_15055,N_8920,N_12319);
and U15056 (N_15056,N_11434,N_10521);
nor U15057 (N_15057,N_9529,N_10000);
nand U15058 (N_15058,N_6357,N_8401);
nand U15059 (N_15059,N_11894,N_6670);
xnor U15060 (N_15060,N_6861,N_7622);
nor U15061 (N_15061,N_11977,N_9409);
and U15062 (N_15062,N_8782,N_8084);
nor U15063 (N_15063,N_8914,N_11619);
nor U15064 (N_15064,N_12240,N_8325);
nor U15065 (N_15065,N_7234,N_7206);
or U15066 (N_15066,N_7794,N_11488);
and U15067 (N_15067,N_10909,N_6832);
nor U15068 (N_15068,N_10086,N_8378);
nor U15069 (N_15069,N_10338,N_11722);
nand U15070 (N_15070,N_8746,N_9781);
and U15071 (N_15071,N_11647,N_10109);
and U15072 (N_15072,N_6570,N_9086);
or U15073 (N_15073,N_7136,N_9370);
or U15074 (N_15074,N_10649,N_8103);
nand U15075 (N_15075,N_7480,N_11308);
nor U15076 (N_15076,N_7910,N_6685);
nor U15077 (N_15077,N_11064,N_10406);
or U15078 (N_15078,N_9729,N_8681);
or U15079 (N_15079,N_8763,N_8708);
nand U15080 (N_15080,N_8416,N_6373);
nand U15081 (N_15081,N_10049,N_11456);
nor U15082 (N_15082,N_9743,N_9728);
and U15083 (N_15083,N_11230,N_7825);
nor U15084 (N_15084,N_6945,N_7914);
or U15085 (N_15085,N_6615,N_9522);
and U15086 (N_15086,N_11207,N_12046);
and U15087 (N_15087,N_8216,N_7890);
and U15088 (N_15088,N_9546,N_7509);
xnor U15089 (N_15089,N_6823,N_8470);
nor U15090 (N_15090,N_10322,N_11309);
nor U15091 (N_15091,N_9767,N_8818);
and U15092 (N_15092,N_11234,N_8446);
or U15093 (N_15093,N_10822,N_10458);
nand U15094 (N_15094,N_9343,N_12464);
or U15095 (N_15095,N_8527,N_9213);
nor U15096 (N_15096,N_12072,N_10634);
xnor U15097 (N_15097,N_6322,N_12296);
or U15098 (N_15098,N_12344,N_9947);
or U15099 (N_15099,N_6598,N_11989);
nand U15100 (N_15100,N_9141,N_10457);
or U15101 (N_15101,N_7591,N_11822);
xor U15102 (N_15102,N_8857,N_11496);
nor U15103 (N_15103,N_11723,N_11631);
and U15104 (N_15104,N_6314,N_10234);
or U15105 (N_15105,N_9596,N_12163);
or U15106 (N_15106,N_10162,N_8456);
or U15107 (N_15107,N_8269,N_12218);
xor U15108 (N_15108,N_11452,N_9427);
and U15109 (N_15109,N_12490,N_7746);
nand U15110 (N_15110,N_10055,N_11022);
or U15111 (N_15111,N_7314,N_10176);
nand U15112 (N_15112,N_6624,N_10421);
and U15113 (N_15113,N_6880,N_7869);
nor U15114 (N_15114,N_11467,N_9502);
or U15115 (N_15115,N_6687,N_11146);
nand U15116 (N_15116,N_11744,N_8098);
or U15117 (N_15117,N_9821,N_7039);
nor U15118 (N_15118,N_6743,N_9978);
and U15119 (N_15119,N_10031,N_6465);
nor U15120 (N_15120,N_7294,N_9407);
or U15121 (N_15121,N_12284,N_11757);
or U15122 (N_15122,N_7467,N_6762);
nand U15123 (N_15123,N_7018,N_8589);
nor U15124 (N_15124,N_8779,N_8321);
or U15125 (N_15125,N_10731,N_12265);
nand U15126 (N_15126,N_12063,N_10459);
or U15127 (N_15127,N_8808,N_10596);
nand U15128 (N_15128,N_6308,N_8219);
nor U15129 (N_15129,N_8473,N_8761);
nor U15130 (N_15130,N_10628,N_9372);
or U15131 (N_15131,N_7512,N_12338);
nor U15132 (N_15132,N_10953,N_7703);
nand U15133 (N_15133,N_8001,N_6882);
and U15134 (N_15134,N_11729,N_6483);
nor U15135 (N_15135,N_9860,N_10090);
or U15136 (N_15136,N_7187,N_9167);
or U15137 (N_15137,N_10522,N_8553);
nand U15138 (N_15138,N_6454,N_8003);
or U15139 (N_15139,N_12134,N_9054);
nor U15140 (N_15140,N_6426,N_7221);
nand U15141 (N_15141,N_10681,N_7236);
and U15142 (N_15142,N_8228,N_9308);
or U15143 (N_15143,N_9214,N_8285);
nand U15144 (N_15144,N_9455,N_11510);
nand U15145 (N_15145,N_10881,N_12136);
xor U15146 (N_15146,N_6840,N_9548);
and U15147 (N_15147,N_9485,N_11554);
nand U15148 (N_15148,N_12305,N_10584);
nand U15149 (N_15149,N_7780,N_10188);
nor U15150 (N_15150,N_11983,N_8075);
nand U15151 (N_15151,N_8143,N_7166);
nor U15152 (N_15152,N_6455,N_9179);
nand U15153 (N_15153,N_10604,N_6544);
nor U15154 (N_15154,N_10206,N_9332);
and U15155 (N_15155,N_10647,N_12104);
and U15156 (N_15156,N_8850,N_7821);
or U15157 (N_15157,N_10134,N_8305);
nand U15158 (N_15158,N_8663,N_7571);
nor U15159 (N_15159,N_9817,N_8594);
xnor U15160 (N_15160,N_12400,N_10385);
or U15161 (N_15161,N_9172,N_6864);
nor U15162 (N_15162,N_6735,N_11321);
and U15163 (N_15163,N_6360,N_8169);
and U15164 (N_15164,N_8010,N_10277);
or U15165 (N_15165,N_8661,N_9575);
nor U15166 (N_15166,N_6856,N_8120);
nand U15167 (N_15167,N_9861,N_9885);
xor U15168 (N_15168,N_7092,N_9992);
or U15169 (N_15169,N_12383,N_10044);
nand U15170 (N_15170,N_10958,N_9206);
nor U15171 (N_15171,N_9121,N_11993);
xnor U15172 (N_15172,N_10369,N_9272);
and U15173 (N_15173,N_10671,N_11477);
nand U15174 (N_15174,N_7860,N_7626);
xnor U15175 (N_15175,N_10706,N_9242);
nor U15176 (N_15176,N_6935,N_9136);
and U15177 (N_15177,N_7982,N_10106);
nor U15178 (N_15178,N_10802,N_9581);
nand U15179 (N_15179,N_9105,N_9503);
and U15180 (N_15180,N_12048,N_11479);
nand U15181 (N_15181,N_11126,N_9699);
nor U15182 (N_15182,N_9380,N_9889);
or U15183 (N_15183,N_6259,N_7995);
xnor U15184 (N_15184,N_11679,N_12135);
or U15185 (N_15185,N_10401,N_9463);
or U15186 (N_15186,N_10312,N_6778);
xor U15187 (N_15187,N_9829,N_12331);
or U15188 (N_15188,N_12391,N_7604);
nand U15189 (N_15189,N_11882,N_11740);
or U15190 (N_15190,N_11120,N_6697);
nor U15191 (N_15191,N_11351,N_8859);
or U15192 (N_15192,N_6294,N_9582);
xor U15193 (N_15193,N_11073,N_10029);
xnor U15194 (N_15194,N_10292,N_11858);
xor U15195 (N_15195,N_7331,N_10295);
or U15196 (N_15196,N_10599,N_10154);
xnor U15197 (N_15197,N_12494,N_7053);
nor U15198 (N_15198,N_11971,N_8509);
and U15199 (N_15199,N_11574,N_8840);
and U15200 (N_15200,N_8395,N_12266);
or U15201 (N_15201,N_6632,N_10307);
nor U15202 (N_15202,N_9900,N_8798);
or U15203 (N_15203,N_7832,N_8595);
nand U15204 (N_15204,N_9450,N_11819);
nor U15205 (N_15205,N_8250,N_6694);
and U15206 (N_15206,N_8809,N_10257);
nor U15207 (N_15207,N_7390,N_12249);
nor U15208 (N_15208,N_10420,N_11941);
and U15209 (N_15209,N_7354,N_6894);
xor U15210 (N_15210,N_9228,N_11171);
nor U15211 (N_15211,N_11541,N_12367);
xnor U15212 (N_15212,N_10935,N_6914);
or U15213 (N_15213,N_7421,N_11437);
nor U15214 (N_15214,N_12016,N_6577);
nor U15215 (N_15215,N_6994,N_8916);
and U15216 (N_15216,N_10361,N_6610);
or U15217 (N_15217,N_10882,N_9721);
nor U15218 (N_15218,N_10513,N_7603);
nor U15219 (N_15219,N_7044,N_10469);
or U15220 (N_15220,N_9235,N_6453);
nor U15221 (N_15221,N_6413,N_11076);
nor U15222 (N_15222,N_6591,N_9788);
xnor U15223 (N_15223,N_7239,N_9000);
or U15224 (N_15224,N_8540,N_8493);
nand U15225 (N_15225,N_9028,N_11125);
nand U15226 (N_15226,N_10752,N_10018);
nand U15227 (N_15227,N_9956,N_10194);
and U15228 (N_15228,N_8554,N_8979);
and U15229 (N_15229,N_7481,N_8545);
or U15230 (N_15230,N_12248,N_8657);
nand U15231 (N_15231,N_7824,N_10135);
xor U15232 (N_15232,N_10386,N_11929);
or U15233 (N_15233,N_6830,N_8053);
xnor U15234 (N_15234,N_10938,N_11031);
or U15235 (N_15235,N_10104,N_7284);
or U15236 (N_15236,N_9634,N_10550);
nand U15237 (N_15237,N_6918,N_11603);
and U15238 (N_15238,N_10690,N_11598);
and U15239 (N_15239,N_10404,N_11192);
xnor U15240 (N_15240,N_10139,N_10435);
or U15241 (N_15241,N_9148,N_9262);
nor U15242 (N_15242,N_12489,N_9628);
and U15243 (N_15243,N_10704,N_12084);
nand U15244 (N_15244,N_11643,N_8516);
nand U15245 (N_15245,N_9461,N_8422);
nor U15246 (N_15246,N_8423,N_10694);
nand U15247 (N_15247,N_11123,N_12474);
xor U15248 (N_15248,N_11310,N_10793);
nor U15249 (N_15249,N_9703,N_9003);
or U15250 (N_15250,N_7425,N_7938);
and U15251 (N_15251,N_11645,N_8834);
nand U15252 (N_15252,N_11027,N_6987);
nand U15253 (N_15253,N_6251,N_10293);
nor U15254 (N_15254,N_9880,N_8178);
nand U15255 (N_15255,N_9717,N_8457);
nor U15256 (N_15256,N_11680,N_7749);
and U15257 (N_15257,N_12117,N_11501);
and U15258 (N_15258,N_12429,N_10174);
or U15259 (N_15259,N_12341,N_9574);
and U15260 (N_15260,N_11005,N_11018);
nor U15261 (N_15261,N_7554,N_10929);
xor U15262 (N_15262,N_9305,N_11112);
nor U15263 (N_15263,N_6661,N_6332);
nor U15264 (N_15264,N_10181,N_6850);
nand U15265 (N_15265,N_8863,N_9959);
and U15266 (N_15266,N_9835,N_9544);
or U15267 (N_15267,N_8613,N_12169);
and U15268 (N_15268,N_12332,N_10590);
nand U15269 (N_15269,N_7370,N_11038);
nand U15270 (N_15270,N_8015,N_9303);
nor U15271 (N_15271,N_9230,N_10434);
nor U15272 (N_15272,N_7449,N_6877);
nor U15273 (N_15273,N_9284,N_7578);
and U15274 (N_15274,N_10214,N_8220);
xnor U15275 (N_15275,N_7519,N_10547);
or U15276 (N_15276,N_11096,N_11402);
nor U15277 (N_15277,N_8670,N_7675);
nor U15278 (N_15278,N_8071,N_10011);
or U15279 (N_15279,N_11410,N_12043);
or U15280 (N_15280,N_8534,N_9630);
nor U15281 (N_15281,N_10448,N_10733);
or U15282 (N_15282,N_8328,N_9061);
nand U15283 (N_15283,N_12285,N_10472);
nor U15284 (N_15284,N_8716,N_11468);
nor U15285 (N_15285,N_11931,N_8153);
or U15286 (N_15286,N_10030,N_6451);
and U15287 (N_15287,N_7443,N_8315);
nand U15288 (N_15288,N_9816,N_8290);
nor U15289 (N_15289,N_10719,N_12010);
nor U15290 (N_15290,N_11877,N_12172);
and U15291 (N_15291,N_10352,N_6758);
nor U15292 (N_15292,N_10225,N_11148);
and U15293 (N_15293,N_11943,N_6316);
nand U15294 (N_15294,N_9336,N_11419);
nand U15295 (N_15295,N_10093,N_9823);
and U15296 (N_15296,N_12182,N_7947);
xnor U15297 (N_15297,N_10715,N_8078);
and U15298 (N_15298,N_8069,N_8551);
xor U15299 (N_15299,N_9334,N_9483);
nor U15300 (N_15300,N_7377,N_11676);
and U15301 (N_15301,N_8109,N_11895);
or U15302 (N_15302,N_12325,N_6275);
nand U15303 (N_15303,N_7050,N_12405);
nand U15304 (N_15304,N_6993,N_11069);
nor U15305 (N_15305,N_10364,N_7195);
and U15306 (N_15306,N_7237,N_11814);
nor U15307 (N_15307,N_12122,N_7809);
nand U15308 (N_15308,N_10395,N_8388);
nand U15309 (N_15309,N_8002,N_10903);
nand U15310 (N_15310,N_6433,N_10167);
nand U15311 (N_15311,N_12165,N_10195);
or U15312 (N_15312,N_12470,N_7888);
and U15313 (N_15313,N_9620,N_9524);
nor U15314 (N_15314,N_7189,N_9477);
xnor U15315 (N_15315,N_8448,N_9369);
nor U15316 (N_15316,N_8065,N_12149);
and U15317 (N_15317,N_9898,N_11489);
nand U15318 (N_15318,N_10315,N_6410);
or U15319 (N_15319,N_11683,N_6296);
or U15320 (N_15320,N_6649,N_12222);
or U15321 (N_15321,N_7605,N_12396);
nand U15322 (N_15322,N_7960,N_11274);
nand U15323 (N_15323,N_10491,N_8987);
nand U15324 (N_15324,N_8340,N_6353);
xor U15325 (N_15325,N_8116,N_11210);
nand U15326 (N_15326,N_7951,N_7227);
and U15327 (N_15327,N_7624,N_10784);
or U15328 (N_15328,N_9404,N_7367);
and U15329 (N_15329,N_9690,N_11773);
nand U15330 (N_15330,N_11616,N_7953);
and U15331 (N_15331,N_12431,N_6569);
or U15332 (N_15332,N_8714,N_9395);
and U15333 (N_15333,N_8405,N_11785);
xor U15334 (N_15334,N_7494,N_10978);
nand U15335 (N_15335,N_9080,N_12150);
nand U15336 (N_15336,N_6295,N_11089);
nor U15337 (N_15337,N_11187,N_10887);
nor U15338 (N_15338,N_7639,N_11850);
and U15339 (N_15339,N_8333,N_6756);
nor U15340 (N_15340,N_9708,N_9641);
nor U15341 (N_15341,N_8060,N_11732);
nand U15342 (N_15342,N_7585,N_11536);
and U15343 (N_15343,N_6961,N_12081);
and U15344 (N_15344,N_10942,N_10623);
nor U15345 (N_15345,N_11232,N_9663);
or U15346 (N_15346,N_7424,N_7305);
nand U15347 (N_15347,N_10444,N_8742);
and U15348 (N_15348,N_6484,N_8582);
or U15349 (N_15349,N_10805,N_8152);
and U15350 (N_15350,N_11135,N_9893);
or U15351 (N_15351,N_8195,N_7652);
or U15352 (N_15352,N_11913,N_8893);
nor U15353 (N_15353,N_11214,N_7719);
nand U15354 (N_15354,N_11372,N_7778);
xor U15355 (N_15355,N_6286,N_9653);
nand U15356 (N_15356,N_11388,N_9283);
xor U15357 (N_15357,N_6297,N_9600);
and U15358 (N_15358,N_10810,N_8052);
nand U15359 (N_15359,N_8284,N_9048);
or U15360 (N_15360,N_7163,N_10613);
nand U15361 (N_15361,N_6302,N_10402);
nor U15362 (N_15362,N_6491,N_10914);
nor U15363 (N_15363,N_10824,N_11926);
nor U15364 (N_15364,N_9624,N_10908);
or U15365 (N_15365,N_9589,N_7008);
or U15366 (N_15366,N_10622,N_9964);
and U15367 (N_15367,N_8025,N_7020);
nor U15368 (N_15368,N_8188,N_10024);
nor U15369 (N_15369,N_9452,N_8191);
and U15370 (N_15370,N_11469,N_9763);
nor U15371 (N_15371,N_9752,N_8999);
xor U15372 (N_15372,N_10682,N_9131);
or U15373 (N_15373,N_8518,N_9223);
nor U15374 (N_15374,N_9239,N_12418);
and U15375 (N_15375,N_8242,N_10568);
and U15376 (N_15376,N_10869,N_10648);
xor U15377 (N_15377,N_6718,N_7676);
and U15378 (N_15378,N_10461,N_6795);
nand U15379 (N_15379,N_12158,N_8728);
nor U15380 (N_15380,N_9613,N_7267);
or U15381 (N_15381,N_7518,N_10242);
xnor U15382 (N_15382,N_8767,N_8127);
and U15383 (N_15383,N_10187,N_7988);
nand U15384 (N_15384,N_9181,N_9879);
nand U15385 (N_15385,N_9593,N_10237);
and U15386 (N_15386,N_7991,N_6621);
nand U15387 (N_15387,N_7495,N_8887);
nand U15388 (N_15388,N_7705,N_7087);
and U15389 (N_15389,N_9445,N_6965);
xnor U15390 (N_15390,N_9480,N_10567);
and U15391 (N_15391,N_12445,N_8891);
nor U15392 (N_15392,N_7010,N_6950);
and U15393 (N_15393,N_9314,N_9815);
nor U15394 (N_15394,N_11907,N_10815);
nand U15395 (N_15395,N_6760,N_11827);
or U15396 (N_15396,N_9625,N_9520);
nor U15397 (N_15397,N_7588,N_11848);
nor U15398 (N_15398,N_7030,N_11666);
or U15399 (N_15399,N_9494,N_8984);
or U15400 (N_15400,N_10732,N_10989);
or U15401 (N_15401,N_7223,N_11322);
or U15402 (N_15402,N_8866,N_8689);
nand U15403 (N_15403,N_10332,N_8097);
nand U15404 (N_15404,N_10310,N_10549);
and U15405 (N_15405,N_10265,N_6390);
nand U15406 (N_15406,N_9878,N_8672);
nand U15407 (N_15407,N_8795,N_6337);
nor U15408 (N_15408,N_7701,N_8506);
nor U15409 (N_15409,N_10460,N_7261);
nand U15410 (N_15410,N_7613,N_12191);
nor U15411 (N_15411,N_8193,N_11461);
or U15412 (N_15412,N_6506,N_12123);
xnor U15413 (N_15413,N_11938,N_11880);
nand U15414 (N_15414,N_10960,N_7882);
nor U15415 (N_15415,N_7802,N_6467);
nor U15416 (N_15416,N_9886,N_6734);
or U15417 (N_15417,N_8123,N_8772);
or U15418 (N_15418,N_6526,N_6951);
and U15419 (N_15419,N_9645,N_6502);
or U15420 (N_15420,N_9306,N_7808);
or U15421 (N_15421,N_11707,N_9134);
or U15422 (N_15422,N_10763,N_10368);
or U15423 (N_15423,N_10507,N_9804);
and U15424 (N_15424,N_9360,N_9656);
and U15425 (N_15425,N_10728,N_7606);
or U15426 (N_15426,N_7312,N_6933);
nand U15427 (N_15427,N_9327,N_7271);
and U15428 (N_15428,N_7477,N_7876);
nand U15429 (N_15429,N_11153,N_6340);
nor U15430 (N_15430,N_7704,N_8323);
nand U15431 (N_15431,N_10761,N_11357);
nand U15432 (N_15432,N_12145,N_7076);
or U15433 (N_15433,N_7559,N_6351);
and U15434 (N_15434,N_10913,N_7617);
nor U15435 (N_15435,N_7317,N_8990);
nand U15436 (N_15436,N_9887,N_10931);
nor U15437 (N_15437,N_9082,N_10249);
or U15438 (N_15438,N_12375,N_9680);
nor U15439 (N_15439,N_11213,N_6800);
nand U15440 (N_15440,N_10058,N_11412);
or U15441 (N_15441,N_11948,N_7762);
nor U15442 (N_15442,N_8390,N_8257);
nand U15443 (N_15443,N_7873,N_10772);
or U15444 (N_15444,N_9644,N_11553);
or U15445 (N_15445,N_9516,N_10175);
and U15446 (N_15446,N_8450,N_12315);
nand U15447 (N_15447,N_11979,N_9598);
nor U15448 (N_15448,N_8083,N_6511);
nor U15449 (N_15449,N_11161,N_9229);
or U15450 (N_15450,N_11637,N_10813);
nand U15451 (N_15451,N_9732,N_10054);
or U15452 (N_15452,N_9777,N_10132);
xor U15453 (N_15453,N_12426,N_7037);
nand U15454 (N_15454,N_10509,N_7408);
nand U15455 (N_15455,N_10962,N_9357);
or U15456 (N_15456,N_7574,N_10009);
nand U15457 (N_15457,N_7123,N_9583);
and U15458 (N_15458,N_11117,N_9871);
nand U15459 (N_15459,N_8977,N_7493);
nor U15460 (N_15460,N_7307,N_8864);
nor U15461 (N_15461,N_12236,N_11652);
nand U15462 (N_15462,N_6395,N_12069);
and U15463 (N_15463,N_7954,N_10082);
or U15464 (N_15464,N_9374,N_8101);
and U15465 (N_15465,N_10281,N_12260);
and U15466 (N_15466,N_7015,N_11247);
or U15467 (N_15467,N_7535,N_6564);
nand U15468 (N_15468,N_12451,N_10357);
nand U15469 (N_15469,N_6962,N_11736);
or U15470 (N_15470,N_9723,N_10708);
xor U15471 (N_15471,N_10925,N_6844);
or U15472 (N_15472,N_9424,N_7709);
nand U15473 (N_15473,N_9715,N_8794);
nand U15474 (N_15474,N_10501,N_7926);
or U15475 (N_15475,N_8512,N_7376);
nand U15476 (N_15476,N_7225,N_11052);
and U15477 (N_15477,N_10923,N_11905);
nand U15478 (N_15478,N_9285,N_8313);
nor U15479 (N_15479,N_10949,N_11399);
and U15480 (N_15480,N_7211,N_10775);
nor U15481 (N_15481,N_8205,N_7804);
or U15482 (N_15482,N_12125,N_7974);
nor U15483 (N_15483,N_7647,N_11799);
nor U15484 (N_15484,N_11211,N_6676);
or U15485 (N_15485,N_10233,N_6609);
and U15486 (N_15486,N_11668,N_9219);
or U15487 (N_15487,N_6857,N_9627);
or U15488 (N_15488,N_10816,N_11846);
or U15489 (N_15489,N_10280,N_11066);
nand U15490 (N_15490,N_11368,N_8430);
or U15491 (N_15491,N_8637,N_9692);
or U15492 (N_15492,N_6488,N_10424);
and U15493 (N_15493,N_7057,N_7172);
or U15494 (N_15494,N_6349,N_8036);
or U15495 (N_15495,N_7826,N_9317);
xnor U15496 (N_15496,N_9446,N_12487);
or U15497 (N_15497,N_11222,N_9759);
nand U15498 (N_15498,N_8806,N_12301);
nor U15499 (N_15499,N_6419,N_10342);
nand U15500 (N_15500,N_8068,N_8058);
nor U15501 (N_15501,N_10674,N_8427);
nand U15502 (N_15502,N_6573,N_12428);
xor U15503 (N_15503,N_7074,N_7330);
and U15504 (N_15504,N_11113,N_12070);
and U15505 (N_15505,N_10517,N_11015);
and U15506 (N_15506,N_7373,N_9010);
nor U15507 (N_15507,N_9406,N_11756);
nand U15508 (N_15508,N_7083,N_9258);
nor U15509 (N_15509,N_11258,N_10884);
and U15510 (N_15510,N_10998,N_11465);
nor U15511 (N_15511,N_7608,N_10019);
nor U15512 (N_15512,N_10495,N_9746);
nor U15513 (N_15513,N_6435,N_10896);
nor U15514 (N_15514,N_12369,N_8263);
xor U15515 (N_15515,N_9011,N_9970);
nor U15516 (N_15516,N_11179,N_10391);
and U15517 (N_15517,N_6814,N_11832);
or U15518 (N_15518,N_9197,N_8549);
and U15519 (N_15519,N_10138,N_7448);
and U15520 (N_15520,N_7689,N_11521);
and U15521 (N_15521,N_9539,N_6347);
xnor U15522 (N_15522,N_11398,N_11967);
nand U15523 (N_15523,N_7096,N_7765);
nor U15524 (N_15524,N_6281,N_7711);
or U15525 (N_15525,N_11075,N_9216);
or U15526 (N_15526,N_9981,N_6388);
xor U15527 (N_15527,N_6507,N_11628);
or U15528 (N_15528,N_8640,N_11105);
nand U15529 (N_15529,N_6730,N_9633);
or U15530 (N_15530,N_9069,N_10559);
nand U15531 (N_15531,N_7659,N_9352);
nor U15532 (N_15532,N_8129,N_7054);
nand U15533 (N_15533,N_11956,N_6528);
or U15534 (N_15534,N_12140,N_12038);
nor U15535 (N_15535,N_6424,N_8602);
or U15536 (N_15536,N_6940,N_12132);
or U15537 (N_15537,N_8231,N_9102);
and U15538 (N_15538,N_10994,N_9836);
or U15539 (N_15539,N_8474,N_6652);
nand U15540 (N_15540,N_12389,N_6575);
nand U15541 (N_15541,N_6745,N_8838);
or U15542 (N_15542,N_9910,N_11455);
nor U15543 (N_15543,N_8181,N_7418);
and U15544 (N_15544,N_10146,N_7492);
nor U15545 (N_15545,N_7867,N_10570);
nand U15546 (N_15546,N_6662,N_6869);
or U15547 (N_15547,N_10770,N_8019);
and U15548 (N_15548,N_11043,N_6717);
or U15549 (N_15549,N_11293,N_7161);
and U15550 (N_15550,N_10276,N_10020);
and U15551 (N_15551,N_9667,N_9129);
xnor U15552 (N_15552,N_11502,N_11528);
nor U15553 (N_15553,N_8770,N_6463);
nand U15554 (N_15554,N_9289,N_12469);
and U15555 (N_15555,N_11292,N_9640);
xor U15556 (N_15556,N_11599,N_10426);
or U15557 (N_15557,N_6464,N_7915);
and U15558 (N_15558,N_7419,N_8603);
nand U15559 (N_15559,N_7966,N_8783);
xor U15560 (N_15560,N_11068,N_8141);
nand U15561 (N_15561,N_9720,N_12045);
and U15562 (N_15562,N_11111,N_9187);
and U15563 (N_15563,N_7090,N_6746);
or U15564 (N_15564,N_7657,N_9444);
nand U15565 (N_15565,N_12384,N_7219);
nor U15566 (N_15566,N_9971,N_10417);
and U15567 (N_15567,N_8725,N_9537);
nand U15568 (N_15568,N_11221,N_9532);
and U15569 (N_15569,N_7673,N_6704);
xor U15570 (N_15570,N_12379,N_10786);
xor U15571 (N_15571,N_11635,N_9066);
nor U15572 (N_15572,N_9361,N_7393);
xor U15573 (N_15573,N_8700,N_12479);
nor U15574 (N_15574,N_10750,N_6660);
and U15575 (N_15575,N_8963,N_6916);
or U15576 (N_15576,N_9779,N_8380);
or U15577 (N_15577,N_10397,N_11133);
and U15578 (N_15578,N_11302,N_10531);
nor U15579 (N_15579,N_11060,N_10667);
nor U15580 (N_15580,N_6973,N_11624);
xor U15581 (N_15581,N_7561,N_8618);
nand U15582 (N_15582,N_10359,N_11611);
and U15583 (N_15583,N_9955,N_8569);
nor U15584 (N_15584,N_11511,N_12271);
nor U15585 (N_15585,N_8356,N_11498);
nand U15586 (N_15586,N_10227,N_10717);
and U15587 (N_15587,N_7321,N_11798);
or U15588 (N_15588,N_9962,N_7062);
or U15589 (N_15589,N_9006,N_11204);
nand U15590 (N_15590,N_8694,N_12173);
nand U15591 (N_15591,N_9555,N_10891);
nand U15592 (N_15592,N_9120,N_6855);
or U15593 (N_15593,N_9397,N_10108);
or U15594 (N_15594,N_10579,N_12124);
or U15595 (N_15595,N_9091,N_10983);
and U15596 (N_15596,N_11007,N_7283);
and U15597 (N_15597,N_11844,N_10716);
or U15598 (N_15598,N_8210,N_8682);
and U15599 (N_15599,N_12339,N_8879);
xnor U15600 (N_15600,N_10917,N_7700);
nand U15601 (N_15601,N_10413,N_12253);
or U15602 (N_15602,N_12324,N_10666);
or U15603 (N_15603,N_10789,N_11472);
nand U15604 (N_15604,N_6925,N_6533);
nor U15605 (N_15605,N_12177,N_6527);
nand U15606 (N_15606,N_8756,N_11688);
nand U15607 (N_15607,N_10259,N_9894);
and U15608 (N_15608,N_7736,N_8968);
or U15609 (N_15609,N_7102,N_9379);
nor U15610 (N_15610,N_7075,N_11594);
nor U15611 (N_15611,N_7127,N_7528);
xor U15612 (N_15612,N_6711,N_8247);
nand U15613 (N_15613,N_10298,N_6804);
nor U15614 (N_15614,N_11700,N_9036);
nand U15615 (N_15615,N_9786,N_7051);
nor U15616 (N_15616,N_10774,N_9749);
nor U15617 (N_15617,N_7727,N_10053);
nand U15618 (N_15618,N_6790,N_11573);
and U15619 (N_15619,N_6968,N_8998);
nor U15620 (N_15620,N_12022,N_8080);
nor U15621 (N_15621,N_9534,N_11656);
nor U15622 (N_15622,N_8392,N_8344);
and U15623 (N_15623,N_8276,N_8110);
nor U15624 (N_15624,N_7874,N_8147);
or U15625 (N_15625,N_12360,N_10378);
xor U15626 (N_15626,N_8360,N_11775);
xnor U15627 (N_15627,N_11721,N_7594);
or U15628 (N_15628,N_11894,N_9783);
nor U15629 (N_15629,N_10331,N_7582);
or U15630 (N_15630,N_11425,N_7697);
and U15631 (N_15631,N_10468,N_7955);
nand U15632 (N_15632,N_7843,N_6710);
xnor U15633 (N_15633,N_10617,N_10962);
nand U15634 (N_15634,N_12071,N_8748);
or U15635 (N_15635,N_7597,N_10014);
nand U15636 (N_15636,N_10608,N_10801);
nand U15637 (N_15637,N_7828,N_7487);
nand U15638 (N_15638,N_10680,N_7461);
nand U15639 (N_15639,N_8232,N_10753);
xnor U15640 (N_15640,N_11776,N_6544);
nor U15641 (N_15641,N_7070,N_11552);
nor U15642 (N_15642,N_11022,N_11773);
and U15643 (N_15643,N_8026,N_8303);
nor U15644 (N_15644,N_8473,N_10251);
nor U15645 (N_15645,N_8962,N_11920);
nor U15646 (N_15646,N_12427,N_9908);
and U15647 (N_15647,N_7560,N_6830);
or U15648 (N_15648,N_8285,N_11539);
or U15649 (N_15649,N_9908,N_10631);
and U15650 (N_15650,N_7338,N_7664);
and U15651 (N_15651,N_11482,N_8612);
xnor U15652 (N_15652,N_11768,N_10544);
nand U15653 (N_15653,N_8699,N_6843);
nand U15654 (N_15654,N_8505,N_11593);
nor U15655 (N_15655,N_6330,N_11730);
or U15656 (N_15656,N_9596,N_11037);
nand U15657 (N_15657,N_9141,N_10191);
or U15658 (N_15658,N_8568,N_11084);
or U15659 (N_15659,N_6590,N_12163);
nand U15660 (N_15660,N_10696,N_9681);
or U15661 (N_15661,N_11475,N_10928);
nand U15662 (N_15662,N_6850,N_8126);
and U15663 (N_15663,N_6694,N_8753);
or U15664 (N_15664,N_6883,N_9214);
nand U15665 (N_15665,N_8141,N_11709);
nor U15666 (N_15666,N_10498,N_11607);
nor U15667 (N_15667,N_11821,N_9097);
nor U15668 (N_15668,N_8706,N_7560);
and U15669 (N_15669,N_10197,N_7126);
nand U15670 (N_15670,N_8162,N_10185);
and U15671 (N_15671,N_11348,N_11561);
or U15672 (N_15672,N_11689,N_9159);
or U15673 (N_15673,N_8111,N_8095);
nand U15674 (N_15674,N_8875,N_8379);
and U15675 (N_15675,N_11106,N_8623);
nand U15676 (N_15676,N_6650,N_9836);
xnor U15677 (N_15677,N_11503,N_11309);
nor U15678 (N_15678,N_12375,N_9209);
or U15679 (N_15679,N_8468,N_7475);
nor U15680 (N_15680,N_8624,N_7063);
nor U15681 (N_15681,N_6992,N_9106);
nor U15682 (N_15682,N_12244,N_6579);
nand U15683 (N_15683,N_6778,N_10210);
and U15684 (N_15684,N_7986,N_11014);
nor U15685 (N_15685,N_6538,N_7843);
xor U15686 (N_15686,N_6789,N_6655);
and U15687 (N_15687,N_7962,N_11355);
or U15688 (N_15688,N_10403,N_11824);
xor U15689 (N_15689,N_8977,N_7708);
or U15690 (N_15690,N_8575,N_9954);
nand U15691 (N_15691,N_8872,N_10130);
or U15692 (N_15692,N_7232,N_9944);
and U15693 (N_15693,N_7712,N_9831);
nand U15694 (N_15694,N_6864,N_10173);
nand U15695 (N_15695,N_7880,N_12265);
and U15696 (N_15696,N_10317,N_6406);
or U15697 (N_15697,N_11388,N_10679);
or U15698 (N_15698,N_11306,N_8664);
nand U15699 (N_15699,N_12194,N_10869);
nand U15700 (N_15700,N_6454,N_10821);
or U15701 (N_15701,N_9255,N_10416);
and U15702 (N_15702,N_7137,N_7410);
and U15703 (N_15703,N_10262,N_10576);
nor U15704 (N_15704,N_11034,N_9093);
nor U15705 (N_15705,N_11545,N_7757);
nand U15706 (N_15706,N_6893,N_8412);
nand U15707 (N_15707,N_6899,N_7643);
nor U15708 (N_15708,N_11789,N_11751);
xnor U15709 (N_15709,N_8564,N_7003);
nor U15710 (N_15710,N_8544,N_10382);
nand U15711 (N_15711,N_7544,N_7316);
nand U15712 (N_15712,N_9514,N_9128);
and U15713 (N_15713,N_11944,N_6288);
nand U15714 (N_15714,N_6439,N_8094);
nand U15715 (N_15715,N_7993,N_11308);
nor U15716 (N_15716,N_12155,N_6495);
nor U15717 (N_15717,N_6715,N_9432);
or U15718 (N_15718,N_8635,N_6350);
and U15719 (N_15719,N_11565,N_8171);
and U15720 (N_15720,N_6922,N_10789);
or U15721 (N_15721,N_11654,N_8907);
nor U15722 (N_15722,N_10615,N_8053);
and U15723 (N_15723,N_8732,N_8930);
or U15724 (N_15724,N_11006,N_9496);
nor U15725 (N_15725,N_7638,N_8181);
nand U15726 (N_15726,N_12389,N_7466);
and U15727 (N_15727,N_11440,N_10032);
nand U15728 (N_15728,N_7997,N_6397);
or U15729 (N_15729,N_6739,N_11397);
xnor U15730 (N_15730,N_7558,N_12354);
nand U15731 (N_15731,N_11535,N_11880);
or U15732 (N_15732,N_10868,N_6337);
xnor U15733 (N_15733,N_11126,N_11597);
nand U15734 (N_15734,N_11337,N_8146);
xnor U15735 (N_15735,N_11883,N_10437);
nor U15736 (N_15736,N_7001,N_6744);
nand U15737 (N_15737,N_6990,N_11771);
or U15738 (N_15738,N_8198,N_8447);
nand U15739 (N_15739,N_10221,N_7850);
nor U15740 (N_15740,N_9660,N_7131);
and U15741 (N_15741,N_9998,N_7475);
or U15742 (N_15742,N_10334,N_10842);
and U15743 (N_15743,N_12232,N_10557);
or U15744 (N_15744,N_8954,N_6553);
or U15745 (N_15745,N_7665,N_12152);
xor U15746 (N_15746,N_9571,N_7449);
nor U15747 (N_15747,N_12225,N_9119);
and U15748 (N_15748,N_11768,N_12446);
and U15749 (N_15749,N_7035,N_11732);
and U15750 (N_15750,N_10451,N_7987);
and U15751 (N_15751,N_7387,N_11080);
or U15752 (N_15752,N_11211,N_8661);
and U15753 (N_15753,N_8469,N_10143);
nand U15754 (N_15754,N_9793,N_11152);
and U15755 (N_15755,N_7549,N_10874);
nand U15756 (N_15756,N_11799,N_8884);
and U15757 (N_15757,N_10643,N_11055);
or U15758 (N_15758,N_6714,N_10863);
and U15759 (N_15759,N_6623,N_10274);
nand U15760 (N_15760,N_8854,N_10926);
nand U15761 (N_15761,N_7799,N_10421);
or U15762 (N_15762,N_11593,N_8347);
and U15763 (N_15763,N_11829,N_10410);
or U15764 (N_15764,N_7485,N_10720);
nor U15765 (N_15765,N_7067,N_6707);
nand U15766 (N_15766,N_12112,N_11953);
nand U15767 (N_15767,N_6619,N_8103);
nor U15768 (N_15768,N_10140,N_6869);
and U15769 (N_15769,N_9268,N_10540);
nor U15770 (N_15770,N_8782,N_9656);
or U15771 (N_15771,N_6349,N_9310);
and U15772 (N_15772,N_11737,N_7345);
xor U15773 (N_15773,N_10834,N_11333);
nor U15774 (N_15774,N_8219,N_9893);
nand U15775 (N_15775,N_10662,N_11821);
xor U15776 (N_15776,N_7200,N_11347);
and U15777 (N_15777,N_10116,N_11130);
xnor U15778 (N_15778,N_6407,N_8783);
and U15779 (N_15779,N_11726,N_10263);
nand U15780 (N_15780,N_9273,N_7299);
nor U15781 (N_15781,N_12197,N_7187);
and U15782 (N_15782,N_11613,N_7088);
xnor U15783 (N_15783,N_7443,N_7178);
or U15784 (N_15784,N_10195,N_7263);
nand U15785 (N_15785,N_10869,N_7368);
nor U15786 (N_15786,N_9114,N_9621);
or U15787 (N_15787,N_8612,N_7198);
nand U15788 (N_15788,N_7809,N_11890);
nand U15789 (N_15789,N_9498,N_12406);
or U15790 (N_15790,N_11504,N_7984);
nand U15791 (N_15791,N_12436,N_12414);
nand U15792 (N_15792,N_12069,N_7688);
and U15793 (N_15793,N_7110,N_11248);
or U15794 (N_15794,N_8797,N_6965);
nand U15795 (N_15795,N_10987,N_7035);
nand U15796 (N_15796,N_6842,N_6318);
nor U15797 (N_15797,N_11190,N_6578);
and U15798 (N_15798,N_6288,N_8062);
nor U15799 (N_15799,N_10445,N_6618);
nor U15800 (N_15800,N_8589,N_7582);
and U15801 (N_15801,N_7249,N_7630);
nand U15802 (N_15802,N_7457,N_9521);
and U15803 (N_15803,N_12309,N_10470);
nand U15804 (N_15804,N_7787,N_11757);
nor U15805 (N_15805,N_8893,N_7775);
and U15806 (N_15806,N_7854,N_10366);
nand U15807 (N_15807,N_7655,N_9483);
nor U15808 (N_15808,N_9002,N_8297);
or U15809 (N_15809,N_6287,N_7311);
nor U15810 (N_15810,N_10459,N_6732);
nor U15811 (N_15811,N_10517,N_6574);
nor U15812 (N_15812,N_8687,N_6395);
nand U15813 (N_15813,N_9789,N_8643);
nand U15814 (N_15814,N_9672,N_12445);
or U15815 (N_15815,N_7965,N_11696);
or U15816 (N_15816,N_12082,N_9196);
nand U15817 (N_15817,N_6744,N_11867);
nand U15818 (N_15818,N_8890,N_8769);
nor U15819 (N_15819,N_10220,N_11032);
nor U15820 (N_15820,N_9374,N_11882);
or U15821 (N_15821,N_7697,N_9856);
nand U15822 (N_15822,N_11727,N_10065);
xor U15823 (N_15823,N_12402,N_9600);
nor U15824 (N_15824,N_11218,N_9545);
nor U15825 (N_15825,N_6289,N_6997);
and U15826 (N_15826,N_10908,N_9288);
nor U15827 (N_15827,N_10196,N_8569);
and U15828 (N_15828,N_8778,N_12297);
nand U15829 (N_15829,N_9049,N_11670);
and U15830 (N_15830,N_6454,N_9304);
nor U15831 (N_15831,N_9688,N_10216);
nor U15832 (N_15832,N_11488,N_11119);
nor U15833 (N_15833,N_10541,N_8711);
or U15834 (N_15834,N_10658,N_11618);
nor U15835 (N_15835,N_6424,N_11208);
and U15836 (N_15836,N_10341,N_10460);
xor U15837 (N_15837,N_11523,N_9578);
nor U15838 (N_15838,N_10261,N_8627);
or U15839 (N_15839,N_10703,N_12400);
xnor U15840 (N_15840,N_8809,N_11912);
and U15841 (N_15841,N_8979,N_7677);
nor U15842 (N_15842,N_6884,N_7039);
nor U15843 (N_15843,N_11178,N_7724);
and U15844 (N_15844,N_9518,N_6924);
or U15845 (N_15845,N_6788,N_6647);
or U15846 (N_15846,N_11391,N_10443);
nor U15847 (N_15847,N_11203,N_6526);
or U15848 (N_15848,N_10707,N_9322);
xor U15849 (N_15849,N_8303,N_10188);
nor U15850 (N_15850,N_9501,N_6438);
nand U15851 (N_15851,N_6436,N_8843);
nand U15852 (N_15852,N_12389,N_12306);
nand U15853 (N_15853,N_10074,N_9323);
nand U15854 (N_15854,N_7570,N_6853);
or U15855 (N_15855,N_11044,N_7865);
xor U15856 (N_15856,N_7022,N_9753);
or U15857 (N_15857,N_8079,N_7463);
or U15858 (N_15858,N_10099,N_7373);
nor U15859 (N_15859,N_12051,N_10733);
nor U15860 (N_15860,N_12299,N_12181);
or U15861 (N_15861,N_7226,N_9381);
xnor U15862 (N_15862,N_11984,N_8232);
or U15863 (N_15863,N_11197,N_8951);
or U15864 (N_15864,N_8473,N_9631);
or U15865 (N_15865,N_8923,N_10215);
and U15866 (N_15866,N_7101,N_10920);
nor U15867 (N_15867,N_10202,N_12353);
nor U15868 (N_15868,N_11194,N_9532);
nor U15869 (N_15869,N_9785,N_7580);
xor U15870 (N_15870,N_6902,N_8605);
and U15871 (N_15871,N_7444,N_6390);
or U15872 (N_15872,N_9669,N_11728);
or U15873 (N_15873,N_10957,N_11305);
xor U15874 (N_15874,N_6993,N_10930);
xnor U15875 (N_15875,N_7809,N_11035);
nand U15876 (N_15876,N_8902,N_9474);
xnor U15877 (N_15877,N_7335,N_9906);
or U15878 (N_15878,N_11768,N_9799);
nor U15879 (N_15879,N_10639,N_11825);
nand U15880 (N_15880,N_8874,N_10300);
or U15881 (N_15881,N_8311,N_10846);
nor U15882 (N_15882,N_8741,N_6532);
xor U15883 (N_15883,N_10549,N_8096);
xnor U15884 (N_15884,N_9348,N_8301);
xnor U15885 (N_15885,N_10141,N_9801);
nor U15886 (N_15886,N_12038,N_8242);
and U15887 (N_15887,N_6828,N_11351);
nor U15888 (N_15888,N_8191,N_10348);
or U15889 (N_15889,N_10141,N_12369);
nand U15890 (N_15890,N_11118,N_6487);
and U15891 (N_15891,N_8427,N_9598);
nand U15892 (N_15892,N_6951,N_10715);
nand U15893 (N_15893,N_10790,N_6575);
or U15894 (N_15894,N_11756,N_12109);
nand U15895 (N_15895,N_10708,N_8880);
or U15896 (N_15896,N_7619,N_9150);
xor U15897 (N_15897,N_7696,N_8857);
nand U15898 (N_15898,N_10763,N_6255);
or U15899 (N_15899,N_7133,N_8232);
and U15900 (N_15900,N_10074,N_7214);
nor U15901 (N_15901,N_8687,N_6929);
nand U15902 (N_15902,N_12259,N_7070);
or U15903 (N_15903,N_11835,N_7348);
and U15904 (N_15904,N_8575,N_6310);
nand U15905 (N_15905,N_8747,N_10863);
or U15906 (N_15906,N_10478,N_6435);
and U15907 (N_15907,N_8772,N_6658);
nand U15908 (N_15908,N_12009,N_11895);
xor U15909 (N_15909,N_6418,N_6680);
nor U15910 (N_15910,N_12266,N_11711);
and U15911 (N_15911,N_11740,N_12198);
or U15912 (N_15912,N_8989,N_9042);
xor U15913 (N_15913,N_9502,N_9618);
or U15914 (N_15914,N_7724,N_8572);
or U15915 (N_15915,N_9182,N_7573);
or U15916 (N_15916,N_8308,N_6553);
and U15917 (N_15917,N_11123,N_6352);
and U15918 (N_15918,N_6748,N_7186);
nor U15919 (N_15919,N_11738,N_10018);
or U15920 (N_15920,N_9058,N_8551);
and U15921 (N_15921,N_8495,N_11729);
nor U15922 (N_15922,N_6278,N_10277);
nor U15923 (N_15923,N_6650,N_11952);
or U15924 (N_15924,N_9903,N_7965);
and U15925 (N_15925,N_10749,N_7203);
or U15926 (N_15926,N_11493,N_11170);
nor U15927 (N_15927,N_9140,N_7267);
or U15928 (N_15928,N_9997,N_7609);
nand U15929 (N_15929,N_6930,N_11805);
and U15930 (N_15930,N_12350,N_10857);
and U15931 (N_15931,N_6623,N_7485);
or U15932 (N_15932,N_8334,N_7014);
xnor U15933 (N_15933,N_12248,N_10227);
nor U15934 (N_15934,N_11020,N_6320);
nor U15935 (N_15935,N_8210,N_10395);
nor U15936 (N_15936,N_7191,N_11795);
nand U15937 (N_15937,N_8333,N_10312);
or U15938 (N_15938,N_7980,N_11046);
nor U15939 (N_15939,N_11128,N_12417);
and U15940 (N_15940,N_11090,N_10376);
xnor U15941 (N_15941,N_11535,N_6820);
or U15942 (N_15942,N_7175,N_8309);
nand U15943 (N_15943,N_6602,N_11261);
or U15944 (N_15944,N_7389,N_10949);
nand U15945 (N_15945,N_10978,N_9996);
or U15946 (N_15946,N_9812,N_7160);
xnor U15947 (N_15947,N_11140,N_9202);
or U15948 (N_15948,N_7058,N_8175);
nand U15949 (N_15949,N_7412,N_10562);
nor U15950 (N_15950,N_8801,N_11999);
nor U15951 (N_15951,N_11898,N_8696);
xnor U15952 (N_15952,N_10660,N_8548);
and U15953 (N_15953,N_12479,N_11986);
nor U15954 (N_15954,N_11844,N_8972);
nand U15955 (N_15955,N_9316,N_9827);
or U15956 (N_15956,N_9141,N_10125);
nor U15957 (N_15957,N_10318,N_9826);
nor U15958 (N_15958,N_8701,N_12493);
or U15959 (N_15959,N_6883,N_11259);
or U15960 (N_15960,N_11470,N_12197);
or U15961 (N_15961,N_12236,N_9488);
nand U15962 (N_15962,N_7122,N_7936);
nand U15963 (N_15963,N_9734,N_7719);
nand U15964 (N_15964,N_8386,N_8589);
nand U15965 (N_15965,N_8907,N_6648);
nand U15966 (N_15966,N_6348,N_9705);
or U15967 (N_15967,N_6748,N_9675);
nand U15968 (N_15968,N_8508,N_10228);
and U15969 (N_15969,N_10273,N_7806);
and U15970 (N_15970,N_6807,N_9183);
and U15971 (N_15971,N_6453,N_11632);
nand U15972 (N_15972,N_7016,N_8108);
xor U15973 (N_15973,N_6404,N_7317);
nor U15974 (N_15974,N_11548,N_10462);
nand U15975 (N_15975,N_7261,N_8827);
and U15976 (N_15976,N_12106,N_10640);
xnor U15977 (N_15977,N_8469,N_10572);
nor U15978 (N_15978,N_11043,N_6301);
xnor U15979 (N_15979,N_9057,N_11623);
or U15980 (N_15980,N_7159,N_11575);
xnor U15981 (N_15981,N_8902,N_11230);
nor U15982 (N_15982,N_10518,N_7019);
or U15983 (N_15983,N_6533,N_6413);
nor U15984 (N_15984,N_7329,N_10867);
or U15985 (N_15985,N_8596,N_8589);
or U15986 (N_15986,N_9664,N_11160);
xnor U15987 (N_15987,N_7242,N_7634);
nor U15988 (N_15988,N_7822,N_11938);
nand U15989 (N_15989,N_8927,N_12404);
and U15990 (N_15990,N_8597,N_8858);
nor U15991 (N_15991,N_8361,N_7910);
and U15992 (N_15992,N_6761,N_11771);
nor U15993 (N_15993,N_6747,N_11669);
nor U15994 (N_15994,N_6803,N_6632);
nor U15995 (N_15995,N_10724,N_8891);
or U15996 (N_15996,N_6978,N_7995);
nand U15997 (N_15997,N_11025,N_10991);
xnor U15998 (N_15998,N_12456,N_10126);
nor U15999 (N_15999,N_12120,N_10914);
nor U16000 (N_16000,N_12141,N_7280);
or U16001 (N_16001,N_7411,N_9777);
nand U16002 (N_16002,N_8753,N_11980);
and U16003 (N_16003,N_7195,N_12258);
nand U16004 (N_16004,N_11029,N_10504);
and U16005 (N_16005,N_6445,N_11233);
or U16006 (N_16006,N_8466,N_11018);
or U16007 (N_16007,N_10763,N_8866);
nor U16008 (N_16008,N_10380,N_11306);
nor U16009 (N_16009,N_12193,N_8564);
nor U16010 (N_16010,N_9672,N_7989);
and U16011 (N_16011,N_11163,N_6526);
and U16012 (N_16012,N_7993,N_6558);
nor U16013 (N_16013,N_10417,N_7978);
nand U16014 (N_16014,N_12380,N_6637);
nand U16015 (N_16015,N_7848,N_12110);
nand U16016 (N_16016,N_10937,N_10436);
and U16017 (N_16017,N_6984,N_9921);
nand U16018 (N_16018,N_9414,N_7139);
xor U16019 (N_16019,N_11465,N_11056);
nand U16020 (N_16020,N_10550,N_9243);
nor U16021 (N_16021,N_10828,N_9443);
nor U16022 (N_16022,N_11147,N_11354);
nor U16023 (N_16023,N_11886,N_12304);
nor U16024 (N_16024,N_11547,N_9560);
and U16025 (N_16025,N_6305,N_8859);
and U16026 (N_16026,N_11117,N_11407);
and U16027 (N_16027,N_7366,N_8821);
or U16028 (N_16028,N_7284,N_12423);
nor U16029 (N_16029,N_11113,N_7694);
or U16030 (N_16030,N_11514,N_8065);
and U16031 (N_16031,N_9086,N_10484);
nor U16032 (N_16032,N_9363,N_11447);
nor U16033 (N_16033,N_7278,N_9099);
xor U16034 (N_16034,N_8509,N_6285);
nor U16035 (N_16035,N_8585,N_9620);
or U16036 (N_16036,N_9665,N_11661);
and U16037 (N_16037,N_8291,N_12012);
and U16038 (N_16038,N_9865,N_7282);
and U16039 (N_16039,N_11533,N_9036);
or U16040 (N_16040,N_10837,N_9900);
nor U16041 (N_16041,N_6973,N_6473);
and U16042 (N_16042,N_10155,N_12307);
and U16043 (N_16043,N_11609,N_7431);
xnor U16044 (N_16044,N_11974,N_10222);
nand U16045 (N_16045,N_6870,N_6999);
and U16046 (N_16046,N_11481,N_8965);
or U16047 (N_16047,N_6797,N_12146);
nand U16048 (N_16048,N_7206,N_11524);
and U16049 (N_16049,N_8777,N_6434);
nor U16050 (N_16050,N_7637,N_8683);
nand U16051 (N_16051,N_7868,N_9341);
or U16052 (N_16052,N_9916,N_10881);
xor U16053 (N_16053,N_10063,N_9287);
or U16054 (N_16054,N_8984,N_7535);
nand U16055 (N_16055,N_7018,N_6614);
nor U16056 (N_16056,N_11581,N_11072);
and U16057 (N_16057,N_6268,N_8603);
nor U16058 (N_16058,N_6809,N_10414);
nand U16059 (N_16059,N_9671,N_8256);
and U16060 (N_16060,N_11491,N_7740);
xnor U16061 (N_16061,N_8767,N_12433);
nand U16062 (N_16062,N_6939,N_7588);
or U16063 (N_16063,N_10159,N_9852);
nand U16064 (N_16064,N_11172,N_8485);
nor U16065 (N_16065,N_6904,N_11260);
xnor U16066 (N_16066,N_6306,N_6517);
and U16067 (N_16067,N_10531,N_10841);
xor U16068 (N_16068,N_11106,N_8514);
and U16069 (N_16069,N_8070,N_11343);
and U16070 (N_16070,N_10116,N_12122);
or U16071 (N_16071,N_10621,N_9539);
or U16072 (N_16072,N_8112,N_8457);
or U16073 (N_16073,N_10521,N_6667);
or U16074 (N_16074,N_8811,N_9682);
or U16075 (N_16075,N_10258,N_12116);
nand U16076 (N_16076,N_6939,N_10252);
and U16077 (N_16077,N_10107,N_7176);
nand U16078 (N_16078,N_8280,N_11928);
or U16079 (N_16079,N_7895,N_7513);
and U16080 (N_16080,N_6524,N_9354);
and U16081 (N_16081,N_12004,N_11781);
xnor U16082 (N_16082,N_6513,N_8925);
or U16083 (N_16083,N_9897,N_6527);
nor U16084 (N_16084,N_8123,N_10347);
and U16085 (N_16085,N_11111,N_6319);
xor U16086 (N_16086,N_9743,N_10718);
and U16087 (N_16087,N_11523,N_6926);
and U16088 (N_16088,N_9819,N_7667);
or U16089 (N_16089,N_11502,N_6471);
nor U16090 (N_16090,N_6772,N_9543);
and U16091 (N_16091,N_10513,N_11459);
and U16092 (N_16092,N_11010,N_11825);
nand U16093 (N_16093,N_9611,N_11647);
xor U16094 (N_16094,N_11383,N_8396);
nand U16095 (N_16095,N_12477,N_7079);
nand U16096 (N_16096,N_10045,N_9386);
xnor U16097 (N_16097,N_6349,N_8266);
and U16098 (N_16098,N_8718,N_7211);
and U16099 (N_16099,N_8810,N_10066);
nor U16100 (N_16100,N_6677,N_8374);
and U16101 (N_16101,N_8442,N_10974);
and U16102 (N_16102,N_12451,N_12080);
nand U16103 (N_16103,N_6749,N_7684);
nand U16104 (N_16104,N_8963,N_6775);
nor U16105 (N_16105,N_11507,N_11187);
and U16106 (N_16106,N_11810,N_8995);
or U16107 (N_16107,N_6645,N_6333);
xor U16108 (N_16108,N_10035,N_9042);
nor U16109 (N_16109,N_7037,N_9379);
xnor U16110 (N_16110,N_8075,N_11577);
nand U16111 (N_16111,N_6304,N_9492);
or U16112 (N_16112,N_10805,N_9782);
nand U16113 (N_16113,N_12265,N_7529);
nand U16114 (N_16114,N_11847,N_12345);
and U16115 (N_16115,N_11269,N_9794);
nor U16116 (N_16116,N_8566,N_9159);
or U16117 (N_16117,N_6545,N_6390);
xnor U16118 (N_16118,N_8949,N_11592);
or U16119 (N_16119,N_10894,N_10448);
xor U16120 (N_16120,N_9594,N_11839);
nor U16121 (N_16121,N_10055,N_7915);
xnor U16122 (N_16122,N_7939,N_6351);
nor U16123 (N_16123,N_10424,N_7044);
nor U16124 (N_16124,N_9248,N_9003);
or U16125 (N_16125,N_8020,N_8580);
nand U16126 (N_16126,N_10458,N_12269);
nand U16127 (N_16127,N_7938,N_12048);
nand U16128 (N_16128,N_11594,N_9760);
or U16129 (N_16129,N_11394,N_8799);
nand U16130 (N_16130,N_7220,N_8105);
and U16131 (N_16131,N_7621,N_9156);
and U16132 (N_16132,N_9326,N_10106);
or U16133 (N_16133,N_11985,N_8981);
and U16134 (N_16134,N_9528,N_12290);
or U16135 (N_16135,N_12335,N_8649);
nor U16136 (N_16136,N_11280,N_6762);
xnor U16137 (N_16137,N_8547,N_11876);
nor U16138 (N_16138,N_6283,N_8442);
and U16139 (N_16139,N_9114,N_10655);
nand U16140 (N_16140,N_6912,N_9287);
nor U16141 (N_16141,N_9330,N_8841);
or U16142 (N_16142,N_7327,N_8481);
or U16143 (N_16143,N_12377,N_8818);
or U16144 (N_16144,N_6399,N_7767);
or U16145 (N_16145,N_10690,N_11964);
nand U16146 (N_16146,N_8822,N_9656);
or U16147 (N_16147,N_9087,N_6354);
or U16148 (N_16148,N_12225,N_10391);
nor U16149 (N_16149,N_11765,N_10336);
and U16150 (N_16150,N_9248,N_7833);
nand U16151 (N_16151,N_11214,N_9400);
or U16152 (N_16152,N_7089,N_10844);
or U16153 (N_16153,N_7503,N_9614);
or U16154 (N_16154,N_12172,N_7836);
xor U16155 (N_16155,N_8501,N_8438);
nand U16156 (N_16156,N_9552,N_11446);
xnor U16157 (N_16157,N_6686,N_9312);
nor U16158 (N_16158,N_6372,N_8708);
or U16159 (N_16159,N_7017,N_8468);
and U16160 (N_16160,N_8303,N_6267);
or U16161 (N_16161,N_8393,N_11147);
nor U16162 (N_16162,N_10348,N_11263);
or U16163 (N_16163,N_8493,N_11591);
and U16164 (N_16164,N_7589,N_11961);
and U16165 (N_16165,N_7521,N_7192);
or U16166 (N_16166,N_10115,N_9892);
nor U16167 (N_16167,N_7636,N_11426);
and U16168 (N_16168,N_11266,N_7399);
or U16169 (N_16169,N_7535,N_11781);
xnor U16170 (N_16170,N_8391,N_9659);
and U16171 (N_16171,N_7198,N_6645);
nand U16172 (N_16172,N_7373,N_9765);
and U16173 (N_16173,N_10310,N_9310);
xor U16174 (N_16174,N_6499,N_10264);
nor U16175 (N_16175,N_9267,N_8461);
or U16176 (N_16176,N_11752,N_6798);
or U16177 (N_16177,N_9940,N_6828);
nand U16178 (N_16178,N_8873,N_8565);
and U16179 (N_16179,N_10459,N_7783);
xor U16180 (N_16180,N_10864,N_9444);
nand U16181 (N_16181,N_7470,N_9891);
and U16182 (N_16182,N_8836,N_7890);
and U16183 (N_16183,N_11327,N_9461);
nand U16184 (N_16184,N_11755,N_7354);
or U16185 (N_16185,N_10111,N_11993);
and U16186 (N_16186,N_11943,N_6494);
xor U16187 (N_16187,N_12387,N_11828);
and U16188 (N_16188,N_6788,N_11905);
and U16189 (N_16189,N_9406,N_12485);
and U16190 (N_16190,N_8466,N_7506);
nand U16191 (N_16191,N_9843,N_6828);
xor U16192 (N_16192,N_7860,N_7602);
or U16193 (N_16193,N_10831,N_7864);
or U16194 (N_16194,N_6306,N_11927);
and U16195 (N_16195,N_9714,N_9854);
nand U16196 (N_16196,N_11525,N_7671);
nor U16197 (N_16197,N_11318,N_11812);
xnor U16198 (N_16198,N_6343,N_7805);
and U16199 (N_16199,N_8411,N_9161);
nor U16200 (N_16200,N_10892,N_7139);
and U16201 (N_16201,N_9115,N_11661);
nand U16202 (N_16202,N_10102,N_10962);
and U16203 (N_16203,N_9642,N_7602);
and U16204 (N_16204,N_7618,N_11905);
nor U16205 (N_16205,N_11926,N_8935);
nor U16206 (N_16206,N_8343,N_6790);
xnor U16207 (N_16207,N_9726,N_6660);
nand U16208 (N_16208,N_6762,N_7207);
or U16209 (N_16209,N_12183,N_11910);
and U16210 (N_16210,N_7200,N_6794);
and U16211 (N_16211,N_8900,N_6752);
and U16212 (N_16212,N_8460,N_10666);
or U16213 (N_16213,N_11152,N_12079);
nand U16214 (N_16214,N_8259,N_10030);
nor U16215 (N_16215,N_9032,N_8457);
xnor U16216 (N_16216,N_7844,N_9965);
nand U16217 (N_16217,N_8165,N_7892);
or U16218 (N_16218,N_7077,N_8952);
and U16219 (N_16219,N_8134,N_9474);
nand U16220 (N_16220,N_9034,N_10119);
xor U16221 (N_16221,N_11564,N_6757);
nand U16222 (N_16222,N_9719,N_7797);
and U16223 (N_16223,N_11695,N_11309);
nor U16224 (N_16224,N_8220,N_10428);
or U16225 (N_16225,N_7999,N_11007);
nand U16226 (N_16226,N_6957,N_6661);
and U16227 (N_16227,N_9716,N_6690);
and U16228 (N_16228,N_9407,N_8403);
or U16229 (N_16229,N_6903,N_10354);
nand U16230 (N_16230,N_10157,N_6355);
nor U16231 (N_16231,N_7327,N_6461);
nand U16232 (N_16232,N_8279,N_10269);
xnor U16233 (N_16233,N_7560,N_11329);
nor U16234 (N_16234,N_7193,N_7444);
nor U16235 (N_16235,N_11687,N_7242);
nand U16236 (N_16236,N_12374,N_8290);
and U16237 (N_16237,N_11700,N_7839);
and U16238 (N_16238,N_10744,N_7147);
nand U16239 (N_16239,N_12443,N_8141);
and U16240 (N_16240,N_11077,N_7861);
and U16241 (N_16241,N_11245,N_6669);
nand U16242 (N_16242,N_7105,N_7841);
and U16243 (N_16243,N_8271,N_10283);
nor U16244 (N_16244,N_7909,N_10941);
and U16245 (N_16245,N_10325,N_10335);
and U16246 (N_16246,N_9602,N_7493);
nand U16247 (N_16247,N_11381,N_6870);
nand U16248 (N_16248,N_10600,N_9365);
or U16249 (N_16249,N_11264,N_8776);
xnor U16250 (N_16250,N_12495,N_6619);
nor U16251 (N_16251,N_7965,N_11714);
nor U16252 (N_16252,N_9521,N_8490);
nand U16253 (N_16253,N_7872,N_10153);
and U16254 (N_16254,N_11727,N_11202);
or U16255 (N_16255,N_9988,N_10820);
nand U16256 (N_16256,N_12294,N_6321);
or U16257 (N_16257,N_6878,N_6460);
nor U16258 (N_16258,N_6381,N_9372);
nand U16259 (N_16259,N_10640,N_11845);
nor U16260 (N_16260,N_9932,N_11460);
and U16261 (N_16261,N_9950,N_8645);
nor U16262 (N_16262,N_7223,N_6547);
nand U16263 (N_16263,N_6254,N_10773);
nor U16264 (N_16264,N_9165,N_12200);
or U16265 (N_16265,N_8143,N_7442);
nand U16266 (N_16266,N_8136,N_8780);
and U16267 (N_16267,N_6283,N_10971);
nor U16268 (N_16268,N_9964,N_10253);
xor U16269 (N_16269,N_6526,N_9577);
nand U16270 (N_16270,N_7280,N_7471);
or U16271 (N_16271,N_9231,N_8752);
or U16272 (N_16272,N_11112,N_6315);
xor U16273 (N_16273,N_12482,N_9746);
xor U16274 (N_16274,N_10844,N_10040);
xor U16275 (N_16275,N_8817,N_6948);
nor U16276 (N_16276,N_8332,N_7056);
nor U16277 (N_16277,N_6303,N_12469);
or U16278 (N_16278,N_9981,N_11691);
or U16279 (N_16279,N_8776,N_7166);
xnor U16280 (N_16280,N_7448,N_9024);
or U16281 (N_16281,N_9192,N_8583);
or U16282 (N_16282,N_12288,N_10134);
xor U16283 (N_16283,N_7676,N_12479);
nand U16284 (N_16284,N_7481,N_7385);
and U16285 (N_16285,N_7898,N_10773);
nand U16286 (N_16286,N_7848,N_12102);
or U16287 (N_16287,N_11707,N_10401);
and U16288 (N_16288,N_6880,N_10396);
and U16289 (N_16289,N_12330,N_11428);
nor U16290 (N_16290,N_11191,N_9811);
and U16291 (N_16291,N_9166,N_10910);
nor U16292 (N_16292,N_7440,N_10909);
nor U16293 (N_16293,N_12495,N_6927);
or U16294 (N_16294,N_9535,N_10629);
nor U16295 (N_16295,N_9676,N_7869);
nor U16296 (N_16296,N_8440,N_8060);
and U16297 (N_16297,N_7637,N_9696);
and U16298 (N_16298,N_7101,N_7507);
and U16299 (N_16299,N_11570,N_9003);
nand U16300 (N_16300,N_11407,N_10099);
nor U16301 (N_16301,N_6467,N_6616);
or U16302 (N_16302,N_7654,N_7858);
nor U16303 (N_16303,N_6306,N_8850);
and U16304 (N_16304,N_7516,N_9879);
nor U16305 (N_16305,N_7049,N_10884);
nand U16306 (N_16306,N_7823,N_10497);
nand U16307 (N_16307,N_8960,N_8549);
and U16308 (N_16308,N_10150,N_7821);
nand U16309 (N_16309,N_7605,N_8358);
xor U16310 (N_16310,N_12395,N_10192);
nand U16311 (N_16311,N_9776,N_10771);
nor U16312 (N_16312,N_10102,N_11460);
or U16313 (N_16313,N_8640,N_11641);
and U16314 (N_16314,N_10768,N_11500);
nor U16315 (N_16315,N_12053,N_10231);
xor U16316 (N_16316,N_8936,N_11756);
nor U16317 (N_16317,N_6427,N_10158);
or U16318 (N_16318,N_9387,N_6435);
or U16319 (N_16319,N_8502,N_9818);
xor U16320 (N_16320,N_11755,N_8156);
nor U16321 (N_16321,N_8866,N_10601);
nand U16322 (N_16322,N_10210,N_10261);
or U16323 (N_16323,N_10538,N_8012);
and U16324 (N_16324,N_10639,N_8366);
xor U16325 (N_16325,N_7684,N_9134);
nand U16326 (N_16326,N_8071,N_11053);
nor U16327 (N_16327,N_8746,N_8226);
xnor U16328 (N_16328,N_8488,N_12414);
or U16329 (N_16329,N_11207,N_10587);
and U16330 (N_16330,N_6995,N_9645);
nand U16331 (N_16331,N_6533,N_11079);
xor U16332 (N_16332,N_10957,N_6483);
xnor U16333 (N_16333,N_9828,N_7280);
nand U16334 (N_16334,N_8693,N_10720);
or U16335 (N_16335,N_6679,N_10497);
and U16336 (N_16336,N_6359,N_11297);
xor U16337 (N_16337,N_9367,N_8976);
or U16338 (N_16338,N_10538,N_8668);
or U16339 (N_16339,N_9948,N_6361);
or U16340 (N_16340,N_11968,N_6500);
nand U16341 (N_16341,N_7624,N_6842);
xnor U16342 (N_16342,N_9437,N_11332);
nand U16343 (N_16343,N_7821,N_12475);
or U16344 (N_16344,N_9196,N_9641);
or U16345 (N_16345,N_11659,N_10781);
xor U16346 (N_16346,N_9728,N_8325);
and U16347 (N_16347,N_6926,N_8810);
and U16348 (N_16348,N_10236,N_9531);
nand U16349 (N_16349,N_8019,N_9924);
nor U16350 (N_16350,N_7008,N_7392);
nand U16351 (N_16351,N_6729,N_9380);
and U16352 (N_16352,N_9010,N_11431);
nand U16353 (N_16353,N_10412,N_6851);
and U16354 (N_16354,N_10031,N_8981);
nor U16355 (N_16355,N_9844,N_11674);
nor U16356 (N_16356,N_10760,N_11093);
and U16357 (N_16357,N_8223,N_8311);
or U16358 (N_16358,N_9007,N_7894);
nand U16359 (N_16359,N_11866,N_10916);
nor U16360 (N_16360,N_7433,N_9589);
xnor U16361 (N_16361,N_12362,N_8138);
or U16362 (N_16362,N_11341,N_9511);
nor U16363 (N_16363,N_9684,N_8232);
or U16364 (N_16364,N_7270,N_11574);
nor U16365 (N_16365,N_11164,N_11246);
or U16366 (N_16366,N_6588,N_6928);
nand U16367 (N_16367,N_6658,N_10632);
nor U16368 (N_16368,N_11792,N_6691);
or U16369 (N_16369,N_12037,N_11797);
and U16370 (N_16370,N_6703,N_7587);
nand U16371 (N_16371,N_11174,N_7062);
nand U16372 (N_16372,N_11135,N_12484);
and U16373 (N_16373,N_10824,N_9822);
xor U16374 (N_16374,N_9080,N_7375);
and U16375 (N_16375,N_11157,N_11608);
and U16376 (N_16376,N_6864,N_6528);
and U16377 (N_16377,N_6822,N_8579);
nor U16378 (N_16378,N_11131,N_10318);
or U16379 (N_16379,N_9906,N_12291);
nor U16380 (N_16380,N_8268,N_12070);
and U16381 (N_16381,N_10502,N_9326);
and U16382 (N_16382,N_7820,N_6813);
and U16383 (N_16383,N_9306,N_12014);
nor U16384 (N_16384,N_10227,N_8158);
xnor U16385 (N_16385,N_11371,N_11739);
or U16386 (N_16386,N_9456,N_6730);
nor U16387 (N_16387,N_10970,N_10843);
xnor U16388 (N_16388,N_12121,N_9429);
nand U16389 (N_16389,N_12139,N_7296);
nor U16390 (N_16390,N_9393,N_7494);
or U16391 (N_16391,N_10881,N_10140);
nor U16392 (N_16392,N_8314,N_8937);
xor U16393 (N_16393,N_11157,N_7324);
nand U16394 (N_16394,N_12372,N_11857);
nand U16395 (N_16395,N_10033,N_9180);
xor U16396 (N_16396,N_11637,N_8006);
and U16397 (N_16397,N_7321,N_8039);
nor U16398 (N_16398,N_9987,N_9521);
and U16399 (N_16399,N_7066,N_8917);
and U16400 (N_16400,N_10108,N_7743);
nor U16401 (N_16401,N_9974,N_12397);
or U16402 (N_16402,N_8714,N_8507);
and U16403 (N_16403,N_10187,N_11288);
or U16404 (N_16404,N_12137,N_10680);
nor U16405 (N_16405,N_10277,N_11657);
and U16406 (N_16406,N_6514,N_8683);
or U16407 (N_16407,N_7575,N_7713);
nand U16408 (N_16408,N_10771,N_11242);
or U16409 (N_16409,N_12233,N_6651);
nor U16410 (N_16410,N_8290,N_10806);
nand U16411 (N_16411,N_9677,N_9012);
or U16412 (N_16412,N_6412,N_8610);
or U16413 (N_16413,N_12109,N_6365);
nor U16414 (N_16414,N_6617,N_10735);
nor U16415 (N_16415,N_8050,N_7483);
and U16416 (N_16416,N_8313,N_6364);
or U16417 (N_16417,N_9886,N_9938);
or U16418 (N_16418,N_8842,N_11025);
or U16419 (N_16419,N_12076,N_8043);
or U16420 (N_16420,N_6374,N_10118);
nand U16421 (N_16421,N_12442,N_9960);
nand U16422 (N_16422,N_8266,N_11719);
nand U16423 (N_16423,N_11754,N_10659);
or U16424 (N_16424,N_11688,N_12055);
nand U16425 (N_16425,N_10729,N_9814);
nor U16426 (N_16426,N_8908,N_6555);
nor U16427 (N_16427,N_11232,N_11814);
and U16428 (N_16428,N_7204,N_9122);
or U16429 (N_16429,N_11273,N_8796);
xor U16430 (N_16430,N_11205,N_10074);
nand U16431 (N_16431,N_9182,N_10703);
or U16432 (N_16432,N_8822,N_12283);
or U16433 (N_16433,N_9870,N_9476);
nor U16434 (N_16434,N_8535,N_10445);
or U16435 (N_16435,N_7655,N_6662);
nand U16436 (N_16436,N_8343,N_6900);
nand U16437 (N_16437,N_12418,N_8835);
nor U16438 (N_16438,N_10794,N_8795);
nand U16439 (N_16439,N_9132,N_11831);
or U16440 (N_16440,N_7773,N_11595);
nand U16441 (N_16441,N_6942,N_7428);
xor U16442 (N_16442,N_8482,N_8711);
nand U16443 (N_16443,N_9539,N_9909);
nor U16444 (N_16444,N_7471,N_10129);
and U16445 (N_16445,N_10768,N_10005);
and U16446 (N_16446,N_8129,N_7949);
and U16447 (N_16447,N_12414,N_8917);
nand U16448 (N_16448,N_6977,N_11067);
xnor U16449 (N_16449,N_11929,N_10876);
or U16450 (N_16450,N_12022,N_10472);
and U16451 (N_16451,N_8895,N_7924);
nor U16452 (N_16452,N_11230,N_7115);
and U16453 (N_16453,N_11308,N_12446);
nor U16454 (N_16454,N_11285,N_11550);
nor U16455 (N_16455,N_9049,N_11595);
nor U16456 (N_16456,N_6251,N_7188);
nor U16457 (N_16457,N_6476,N_11697);
nor U16458 (N_16458,N_10207,N_9048);
and U16459 (N_16459,N_10968,N_9187);
or U16460 (N_16460,N_7841,N_9690);
nor U16461 (N_16461,N_6420,N_10237);
and U16462 (N_16462,N_9095,N_10678);
and U16463 (N_16463,N_7218,N_12042);
or U16464 (N_16464,N_9866,N_11615);
nor U16465 (N_16465,N_7745,N_10589);
and U16466 (N_16466,N_11086,N_11511);
nor U16467 (N_16467,N_8170,N_7257);
or U16468 (N_16468,N_7600,N_11839);
nand U16469 (N_16469,N_6633,N_10239);
nand U16470 (N_16470,N_7497,N_10046);
nor U16471 (N_16471,N_7773,N_11501);
nor U16472 (N_16472,N_9822,N_6263);
or U16473 (N_16473,N_8324,N_10941);
nand U16474 (N_16474,N_7755,N_6973);
or U16475 (N_16475,N_6760,N_11873);
nor U16476 (N_16476,N_9036,N_7826);
nor U16477 (N_16477,N_11529,N_10777);
nor U16478 (N_16478,N_10684,N_8913);
and U16479 (N_16479,N_10304,N_7554);
nand U16480 (N_16480,N_11280,N_6686);
nand U16481 (N_16481,N_11976,N_7550);
or U16482 (N_16482,N_9511,N_10820);
or U16483 (N_16483,N_7179,N_12014);
or U16484 (N_16484,N_7003,N_6329);
and U16485 (N_16485,N_7718,N_8683);
nor U16486 (N_16486,N_7398,N_8604);
nand U16487 (N_16487,N_10278,N_9089);
xor U16488 (N_16488,N_10276,N_6730);
or U16489 (N_16489,N_10408,N_7757);
nand U16490 (N_16490,N_7836,N_8473);
or U16491 (N_16491,N_9168,N_11489);
and U16492 (N_16492,N_12225,N_7491);
nor U16493 (N_16493,N_11195,N_6985);
nand U16494 (N_16494,N_6660,N_7409);
nand U16495 (N_16495,N_7227,N_10080);
or U16496 (N_16496,N_7490,N_11276);
and U16497 (N_16497,N_11813,N_7700);
and U16498 (N_16498,N_8121,N_7740);
nand U16499 (N_16499,N_11211,N_12470);
and U16500 (N_16500,N_6373,N_9253);
and U16501 (N_16501,N_8134,N_10115);
or U16502 (N_16502,N_7249,N_9794);
nand U16503 (N_16503,N_9399,N_6678);
nand U16504 (N_16504,N_12364,N_8930);
nand U16505 (N_16505,N_8510,N_9750);
and U16506 (N_16506,N_11091,N_11822);
or U16507 (N_16507,N_6525,N_8986);
nand U16508 (N_16508,N_9131,N_10026);
nor U16509 (N_16509,N_8947,N_9256);
nor U16510 (N_16510,N_8865,N_8170);
xor U16511 (N_16511,N_9476,N_6371);
and U16512 (N_16512,N_9269,N_10903);
nand U16513 (N_16513,N_11055,N_12212);
and U16514 (N_16514,N_6686,N_6885);
and U16515 (N_16515,N_9997,N_8318);
nor U16516 (N_16516,N_9029,N_11627);
and U16517 (N_16517,N_9000,N_9888);
and U16518 (N_16518,N_7988,N_6878);
or U16519 (N_16519,N_6351,N_11534);
nor U16520 (N_16520,N_12230,N_10125);
nor U16521 (N_16521,N_10900,N_7704);
nor U16522 (N_16522,N_8004,N_10429);
nor U16523 (N_16523,N_9072,N_9227);
nor U16524 (N_16524,N_10054,N_12142);
nand U16525 (N_16525,N_8584,N_11508);
nor U16526 (N_16526,N_6551,N_7664);
or U16527 (N_16527,N_8714,N_6518);
nor U16528 (N_16528,N_9446,N_11552);
and U16529 (N_16529,N_6720,N_10852);
nand U16530 (N_16530,N_8744,N_6616);
nand U16531 (N_16531,N_11819,N_7414);
or U16532 (N_16532,N_8569,N_9971);
nand U16533 (N_16533,N_8201,N_11727);
nor U16534 (N_16534,N_8802,N_11713);
nor U16535 (N_16535,N_8108,N_10341);
nor U16536 (N_16536,N_7502,N_11609);
or U16537 (N_16537,N_12289,N_8454);
or U16538 (N_16538,N_9998,N_8687);
xor U16539 (N_16539,N_11410,N_11479);
nor U16540 (N_16540,N_12204,N_8437);
nor U16541 (N_16541,N_11194,N_8286);
nor U16542 (N_16542,N_9126,N_8931);
nand U16543 (N_16543,N_9167,N_10586);
nand U16544 (N_16544,N_7766,N_11760);
nand U16545 (N_16545,N_10066,N_10977);
nand U16546 (N_16546,N_6588,N_6969);
and U16547 (N_16547,N_7470,N_10561);
or U16548 (N_16548,N_12408,N_8166);
or U16549 (N_16549,N_6830,N_7403);
xor U16550 (N_16550,N_9993,N_10772);
or U16551 (N_16551,N_11142,N_10625);
nor U16552 (N_16552,N_12115,N_10998);
and U16553 (N_16553,N_7159,N_10728);
nand U16554 (N_16554,N_7569,N_7375);
or U16555 (N_16555,N_11464,N_9475);
xor U16556 (N_16556,N_7522,N_7726);
nor U16557 (N_16557,N_10010,N_10793);
and U16558 (N_16558,N_7160,N_9270);
or U16559 (N_16559,N_11018,N_8352);
xor U16560 (N_16560,N_8233,N_10114);
or U16561 (N_16561,N_6287,N_7935);
nand U16562 (N_16562,N_10338,N_12058);
nor U16563 (N_16563,N_12476,N_7260);
nand U16564 (N_16564,N_7652,N_10078);
xnor U16565 (N_16565,N_8567,N_10490);
nand U16566 (N_16566,N_8491,N_8719);
xnor U16567 (N_16567,N_9553,N_12234);
and U16568 (N_16568,N_9707,N_9655);
and U16569 (N_16569,N_11783,N_6598);
nor U16570 (N_16570,N_7214,N_8655);
and U16571 (N_16571,N_11800,N_8569);
or U16572 (N_16572,N_11772,N_11680);
xor U16573 (N_16573,N_10029,N_8683);
and U16574 (N_16574,N_9829,N_7475);
or U16575 (N_16575,N_6403,N_10844);
nand U16576 (N_16576,N_8164,N_12134);
and U16577 (N_16577,N_7689,N_12349);
nor U16578 (N_16578,N_9279,N_8299);
nor U16579 (N_16579,N_8000,N_11407);
or U16580 (N_16580,N_11332,N_10211);
and U16581 (N_16581,N_11879,N_6654);
nor U16582 (N_16582,N_9646,N_10487);
nor U16583 (N_16583,N_9188,N_11182);
nor U16584 (N_16584,N_12062,N_10200);
nor U16585 (N_16585,N_6586,N_10261);
nor U16586 (N_16586,N_6811,N_10454);
or U16587 (N_16587,N_7710,N_9569);
nor U16588 (N_16588,N_9618,N_7031);
and U16589 (N_16589,N_7065,N_10986);
and U16590 (N_16590,N_11430,N_10895);
and U16591 (N_16591,N_9735,N_10452);
or U16592 (N_16592,N_11772,N_9719);
or U16593 (N_16593,N_9318,N_9862);
nor U16594 (N_16594,N_6884,N_12124);
or U16595 (N_16595,N_10923,N_9451);
nand U16596 (N_16596,N_7192,N_10631);
or U16597 (N_16597,N_7042,N_9790);
xnor U16598 (N_16598,N_11001,N_7431);
nand U16599 (N_16599,N_6879,N_11855);
nor U16600 (N_16600,N_8412,N_10494);
or U16601 (N_16601,N_6919,N_11396);
and U16602 (N_16602,N_7860,N_12279);
nor U16603 (N_16603,N_9175,N_8855);
or U16604 (N_16604,N_6822,N_12266);
nand U16605 (N_16605,N_12089,N_8858);
or U16606 (N_16606,N_10757,N_12070);
and U16607 (N_16607,N_10395,N_9274);
and U16608 (N_16608,N_10721,N_11890);
and U16609 (N_16609,N_9262,N_11619);
nor U16610 (N_16610,N_12498,N_10265);
nor U16611 (N_16611,N_9415,N_7413);
xor U16612 (N_16612,N_10080,N_8753);
and U16613 (N_16613,N_10920,N_10528);
nor U16614 (N_16614,N_6432,N_10743);
nand U16615 (N_16615,N_8200,N_7475);
or U16616 (N_16616,N_9753,N_12495);
nand U16617 (N_16617,N_7816,N_10528);
xor U16618 (N_16618,N_8031,N_6895);
and U16619 (N_16619,N_11678,N_11763);
nand U16620 (N_16620,N_11083,N_11559);
and U16621 (N_16621,N_9326,N_10461);
nand U16622 (N_16622,N_8124,N_8928);
or U16623 (N_16623,N_10017,N_8215);
nor U16624 (N_16624,N_6998,N_7327);
or U16625 (N_16625,N_6743,N_8236);
nor U16626 (N_16626,N_8204,N_7338);
xor U16627 (N_16627,N_11356,N_9803);
or U16628 (N_16628,N_8412,N_10977);
and U16629 (N_16629,N_10965,N_11999);
and U16630 (N_16630,N_7219,N_11115);
nor U16631 (N_16631,N_10337,N_11605);
xnor U16632 (N_16632,N_11447,N_12295);
or U16633 (N_16633,N_7266,N_8959);
nand U16634 (N_16634,N_8700,N_10031);
nor U16635 (N_16635,N_11800,N_6793);
nand U16636 (N_16636,N_8752,N_8196);
nand U16637 (N_16637,N_11744,N_12237);
nand U16638 (N_16638,N_9604,N_9309);
or U16639 (N_16639,N_12265,N_9685);
xnor U16640 (N_16640,N_7768,N_9463);
or U16641 (N_16641,N_6692,N_9465);
nand U16642 (N_16642,N_7415,N_7577);
and U16643 (N_16643,N_7155,N_10218);
nand U16644 (N_16644,N_10882,N_8578);
xnor U16645 (N_16645,N_7052,N_8568);
nand U16646 (N_16646,N_10112,N_10733);
or U16647 (N_16647,N_11926,N_8647);
and U16648 (N_16648,N_6646,N_10266);
nor U16649 (N_16649,N_7197,N_10217);
or U16650 (N_16650,N_12344,N_7817);
xor U16651 (N_16651,N_10079,N_7250);
and U16652 (N_16652,N_11439,N_10665);
and U16653 (N_16653,N_11509,N_7662);
nor U16654 (N_16654,N_6723,N_7986);
or U16655 (N_16655,N_8239,N_6904);
nor U16656 (N_16656,N_6612,N_7544);
or U16657 (N_16657,N_11304,N_11395);
nor U16658 (N_16658,N_8820,N_12416);
and U16659 (N_16659,N_11799,N_6322);
or U16660 (N_16660,N_8473,N_11288);
or U16661 (N_16661,N_6605,N_10038);
nor U16662 (N_16662,N_6525,N_9500);
nand U16663 (N_16663,N_6781,N_9693);
nor U16664 (N_16664,N_6720,N_8917);
nand U16665 (N_16665,N_12009,N_11488);
or U16666 (N_16666,N_7980,N_8812);
nor U16667 (N_16667,N_7047,N_11262);
nand U16668 (N_16668,N_11223,N_6316);
nand U16669 (N_16669,N_9717,N_9032);
and U16670 (N_16670,N_11454,N_6791);
and U16671 (N_16671,N_7752,N_7654);
or U16672 (N_16672,N_7387,N_9109);
and U16673 (N_16673,N_11885,N_11582);
nor U16674 (N_16674,N_6794,N_8279);
and U16675 (N_16675,N_12131,N_9981);
and U16676 (N_16676,N_8384,N_8394);
and U16677 (N_16677,N_10662,N_8643);
and U16678 (N_16678,N_10227,N_7506);
xnor U16679 (N_16679,N_11814,N_10058);
nand U16680 (N_16680,N_8886,N_12396);
nor U16681 (N_16681,N_12317,N_12065);
and U16682 (N_16682,N_6713,N_12337);
or U16683 (N_16683,N_6720,N_10740);
and U16684 (N_16684,N_8478,N_12298);
and U16685 (N_16685,N_7207,N_7511);
nor U16686 (N_16686,N_6753,N_9709);
nand U16687 (N_16687,N_7827,N_9419);
nand U16688 (N_16688,N_9564,N_11820);
and U16689 (N_16689,N_9832,N_8339);
xor U16690 (N_16690,N_6703,N_7215);
and U16691 (N_16691,N_10147,N_8237);
nor U16692 (N_16692,N_9712,N_12173);
and U16693 (N_16693,N_8514,N_9187);
or U16694 (N_16694,N_11906,N_9097);
xor U16695 (N_16695,N_11404,N_8269);
nand U16696 (N_16696,N_7118,N_8020);
or U16697 (N_16697,N_8737,N_7260);
nand U16698 (N_16698,N_6623,N_7715);
nor U16699 (N_16699,N_11440,N_9372);
nor U16700 (N_16700,N_11048,N_8224);
nand U16701 (N_16701,N_9725,N_7049);
nand U16702 (N_16702,N_7789,N_11965);
and U16703 (N_16703,N_12447,N_12064);
and U16704 (N_16704,N_6742,N_7095);
nand U16705 (N_16705,N_6779,N_8428);
and U16706 (N_16706,N_10428,N_12201);
nand U16707 (N_16707,N_10562,N_6816);
nand U16708 (N_16708,N_8163,N_9925);
and U16709 (N_16709,N_11226,N_7946);
and U16710 (N_16710,N_12224,N_12219);
and U16711 (N_16711,N_12254,N_9396);
nor U16712 (N_16712,N_9971,N_7814);
nor U16713 (N_16713,N_10909,N_10674);
nor U16714 (N_16714,N_9636,N_7282);
nand U16715 (N_16715,N_8485,N_10700);
nand U16716 (N_16716,N_12139,N_12407);
and U16717 (N_16717,N_11808,N_8063);
nand U16718 (N_16718,N_6976,N_12169);
or U16719 (N_16719,N_6307,N_11107);
or U16720 (N_16720,N_6901,N_7719);
or U16721 (N_16721,N_10858,N_8204);
and U16722 (N_16722,N_9674,N_8705);
or U16723 (N_16723,N_6358,N_9200);
or U16724 (N_16724,N_9024,N_7479);
nor U16725 (N_16725,N_9865,N_7592);
nor U16726 (N_16726,N_10157,N_7693);
xnor U16727 (N_16727,N_7438,N_8407);
nand U16728 (N_16728,N_6329,N_8902);
nand U16729 (N_16729,N_9180,N_11902);
xor U16730 (N_16730,N_6622,N_10563);
or U16731 (N_16731,N_6988,N_7956);
and U16732 (N_16732,N_8272,N_10829);
nand U16733 (N_16733,N_11363,N_11120);
nand U16734 (N_16734,N_9550,N_10930);
xor U16735 (N_16735,N_9346,N_11369);
or U16736 (N_16736,N_10034,N_9641);
or U16737 (N_16737,N_11773,N_8387);
and U16738 (N_16738,N_8023,N_9253);
xor U16739 (N_16739,N_11163,N_10789);
and U16740 (N_16740,N_10032,N_7589);
nor U16741 (N_16741,N_7618,N_8028);
and U16742 (N_16742,N_7886,N_12218);
nand U16743 (N_16743,N_8001,N_9627);
or U16744 (N_16744,N_7988,N_9122);
nand U16745 (N_16745,N_8786,N_11639);
nor U16746 (N_16746,N_6865,N_12016);
and U16747 (N_16747,N_8184,N_11472);
nand U16748 (N_16748,N_7331,N_11303);
and U16749 (N_16749,N_7032,N_7739);
nand U16750 (N_16750,N_6263,N_8695);
nor U16751 (N_16751,N_9419,N_8722);
nand U16752 (N_16752,N_7580,N_7402);
nand U16753 (N_16753,N_10891,N_8821);
nand U16754 (N_16754,N_7456,N_6587);
or U16755 (N_16755,N_12142,N_8723);
and U16756 (N_16756,N_10996,N_12283);
and U16757 (N_16757,N_10319,N_9908);
or U16758 (N_16758,N_9560,N_6748);
and U16759 (N_16759,N_11514,N_11499);
nor U16760 (N_16760,N_12066,N_10803);
or U16761 (N_16761,N_10430,N_9092);
nand U16762 (N_16762,N_10253,N_7058);
nor U16763 (N_16763,N_11493,N_7816);
and U16764 (N_16764,N_10239,N_7397);
nor U16765 (N_16765,N_10087,N_8411);
and U16766 (N_16766,N_7179,N_6978);
nand U16767 (N_16767,N_9449,N_10049);
xnor U16768 (N_16768,N_7044,N_8524);
nor U16769 (N_16769,N_6704,N_8463);
or U16770 (N_16770,N_6318,N_7331);
and U16771 (N_16771,N_10943,N_11509);
and U16772 (N_16772,N_9125,N_9994);
and U16773 (N_16773,N_7615,N_10723);
xnor U16774 (N_16774,N_8618,N_6400);
nand U16775 (N_16775,N_10158,N_10725);
nand U16776 (N_16776,N_9400,N_10194);
and U16777 (N_16777,N_9567,N_7837);
or U16778 (N_16778,N_7762,N_10322);
or U16779 (N_16779,N_10396,N_11501);
or U16780 (N_16780,N_11074,N_10441);
or U16781 (N_16781,N_9384,N_6374);
or U16782 (N_16782,N_8924,N_11943);
or U16783 (N_16783,N_10047,N_6802);
nand U16784 (N_16784,N_7434,N_9352);
or U16785 (N_16785,N_6870,N_7394);
nand U16786 (N_16786,N_11030,N_10576);
and U16787 (N_16787,N_8797,N_12246);
xnor U16788 (N_16788,N_12219,N_6336);
nor U16789 (N_16789,N_6673,N_7287);
nor U16790 (N_16790,N_9778,N_6765);
nand U16791 (N_16791,N_6652,N_8845);
xnor U16792 (N_16792,N_7316,N_12375);
xor U16793 (N_16793,N_7276,N_8262);
or U16794 (N_16794,N_11042,N_6433);
and U16795 (N_16795,N_11784,N_11961);
nand U16796 (N_16796,N_8393,N_10659);
xor U16797 (N_16797,N_9917,N_8575);
nor U16798 (N_16798,N_6362,N_7329);
nand U16799 (N_16799,N_10917,N_12130);
and U16800 (N_16800,N_10863,N_9252);
nand U16801 (N_16801,N_11571,N_7694);
and U16802 (N_16802,N_7702,N_7015);
and U16803 (N_16803,N_11428,N_9710);
nand U16804 (N_16804,N_11388,N_10594);
nand U16805 (N_16805,N_8631,N_8713);
or U16806 (N_16806,N_10317,N_12157);
nand U16807 (N_16807,N_12130,N_9621);
or U16808 (N_16808,N_10844,N_8714);
or U16809 (N_16809,N_9295,N_8639);
and U16810 (N_16810,N_11625,N_7723);
or U16811 (N_16811,N_11229,N_6333);
or U16812 (N_16812,N_11496,N_10661);
or U16813 (N_16813,N_9292,N_9982);
or U16814 (N_16814,N_9129,N_7525);
xor U16815 (N_16815,N_9636,N_10753);
or U16816 (N_16816,N_10731,N_6866);
or U16817 (N_16817,N_9151,N_8895);
nand U16818 (N_16818,N_6757,N_6535);
nand U16819 (N_16819,N_8459,N_12231);
xnor U16820 (N_16820,N_11595,N_8017);
xor U16821 (N_16821,N_12142,N_8667);
nand U16822 (N_16822,N_9530,N_7320);
and U16823 (N_16823,N_10619,N_9332);
and U16824 (N_16824,N_9407,N_7589);
xnor U16825 (N_16825,N_6701,N_7608);
or U16826 (N_16826,N_8387,N_8873);
nand U16827 (N_16827,N_9508,N_11941);
nor U16828 (N_16828,N_10516,N_11061);
and U16829 (N_16829,N_7803,N_7142);
nand U16830 (N_16830,N_7856,N_10542);
nand U16831 (N_16831,N_11397,N_7395);
or U16832 (N_16832,N_9317,N_7286);
or U16833 (N_16833,N_8470,N_11782);
and U16834 (N_16834,N_7270,N_7422);
or U16835 (N_16835,N_8999,N_9373);
xnor U16836 (N_16836,N_12364,N_6363);
nand U16837 (N_16837,N_7484,N_11544);
and U16838 (N_16838,N_9249,N_7889);
nand U16839 (N_16839,N_6449,N_8478);
and U16840 (N_16840,N_11555,N_8493);
or U16841 (N_16841,N_6354,N_6813);
or U16842 (N_16842,N_10198,N_8558);
nand U16843 (N_16843,N_11926,N_8960);
nand U16844 (N_16844,N_10053,N_6954);
or U16845 (N_16845,N_6798,N_10371);
and U16846 (N_16846,N_8581,N_11209);
nand U16847 (N_16847,N_10609,N_7859);
nor U16848 (N_16848,N_6705,N_11752);
nor U16849 (N_16849,N_7610,N_6546);
and U16850 (N_16850,N_10706,N_8104);
or U16851 (N_16851,N_10424,N_7625);
xnor U16852 (N_16852,N_7232,N_7247);
or U16853 (N_16853,N_10105,N_6297);
nand U16854 (N_16854,N_10067,N_8867);
or U16855 (N_16855,N_8912,N_11330);
nand U16856 (N_16856,N_7628,N_11314);
nor U16857 (N_16857,N_10756,N_7088);
or U16858 (N_16858,N_10510,N_7558);
or U16859 (N_16859,N_10793,N_9756);
nand U16860 (N_16860,N_9445,N_8442);
xnor U16861 (N_16861,N_7527,N_6559);
nor U16862 (N_16862,N_6721,N_12198);
nand U16863 (N_16863,N_8002,N_8944);
nor U16864 (N_16864,N_8851,N_6837);
and U16865 (N_16865,N_11382,N_12430);
nor U16866 (N_16866,N_8696,N_9033);
and U16867 (N_16867,N_10995,N_10355);
or U16868 (N_16868,N_9238,N_6712);
and U16869 (N_16869,N_6478,N_9219);
or U16870 (N_16870,N_11947,N_6344);
xnor U16871 (N_16871,N_10784,N_6537);
nand U16872 (N_16872,N_12062,N_10929);
and U16873 (N_16873,N_10879,N_9659);
nand U16874 (N_16874,N_11497,N_11575);
nor U16875 (N_16875,N_11839,N_7856);
or U16876 (N_16876,N_6586,N_9316);
nand U16877 (N_16877,N_6383,N_11054);
nand U16878 (N_16878,N_7977,N_10738);
nor U16879 (N_16879,N_11013,N_8115);
xnor U16880 (N_16880,N_8940,N_11498);
nand U16881 (N_16881,N_6957,N_8276);
or U16882 (N_16882,N_10399,N_9252);
and U16883 (N_16883,N_6260,N_7686);
or U16884 (N_16884,N_7091,N_9607);
nand U16885 (N_16885,N_7425,N_7790);
xnor U16886 (N_16886,N_11532,N_11290);
nor U16887 (N_16887,N_10340,N_7196);
nand U16888 (N_16888,N_6801,N_7662);
nand U16889 (N_16889,N_11469,N_7097);
nand U16890 (N_16890,N_6504,N_11714);
and U16891 (N_16891,N_10215,N_10254);
and U16892 (N_16892,N_9086,N_8142);
or U16893 (N_16893,N_12415,N_7795);
nor U16894 (N_16894,N_9123,N_10171);
nand U16895 (N_16895,N_7416,N_7747);
nor U16896 (N_16896,N_7890,N_8869);
nand U16897 (N_16897,N_9977,N_7520);
xnor U16898 (N_16898,N_11690,N_9058);
and U16899 (N_16899,N_10344,N_8686);
or U16900 (N_16900,N_7699,N_10776);
or U16901 (N_16901,N_6686,N_11625);
and U16902 (N_16902,N_11416,N_8136);
or U16903 (N_16903,N_7063,N_6814);
or U16904 (N_16904,N_12072,N_9245);
nand U16905 (N_16905,N_10719,N_12009);
xnor U16906 (N_16906,N_8520,N_8247);
or U16907 (N_16907,N_6803,N_9144);
xnor U16908 (N_16908,N_12333,N_10790);
and U16909 (N_16909,N_7815,N_7963);
nor U16910 (N_16910,N_9012,N_9048);
nand U16911 (N_16911,N_8899,N_8499);
or U16912 (N_16912,N_7415,N_7382);
or U16913 (N_16913,N_10060,N_11118);
nand U16914 (N_16914,N_9607,N_10946);
xor U16915 (N_16915,N_6447,N_11253);
nand U16916 (N_16916,N_7325,N_10530);
xnor U16917 (N_16917,N_12267,N_8750);
nor U16918 (N_16918,N_8759,N_12224);
or U16919 (N_16919,N_6315,N_9067);
nor U16920 (N_16920,N_9802,N_10869);
nand U16921 (N_16921,N_9528,N_12039);
nor U16922 (N_16922,N_8264,N_11103);
or U16923 (N_16923,N_9297,N_6354);
nor U16924 (N_16924,N_6306,N_11201);
or U16925 (N_16925,N_10969,N_8384);
or U16926 (N_16926,N_9362,N_10388);
nand U16927 (N_16927,N_8592,N_9942);
or U16928 (N_16928,N_8923,N_8222);
nand U16929 (N_16929,N_9706,N_10143);
or U16930 (N_16930,N_9358,N_8527);
or U16931 (N_16931,N_9195,N_6484);
nand U16932 (N_16932,N_6933,N_6542);
and U16933 (N_16933,N_12184,N_9191);
or U16934 (N_16934,N_10756,N_9542);
nor U16935 (N_16935,N_8985,N_7584);
nor U16936 (N_16936,N_8457,N_12011);
nand U16937 (N_16937,N_10156,N_9813);
nand U16938 (N_16938,N_11196,N_7803);
and U16939 (N_16939,N_11521,N_12333);
or U16940 (N_16940,N_11666,N_9019);
or U16941 (N_16941,N_10255,N_8356);
nand U16942 (N_16942,N_8638,N_6645);
xnor U16943 (N_16943,N_10487,N_6659);
and U16944 (N_16944,N_11935,N_6745);
and U16945 (N_16945,N_11065,N_11153);
and U16946 (N_16946,N_10330,N_7534);
nand U16947 (N_16947,N_6910,N_9815);
nand U16948 (N_16948,N_10944,N_7901);
or U16949 (N_16949,N_11187,N_7896);
nand U16950 (N_16950,N_7709,N_8251);
and U16951 (N_16951,N_12174,N_6727);
and U16952 (N_16952,N_11651,N_8567);
nand U16953 (N_16953,N_9533,N_9074);
nand U16954 (N_16954,N_7024,N_8062);
nor U16955 (N_16955,N_9884,N_12204);
nor U16956 (N_16956,N_10581,N_7589);
and U16957 (N_16957,N_7580,N_7066);
nor U16958 (N_16958,N_9632,N_6311);
and U16959 (N_16959,N_9808,N_7236);
or U16960 (N_16960,N_10571,N_6846);
nor U16961 (N_16961,N_9244,N_12218);
and U16962 (N_16962,N_10361,N_12175);
or U16963 (N_16963,N_9427,N_10629);
and U16964 (N_16964,N_10570,N_11641);
and U16965 (N_16965,N_7000,N_10868);
and U16966 (N_16966,N_6604,N_8657);
nor U16967 (N_16967,N_8292,N_9789);
or U16968 (N_16968,N_7136,N_9767);
xor U16969 (N_16969,N_10074,N_7513);
xnor U16970 (N_16970,N_10483,N_6472);
and U16971 (N_16971,N_11991,N_9719);
xor U16972 (N_16972,N_10795,N_10264);
or U16973 (N_16973,N_11560,N_8267);
or U16974 (N_16974,N_6450,N_8963);
and U16975 (N_16975,N_7497,N_11285);
and U16976 (N_16976,N_11723,N_6321);
nand U16977 (N_16977,N_8946,N_10258);
nand U16978 (N_16978,N_6947,N_7987);
or U16979 (N_16979,N_8413,N_9199);
nand U16980 (N_16980,N_7149,N_8640);
or U16981 (N_16981,N_11274,N_8394);
and U16982 (N_16982,N_7678,N_6733);
nor U16983 (N_16983,N_11381,N_8077);
and U16984 (N_16984,N_12117,N_12213);
nor U16985 (N_16985,N_11448,N_11438);
and U16986 (N_16986,N_8233,N_10058);
nand U16987 (N_16987,N_9275,N_7188);
xnor U16988 (N_16988,N_9908,N_8737);
nand U16989 (N_16989,N_11416,N_6304);
xnor U16990 (N_16990,N_8665,N_11007);
and U16991 (N_16991,N_12078,N_12147);
nor U16992 (N_16992,N_11759,N_12449);
or U16993 (N_16993,N_11863,N_6576);
nand U16994 (N_16994,N_7058,N_7998);
or U16995 (N_16995,N_7638,N_10109);
nor U16996 (N_16996,N_6735,N_9651);
and U16997 (N_16997,N_6725,N_10685);
or U16998 (N_16998,N_9804,N_10627);
nand U16999 (N_16999,N_9866,N_6982);
nand U17000 (N_17000,N_12255,N_8514);
nor U17001 (N_17001,N_11114,N_12063);
and U17002 (N_17002,N_11924,N_6911);
nand U17003 (N_17003,N_12359,N_11536);
nor U17004 (N_17004,N_11524,N_9809);
nand U17005 (N_17005,N_11248,N_8863);
nand U17006 (N_17006,N_6884,N_12344);
or U17007 (N_17007,N_7307,N_10712);
xnor U17008 (N_17008,N_11194,N_7883);
and U17009 (N_17009,N_6654,N_6423);
xor U17010 (N_17010,N_6858,N_7220);
and U17011 (N_17011,N_10347,N_9591);
xor U17012 (N_17012,N_8840,N_8799);
nor U17013 (N_17013,N_8512,N_7700);
nand U17014 (N_17014,N_12100,N_7467);
and U17015 (N_17015,N_9773,N_11129);
or U17016 (N_17016,N_7668,N_8902);
and U17017 (N_17017,N_8235,N_10229);
or U17018 (N_17018,N_7943,N_10707);
nor U17019 (N_17019,N_10338,N_11350);
and U17020 (N_17020,N_11153,N_7929);
nand U17021 (N_17021,N_11126,N_10192);
nor U17022 (N_17022,N_11413,N_11204);
nor U17023 (N_17023,N_6493,N_7296);
or U17024 (N_17024,N_10618,N_11156);
nor U17025 (N_17025,N_8964,N_7948);
and U17026 (N_17026,N_10014,N_10362);
and U17027 (N_17027,N_8214,N_8691);
nor U17028 (N_17028,N_11334,N_11504);
and U17029 (N_17029,N_12145,N_7322);
xor U17030 (N_17030,N_10323,N_8048);
and U17031 (N_17031,N_10493,N_6341);
nand U17032 (N_17032,N_10575,N_12407);
or U17033 (N_17033,N_7275,N_8477);
and U17034 (N_17034,N_12426,N_11880);
and U17035 (N_17035,N_11949,N_7088);
or U17036 (N_17036,N_11313,N_7166);
and U17037 (N_17037,N_8986,N_7360);
nand U17038 (N_17038,N_11832,N_9280);
nor U17039 (N_17039,N_10245,N_8143);
nand U17040 (N_17040,N_10944,N_8776);
nand U17041 (N_17041,N_11875,N_6864);
nor U17042 (N_17042,N_12184,N_10761);
nor U17043 (N_17043,N_11436,N_12138);
nor U17044 (N_17044,N_10873,N_11098);
xnor U17045 (N_17045,N_12472,N_11620);
nand U17046 (N_17046,N_6919,N_12327);
nand U17047 (N_17047,N_7209,N_7935);
or U17048 (N_17048,N_8241,N_6411);
and U17049 (N_17049,N_8891,N_6822);
and U17050 (N_17050,N_8794,N_11777);
or U17051 (N_17051,N_11358,N_8868);
and U17052 (N_17052,N_9403,N_9874);
nor U17053 (N_17053,N_9745,N_10771);
or U17054 (N_17054,N_11986,N_12460);
or U17055 (N_17055,N_10472,N_7416);
nor U17056 (N_17056,N_9564,N_7591);
nand U17057 (N_17057,N_7390,N_10314);
nand U17058 (N_17058,N_8179,N_7271);
and U17059 (N_17059,N_8068,N_7309);
nor U17060 (N_17060,N_11523,N_7944);
nand U17061 (N_17061,N_9914,N_10156);
or U17062 (N_17062,N_9579,N_7130);
or U17063 (N_17063,N_12421,N_7751);
or U17064 (N_17064,N_7450,N_11249);
nand U17065 (N_17065,N_7719,N_11640);
nand U17066 (N_17066,N_12320,N_12149);
nand U17067 (N_17067,N_11298,N_9140);
or U17068 (N_17068,N_8756,N_8376);
nor U17069 (N_17069,N_8253,N_9715);
nor U17070 (N_17070,N_12313,N_8952);
nand U17071 (N_17071,N_9085,N_7600);
and U17072 (N_17072,N_10456,N_10220);
nor U17073 (N_17073,N_7247,N_7860);
and U17074 (N_17074,N_12031,N_10226);
or U17075 (N_17075,N_12442,N_9931);
nand U17076 (N_17076,N_6547,N_8941);
and U17077 (N_17077,N_11287,N_12131);
nand U17078 (N_17078,N_11422,N_7795);
nand U17079 (N_17079,N_7782,N_7674);
and U17080 (N_17080,N_11483,N_7268);
and U17081 (N_17081,N_11224,N_6464);
and U17082 (N_17082,N_7283,N_8463);
nand U17083 (N_17083,N_6943,N_6760);
nor U17084 (N_17084,N_11376,N_7077);
nor U17085 (N_17085,N_11409,N_10014);
or U17086 (N_17086,N_7929,N_8331);
nand U17087 (N_17087,N_8419,N_12389);
or U17088 (N_17088,N_10550,N_12436);
nand U17089 (N_17089,N_7632,N_7828);
nor U17090 (N_17090,N_11223,N_9250);
or U17091 (N_17091,N_7205,N_10719);
xnor U17092 (N_17092,N_7312,N_6392);
nand U17093 (N_17093,N_12399,N_11734);
nor U17094 (N_17094,N_10383,N_8732);
and U17095 (N_17095,N_11463,N_10887);
or U17096 (N_17096,N_10736,N_6560);
or U17097 (N_17097,N_9819,N_7989);
nor U17098 (N_17098,N_11061,N_11039);
or U17099 (N_17099,N_9153,N_12241);
and U17100 (N_17100,N_8957,N_7088);
nand U17101 (N_17101,N_11882,N_9699);
or U17102 (N_17102,N_6547,N_7554);
or U17103 (N_17103,N_11347,N_7196);
or U17104 (N_17104,N_10397,N_8796);
or U17105 (N_17105,N_10069,N_11366);
nand U17106 (N_17106,N_11978,N_9389);
and U17107 (N_17107,N_6375,N_9614);
nor U17108 (N_17108,N_10683,N_9170);
or U17109 (N_17109,N_10953,N_6519);
nor U17110 (N_17110,N_8570,N_8670);
xor U17111 (N_17111,N_10527,N_10199);
nor U17112 (N_17112,N_10468,N_6478);
nor U17113 (N_17113,N_6427,N_11949);
nor U17114 (N_17114,N_9458,N_10308);
nor U17115 (N_17115,N_8691,N_10552);
nand U17116 (N_17116,N_6756,N_11964);
nor U17117 (N_17117,N_10627,N_8968);
and U17118 (N_17118,N_7063,N_12407);
nand U17119 (N_17119,N_11770,N_12445);
and U17120 (N_17120,N_8455,N_10260);
or U17121 (N_17121,N_12442,N_8660);
or U17122 (N_17122,N_7835,N_7491);
and U17123 (N_17123,N_11437,N_9492);
and U17124 (N_17124,N_11380,N_10328);
nand U17125 (N_17125,N_7286,N_12314);
xnor U17126 (N_17126,N_9455,N_7469);
or U17127 (N_17127,N_8904,N_7751);
and U17128 (N_17128,N_6749,N_6588);
and U17129 (N_17129,N_10953,N_7865);
and U17130 (N_17130,N_9186,N_11879);
and U17131 (N_17131,N_10104,N_6613);
and U17132 (N_17132,N_6611,N_6975);
and U17133 (N_17133,N_8290,N_7384);
nand U17134 (N_17134,N_11041,N_11072);
and U17135 (N_17135,N_10508,N_7208);
or U17136 (N_17136,N_6952,N_9424);
nand U17137 (N_17137,N_7026,N_11763);
nor U17138 (N_17138,N_11412,N_8098);
and U17139 (N_17139,N_7947,N_11584);
or U17140 (N_17140,N_9924,N_10875);
nand U17141 (N_17141,N_7991,N_7800);
nand U17142 (N_17142,N_10950,N_7693);
xnor U17143 (N_17143,N_9799,N_8649);
nor U17144 (N_17144,N_10479,N_10865);
and U17145 (N_17145,N_11754,N_11369);
or U17146 (N_17146,N_9195,N_8720);
xnor U17147 (N_17147,N_9387,N_9984);
nor U17148 (N_17148,N_9067,N_6879);
xor U17149 (N_17149,N_9862,N_10362);
or U17150 (N_17150,N_8160,N_9178);
nor U17151 (N_17151,N_8147,N_9276);
nand U17152 (N_17152,N_11684,N_11725);
and U17153 (N_17153,N_8301,N_10978);
or U17154 (N_17154,N_8021,N_10137);
nand U17155 (N_17155,N_10912,N_7882);
nor U17156 (N_17156,N_11709,N_8410);
or U17157 (N_17157,N_8020,N_9784);
nand U17158 (N_17158,N_12000,N_7620);
and U17159 (N_17159,N_10155,N_8641);
nand U17160 (N_17160,N_6733,N_7316);
or U17161 (N_17161,N_6687,N_8092);
and U17162 (N_17162,N_10689,N_12246);
or U17163 (N_17163,N_9562,N_9960);
nor U17164 (N_17164,N_10561,N_11171);
or U17165 (N_17165,N_6557,N_9891);
and U17166 (N_17166,N_6510,N_12125);
or U17167 (N_17167,N_7603,N_6799);
or U17168 (N_17168,N_8442,N_11775);
nor U17169 (N_17169,N_11977,N_6599);
nor U17170 (N_17170,N_8298,N_6444);
nor U17171 (N_17171,N_10525,N_12470);
and U17172 (N_17172,N_11714,N_9277);
or U17173 (N_17173,N_11052,N_9434);
and U17174 (N_17174,N_11225,N_10616);
nor U17175 (N_17175,N_10038,N_10362);
nor U17176 (N_17176,N_11881,N_8367);
and U17177 (N_17177,N_9207,N_6946);
and U17178 (N_17178,N_12238,N_9039);
nor U17179 (N_17179,N_9855,N_11602);
nor U17180 (N_17180,N_10488,N_10305);
nand U17181 (N_17181,N_10148,N_7273);
or U17182 (N_17182,N_10988,N_7976);
nor U17183 (N_17183,N_8801,N_7817);
nand U17184 (N_17184,N_9907,N_7603);
nor U17185 (N_17185,N_10218,N_6497);
nand U17186 (N_17186,N_8261,N_6961);
nand U17187 (N_17187,N_8145,N_8068);
and U17188 (N_17188,N_8042,N_12092);
and U17189 (N_17189,N_7714,N_11312);
xnor U17190 (N_17190,N_8397,N_9361);
nor U17191 (N_17191,N_10981,N_11225);
or U17192 (N_17192,N_8599,N_7173);
and U17193 (N_17193,N_8184,N_8984);
xor U17194 (N_17194,N_7401,N_8355);
nor U17195 (N_17195,N_10574,N_9881);
or U17196 (N_17196,N_6438,N_11506);
nand U17197 (N_17197,N_10954,N_10961);
and U17198 (N_17198,N_9350,N_10152);
and U17199 (N_17199,N_8287,N_7375);
and U17200 (N_17200,N_6891,N_10625);
nor U17201 (N_17201,N_8214,N_10199);
nor U17202 (N_17202,N_11117,N_7053);
nand U17203 (N_17203,N_7801,N_7254);
nor U17204 (N_17204,N_11758,N_10287);
nand U17205 (N_17205,N_8637,N_6430);
and U17206 (N_17206,N_9799,N_6542);
nor U17207 (N_17207,N_11816,N_12188);
and U17208 (N_17208,N_8036,N_8429);
or U17209 (N_17209,N_9819,N_8274);
nor U17210 (N_17210,N_7878,N_12016);
and U17211 (N_17211,N_9962,N_6990);
and U17212 (N_17212,N_7088,N_10898);
nor U17213 (N_17213,N_10448,N_9698);
nor U17214 (N_17214,N_7413,N_7726);
nand U17215 (N_17215,N_7389,N_7362);
nand U17216 (N_17216,N_11384,N_6851);
nand U17217 (N_17217,N_9571,N_10237);
nor U17218 (N_17218,N_10401,N_9895);
or U17219 (N_17219,N_8284,N_9544);
or U17220 (N_17220,N_9733,N_8709);
nand U17221 (N_17221,N_11432,N_11168);
or U17222 (N_17222,N_6362,N_8300);
and U17223 (N_17223,N_9263,N_12066);
xnor U17224 (N_17224,N_12165,N_8698);
and U17225 (N_17225,N_7339,N_10298);
and U17226 (N_17226,N_12286,N_7136);
nand U17227 (N_17227,N_8747,N_8975);
and U17228 (N_17228,N_11424,N_7415);
nand U17229 (N_17229,N_7790,N_7805);
and U17230 (N_17230,N_10607,N_9156);
nand U17231 (N_17231,N_12339,N_8990);
and U17232 (N_17232,N_8417,N_7495);
and U17233 (N_17233,N_10082,N_6625);
or U17234 (N_17234,N_8797,N_7221);
nand U17235 (N_17235,N_6989,N_7109);
or U17236 (N_17236,N_12405,N_6771);
nand U17237 (N_17237,N_12374,N_8641);
nor U17238 (N_17238,N_7254,N_6624);
or U17239 (N_17239,N_11648,N_11307);
and U17240 (N_17240,N_8167,N_10040);
nand U17241 (N_17241,N_6629,N_7946);
or U17242 (N_17242,N_12205,N_8109);
and U17243 (N_17243,N_10838,N_8989);
nand U17244 (N_17244,N_10440,N_7154);
xnor U17245 (N_17245,N_8749,N_10402);
nor U17246 (N_17246,N_7262,N_11711);
or U17247 (N_17247,N_6387,N_10333);
or U17248 (N_17248,N_12326,N_9195);
nor U17249 (N_17249,N_6648,N_7549);
and U17250 (N_17250,N_7269,N_9684);
nor U17251 (N_17251,N_9515,N_7306);
nor U17252 (N_17252,N_7633,N_12451);
or U17253 (N_17253,N_10994,N_6685);
and U17254 (N_17254,N_12146,N_11048);
or U17255 (N_17255,N_8500,N_7709);
nand U17256 (N_17256,N_8831,N_9249);
or U17257 (N_17257,N_10739,N_10351);
or U17258 (N_17258,N_10604,N_11964);
and U17259 (N_17259,N_12034,N_12433);
nand U17260 (N_17260,N_11489,N_9862);
and U17261 (N_17261,N_8245,N_12270);
nor U17262 (N_17262,N_12172,N_7065);
nand U17263 (N_17263,N_10750,N_10905);
nor U17264 (N_17264,N_8217,N_12059);
nand U17265 (N_17265,N_7527,N_8694);
and U17266 (N_17266,N_10472,N_11439);
and U17267 (N_17267,N_10359,N_8816);
nand U17268 (N_17268,N_11181,N_8109);
or U17269 (N_17269,N_6964,N_6852);
or U17270 (N_17270,N_10950,N_9520);
and U17271 (N_17271,N_10123,N_10039);
and U17272 (N_17272,N_7949,N_10931);
and U17273 (N_17273,N_9237,N_10611);
nor U17274 (N_17274,N_6454,N_8122);
and U17275 (N_17275,N_8911,N_10537);
or U17276 (N_17276,N_6380,N_7465);
nand U17277 (N_17277,N_9258,N_10489);
nor U17278 (N_17278,N_7866,N_9131);
and U17279 (N_17279,N_7345,N_6822);
xnor U17280 (N_17280,N_6914,N_7044);
and U17281 (N_17281,N_10975,N_8339);
and U17282 (N_17282,N_10222,N_12079);
nor U17283 (N_17283,N_8466,N_8146);
nand U17284 (N_17284,N_11226,N_8623);
and U17285 (N_17285,N_11119,N_8243);
nand U17286 (N_17286,N_8704,N_11986);
nand U17287 (N_17287,N_7757,N_6459);
or U17288 (N_17288,N_12048,N_12200);
and U17289 (N_17289,N_9832,N_10860);
nor U17290 (N_17290,N_10564,N_7029);
and U17291 (N_17291,N_12022,N_9517);
xnor U17292 (N_17292,N_10188,N_10116);
nor U17293 (N_17293,N_8165,N_9527);
nor U17294 (N_17294,N_9299,N_9237);
nor U17295 (N_17295,N_11985,N_7849);
and U17296 (N_17296,N_7280,N_7296);
nand U17297 (N_17297,N_12055,N_11874);
xor U17298 (N_17298,N_6929,N_7419);
and U17299 (N_17299,N_8990,N_8522);
nor U17300 (N_17300,N_6492,N_8972);
and U17301 (N_17301,N_6418,N_8420);
nor U17302 (N_17302,N_6832,N_9678);
and U17303 (N_17303,N_10618,N_11259);
or U17304 (N_17304,N_6980,N_8263);
and U17305 (N_17305,N_8305,N_10260);
or U17306 (N_17306,N_8789,N_7106);
nand U17307 (N_17307,N_10727,N_11686);
and U17308 (N_17308,N_7512,N_9972);
nor U17309 (N_17309,N_7031,N_12329);
nor U17310 (N_17310,N_9672,N_11970);
and U17311 (N_17311,N_6737,N_9732);
nor U17312 (N_17312,N_7742,N_11452);
nand U17313 (N_17313,N_8862,N_7234);
and U17314 (N_17314,N_9877,N_10798);
xor U17315 (N_17315,N_8083,N_12374);
xnor U17316 (N_17316,N_8607,N_8975);
nor U17317 (N_17317,N_10657,N_8745);
nor U17318 (N_17318,N_9664,N_7475);
and U17319 (N_17319,N_9413,N_6717);
xnor U17320 (N_17320,N_8864,N_8563);
nand U17321 (N_17321,N_11533,N_11674);
nor U17322 (N_17322,N_8710,N_8668);
nand U17323 (N_17323,N_11140,N_8273);
and U17324 (N_17324,N_6255,N_8867);
nand U17325 (N_17325,N_6426,N_8120);
or U17326 (N_17326,N_7525,N_10285);
nor U17327 (N_17327,N_6458,N_7265);
or U17328 (N_17328,N_6986,N_6469);
and U17329 (N_17329,N_9640,N_11432);
or U17330 (N_17330,N_6524,N_7665);
nor U17331 (N_17331,N_6943,N_8979);
nor U17332 (N_17332,N_11419,N_11947);
and U17333 (N_17333,N_10150,N_10750);
or U17334 (N_17334,N_6413,N_8018);
and U17335 (N_17335,N_10544,N_8313);
or U17336 (N_17336,N_12282,N_6714);
and U17337 (N_17337,N_11072,N_11256);
nor U17338 (N_17338,N_9225,N_11100);
nand U17339 (N_17339,N_7504,N_11564);
nor U17340 (N_17340,N_9740,N_10700);
and U17341 (N_17341,N_8646,N_9654);
and U17342 (N_17342,N_10786,N_12120);
nand U17343 (N_17343,N_10521,N_9378);
nand U17344 (N_17344,N_7661,N_10199);
and U17345 (N_17345,N_7225,N_9888);
nor U17346 (N_17346,N_10638,N_6261);
nor U17347 (N_17347,N_11816,N_10076);
nor U17348 (N_17348,N_8300,N_10266);
xnor U17349 (N_17349,N_11633,N_9328);
or U17350 (N_17350,N_10479,N_8331);
nor U17351 (N_17351,N_11437,N_7183);
nand U17352 (N_17352,N_8566,N_8446);
or U17353 (N_17353,N_8288,N_8313);
or U17354 (N_17354,N_7082,N_7626);
and U17355 (N_17355,N_9287,N_7167);
and U17356 (N_17356,N_12258,N_7448);
or U17357 (N_17357,N_8508,N_7079);
and U17358 (N_17358,N_8350,N_8798);
xnor U17359 (N_17359,N_10488,N_8328);
nand U17360 (N_17360,N_11798,N_9974);
nor U17361 (N_17361,N_8775,N_8691);
or U17362 (N_17362,N_9406,N_7670);
xnor U17363 (N_17363,N_10924,N_7861);
or U17364 (N_17364,N_12252,N_12072);
or U17365 (N_17365,N_12352,N_10614);
or U17366 (N_17366,N_10432,N_8852);
nor U17367 (N_17367,N_11998,N_7578);
nor U17368 (N_17368,N_12418,N_7426);
nor U17369 (N_17369,N_11069,N_7889);
nand U17370 (N_17370,N_10667,N_11984);
and U17371 (N_17371,N_8578,N_11479);
or U17372 (N_17372,N_12464,N_6507);
or U17373 (N_17373,N_8219,N_10329);
or U17374 (N_17374,N_6268,N_7061);
nand U17375 (N_17375,N_10036,N_7470);
nor U17376 (N_17376,N_7247,N_10098);
nand U17377 (N_17377,N_10759,N_6480);
nand U17378 (N_17378,N_7939,N_8512);
or U17379 (N_17379,N_11363,N_8604);
and U17380 (N_17380,N_6512,N_10014);
or U17381 (N_17381,N_10823,N_7337);
or U17382 (N_17382,N_9543,N_9859);
or U17383 (N_17383,N_7425,N_6980);
or U17384 (N_17384,N_9018,N_8492);
nor U17385 (N_17385,N_7916,N_10679);
and U17386 (N_17386,N_9149,N_11748);
or U17387 (N_17387,N_11770,N_7667);
and U17388 (N_17388,N_6445,N_10579);
nand U17389 (N_17389,N_12485,N_11748);
or U17390 (N_17390,N_11116,N_10133);
xnor U17391 (N_17391,N_6993,N_8508);
or U17392 (N_17392,N_8902,N_11444);
nor U17393 (N_17393,N_11361,N_7152);
xnor U17394 (N_17394,N_8323,N_7274);
and U17395 (N_17395,N_9629,N_6260);
and U17396 (N_17396,N_10199,N_8948);
nor U17397 (N_17397,N_7618,N_10918);
nand U17398 (N_17398,N_7746,N_11222);
nand U17399 (N_17399,N_9183,N_8312);
and U17400 (N_17400,N_9422,N_7726);
xor U17401 (N_17401,N_11702,N_10443);
nand U17402 (N_17402,N_7981,N_10657);
xor U17403 (N_17403,N_6316,N_6320);
xor U17404 (N_17404,N_6297,N_12163);
nand U17405 (N_17405,N_9664,N_8199);
nor U17406 (N_17406,N_11542,N_9781);
nand U17407 (N_17407,N_9209,N_7277);
and U17408 (N_17408,N_10040,N_9042);
nor U17409 (N_17409,N_10208,N_6953);
or U17410 (N_17410,N_8249,N_8868);
nand U17411 (N_17411,N_7100,N_7413);
nor U17412 (N_17412,N_11635,N_10129);
or U17413 (N_17413,N_9361,N_10996);
xor U17414 (N_17414,N_8374,N_11552);
xor U17415 (N_17415,N_11896,N_6526);
nand U17416 (N_17416,N_9630,N_10480);
nor U17417 (N_17417,N_8947,N_11001);
xor U17418 (N_17418,N_9160,N_6727);
nor U17419 (N_17419,N_9749,N_10215);
and U17420 (N_17420,N_7644,N_8282);
and U17421 (N_17421,N_12089,N_6637);
or U17422 (N_17422,N_10564,N_8119);
or U17423 (N_17423,N_9264,N_6363);
or U17424 (N_17424,N_9072,N_10544);
nand U17425 (N_17425,N_11054,N_12124);
or U17426 (N_17426,N_10336,N_9678);
and U17427 (N_17427,N_10818,N_7170);
nor U17428 (N_17428,N_6855,N_7967);
or U17429 (N_17429,N_8314,N_10711);
nor U17430 (N_17430,N_10725,N_9072);
and U17431 (N_17431,N_7775,N_8845);
nand U17432 (N_17432,N_8101,N_9833);
nor U17433 (N_17433,N_10879,N_9761);
and U17434 (N_17434,N_11253,N_6301);
nand U17435 (N_17435,N_10246,N_11801);
nor U17436 (N_17436,N_6801,N_6638);
xor U17437 (N_17437,N_9410,N_6965);
nand U17438 (N_17438,N_9238,N_8150);
or U17439 (N_17439,N_9446,N_10890);
nand U17440 (N_17440,N_10334,N_9847);
nand U17441 (N_17441,N_7421,N_9106);
nor U17442 (N_17442,N_8698,N_10933);
nor U17443 (N_17443,N_7211,N_11554);
or U17444 (N_17444,N_10333,N_9178);
nor U17445 (N_17445,N_11680,N_9354);
nor U17446 (N_17446,N_8998,N_11543);
or U17447 (N_17447,N_6470,N_10979);
nand U17448 (N_17448,N_9507,N_11536);
nor U17449 (N_17449,N_7285,N_9582);
or U17450 (N_17450,N_6327,N_12113);
nor U17451 (N_17451,N_12252,N_11609);
nand U17452 (N_17452,N_8551,N_6533);
nand U17453 (N_17453,N_8926,N_7258);
nor U17454 (N_17454,N_12262,N_11114);
nor U17455 (N_17455,N_8269,N_12415);
nor U17456 (N_17456,N_10451,N_12315);
nor U17457 (N_17457,N_11093,N_9921);
nor U17458 (N_17458,N_12212,N_9438);
and U17459 (N_17459,N_9930,N_9620);
nand U17460 (N_17460,N_8288,N_6417);
and U17461 (N_17461,N_8024,N_9105);
nor U17462 (N_17462,N_9480,N_11368);
and U17463 (N_17463,N_9084,N_7596);
nor U17464 (N_17464,N_8228,N_7724);
nor U17465 (N_17465,N_9462,N_6719);
nor U17466 (N_17466,N_7621,N_8000);
or U17467 (N_17467,N_6738,N_11034);
and U17468 (N_17468,N_11738,N_8361);
or U17469 (N_17469,N_10652,N_9565);
xor U17470 (N_17470,N_10515,N_7051);
xnor U17471 (N_17471,N_11402,N_8522);
nor U17472 (N_17472,N_6503,N_12299);
or U17473 (N_17473,N_8778,N_6516);
or U17474 (N_17474,N_8466,N_10667);
nand U17475 (N_17475,N_10540,N_6835);
nor U17476 (N_17476,N_11086,N_8725);
nand U17477 (N_17477,N_9560,N_11707);
or U17478 (N_17478,N_6601,N_7371);
or U17479 (N_17479,N_7812,N_11780);
or U17480 (N_17480,N_9268,N_11609);
nand U17481 (N_17481,N_11731,N_11100);
or U17482 (N_17482,N_7322,N_11172);
and U17483 (N_17483,N_11467,N_8206);
nor U17484 (N_17484,N_7881,N_7826);
xor U17485 (N_17485,N_11616,N_7577);
or U17486 (N_17486,N_11035,N_8089);
xnor U17487 (N_17487,N_9507,N_8081);
nor U17488 (N_17488,N_8226,N_10434);
nor U17489 (N_17489,N_7208,N_8275);
xor U17490 (N_17490,N_9564,N_11270);
nor U17491 (N_17491,N_6351,N_10699);
and U17492 (N_17492,N_6418,N_6475);
and U17493 (N_17493,N_11062,N_7150);
or U17494 (N_17494,N_12274,N_7472);
and U17495 (N_17495,N_7826,N_7705);
and U17496 (N_17496,N_8082,N_7620);
nand U17497 (N_17497,N_7642,N_11571);
and U17498 (N_17498,N_6669,N_8840);
nor U17499 (N_17499,N_10599,N_6440);
or U17500 (N_17500,N_10484,N_10268);
xnor U17501 (N_17501,N_6872,N_10218);
or U17502 (N_17502,N_7886,N_8139);
nand U17503 (N_17503,N_8536,N_9915);
nor U17504 (N_17504,N_7223,N_12475);
xnor U17505 (N_17505,N_7619,N_6687);
nand U17506 (N_17506,N_12011,N_10279);
and U17507 (N_17507,N_10274,N_10731);
and U17508 (N_17508,N_11213,N_7752);
and U17509 (N_17509,N_6580,N_9602);
nor U17510 (N_17510,N_11261,N_7528);
or U17511 (N_17511,N_6977,N_11064);
nor U17512 (N_17512,N_11708,N_6286);
nor U17513 (N_17513,N_8543,N_6292);
nand U17514 (N_17514,N_9193,N_9512);
xnor U17515 (N_17515,N_10368,N_9660);
nand U17516 (N_17516,N_10040,N_8911);
nand U17517 (N_17517,N_6994,N_9048);
nor U17518 (N_17518,N_7601,N_11761);
or U17519 (N_17519,N_8588,N_10812);
and U17520 (N_17520,N_11629,N_9600);
nand U17521 (N_17521,N_10971,N_8366);
and U17522 (N_17522,N_9956,N_10775);
nor U17523 (N_17523,N_11534,N_10131);
and U17524 (N_17524,N_8767,N_8378);
or U17525 (N_17525,N_8751,N_8155);
and U17526 (N_17526,N_9879,N_9696);
nor U17527 (N_17527,N_9441,N_11386);
nand U17528 (N_17528,N_6492,N_6530);
or U17529 (N_17529,N_11654,N_11074);
and U17530 (N_17530,N_8319,N_7056);
xnor U17531 (N_17531,N_6293,N_11924);
and U17532 (N_17532,N_7674,N_9491);
nand U17533 (N_17533,N_6376,N_11732);
nor U17534 (N_17534,N_11792,N_6547);
or U17535 (N_17535,N_9031,N_9552);
nand U17536 (N_17536,N_8874,N_8817);
nor U17537 (N_17537,N_11301,N_9165);
and U17538 (N_17538,N_8412,N_7643);
xnor U17539 (N_17539,N_7067,N_7095);
nand U17540 (N_17540,N_11967,N_8574);
nor U17541 (N_17541,N_6978,N_8716);
nor U17542 (N_17542,N_6366,N_10067);
and U17543 (N_17543,N_12337,N_11722);
or U17544 (N_17544,N_11275,N_10399);
nor U17545 (N_17545,N_6753,N_9764);
nor U17546 (N_17546,N_9183,N_8197);
nand U17547 (N_17547,N_8099,N_9124);
or U17548 (N_17548,N_7407,N_12359);
nand U17549 (N_17549,N_11358,N_11475);
and U17550 (N_17550,N_11793,N_6787);
and U17551 (N_17551,N_11270,N_11225);
nor U17552 (N_17552,N_8686,N_7502);
nand U17553 (N_17553,N_11332,N_7325);
and U17554 (N_17554,N_8278,N_10554);
and U17555 (N_17555,N_11880,N_10058);
and U17556 (N_17556,N_9196,N_11671);
nand U17557 (N_17557,N_11853,N_11730);
xor U17558 (N_17558,N_11388,N_12498);
nand U17559 (N_17559,N_10057,N_7831);
and U17560 (N_17560,N_11443,N_10800);
nor U17561 (N_17561,N_9396,N_8111);
nand U17562 (N_17562,N_8703,N_11889);
nor U17563 (N_17563,N_8368,N_9563);
xnor U17564 (N_17564,N_12329,N_7654);
nor U17565 (N_17565,N_9416,N_6988);
or U17566 (N_17566,N_6551,N_11080);
nand U17567 (N_17567,N_8743,N_12415);
xor U17568 (N_17568,N_7349,N_6421);
or U17569 (N_17569,N_7302,N_6876);
and U17570 (N_17570,N_10343,N_11052);
or U17571 (N_17571,N_7770,N_9327);
nor U17572 (N_17572,N_8863,N_7802);
or U17573 (N_17573,N_7269,N_6733);
nor U17574 (N_17574,N_7087,N_12422);
nand U17575 (N_17575,N_10107,N_12067);
or U17576 (N_17576,N_6658,N_9132);
and U17577 (N_17577,N_9439,N_7409);
nand U17578 (N_17578,N_10707,N_8880);
nand U17579 (N_17579,N_11599,N_10309);
nor U17580 (N_17580,N_10008,N_7139);
or U17581 (N_17581,N_10570,N_8238);
nor U17582 (N_17582,N_10798,N_6616);
or U17583 (N_17583,N_11965,N_10206);
or U17584 (N_17584,N_9712,N_9189);
or U17585 (N_17585,N_9792,N_8328);
and U17586 (N_17586,N_11856,N_8106);
nand U17587 (N_17587,N_11890,N_9837);
xnor U17588 (N_17588,N_12349,N_10720);
and U17589 (N_17589,N_10503,N_6661);
and U17590 (N_17590,N_7921,N_10750);
nand U17591 (N_17591,N_9674,N_7869);
nor U17592 (N_17592,N_11653,N_7816);
and U17593 (N_17593,N_11420,N_10304);
nand U17594 (N_17594,N_10986,N_7026);
nor U17595 (N_17595,N_11292,N_10526);
xor U17596 (N_17596,N_10780,N_6620);
and U17597 (N_17597,N_6901,N_9021);
xnor U17598 (N_17598,N_7705,N_9978);
nor U17599 (N_17599,N_6646,N_11900);
nand U17600 (N_17600,N_9733,N_10433);
nand U17601 (N_17601,N_12152,N_11338);
or U17602 (N_17602,N_8333,N_6722);
or U17603 (N_17603,N_11683,N_11455);
or U17604 (N_17604,N_8090,N_8642);
nand U17605 (N_17605,N_8329,N_9292);
nand U17606 (N_17606,N_10725,N_11809);
and U17607 (N_17607,N_10894,N_7682);
nand U17608 (N_17608,N_10827,N_7867);
or U17609 (N_17609,N_8770,N_12328);
and U17610 (N_17610,N_8950,N_7950);
and U17611 (N_17611,N_11854,N_11990);
xnor U17612 (N_17612,N_8650,N_11431);
nor U17613 (N_17613,N_9585,N_7402);
nor U17614 (N_17614,N_6625,N_12085);
or U17615 (N_17615,N_7651,N_11091);
and U17616 (N_17616,N_11458,N_12115);
xor U17617 (N_17617,N_9017,N_8214);
and U17618 (N_17618,N_10656,N_8936);
nor U17619 (N_17619,N_6265,N_6349);
xor U17620 (N_17620,N_9984,N_7190);
xnor U17621 (N_17621,N_7448,N_9275);
or U17622 (N_17622,N_11893,N_6952);
or U17623 (N_17623,N_6649,N_8592);
or U17624 (N_17624,N_9865,N_6542);
xor U17625 (N_17625,N_8753,N_11995);
and U17626 (N_17626,N_11257,N_10705);
nor U17627 (N_17627,N_12416,N_11518);
and U17628 (N_17628,N_7075,N_10338);
and U17629 (N_17629,N_12022,N_8787);
or U17630 (N_17630,N_10226,N_7840);
or U17631 (N_17631,N_10841,N_7372);
xnor U17632 (N_17632,N_11308,N_6445);
nor U17633 (N_17633,N_9868,N_8732);
nand U17634 (N_17634,N_10017,N_12204);
nor U17635 (N_17635,N_9244,N_9009);
nor U17636 (N_17636,N_10819,N_7139);
nand U17637 (N_17637,N_11369,N_8971);
nand U17638 (N_17638,N_12127,N_8902);
nand U17639 (N_17639,N_12490,N_6291);
nand U17640 (N_17640,N_8875,N_10940);
or U17641 (N_17641,N_10405,N_12102);
nor U17642 (N_17642,N_9141,N_8802);
and U17643 (N_17643,N_10260,N_7039);
nor U17644 (N_17644,N_10171,N_10987);
nor U17645 (N_17645,N_8810,N_10560);
and U17646 (N_17646,N_9721,N_8146);
nand U17647 (N_17647,N_8929,N_8264);
nor U17648 (N_17648,N_11980,N_6490);
or U17649 (N_17649,N_12266,N_10007);
nor U17650 (N_17650,N_11958,N_7059);
and U17651 (N_17651,N_10278,N_10006);
nand U17652 (N_17652,N_7646,N_10409);
nor U17653 (N_17653,N_10772,N_11337);
nor U17654 (N_17654,N_10893,N_7449);
or U17655 (N_17655,N_12353,N_7073);
or U17656 (N_17656,N_8971,N_9377);
nor U17657 (N_17657,N_6281,N_11188);
nand U17658 (N_17658,N_8559,N_7420);
nor U17659 (N_17659,N_8544,N_12384);
or U17660 (N_17660,N_11878,N_8721);
and U17661 (N_17661,N_6760,N_12468);
and U17662 (N_17662,N_8425,N_9142);
or U17663 (N_17663,N_8011,N_7968);
xnor U17664 (N_17664,N_9899,N_11930);
nor U17665 (N_17665,N_10192,N_10644);
nor U17666 (N_17666,N_7074,N_6814);
and U17667 (N_17667,N_7652,N_8431);
nor U17668 (N_17668,N_8129,N_7389);
nor U17669 (N_17669,N_11878,N_10373);
or U17670 (N_17670,N_7409,N_9109);
nand U17671 (N_17671,N_6313,N_7919);
nand U17672 (N_17672,N_9215,N_11215);
or U17673 (N_17673,N_6315,N_6744);
and U17674 (N_17674,N_9842,N_6710);
and U17675 (N_17675,N_9038,N_7228);
and U17676 (N_17676,N_7578,N_6376);
and U17677 (N_17677,N_7099,N_9758);
or U17678 (N_17678,N_9194,N_7396);
and U17679 (N_17679,N_8478,N_7473);
nor U17680 (N_17680,N_6511,N_12101);
or U17681 (N_17681,N_7121,N_8982);
nand U17682 (N_17682,N_9810,N_11922);
nand U17683 (N_17683,N_6638,N_11116);
or U17684 (N_17684,N_6629,N_6828);
nor U17685 (N_17685,N_12483,N_11570);
nand U17686 (N_17686,N_8948,N_10959);
xor U17687 (N_17687,N_9684,N_7678);
and U17688 (N_17688,N_8323,N_12220);
or U17689 (N_17689,N_7984,N_8491);
nand U17690 (N_17690,N_9958,N_9989);
xor U17691 (N_17691,N_11974,N_10386);
nor U17692 (N_17692,N_8598,N_7844);
or U17693 (N_17693,N_8197,N_8416);
and U17694 (N_17694,N_8919,N_10445);
nor U17695 (N_17695,N_10316,N_6720);
and U17696 (N_17696,N_10892,N_10858);
or U17697 (N_17697,N_9338,N_11613);
and U17698 (N_17698,N_6985,N_10887);
nand U17699 (N_17699,N_6884,N_11636);
and U17700 (N_17700,N_12352,N_10183);
nand U17701 (N_17701,N_11202,N_7938);
or U17702 (N_17702,N_6652,N_8910);
nor U17703 (N_17703,N_9281,N_6511);
nand U17704 (N_17704,N_11196,N_10001);
or U17705 (N_17705,N_10999,N_10284);
nand U17706 (N_17706,N_10603,N_10375);
nor U17707 (N_17707,N_11792,N_12387);
nand U17708 (N_17708,N_8708,N_12468);
or U17709 (N_17709,N_8013,N_7470);
or U17710 (N_17710,N_9293,N_10941);
nor U17711 (N_17711,N_11547,N_7860);
or U17712 (N_17712,N_12339,N_9087);
nor U17713 (N_17713,N_6557,N_8814);
and U17714 (N_17714,N_9281,N_8023);
nand U17715 (N_17715,N_11296,N_6251);
or U17716 (N_17716,N_9424,N_9471);
xor U17717 (N_17717,N_10846,N_8522);
nand U17718 (N_17718,N_6562,N_6261);
or U17719 (N_17719,N_7553,N_6357);
and U17720 (N_17720,N_6410,N_10364);
nand U17721 (N_17721,N_9539,N_6811);
and U17722 (N_17722,N_6989,N_9445);
nand U17723 (N_17723,N_11010,N_9667);
nand U17724 (N_17724,N_7396,N_11713);
or U17725 (N_17725,N_9473,N_7436);
or U17726 (N_17726,N_9599,N_7088);
nand U17727 (N_17727,N_11396,N_6895);
or U17728 (N_17728,N_9752,N_9618);
nand U17729 (N_17729,N_7473,N_9648);
and U17730 (N_17730,N_11694,N_7112);
nor U17731 (N_17731,N_10821,N_11835);
and U17732 (N_17732,N_11999,N_9219);
nand U17733 (N_17733,N_7145,N_11569);
or U17734 (N_17734,N_7378,N_7360);
nor U17735 (N_17735,N_9452,N_6461);
nor U17736 (N_17736,N_8928,N_8198);
nand U17737 (N_17737,N_8781,N_12438);
nor U17738 (N_17738,N_7647,N_11301);
nor U17739 (N_17739,N_7170,N_7784);
nor U17740 (N_17740,N_12477,N_9749);
nor U17741 (N_17741,N_6346,N_11497);
and U17742 (N_17742,N_12256,N_11841);
nor U17743 (N_17743,N_7877,N_7306);
nand U17744 (N_17744,N_8625,N_10894);
nor U17745 (N_17745,N_8353,N_10247);
nand U17746 (N_17746,N_12300,N_7868);
and U17747 (N_17747,N_11223,N_7036);
nor U17748 (N_17748,N_8258,N_9486);
nor U17749 (N_17749,N_9094,N_11820);
or U17750 (N_17750,N_8470,N_12036);
nor U17751 (N_17751,N_6591,N_10121);
nor U17752 (N_17752,N_12240,N_10622);
and U17753 (N_17753,N_9635,N_9540);
nand U17754 (N_17754,N_6821,N_10501);
and U17755 (N_17755,N_11290,N_7252);
or U17756 (N_17756,N_9682,N_11722);
or U17757 (N_17757,N_6962,N_7196);
xnor U17758 (N_17758,N_11559,N_8159);
nor U17759 (N_17759,N_9716,N_11903);
or U17760 (N_17760,N_10108,N_6445);
nor U17761 (N_17761,N_7525,N_8114);
or U17762 (N_17762,N_11061,N_8958);
nor U17763 (N_17763,N_7638,N_11689);
nand U17764 (N_17764,N_11475,N_7563);
and U17765 (N_17765,N_9266,N_8297);
and U17766 (N_17766,N_9488,N_11184);
and U17767 (N_17767,N_9826,N_10353);
or U17768 (N_17768,N_12269,N_7643);
nor U17769 (N_17769,N_11846,N_7500);
and U17770 (N_17770,N_7438,N_10101);
nor U17771 (N_17771,N_7136,N_8705);
nor U17772 (N_17772,N_7035,N_6826);
nand U17773 (N_17773,N_11798,N_6680);
nand U17774 (N_17774,N_11846,N_10939);
nand U17775 (N_17775,N_7891,N_10836);
nor U17776 (N_17776,N_11165,N_10107);
nor U17777 (N_17777,N_8217,N_9606);
and U17778 (N_17778,N_6740,N_9629);
or U17779 (N_17779,N_7506,N_8398);
nor U17780 (N_17780,N_9551,N_9733);
and U17781 (N_17781,N_11525,N_9380);
nand U17782 (N_17782,N_6708,N_11408);
xnor U17783 (N_17783,N_8859,N_9101);
or U17784 (N_17784,N_10944,N_11306);
xnor U17785 (N_17785,N_7676,N_7760);
xnor U17786 (N_17786,N_12050,N_12481);
and U17787 (N_17787,N_9513,N_11444);
nor U17788 (N_17788,N_12078,N_6725);
nor U17789 (N_17789,N_10085,N_12234);
and U17790 (N_17790,N_6596,N_10433);
or U17791 (N_17791,N_11920,N_9905);
or U17792 (N_17792,N_9627,N_10106);
nand U17793 (N_17793,N_11201,N_9157);
or U17794 (N_17794,N_8684,N_11966);
nor U17795 (N_17795,N_12263,N_7964);
or U17796 (N_17796,N_10039,N_10986);
nand U17797 (N_17797,N_9626,N_9569);
and U17798 (N_17798,N_10929,N_12265);
or U17799 (N_17799,N_9229,N_6779);
or U17800 (N_17800,N_8241,N_7781);
and U17801 (N_17801,N_8863,N_8292);
nor U17802 (N_17802,N_6638,N_8090);
nand U17803 (N_17803,N_9737,N_6256);
nand U17804 (N_17804,N_11773,N_9534);
xor U17805 (N_17805,N_10152,N_12342);
or U17806 (N_17806,N_7827,N_8320);
or U17807 (N_17807,N_8758,N_8491);
and U17808 (N_17808,N_10498,N_7259);
and U17809 (N_17809,N_10984,N_10674);
nand U17810 (N_17810,N_6864,N_10675);
and U17811 (N_17811,N_10558,N_8179);
nand U17812 (N_17812,N_8896,N_10225);
or U17813 (N_17813,N_11388,N_8034);
or U17814 (N_17814,N_6679,N_6730);
or U17815 (N_17815,N_11271,N_6708);
xnor U17816 (N_17816,N_8604,N_9888);
or U17817 (N_17817,N_12140,N_8211);
nand U17818 (N_17818,N_8755,N_12388);
or U17819 (N_17819,N_6306,N_10468);
nand U17820 (N_17820,N_8733,N_10989);
xnor U17821 (N_17821,N_10908,N_12036);
nand U17822 (N_17822,N_8829,N_7677);
nand U17823 (N_17823,N_10243,N_6737);
nand U17824 (N_17824,N_7205,N_11928);
and U17825 (N_17825,N_10588,N_10301);
nand U17826 (N_17826,N_10728,N_9201);
xnor U17827 (N_17827,N_12369,N_10095);
nand U17828 (N_17828,N_11723,N_7129);
nor U17829 (N_17829,N_10357,N_10813);
or U17830 (N_17830,N_9966,N_11160);
nor U17831 (N_17831,N_6718,N_10894);
xor U17832 (N_17832,N_8247,N_11383);
or U17833 (N_17833,N_9243,N_8289);
nand U17834 (N_17834,N_9122,N_7948);
and U17835 (N_17835,N_9340,N_11998);
or U17836 (N_17836,N_11556,N_7160);
and U17837 (N_17837,N_10500,N_10760);
or U17838 (N_17838,N_8355,N_9137);
or U17839 (N_17839,N_10089,N_7796);
nor U17840 (N_17840,N_9995,N_11419);
or U17841 (N_17841,N_9450,N_10998);
nand U17842 (N_17842,N_9809,N_8123);
nand U17843 (N_17843,N_10176,N_11868);
xor U17844 (N_17844,N_11882,N_7362);
or U17845 (N_17845,N_9090,N_8735);
and U17846 (N_17846,N_11772,N_11958);
and U17847 (N_17847,N_7496,N_10913);
nand U17848 (N_17848,N_12181,N_9516);
or U17849 (N_17849,N_7849,N_8802);
nor U17850 (N_17850,N_9367,N_8231);
nor U17851 (N_17851,N_11252,N_9250);
nor U17852 (N_17852,N_9779,N_7700);
nand U17853 (N_17853,N_11942,N_9334);
and U17854 (N_17854,N_10848,N_7699);
and U17855 (N_17855,N_10406,N_8371);
nand U17856 (N_17856,N_7013,N_12422);
or U17857 (N_17857,N_6995,N_7817);
or U17858 (N_17858,N_8264,N_8392);
nor U17859 (N_17859,N_6259,N_7208);
nor U17860 (N_17860,N_11637,N_11457);
and U17861 (N_17861,N_11904,N_11969);
nor U17862 (N_17862,N_8017,N_8516);
nor U17863 (N_17863,N_9418,N_10308);
nor U17864 (N_17864,N_9282,N_11489);
or U17865 (N_17865,N_8121,N_11785);
or U17866 (N_17866,N_6463,N_8688);
and U17867 (N_17867,N_7701,N_6698);
xor U17868 (N_17868,N_7709,N_7918);
or U17869 (N_17869,N_10548,N_9811);
nand U17870 (N_17870,N_10037,N_10273);
and U17871 (N_17871,N_9537,N_9572);
and U17872 (N_17872,N_10505,N_8925);
nor U17873 (N_17873,N_9324,N_7495);
or U17874 (N_17874,N_9765,N_10961);
nor U17875 (N_17875,N_11174,N_8984);
and U17876 (N_17876,N_7335,N_8761);
nor U17877 (N_17877,N_10229,N_8295);
and U17878 (N_17878,N_10341,N_8459);
or U17879 (N_17879,N_10515,N_11007);
nor U17880 (N_17880,N_9338,N_8707);
and U17881 (N_17881,N_9602,N_7516);
and U17882 (N_17882,N_10063,N_10654);
and U17883 (N_17883,N_8138,N_7078);
nand U17884 (N_17884,N_11225,N_10008);
and U17885 (N_17885,N_11632,N_9309);
or U17886 (N_17886,N_8125,N_7984);
nand U17887 (N_17887,N_11200,N_10637);
nand U17888 (N_17888,N_8868,N_9738);
and U17889 (N_17889,N_12332,N_11364);
nand U17890 (N_17890,N_8449,N_6528);
and U17891 (N_17891,N_11098,N_11930);
nor U17892 (N_17892,N_10396,N_12182);
nor U17893 (N_17893,N_11498,N_9894);
and U17894 (N_17894,N_10129,N_9678);
nor U17895 (N_17895,N_8200,N_9112);
nor U17896 (N_17896,N_10699,N_9563);
nor U17897 (N_17897,N_10769,N_11028);
xor U17898 (N_17898,N_7271,N_11864);
nand U17899 (N_17899,N_11411,N_10268);
nor U17900 (N_17900,N_6270,N_8431);
nand U17901 (N_17901,N_8849,N_10119);
or U17902 (N_17902,N_11965,N_12489);
nor U17903 (N_17903,N_10903,N_12177);
or U17904 (N_17904,N_11962,N_10946);
or U17905 (N_17905,N_10467,N_10540);
nand U17906 (N_17906,N_9080,N_6976);
xnor U17907 (N_17907,N_9300,N_9161);
and U17908 (N_17908,N_8632,N_10266);
nor U17909 (N_17909,N_12352,N_11994);
nand U17910 (N_17910,N_8288,N_10349);
nand U17911 (N_17911,N_11355,N_7555);
xnor U17912 (N_17912,N_8272,N_8831);
nand U17913 (N_17913,N_12439,N_7214);
nor U17914 (N_17914,N_10482,N_7703);
and U17915 (N_17915,N_6674,N_8520);
or U17916 (N_17916,N_10733,N_8449);
and U17917 (N_17917,N_8161,N_9990);
nand U17918 (N_17918,N_7912,N_7506);
nand U17919 (N_17919,N_6751,N_8570);
nand U17920 (N_17920,N_10855,N_8406);
nor U17921 (N_17921,N_7055,N_7145);
nor U17922 (N_17922,N_8984,N_6540);
and U17923 (N_17923,N_9379,N_7444);
or U17924 (N_17924,N_8216,N_9426);
nand U17925 (N_17925,N_8203,N_11437);
nor U17926 (N_17926,N_12047,N_11553);
nand U17927 (N_17927,N_8624,N_8235);
nor U17928 (N_17928,N_9607,N_9693);
or U17929 (N_17929,N_9098,N_8846);
nand U17930 (N_17930,N_10763,N_8292);
and U17931 (N_17931,N_12117,N_7602);
xor U17932 (N_17932,N_11872,N_10470);
or U17933 (N_17933,N_11309,N_10897);
or U17934 (N_17934,N_9572,N_9947);
nand U17935 (N_17935,N_11904,N_8354);
nor U17936 (N_17936,N_8622,N_10488);
nor U17937 (N_17937,N_11684,N_11617);
or U17938 (N_17938,N_11262,N_11314);
and U17939 (N_17939,N_12262,N_6965);
or U17940 (N_17940,N_11685,N_8910);
xor U17941 (N_17941,N_9903,N_10562);
or U17942 (N_17942,N_9388,N_8548);
xor U17943 (N_17943,N_11860,N_8809);
and U17944 (N_17944,N_10728,N_7373);
nand U17945 (N_17945,N_8779,N_8352);
and U17946 (N_17946,N_6722,N_8451);
or U17947 (N_17947,N_9847,N_6322);
nor U17948 (N_17948,N_8038,N_10503);
nor U17949 (N_17949,N_8149,N_11726);
nor U17950 (N_17950,N_7460,N_7291);
xor U17951 (N_17951,N_10491,N_10673);
and U17952 (N_17952,N_10153,N_9785);
or U17953 (N_17953,N_10979,N_11130);
or U17954 (N_17954,N_10852,N_9203);
nand U17955 (N_17955,N_10183,N_7434);
and U17956 (N_17956,N_7108,N_9624);
and U17957 (N_17957,N_6789,N_9741);
nand U17958 (N_17958,N_12345,N_12062);
and U17959 (N_17959,N_7812,N_8946);
xor U17960 (N_17960,N_6283,N_7012);
nor U17961 (N_17961,N_6789,N_8129);
and U17962 (N_17962,N_10716,N_9899);
nand U17963 (N_17963,N_9734,N_8278);
or U17964 (N_17964,N_9269,N_6505);
nand U17965 (N_17965,N_11503,N_10188);
nand U17966 (N_17966,N_7535,N_10214);
xnor U17967 (N_17967,N_9826,N_6916);
or U17968 (N_17968,N_6788,N_10510);
and U17969 (N_17969,N_9100,N_9306);
nand U17970 (N_17970,N_10394,N_11763);
and U17971 (N_17971,N_12219,N_7928);
nand U17972 (N_17972,N_7940,N_9374);
and U17973 (N_17973,N_8360,N_6568);
nor U17974 (N_17974,N_9814,N_8764);
or U17975 (N_17975,N_9089,N_12063);
or U17976 (N_17976,N_11758,N_12224);
nor U17977 (N_17977,N_9639,N_7912);
nand U17978 (N_17978,N_7890,N_8431);
nor U17979 (N_17979,N_6264,N_8448);
and U17980 (N_17980,N_6294,N_9714);
and U17981 (N_17981,N_12371,N_6287);
and U17982 (N_17982,N_10297,N_11157);
nor U17983 (N_17983,N_11550,N_7188);
nor U17984 (N_17984,N_8064,N_11614);
and U17985 (N_17985,N_7963,N_7395);
or U17986 (N_17986,N_11964,N_11302);
nor U17987 (N_17987,N_11517,N_8236);
nor U17988 (N_17988,N_10440,N_8109);
nor U17989 (N_17989,N_8280,N_9481);
or U17990 (N_17990,N_10587,N_10326);
xor U17991 (N_17991,N_8986,N_7170);
xnor U17992 (N_17992,N_8388,N_12454);
and U17993 (N_17993,N_10082,N_6297);
nor U17994 (N_17994,N_9770,N_9790);
and U17995 (N_17995,N_6420,N_12228);
nand U17996 (N_17996,N_9611,N_9097);
and U17997 (N_17997,N_11490,N_9710);
xnor U17998 (N_17998,N_10559,N_10543);
xnor U17999 (N_17999,N_10096,N_8261);
and U18000 (N_18000,N_11452,N_7826);
nand U18001 (N_18001,N_11363,N_6373);
and U18002 (N_18002,N_10207,N_12462);
nor U18003 (N_18003,N_8341,N_9169);
and U18004 (N_18004,N_9717,N_10517);
and U18005 (N_18005,N_12339,N_9045);
nand U18006 (N_18006,N_7472,N_9821);
nand U18007 (N_18007,N_7453,N_11274);
nor U18008 (N_18008,N_11805,N_10492);
nand U18009 (N_18009,N_7525,N_6472);
xor U18010 (N_18010,N_8501,N_6551);
nor U18011 (N_18011,N_7666,N_8502);
nor U18012 (N_18012,N_10215,N_11026);
and U18013 (N_18013,N_11932,N_10935);
and U18014 (N_18014,N_10232,N_6925);
or U18015 (N_18015,N_9095,N_10027);
and U18016 (N_18016,N_8308,N_12253);
or U18017 (N_18017,N_10858,N_10052);
xnor U18018 (N_18018,N_9509,N_7497);
xnor U18019 (N_18019,N_9452,N_10555);
nor U18020 (N_18020,N_9821,N_11254);
nor U18021 (N_18021,N_6870,N_8412);
or U18022 (N_18022,N_8738,N_8656);
or U18023 (N_18023,N_9607,N_10870);
nor U18024 (N_18024,N_7140,N_10590);
nand U18025 (N_18025,N_9454,N_7223);
and U18026 (N_18026,N_12299,N_7119);
xnor U18027 (N_18027,N_9468,N_8404);
or U18028 (N_18028,N_12178,N_11822);
xnor U18029 (N_18029,N_9035,N_7865);
or U18030 (N_18030,N_7950,N_11241);
or U18031 (N_18031,N_8365,N_8599);
or U18032 (N_18032,N_8956,N_8349);
xor U18033 (N_18033,N_10031,N_10640);
and U18034 (N_18034,N_7508,N_11552);
nor U18035 (N_18035,N_10337,N_7398);
nor U18036 (N_18036,N_7616,N_9458);
and U18037 (N_18037,N_12354,N_11017);
or U18038 (N_18038,N_8781,N_11441);
nand U18039 (N_18039,N_9865,N_7780);
nand U18040 (N_18040,N_9844,N_7315);
xor U18041 (N_18041,N_8076,N_9129);
nand U18042 (N_18042,N_10590,N_6764);
and U18043 (N_18043,N_12335,N_6726);
and U18044 (N_18044,N_10145,N_8934);
nor U18045 (N_18045,N_8771,N_11001);
or U18046 (N_18046,N_11129,N_7435);
nand U18047 (N_18047,N_6363,N_11655);
nand U18048 (N_18048,N_8096,N_11199);
nand U18049 (N_18049,N_7705,N_11572);
and U18050 (N_18050,N_7923,N_12304);
and U18051 (N_18051,N_9308,N_6912);
or U18052 (N_18052,N_9449,N_6966);
and U18053 (N_18053,N_8589,N_7724);
nor U18054 (N_18054,N_6703,N_8196);
nand U18055 (N_18055,N_11077,N_10735);
or U18056 (N_18056,N_8019,N_8277);
or U18057 (N_18057,N_9062,N_8341);
nor U18058 (N_18058,N_10622,N_10564);
xnor U18059 (N_18059,N_6585,N_8638);
and U18060 (N_18060,N_8177,N_9307);
nand U18061 (N_18061,N_9778,N_10745);
and U18062 (N_18062,N_9179,N_9653);
or U18063 (N_18063,N_6943,N_11842);
nand U18064 (N_18064,N_8156,N_8250);
and U18065 (N_18065,N_7837,N_11324);
nor U18066 (N_18066,N_10713,N_8899);
and U18067 (N_18067,N_10989,N_11821);
nand U18068 (N_18068,N_10638,N_12482);
nor U18069 (N_18069,N_11877,N_11198);
nor U18070 (N_18070,N_9507,N_6816);
xor U18071 (N_18071,N_9103,N_8495);
nand U18072 (N_18072,N_10353,N_6538);
or U18073 (N_18073,N_7409,N_6772);
nor U18074 (N_18074,N_7485,N_8979);
nand U18075 (N_18075,N_7641,N_9804);
nor U18076 (N_18076,N_6427,N_10985);
nand U18077 (N_18077,N_6330,N_9180);
and U18078 (N_18078,N_9191,N_8805);
nand U18079 (N_18079,N_7576,N_12344);
or U18080 (N_18080,N_11862,N_10254);
xnor U18081 (N_18081,N_9500,N_10770);
xnor U18082 (N_18082,N_7980,N_10397);
and U18083 (N_18083,N_6748,N_11685);
nor U18084 (N_18084,N_7192,N_12376);
and U18085 (N_18085,N_9711,N_9349);
or U18086 (N_18086,N_10381,N_8220);
and U18087 (N_18087,N_12041,N_8296);
or U18088 (N_18088,N_7891,N_9773);
and U18089 (N_18089,N_10225,N_6903);
nor U18090 (N_18090,N_11354,N_7703);
or U18091 (N_18091,N_12242,N_8666);
xor U18092 (N_18092,N_7774,N_6495);
and U18093 (N_18093,N_12155,N_9571);
nor U18094 (N_18094,N_7136,N_8248);
nand U18095 (N_18095,N_7801,N_8615);
nor U18096 (N_18096,N_9238,N_10164);
xor U18097 (N_18097,N_6802,N_8343);
xnor U18098 (N_18098,N_11713,N_6265);
and U18099 (N_18099,N_10686,N_9259);
nand U18100 (N_18100,N_10772,N_10144);
nand U18101 (N_18101,N_10912,N_9663);
or U18102 (N_18102,N_10857,N_10011);
nor U18103 (N_18103,N_8630,N_9203);
nand U18104 (N_18104,N_10013,N_6698);
or U18105 (N_18105,N_8507,N_10581);
nor U18106 (N_18106,N_12190,N_12111);
or U18107 (N_18107,N_10878,N_9665);
nor U18108 (N_18108,N_10493,N_7516);
and U18109 (N_18109,N_8368,N_10465);
and U18110 (N_18110,N_6766,N_11898);
nand U18111 (N_18111,N_12038,N_9630);
and U18112 (N_18112,N_12463,N_12462);
and U18113 (N_18113,N_9152,N_11554);
nand U18114 (N_18114,N_11166,N_8512);
or U18115 (N_18115,N_12265,N_7977);
nor U18116 (N_18116,N_7259,N_9147);
or U18117 (N_18117,N_7898,N_6446);
and U18118 (N_18118,N_12092,N_7809);
or U18119 (N_18119,N_8973,N_9651);
or U18120 (N_18120,N_7185,N_11384);
or U18121 (N_18121,N_10280,N_10596);
nand U18122 (N_18122,N_12228,N_10659);
or U18123 (N_18123,N_9045,N_8673);
nand U18124 (N_18124,N_7948,N_11892);
nor U18125 (N_18125,N_8662,N_6692);
nor U18126 (N_18126,N_11281,N_6610);
nand U18127 (N_18127,N_7385,N_7914);
and U18128 (N_18128,N_11929,N_9562);
or U18129 (N_18129,N_11260,N_12338);
or U18130 (N_18130,N_11576,N_11367);
xnor U18131 (N_18131,N_8362,N_9863);
nor U18132 (N_18132,N_10392,N_10163);
or U18133 (N_18133,N_9088,N_8554);
or U18134 (N_18134,N_8478,N_10793);
or U18135 (N_18135,N_11696,N_10164);
nor U18136 (N_18136,N_7914,N_9457);
nand U18137 (N_18137,N_8586,N_12010);
nor U18138 (N_18138,N_6280,N_9084);
nor U18139 (N_18139,N_6415,N_7615);
or U18140 (N_18140,N_11611,N_8794);
and U18141 (N_18141,N_8790,N_8990);
nor U18142 (N_18142,N_12079,N_6390);
nor U18143 (N_18143,N_11085,N_6394);
and U18144 (N_18144,N_9088,N_12491);
nand U18145 (N_18145,N_12369,N_8930);
and U18146 (N_18146,N_9805,N_9424);
and U18147 (N_18147,N_8243,N_11822);
or U18148 (N_18148,N_11871,N_11407);
or U18149 (N_18149,N_11805,N_7820);
nor U18150 (N_18150,N_7103,N_6882);
or U18151 (N_18151,N_11507,N_7819);
and U18152 (N_18152,N_6905,N_10064);
and U18153 (N_18153,N_10974,N_7905);
nand U18154 (N_18154,N_10308,N_8768);
and U18155 (N_18155,N_12007,N_10316);
and U18156 (N_18156,N_11326,N_9640);
nand U18157 (N_18157,N_9911,N_10525);
nor U18158 (N_18158,N_7009,N_10627);
nor U18159 (N_18159,N_10296,N_6698);
nand U18160 (N_18160,N_9394,N_8264);
nand U18161 (N_18161,N_9358,N_11456);
or U18162 (N_18162,N_7031,N_10137);
and U18163 (N_18163,N_8192,N_9182);
and U18164 (N_18164,N_6859,N_9963);
or U18165 (N_18165,N_6601,N_9132);
or U18166 (N_18166,N_10105,N_9880);
nor U18167 (N_18167,N_10237,N_8527);
or U18168 (N_18168,N_6411,N_7681);
nand U18169 (N_18169,N_6329,N_10327);
or U18170 (N_18170,N_11226,N_9484);
or U18171 (N_18171,N_8607,N_8540);
nand U18172 (N_18172,N_12414,N_11897);
nor U18173 (N_18173,N_8968,N_7691);
nand U18174 (N_18174,N_8612,N_9285);
nand U18175 (N_18175,N_12034,N_11054);
xor U18176 (N_18176,N_9480,N_8417);
or U18177 (N_18177,N_6719,N_12331);
or U18178 (N_18178,N_9741,N_10827);
xor U18179 (N_18179,N_9385,N_6599);
xnor U18180 (N_18180,N_11943,N_9772);
nor U18181 (N_18181,N_11515,N_7724);
nand U18182 (N_18182,N_8541,N_6861);
xor U18183 (N_18183,N_10638,N_9201);
nor U18184 (N_18184,N_7320,N_7140);
nor U18185 (N_18185,N_8841,N_6702);
and U18186 (N_18186,N_9926,N_9703);
or U18187 (N_18187,N_8445,N_11075);
or U18188 (N_18188,N_7603,N_11415);
nand U18189 (N_18189,N_6780,N_9574);
or U18190 (N_18190,N_7134,N_12277);
or U18191 (N_18191,N_10307,N_12403);
nand U18192 (N_18192,N_7815,N_8782);
and U18193 (N_18193,N_11453,N_8148);
nor U18194 (N_18194,N_11404,N_12269);
nor U18195 (N_18195,N_6622,N_7008);
and U18196 (N_18196,N_10579,N_7193);
and U18197 (N_18197,N_10350,N_9351);
nand U18198 (N_18198,N_6864,N_9478);
nand U18199 (N_18199,N_11698,N_6531);
nand U18200 (N_18200,N_11963,N_11203);
xor U18201 (N_18201,N_9745,N_7979);
nor U18202 (N_18202,N_10310,N_10195);
nand U18203 (N_18203,N_10493,N_11358);
or U18204 (N_18204,N_8512,N_12046);
nor U18205 (N_18205,N_9471,N_9839);
nor U18206 (N_18206,N_6452,N_7425);
and U18207 (N_18207,N_11045,N_11595);
or U18208 (N_18208,N_12333,N_6456);
and U18209 (N_18209,N_7384,N_8656);
nand U18210 (N_18210,N_8155,N_8529);
nand U18211 (N_18211,N_7726,N_8108);
or U18212 (N_18212,N_7631,N_8799);
nand U18213 (N_18213,N_9992,N_9609);
and U18214 (N_18214,N_9824,N_10283);
or U18215 (N_18215,N_6436,N_12036);
nor U18216 (N_18216,N_7392,N_10482);
nor U18217 (N_18217,N_8933,N_8547);
nor U18218 (N_18218,N_7504,N_9238);
xor U18219 (N_18219,N_6679,N_8629);
xor U18220 (N_18220,N_11570,N_7536);
and U18221 (N_18221,N_8791,N_11638);
or U18222 (N_18222,N_9213,N_7725);
nor U18223 (N_18223,N_6504,N_7825);
nor U18224 (N_18224,N_11078,N_9899);
and U18225 (N_18225,N_8478,N_6603);
or U18226 (N_18226,N_10432,N_8289);
nand U18227 (N_18227,N_10554,N_7581);
nand U18228 (N_18228,N_11440,N_8824);
nor U18229 (N_18229,N_11393,N_10021);
nor U18230 (N_18230,N_8960,N_10079);
nand U18231 (N_18231,N_8212,N_10359);
nor U18232 (N_18232,N_10694,N_6846);
nor U18233 (N_18233,N_6486,N_8485);
xor U18234 (N_18234,N_12353,N_7917);
nand U18235 (N_18235,N_7642,N_6942);
or U18236 (N_18236,N_9117,N_7297);
nand U18237 (N_18237,N_12455,N_6388);
and U18238 (N_18238,N_6854,N_9716);
or U18239 (N_18239,N_11725,N_10247);
and U18240 (N_18240,N_7327,N_10908);
nand U18241 (N_18241,N_8669,N_8464);
and U18242 (N_18242,N_11732,N_10767);
nor U18243 (N_18243,N_6805,N_8162);
or U18244 (N_18244,N_11850,N_12164);
or U18245 (N_18245,N_8934,N_6516);
and U18246 (N_18246,N_10718,N_8788);
nand U18247 (N_18247,N_8660,N_12377);
and U18248 (N_18248,N_10946,N_7511);
nand U18249 (N_18249,N_11682,N_11948);
nand U18250 (N_18250,N_11660,N_12361);
or U18251 (N_18251,N_7587,N_8503);
nor U18252 (N_18252,N_7452,N_6277);
nor U18253 (N_18253,N_11780,N_7710);
or U18254 (N_18254,N_9206,N_10648);
or U18255 (N_18255,N_10851,N_9658);
or U18256 (N_18256,N_7286,N_12202);
or U18257 (N_18257,N_8074,N_9930);
nand U18258 (N_18258,N_7676,N_10056);
nand U18259 (N_18259,N_7189,N_12340);
and U18260 (N_18260,N_6921,N_11774);
or U18261 (N_18261,N_8906,N_6573);
and U18262 (N_18262,N_10678,N_9475);
and U18263 (N_18263,N_9424,N_12353);
or U18264 (N_18264,N_6252,N_9277);
and U18265 (N_18265,N_8547,N_9366);
and U18266 (N_18266,N_11767,N_9807);
nor U18267 (N_18267,N_12476,N_7791);
xnor U18268 (N_18268,N_8894,N_7086);
nand U18269 (N_18269,N_9705,N_8194);
and U18270 (N_18270,N_6464,N_10397);
xor U18271 (N_18271,N_11047,N_10815);
nor U18272 (N_18272,N_11189,N_7462);
nand U18273 (N_18273,N_10196,N_7460);
nor U18274 (N_18274,N_12411,N_8649);
and U18275 (N_18275,N_7471,N_8760);
xor U18276 (N_18276,N_8002,N_11599);
or U18277 (N_18277,N_10679,N_10824);
nand U18278 (N_18278,N_6512,N_8515);
or U18279 (N_18279,N_7122,N_10400);
and U18280 (N_18280,N_12306,N_6541);
nor U18281 (N_18281,N_11799,N_10109);
xor U18282 (N_18282,N_10930,N_11404);
and U18283 (N_18283,N_12002,N_8283);
nor U18284 (N_18284,N_12170,N_6486);
nand U18285 (N_18285,N_9677,N_9647);
nor U18286 (N_18286,N_7891,N_9571);
nand U18287 (N_18287,N_9194,N_9114);
or U18288 (N_18288,N_7333,N_12088);
or U18289 (N_18289,N_10151,N_8505);
nand U18290 (N_18290,N_10129,N_8094);
nand U18291 (N_18291,N_7611,N_11098);
nand U18292 (N_18292,N_7355,N_12327);
and U18293 (N_18293,N_11726,N_10014);
or U18294 (N_18294,N_12452,N_12344);
nor U18295 (N_18295,N_7489,N_7209);
xnor U18296 (N_18296,N_9756,N_9181);
nand U18297 (N_18297,N_7834,N_11089);
or U18298 (N_18298,N_11379,N_6313);
nand U18299 (N_18299,N_7487,N_7182);
nand U18300 (N_18300,N_9515,N_10973);
and U18301 (N_18301,N_7559,N_9427);
nand U18302 (N_18302,N_10487,N_9190);
and U18303 (N_18303,N_11840,N_6261);
nand U18304 (N_18304,N_11958,N_11749);
and U18305 (N_18305,N_11022,N_12093);
and U18306 (N_18306,N_6252,N_12298);
nor U18307 (N_18307,N_9082,N_11492);
and U18308 (N_18308,N_8744,N_7683);
or U18309 (N_18309,N_6633,N_6714);
nor U18310 (N_18310,N_9054,N_10290);
xnor U18311 (N_18311,N_7106,N_8844);
nor U18312 (N_18312,N_6570,N_9136);
nand U18313 (N_18313,N_9401,N_7440);
xnor U18314 (N_18314,N_8135,N_6661);
nor U18315 (N_18315,N_12342,N_6807);
or U18316 (N_18316,N_7041,N_11554);
nand U18317 (N_18317,N_10653,N_7854);
or U18318 (N_18318,N_7333,N_9015);
xnor U18319 (N_18319,N_6744,N_8652);
nor U18320 (N_18320,N_8635,N_7897);
nand U18321 (N_18321,N_10731,N_12077);
xor U18322 (N_18322,N_11832,N_7682);
xnor U18323 (N_18323,N_9313,N_9084);
and U18324 (N_18324,N_7574,N_10157);
nor U18325 (N_18325,N_9839,N_10262);
xor U18326 (N_18326,N_12131,N_6796);
nor U18327 (N_18327,N_10319,N_7347);
nand U18328 (N_18328,N_9393,N_8957);
nand U18329 (N_18329,N_6343,N_9272);
xor U18330 (N_18330,N_8290,N_11661);
nor U18331 (N_18331,N_12144,N_6684);
or U18332 (N_18332,N_10531,N_8684);
or U18333 (N_18333,N_12037,N_9802);
nand U18334 (N_18334,N_7169,N_11069);
and U18335 (N_18335,N_11501,N_11707);
nor U18336 (N_18336,N_6999,N_10433);
nand U18337 (N_18337,N_11800,N_10256);
or U18338 (N_18338,N_9261,N_6828);
and U18339 (N_18339,N_8916,N_9091);
and U18340 (N_18340,N_6382,N_7450);
nor U18341 (N_18341,N_6909,N_10058);
nor U18342 (N_18342,N_11220,N_6865);
nor U18343 (N_18343,N_12202,N_8816);
nand U18344 (N_18344,N_9076,N_8899);
nor U18345 (N_18345,N_7694,N_10939);
nor U18346 (N_18346,N_11817,N_10790);
or U18347 (N_18347,N_12321,N_10228);
and U18348 (N_18348,N_11458,N_9285);
or U18349 (N_18349,N_7562,N_7350);
and U18350 (N_18350,N_11133,N_10416);
and U18351 (N_18351,N_6792,N_7540);
nor U18352 (N_18352,N_10692,N_10006);
nand U18353 (N_18353,N_11222,N_12456);
nor U18354 (N_18354,N_6677,N_8729);
and U18355 (N_18355,N_6750,N_7783);
nor U18356 (N_18356,N_11386,N_10951);
nand U18357 (N_18357,N_11699,N_10617);
and U18358 (N_18358,N_11691,N_11377);
and U18359 (N_18359,N_8238,N_11872);
and U18360 (N_18360,N_10844,N_11190);
nor U18361 (N_18361,N_11886,N_12421);
and U18362 (N_18362,N_11526,N_9492);
nand U18363 (N_18363,N_6613,N_9224);
nand U18364 (N_18364,N_8372,N_6991);
nand U18365 (N_18365,N_10590,N_8116);
nor U18366 (N_18366,N_10821,N_9203);
nor U18367 (N_18367,N_6881,N_8159);
xor U18368 (N_18368,N_7206,N_7618);
xnor U18369 (N_18369,N_6634,N_12279);
nand U18370 (N_18370,N_8893,N_12045);
and U18371 (N_18371,N_8951,N_6788);
and U18372 (N_18372,N_8071,N_8023);
and U18373 (N_18373,N_7603,N_6844);
or U18374 (N_18374,N_9903,N_8149);
and U18375 (N_18375,N_8670,N_11881);
xnor U18376 (N_18376,N_11388,N_6633);
nand U18377 (N_18377,N_11972,N_10418);
or U18378 (N_18378,N_9006,N_10556);
and U18379 (N_18379,N_9744,N_7252);
or U18380 (N_18380,N_11915,N_6300);
or U18381 (N_18381,N_12453,N_10920);
nand U18382 (N_18382,N_12137,N_8334);
and U18383 (N_18383,N_10763,N_10747);
nor U18384 (N_18384,N_10261,N_7523);
nand U18385 (N_18385,N_8318,N_8735);
nand U18386 (N_18386,N_11280,N_8038);
or U18387 (N_18387,N_7949,N_10587);
nor U18388 (N_18388,N_10349,N_6892);
nor U18389 (N_18389,N_11820,N_8714);
or U18390 (N_18390,N_8357,N_7808);
nor U18391 (N_18391,N_11525,N_9242);
xor U18392 (N_18392,N_8430,N_7497);
nor U18393 (N_18393,N_6425,N_10336);
and U18394 (N_18394,N_9452,N_8347);
or U18395 (N_18395,N_11521,N_6455);
and U18396 (N_18396,N_8869,N_9085);
or U18397 (N_18397,N_10534,N_6543);
nor U18398 (N_18398,N_10664,N_11347);
nand U18399 (N_18399,N_10014,N_8082);
nand U18400 (N_18400,N_11440,N_7239);
or U18401 (N_18401,N_10483,N_8657);
and U18402 (N_18402,N_8983,N_9060);
nand U18403 (N_18403,N_6665,N_11084);
and U18404 (N_18404,N_6933,N_6863);
nor U18405 (N_18405,N_10194,N_9128);
and U18406 (N_18406,N_9979,N_7534);
nand U18407 (N_18407,N_8776,N_11448);
nand U18408 (N_18408,N_7353,N_10445);
or U18409 (N_18409,N_9242,N_7597);
or U18410 (N_18410,N_10009,N_10514);
nor U18411 (N_18411,N_10291,N_9175);
or U18412 (N_18412,N_10332,N_11979);
nor U18413 (N_18413,N_12449,N_11053);
and U18414 (N_18414,N_7407,N_11555);
and U18415 (N_18415,N_11349,N_8202);
nand U18416 (N_18416,N_10140,N_11075);
nor U18417 (N_18417,N_11078,N_9977);
or U18418 (N_18418,N_11196,N_6637);
and U18419 (N_18419,N_11296,N_7273);
nand U18420 (N_18420,N_7764,N_8701);
xnor U18421 (N_18421,N_9291,N_12390);
and U18422 (N_18422,N_12473,N_9296);
nor U18423 (N_18423,N_10540,N_7129);
xnor U18424 (N_18424,N_7907,N_9709);
and U18425 (N_18425,N_11361,N_8105);
and U18426 (N_18426,N_8948,N_9270);
nor U18427 (N_18427,N_11487,N_6737);
and U18428 (N_18428,N_9224,N_10017);
xnor U18429 (N_18429,N_11351,N_11874);
nand U18430 (N_18430,N_8853,N_7480);
xor U18431 (N_18431,N_8582,N_10247);
xor U18432 (N_18432,N_7212,N_11787);
nand U18433 (N_18433,N_9145,N_10581);
or U18434 (N_18434,N_7111,N_11375);
nand U18435 (N_18435,N_6563,N_9888);
nand U18436 (N_18436,N_10113,N_12485);
and U18437 (N_18437,N_10876,N_8721);
xor U18438 (N_18438,N_11842,N_11391);
and U18439 (N_18439,N_7119,N_8933);
nand U18440 (N_18440,N_8861,N_8652);
nor U18441 (N_18441,N_6458,N_12222);
nand U18442 (N_18442,N_12129,N_9643);
or U18443 (N_18443,N_9995,N_9806);
or U18444 (N_18444,N_10036,N_12105);
or U18445 (N_18445,N_10068,N_9007);
nor U18446 (N_18446,N_6260,N_10886);
nor U18447 (N_18447,N_12093,N_12358);
nand U18448 (N_18448,N_12062,N_6813);
nand U18449 (N_18449,N_11311,N_10314);
nor U18450 (N_18450,N_7882,N_7398);
or U18451 (N_18451,N_6303,N_9546);
or U18452 (N_18452,N_8492,N_10151);
or U18453 (N_18453,N_7806,N_9100);
nand U18454 (N_18454,N_11840,N_10521);
and U18455 (N_18455,N_6977,N_9523);
nand U18456 (N_18456,N_8382,N_6378);
or U18457 (N_18457,N_6579,N_9535);
nand U18458 (N_18458,N_7869,N_6858);
nor U18459 (N_18459,N_9663,N_6767);
nand U18460 (N_18460,N_6924,N_12207);
nand U18461 (N_18461,N_7727,N_8740);
and U18462 (N_18462,N_12393,N_9431);
nor U18463 (N_18463,N_12068,N_10117);
xor U18464 (N_18464,N_10101,N_6328);
or U18465 (N_18465,N_10604,N_7878);
and U18466 (N_18466,N_7639,N_11156);
and U18467 (N_18467,N_7321,N_11953);
and U18468 (N_18468,N_6938,N_8644);
and U18469 (N_18469,N_8221,N_10844);
nand U18470 (N_18470,N_12037,N_10932);
nand U18471 (N_18471,N_11731,N_7755);
xnor U18472 (N_18472,N_8409,N_11472);
or U18473 (N_18473,N_8196,N_10669);
xor U18474 (N_18474,N_7544,N_8777);
nand U18475 (N_18475,N_9691,N_9272);
nor U18476 (N_18476,N_11054,N_6746);
and U18477 (N_18477,N_12226,N_6433);
nor U18478 (N_18478,N_8422,N_8027);
or U18479 (N_18479,N_12150,N_9375);
nor U18480 (N_18480,N_9441,N_9896);
nor U18481 (N_18481,N_9507,N_10393);
nand U18482 (N_18482,N_12436,N_8421);
nor U18483 (N_18483,N_8773,N_6597);
nor U18484 (N_18484,N_11824,N_9368);
and U18485 (N_18485,N_11709,N_7564);
nand U18486 (N_18486,N_12090,N_7190);
nand U18487 (N_18487,N_8137,N_9787);
nand U18488 (N_18488,N_8066,N_9806);
and U18489 (N_18489,N_11182,N_8993);
nand U18490 (N_18490,N_7706,N_11737);
and U18491 (N_18491,N_7855,N_11747);
nand U18492 (N_18492,N_6566,N_8099);
and U18493 (N_18493,N_9034,N_9773);
nand U18494 (N_18494,N_9636,N_8943);
or U18495 (N_18495,N_8881,N_8462);
nand U18496 (N_18496,N_6608,N_9590);
nor U18497 (N_18497,N_10078,N_9418);
or U18498 (N_18498,N_11847,N_10338);
nor U18499 (N_18499,N_6759,N_10181);
or U18500 (N_18500,N_6734,N_9287);
and U18501 (N_18501,N_8719,N_12287);
or U18502 (N_18502,N_10120,N_8620);
and U18503 (N_18503,N_11268,N_8312);
nand U18504 (N_18504,N_9886,N_7253);
xor U18505 (N_18505,N_11799,N_8993);
nand U18506 (N_18506,N_11143,N_7631);
or U18507 (N_18507,N_12253,N_7438);
nor U18508 (N_18508,N_7540,N_8859);
and U18509 (N_18509,N_8516,N_7733);
nor U18510 (N_18510,N_8049,N_9159);
or U18511 (N_18511,N_9213,N_11675);
and U18512 (N_18512,N_8706,N_8779);
and U18513 (N_18513,N_9418,N_8074);
or U18514 (N_18514,N_6806,N_9437);
nand U18515 (N_18515,N_11513,N_8819);
nand U18516 (N_18516,N_9394,N_7987);
or U18517 (N_18517,N_9000,N_6543);
or U18518 (N_18518,N_11365,N_8833);
nand U18519 (N_18519,N_10075,N_8225);
nand U18520 (N_18520,N_12360,N_11097);
nand U18521 (N_18521,N_11687,N_8849);
and U18522 (N_18522,N_9540,N_11895);
and U18523 (N_18523,N_10416,N_11733);
or U18524 (N_18524,N_10618,N_11700);
and U18525 (N_18525,N_8912,N_9386);
nor U18526 (N_18526,N_9283,N_10931);
nor U18527 (N_18527,N_9965,N_6802);
or U18528 (N_18528,N_9261,N_7458);
and U18529 (N_18529,N_12377,N_12427);
or U18530 (N_18530,N_6565,N_6687);
and U18531 (N_18531,N_10389,N_9664);
and U18532 (N_18532,N_6294,N_10438);
nor U18533 (N_18533,N_8488,N_6938);
xnor U18534 (N_18534,N_7721,N_10432);
or U18535 (N_18535,N_9265,N_9644);
or U18536 (N_18536,N_8405,N_10553);
or U18537 (N_18537,N_11735,N_8808);
xor U18538 (N_18538,N_12281,N_8317);
or U18539 (N_18539,N_10992,N_6826);
nand U18540 (N_18540,N_9344,N_11929);
and U18541 (N_18541,N_6341,N_10877);
or U18542 (N_18542,N_11779,N_9050);
and U18543 (N_18543,N_11329,N_6576);
nor U18544 (N_18544,N_12329,N_11389);
nor U18545 (N_18545,N_11011,N_10053);
nand U18546 (N_18546,N_8604,N_6578);
xnor U18547 (N_18547,N_8590,N_7478);
xnor U18548 (N_18548,N_7905,N_7506);
nand U18549 (N_18549,N_9934,N_7287);
xor U18550 (N_18550,N_11815,N_10559);
and U18551 (N_18551,N_11156,N_8509);
nor U18552 (N_18552,N_12059,N_6785);
xnor U18553 (N_18553,N_11086,N_9226);
nand U18554 (N_18554,N_6867,N_9770);
nand U18555 (N_18555,N_8873,N_8867);
nand U18556 (N_18556,N_10949,N_9042);
and U18557 (N_18557,N_8071,N_10200);
or U18558 (N_18558,N_12185,N_10359);
or U18559 (N_18559,N_8196,N_10454);
and U18560 (N_18560,N_10893,N_10621);
nor U18561 (N_18561,N_7817,N_7929);
xnor U18562 (N_18562,N_8282,N_9302);
nand U18563 (N_18563,N_10585,N_12066);
or U18564 (N_18564,N_7291,N_8841);
nor U18565 (N_18565,N_10071,N_10301);
and U18566 (N_18566,N_8043,N_12309);
nand U18567 (N_18567,N_7335,N_8588);
or U18568 (N_18568,N_9768,N_6260);
and U18569 (N_18569,N_6989,N_10088);
and U18570 (N_18570,N_9940,N_9015);
or U18571 (N_18571,N_8000,N_12163);
xnor U18572 (N_18572,N_10104,N_6876);
xor U18573 (N_18573,N_10373,N_9232);
and U18574 (N_18574,N_11230,N_7537);
nand U18575 (N_18575,N_9072,N_7556);
and U18576 (N_18576,N_10459,N_8252);
xor U18577 (N_18577,N_6357,N_9125);
nor U18578 (N_18578,N_8853,N_10531);
or U18579 (N_18579,N_7827,N_8993);
nand U18580 (N_18580,N_6574,N_6652);
nor U18581 (N_18581,N_6853,N_10121);
xnor U18582 (N_18582,N_11694,N_9307);
nor U18583 (N_18583,N_10904,N_6805);
and U18584 (N_18584,N_7505,N_9711);
nand U18585 (N_18585,N_7166,N_12308);
nor U18586 (N_18586,N_7106,N_8875);
and U18587 (N_18587,N_11779,N_7468);
nand U18588 (N_18588,N_10918,N_8785);
nor U18589 (N_18589,N_8059,N_11247);
or U18590 (N_18590,N_7838,N_9070);
and U18591 (N_18591,N_6622,N_10954);
nor U18592 (N_18592,N_11319,N_11344);
nor U18593 (N_18593,N_7409,N_8228);
xor U18594 (N_18594,N_11750,N_10214);
nand U18595 (N_18595,N_7986,N_11517);
or U18596 (N_18596,N_9759,N_8408);
nand U18597 (N_18597,N_9100,N_6652);
nand U18598 (N_18598,N_11468,N_9893);
nor U18599 (N_18599,N_6898,N_12366);
nor U18600 (N_18600,N_7026,N_8113);
or U18601 (N_18601,N_8950,N_11694);
nor U18602 (N_18602,N_11826,N_11490);
and U18603 (N_18603,N_8620,N_8340);
and U18604 (N_18604,N_10559,N_11088);
and U18605 (N_18605,N_10544,N_8817);
nor U18606 (N_18606,N_7865,N_6961);
and U18607 (N_18607,N_7682,N_7659);
xnor U18608 (N_18608,N_9672,N_9902);
and U18609 (N_18609,N_9864,N_9538);
nand U18610 (N_18610,N_9700,N_7700);
or U18611 (N_18611,N_7533,N_8346);
and U18612 (N_18612,N_11700,N_10413);
nor U18613 (N_18613,N_6621,N_9217);
or U18614 (N_18614,N_10214,N_7567);
or U18615 (N_18615,N_8703,N_6463);
nor U18616 (N_18616,N_11786,N_7307);
nor U18617 (N_18617,N_7565,N_7476);
nor U18618 (N_18618,N_9121,N_7100);
and U18619 (N_18619,N_7813,N_6855);
nand U18620 (N_18620,N_7745,N_7277);
nand U18621 (N_18621,N_9500,N_7271);
nand U18622 (N_18622,N_8329,N_6903);
nand U18623 (N_18623,N_7554,N_11774);
or U18624 (N_18624,N_10811,N_10247);
or U18625 (N_18625,N_8929,N_7162);
xnor U18626 (N_18626,N_9820,N_6906);
nor U18627 (N_18627,N_8849,N_8845);
nand U18628 (N_18628,N_8988,N_9097);
nor U18629 (N_18629,N_11271,N_9357);
xor U18630 (N_18630,N_7060,N_8356);
nor U18631 (N_18631,N_8476,N_9964);
nand U18632 (N_18632,N_12448,N_11001);
xor U18633 (N_18633,N_8564,N_10977);
nand U18634 (N_18634,N_9292,N_6846);
and U18635 (N_18635,N_12415,N_10031);
and U18636 (N_18636,N_8371,N_8118);
and U18637 (N_18637,N_6649,N_9563);
nor U18638 (N_18638,N_9304,N_10364);
and U18639 (N_18639,N_7646,N_8677);
and U18640 (N_18640,N_9783,N_10781);
and U18641 (N_18641,N_9991,N_7655);
and U18642 (N_18642,N_8529,N_11806);
xor U18643 (N_18643,N_9136,N_7396);
or U18644 (N_18644,N_9577,N_11729);
and U18645 (N_18645,N_9697,N_7603);
nor U18646 (N_18646,N_8817,N_9546);
or U18647 (N_18647,N_10340,N_8601);
or U18648 (N_18648,N_11265,N_10600);
nand U18649 (N_18649,N_9679,N_9965);
or U18650 (N_18650,N_10499,N_7079);
nand U18651 (N_18651,N_9797,N_11678);
nand U18652 (N_18652,N_7860,N_7850);
nand U18653 (N_18653,N_10487,N_11035);
nand U18654 (N_18654,N_11506,N_8120);
and U18655 (N_18655,N_9619,N_7824);
nand U18656 (N_18656,N_7919,N_6398);
and U18657 (N_18657,N_9499,N_12258);
or U18658 (N_18658,N_8243,N_6497);
or U18659 (N_18659,N_12156,N_6958);
nor U18660 (N_18660,N_10280,N_8394);
nor U18661 (N_18661,N_6606,N_10959);
and U18662 (N_18662,N_11924,N_7787);
nor U18663 (N_18663,N_6858,N_8502);
and U18664 (N_18664,N_8341,N_6698);
nand U18665 (N_18665,N_7263,N_6869);
and U18666 (N_18666,N_11815,N_11891);
nor U18667 (N_18667,N_7975,N_8828);
nand U18668 (N_18668,N_8721,N_7559);
xnor U18669 (N_18669,N_9216,N_12131);
xor U18670 (N_18670,N_6733,N_8013);
and U18671 (N_18671,N_9400,N_11844);
nand U18672 (N_18672,N_8938,N_7746);
and U18673 (N_18673,N_7785,N_12277);
or U18674 (N_18674,N_12147,N_6561);
or U18675 (N_18675,N_9708,N_7191);
xnor U18676 (N_18676,N_12043,N_10784);
nor U18677 (N_18677,N_7295,N_10873);
nor U18678 (N_18678,N_11930,N_11304);
and U18679 (N_18679,N_9050,N_10720);
or U18680 (N_18680,N_6523,N_9568);
or U18681 (N_18681,N_7885,N_9100);
and U18682 (N_18682,N_6862,N_8891);
or U18683 (N_18683,N_6723,N_6902);
nor U18684 (N_18684,N_8473,N_8762);
and U18685 (N_18685,N_12472,N_12228);
xnor U18686 (N_18686,N_9162,N_6672);
or U18687 (N_18687,N_10807,N_7341);
and U18688 (N_18688,N_6337,N_9951);
nand U18689 (N_18689,N_11342,N_9006);
nand U18690 (N_18690,N_7821,N_6754);
nor U18691 (N_18691,N_9178,N_7669);
nand U18692 (N_18692,N_6923,N_10048);
nand U18693 (N_18693,N_9890,N_7492);
nand U18694 (N_18694,N_9889,N_10816);
or U18695 (N_18695,N_7900,N_10878);
nand U18696 (N_18696,N_9483,N_11105);
or U18697 (N_18697,N_6501,N_6643);
xnor U18698 (N_18698,N_12034,N_7221);
nand U18699 (N_18699,N_11638,N_8213);
or U18700 (N_18700,N_8824,N_9346);
xnor U18701 (N_18701,N_9773,N_6289);
nand U18702 (N_18702,N_8354,N_11762);
nor U18703 (N_18703,N_11941,N_10177);
nand U18704 (N_18704,N_8554,N_7321);
nand U18705 (N_18705,N_10756,N_12170);
nor U18706 (N_18706,N_9598,N_10515);
nand U18707 (N_18707,N_6299,N_8640);
or U18708 (N_18708,N_9813,N_11237);
and U18709 (N_18709,N_8839,N_11309);
nor U18710 (N_18710,N_6419,N_9350);
or U18711 (N_18711,N_8801,N_8092);
nand U18712 (N_18712,N_7071,N_11548);
nor U18713 (N_18713,N_9240,N_10452);
nor U18714 (N_18714,N_9823,N_11732);
nor U18715 (N_18715,N_8936,N_6449);
or U18716 (N_18716,N_9146,N_11865);
nor U18717 (N_18717,N_12477,N_7816);
or U18718 (N_18718,N_11559,N_8713);
nand U18719 (N_18719,N_10423,N_10163);
nor U18720 (N_18720,N_7723,N_8559);
or U18721 (N_18721,N_10247,N_11365);
and U18722 (N_18722,N_7229,N_12119);
nor U18723 (N_18723,N_8600,N_11034);
and U18724 (N_18724,N_12026,N_9327);
xor U18725 (N_18725,N_12462,N_12370);
or U18726 (N_18726,N_9351,N_8642);
nor U18727 (N_18727,N_10109,N_7929);
and U18728 (N_18728,N_6989,N_7207);
nor U18729 (N_18729,N_6576,N_10160);
or U18730 (N_18730,N_7565,N_10751);
and U18731 (N_18731,N_11553,N_7695);
and U18732 (N_18732,N_9779,N_9278);
and U18733 (N_18733,N_8495,N_10064);
nor U18734 (N_18734,N_10637,N_8819);
nand U18735 (N_18735,N_11523,N_11613);
nor U18736 (N_18736,N_6410,N_6481);
nand U18737 (N_18737,N_8673,N_7171);
or U18738 (N_18738,N_10333,N_9750);
xnor U18739 (N_18739,N_9457,N_6871);
xnor U18740 (N_18740,N_8782,N_10466);
and U18741 (N_18741,N_11866,N_9532);
nand U18742 (N_18742,N_9272,N_12096);
and U18743 (N_18743,N_7184,N_11051);
and U18744 (N_18744,N_9811,N_10289);
nand U18745 (N_18745,N_9347,N_8534);
nor U18746 (N_18746,N_8915,N_10576);
nand U18747 (N_18747,N_11039,N_9880);
or U18748 (N_18748,N_7526,N_7450);
and U18749 (N_18749,N_8903,N_10919);
and U18750 (N_18750,N_13374,N_16540);
and U18751 (N_18751,N_16296,N_15023);
nor U18752 (N_18752,N_14336,N_13730);
and U18753 (N_18753,N_17697,N_12573);
and U18754 (N_18754,N_16232,N_12793);
and U18755 (N_18755,N_13464,N_13042);
and U18756 (N_18756,N_17538,N_13302);
nand U18757 (N_18757,N_17474,N_13776);
or U18758 (N_18758,N_13455,N_14632);
nor U18759 (N_18759,N_15606,N_13153);
and U18760 (N_18760,N_14316,N_14181);
nand U18761 (N_18761,N_15855,N_17950);
xnor U18762 (N_18762,N_13401,N_14600);
nand U18763 (N_18763,N_18130,N_16925);
and U18764 (N_18764,N_15942,N_14379);
nor U18765 (N_18765,N_12665,N_17267);
or U18766 (N_18766,N_18282,N_14978);
xnor U18767 (N_18767,N_16693,N_17013);
xor U18768 (N_18768,N_12757,N_18656);
or U18769 (N_18769,N_16533,N_16317);
or U18770 (N_18770,N_18342,N_17226);
or U18771 (N_18771,N_12918,N_18539);
nor U18772 (N_18772,N_13486,N_17814);
nand U18773 (N_18773,N_16749,N_12820);
xor U18774 (N_18774,N_16347,N_14505);
nor U18775 (N_18775,N_17532,N_15796);
or U18776 (N_18776,N_13770,N_14271);
and U18777 (N_18777,N_18525,N_13540);
nor U18778 (N_18778,N_16730,N_17109);
or U18779 (N_18779,N_18194,N_18346);
nor U18780 (N_18780,N_12522,N_15823);
or U18781 (N_18781,N_15920,N_15253);
or U18782 (N_18782,N_18232,N_12632);
and U18783 (N_18783,N_13750,N_13121);
xnor U18784 (N_18784,N_16816,N_18544);
nand U18785 (N_18785,N_15757,N_15870);
or U18786 (N_18786,N_17142,N_18457);
and U18787 (N_18787,N_15625,N_15104);
nand U18788 (N_18788,N_18448,N_16947);
nand U18789 (N_18789,N_12727,N_15396);
and U18790 (N_18790,N_13838,N_12525);
nand U18791 (N_18791,N_18423,N_17342);
and U18792 (N_18792,N_18545,N_14279);
or U18793 (N_18793,N_12978,N_14936);
or U18794 (N_18794,N_14390,N_17012);
xnor U18795 (N_18795,N_16879,N_17736);
nand U18796 (N_18796,N_14631,N_18308);
nand U18797 (N_18797,N_14592,N_14244);
nor U18798 (N_18798,N_13938,N_15360);
or U18799 (N_18799,N_14014,N_14441);
nor U18800 (N_18800,N_15410,N_14041);
and U18801 (N_18801,N_13708,N_15677);
or U18802 (N_18802,N_12566,N_13545);
or U18803 (N_18803,N_14167,N_13445);
or U18804 (N_18804,N_16885,N_16256);
xor U18805 (N_18805,N_16843,N_14677);
and U18806 (N_18806,N_15466,N_16475);
nand U18807 (N_18807,N_16532,N_16093);
nor U18808 (N_18808,N_15668,N_13483);
and U18809 (N_18809,N_16417,N_14026);
nor U18810 (N_18810,N_13740,N_14469);
xor U18811 (N_18811,N_12840,N_15672);
or U18812 (N_18812,N_17333,N_13339);
or U18813 (N_18813,N_16293,N_17786);
nor U18814 (N_18814,N_12680,N_16601);
nor U18815 (N_18815,N_12723,N_14446);
xnor U18816 (N_18816,N_15972,N_16724);
nor U18817 (N_18817,N_16725,N_15459);
or U18818 (N_18818,N_13217,N_15358);
nor U18819 (N_18819,N_17447,N_18198);
nor U18820 (N_18820,N_13356,N_18616);
nand U18821 (N_18821,N_16252,N_13381);
or U18822 (N_18822,N_15762,N_18007);
or U18823 (N_18823,N_12587,N_17312);
nand U18824 (N_18824,N_16991,N_14928);
and U18825 (N_18825,N_14879,N_13937);
nor U18826 (N_18826,N_17325,N_14752);
or U18827 (N_18827,N_15804,N_18627);
nor U18828 (N_18828,N_16972,N_13078);
nor U18829 (N_18829,N_15968,N_16710);
and U18830 (N_18830,N_15304,N_16624);
nand U18831 (N_18831,N_16770,N_13604);
or U18832 (N_18832,N_14957,N_13594);
and U18833 (N_18833,N_13961,N_16344);
and U18834 (N_18834,N_15062,N_18623);
and U18835 (N_18835,N_18048,N_13705);
nor U18836 (N_18836,N_12906,N_13942);
xnor U18837 (N_18837,N_18648,N_15722);
xnor U18838 (N_18838,N_17866,N_16203);
nand U18839 (N_18839,N_15875,N_13935);
nor U18840 (N_18840,N_12790,N_17323);
nor U18841 (N_18841,N_17420,N_17236);
and U18842 (N_18842,N_14912,N_15335);
or U18843 (N_18843,N_17263,N_16267);
xor U18844 (N_18844,N_12631,N_14163);
nor U18845 (N_18845,N_16445,N_12744);
nor U18846 (N_18846,N_16513,N_13627);
nand U18847 (N_18847,N_13715,N_14411);
xor U18848 (N_18848,N_16893,N_12877);
nor U18849 (N_18849,N_17023,N_16968);
nor U18850 (N_18850,N_14251,N_13314);
nor U18851 (N_18851,N_14777,N_16786);
or U18852 (N_18852,N_17001,N_13008);
and U18853 (N_18853,N_16735,N_13949);
xnor U18854 (N_18854,N_15128,N_14521);
nor U18855 (N_18855,N_16509,N_12677);
and U18856 (N_18856,N_13391,N_14385);
and U18857 (N_18857,N_15597,N_13492);
and U18858 (N_18858,N_16107,N_17178);
or U18859 (N_18859,N_14975,N_13116);
nand U18860 (N_18860,N_17644,N_15257);
or U18861 (N_18861,N_12964,N_12528);
nor U18862 (N_18862,N_13568,N_17443);
nor U18863 (N_18863,N_16425,N_16605);
or U18864 (N_18864,N_18298,N_12944);
and U18865 (N_18865,N_16916,N_15027);
xnor U18866 (N_18866,N_16635,N_14992);
nor U18867 (N_18867,N_17617,N_17303);
nand U18868 (N_18868,N_14878,N_16384);
or U18869 (N_18869,N_16497,N_18182);
nor U18870 (N_18870,N_17689,N_18235);
nand U18871 (N_18871,N_15789,N_14257);
nand U18872 (N_18872,N_12618,N_17275);
nand U18873 (N_18873,N_14546,N_18725);
and U18874 (N_18874,N_18701,N_16415);
and U18875 (N_18875,N_15526,N_16284);
or U18876 (N_18876,N_15500,N_17609);
or U18877 (N_18877,N_18234,N_16414);
or U18878 (N_18878,N_15109,N_14525);
nor U18879 (N_18879,N_18599,N_18651);
nand U18880 (N_18880,N_17147,N_13056);
nand U18881 (N_18881,N_15498,N_13058);
or U18882 (N_18882,N_17534,N_15317);
nor U18883 (N_18883,N_16453,N_13647);
nor U18884 (N_18884,N_13433,N_12611);
nor U18885 (N_18885,N_17189,N_16997);
and U18886 (N_18886,N_16768,N_15822);
or U18887 (N_18887,N_17788,N_14341);
and U18888 (N_18888,N_16652,N_13046);
nor U18889 (N_18889,N_16423,N_14935);
nand U18890 (N_18890,N_15996,N_14863);
or U18891 (N_18891,N_16887,N_14808);
nor U18892 (N_18892,N_15457,N_13890);
nand U18893 (N_18893,N_18091,N_17586);
nor U18894 (N_18894,N_15921,N_15352);
or U18895 (N_18895,N_16457,N_13425);
nor U18896 (N_18896,N_16389,N_15419);
or U18897 (N_18897,N_12546,N_14304);
nor U18898 (N_18898,N_16313,N_13535);
and U18899 (N_18899,N_17005,N_15977);
nor U18900 (N_18900,N_18345,N_14328);
and U18901 (N_18901,N_14780,N_14261);
or U18902 (N_18902,N_14319,N_12841);
or U18903 (N_18903,N_14644,N_13621);
and U18904 (N_18904,N_18507,N_15928);
nor U18905 (N_18905,N_13885,N_12803);
and U18906 (N_18906,N_17569,N_18550);
and U18907 (N_18907,N_17799,N_13585);
nor U18908 (N_18908,N_18491,N_15514);
nor U18909 (N_18909,N_18053,N_13934);
and U18910 (N_18910,N_18426,N_13189);
and U18911 (N_18911,N_18337,N_15980);
and U18912 (N_18912,N_12670,N_17271);
and U18913 (N_18913,N_17336,N_14413);
nand U18914 (N_18914,N_18558,N_16867);
or U18915 (N_18915,N_15448,N_16630);
nand U18916 (N_18916,N_15603,N_16585);
nand U18917 (N_18917,N_14009,N_13923);
nand U18918 (N_18918,N_13476,N_16574);
nand U18919 (N_18919,N_14587,N_14637);
nand U18920 (N_18920,N_16969,N_12696);
and U18921 (N_18921,N_14060,N_15879);
or U18922 (N_18922,N_12802,N_18127);
and U18923 (N_18923,N_15661,N_18025);
and U18924 (N_18924,N_13139,N_14406);
and U18925 (N_18925,N_12997,N_13419);
nand U18926 (N_18926,N_13519,N_18196);
nor U18927 (N_18927,N_16748,N_15101);
nand U18928 (N_18928,N_18398,N_14507);
nor U18929 (N_18929,N_18528,N_14554);
and U18930 (N_18930,N_13623,N_15848);
nor U18931 (N_18931,N_16923,N_12876);
or U18932 (N_18932,N_14360,N_12507);
nor U18933 (N_18933,N_17165,N_18236);
xor U18934 (N_18934,N_17824,N_18208);
or U18935 (N_18935,N_15562,N_14420);
nor U18936 (N_18936,N_14877,N_14841);
nor U18937 (N_18937,N_16642,N_13872);
and U18938 (N_18938,N_13548,N_16266);
nor U18939 (N_18939,N_15647,N_15389);
or U18940 (N_18940,N_18051,N_13992);
nor U18941 (N_18941,N_14461,N_14388);
xor U18942 (N_18942,N_15939,N_18187);
nand U18943 (N_18943,N_17287,N_16122);
and U18944 (N_18944,N_16699,N_13734);
nand U18945 (N_18945,N_13493,N_13063);
or U18946 (N_18946,N_18008,N_14905);
nand U18947 (N_18947,N_17953,N_13386);
nor U18948 (N_18948,N_14933,N_13372);
or U18949 (N_18949,N_13466,N_12594);
or U18950 (N_18950,N_15041,N_15851);
nor U18951 (N_18951,N_16025,N_17429);
and U18952 (N_18952,N_15753,N_18253);
or U18953 (N_18953,N_18071,N_13598);
or U18954 (N_18954,N_12725,N_17505);
and U18955 (N_18955,N_15281,N_17311);
and U18956 (N_18956,N_17280,N_15657);
and U18957 (N_18957,N_15014,N_16162);
nand U18958 (N_18958,N_18445,N_17565);
and U18959 (N_18959,N_12954,N_15692);
nor U18960 (N_18960,N_15797,N_15127);
and U18961 (N_18961,N_13323,N_14395);
nor U18962 (N_18962,N_15948,N_12502);
and U18963 (N_18963,N_13000,N_13773);
nand U18964 (N_18964,N_16449,N_17868);
nand U18965 (N_18965,N_16094,N_12628);
nand U18966 (N_18966,N_15084,N_12729);
and U18967 (N_18967,N_14019,N_16557);
nand U18968 (N_18968,N_12728,N_15213);
and U18969 (N_18969,N_14410,N_16620);
nand U18970 (N_18970,N_15286,N_15428);
or U18971 (N_18971,N_14083,N_15516);
or U18972 (N_18972,N_16776,N_18710);
nand U18973 (N_18973,N_16712,N_13043);
or U18974 (N_18974,N_17640,N_13470);
xor U18975 (N_18975,N_13211,N_16657);
xor U18976 (N_18976,N_18425,N_17625);
and U18977 (N_18977,N_18715,N_12578);
nor U18978 (N_18978,N_13093,N_13396);
and U18979 (N_18979,N_15187,N_17401);
nor U18980 (N_18980,N_17873,N_14909);
and U18981 (N_18981,N_15145,N_14913);
nor U18982 (N_18982,N_13659,N_18180);
and U18983 (N_18983,N_17428,N_14378);
nand U18984 (N_18984,N_15015,N_17975);
or U18985 (N_18985,N_13031,N_15832);
nand U18986 (N_18986,N_13276,N_18277);
nor U18987 (N_18987,N_14591,N_15946);
and U18988 (N_18988,N_15739,N_18576);
nand U18989 (N_18989,N_15566,N_15183);
or U18990 (N_18990,N_13275,N_14571);
and U18991 (N_18991,N_17934,N_14775);
and U18992 (N_18992,N_17389,N_14498);
and U18993 (N_18993,N_17997,N_15475);
nor U18994 (N_18994,N_16790,N_12779);
and U18995 (N_18995,N_13791,N_16520);
nor U18996 (N_18996,N_18063,N_18359);
and U18997 (N_18997,N_14674,N_14856);
or U18998 (N_18998,N_13956,N_15313);
nor U18999 (N_18999,N_15278,N_18114);
nor U19000 (N_19000,N_13216,N_13224);
and U19001 (N_19001,N_16376,N_15510);
or U19002 (N_19002,N_13634,N_14621);
nand U19003 (N_19003,N_17986,N_15857);
and U19004 (N_19004,N_12610,N_18205);
nand U19005 (N_19005,N_14986,N_17525);
nand U19006 (N_19006,N_12821,N_13782);
xor U19007 (N_19007,N_13729,N_13907);
nand U19008 (N_19008,N_18289,N_16292);
and U19009 (N_19009,N_14002,N_14593);
xnor U19010 (N_19010,N_14307,N_17916);
or U19011 (N_19011,N_17437,N_18142);
nand U19012 (N_19012,N_18256,N_12915);
nor U19013 (N_19013,N_14065,N_18642);
and U19014 (N_19014,N_16694,N_13716);
or U19015 (N_19015,N_14810,N_18296);
nor U19016 (N_19016,N_14444,N_13501);
nand U19017 (N_19017,N_18744,N_14246);
and U19018 (N_19018,N_12942,N_14322);
or U19019 (N_19019,N_15247,N_14838);
and U19020 (N_19020,N_15890,N_17466);
or U19021 (N_19021,N_16764,N_13354);
and U19022 (N_19022,N_14764,N_12734);
nand U19023 (N_19023,N_18489,N_13979);
nand U19024 (N_19024,N_12601,N_17821);
nand U19025 (N_19025,N_16807,N_15530);
nand U19026 (N_19026,N_16402,N_14500);
nor U19027 (N_19027,N_14721,N_18462);
nand U19028 (N_19028,N_12605,N_16200);
nor U19029 (N_19029,N_18559,N_16371);
and U19030 (N_19030,N_18242,N_13377);
or U19031 (N_19031,N_13289,N_14459);
and U19032 (N_19032,N_18252,N_13030);
nand U19033 (N_19033,N_13766,N_17996);
and U19034 (N_19034,N_13193,N_15019);
nor U19035 (N_19035,N_15158,N_17862);
or U19036 (N_19036,N_15214,N_15095);
or U19037 (N_19037,N_15649,N_18742);
nand U19038 (N_19038,N_15151,N_18211);
nor U19039 (N_19039,N_13691,N_14214);
nor U19040 (N_19040,N_13821,N_17239);
xnor U19041 (N_19041,N_17203,N_13165);
and U19042 (N_19042,N_13950,N_16424);
nand U19043 (N_19043,N_17943,N_16028);
or U19044 (N_19044,N_17208,N_14747);
nor U19045 (N_19045,N_14127,N_18221);
or U19046 (N_19046,N_15163,N_13188);
and U19047 (N_19047,N_15591,N_13565);
nor U19048 (N_19048,N_17710,N_15346);
or U19049 (N_19049,N_15297,N_14303);
nand U19050 (N_19050,N_16610,N_15340);
or U19051 (N_19051,N_15424,N_16476);
and U19052 (N_19052,N_15669,N_17702);
nor U19053 (N_19053,N_12787,N_17000);
or U19054 (N_19054,N_15758,N_16942);
xnor U19055 (N_19055,N_18708,N_14132);
and U19056 (N_19056,N_16335,N_13728);
and U19057 (N_19057,N_18158,N_13665);
or U19058 (N_19058,N_13184,N_13334);
and U19059 (N_19059,N_17610,N_15940);
nand U19060 (N_19060,N_16840,N_14831);
nand U19061 (N_19061,N_17936,N_17364);
nand U19062 (N_19062,N_16922,N_15152);
nand U19063 (N_19063,N_14087,N_18229);
and U19064 (N_19064,N_16368,N_14397);
and U19065 (N_19065,N_13410,N_13688);
nand U19066 (N_19066,N_16491,N_15755);
or U19067 (N_19067,N_16789,N_14815);
xor U19068 (N_19068,N_15232,N_16303);
nor U19069 (N_19069,N_13235,N_14842);
or U19070 (N_19070,N_14911,N_16332);
or U19071 (N_19071,N_16103,N_14197);
nor U19072 (N_19072,N_18199,N_16006);
nor U19073 (N_19073,N_16035,N_12887);
and U19074 (N_19074,N_16007,N_18514);
and U19075 (N_19075,N_18458,N_15174);
xor U19076 (N_19076,N_15901,N_14769);
or U19077 (N_19077,N_15421,N_13957);
xnor U19078 (N_19078,N_17921,N_16206);
and U19079 (N_19079,N_13051,N_13457);
or U19080 (N_19080,N_14596,N_17794);
or U19081 (N_19081,N_13577,N_13075);
and U19082 (N_19082,N_15464,N_14787);
nor U19083 (N_19083,N_13984,N_18119);
or U19084 (N_19084,N_13684,N_16788);
and U19085 (N_19085,N_17745,N_16331);
or U19086 (N_19086,N_15844,N_12742);
nor U19087 (N_19087,N_18052,N_16091);
or U19088 (N_19088,N_18748,N_14514);
nand U19089 (N_19089,N_15058,N_17260);
and U19090 (N_19090,N_18029,N_16003);
nand U19091 (N_19091,N_17070,N_18269);
and U19092 (N_19092,N_13972,N_15406);
nor U19093 (N_19093,N_18064,N_14695);
or U19094 (N_19094,N_15502,N_12773);
nor U19095 (N_19095,N_16121,N_12564);
nand U19096 (N_19096,N_12570,N_16729);
and U19097 (N_19097,N_13028,N_16911);
xor U19098 (N_19098,N_17549,N_18351);
nor U19099 (N_19099,N_15215,N_17818);
or U19100 (N_19100,N_17110,N_17011);
nor U19101 (N_19101,N_14872,N_14997);
and U19102 (N_19102,N_16286,N_14458);
or U19103 (N_19103,N_15916,N_17557);
and U19104 (N_19104,N_16343,N_17202);
nor U19105 (N_19105,N_13079,N_15981);
xnor U19106 (N_19106,N_16551,N_12881);
nand U19107 (N_19107,N_15721,N_14979);
nand U19108 (N_19108,N_13111,N_14742);
xnor U19109 (N_19109,N_12555,N_12731);
nand U19110 (N_19110,N_16707,N_18446);
and U19111 (N_19111,N_16282,N_15644);
nor U19112 (N_19112,N_13567,N_17732);
nor U19113 (N_19113,N_18303,N_13270);
or U19114 (N_19114,N_17167,N_14727);
or U19115 (N_19115,N_18455,N_12925);
and U19116 (N_19116,N_14106,N_13722);
xor U19117 (N_19117,N_12855,N_12625);
or U19118 (N_19118,N_16291,N_14823);
xnor U19119 (N_19119,N_16116,N_17891);
nand U19120 (N_19120,N_15840,N_15455);
xor U19121 (N_19121,N_16677,N_17805);
and U19122 (N_19122,N_12844,N_15306);
or U19123 (N_19123,N_12621,N_12682);
nor U19124 (N_19124,N_13544,N_17845);
nor U19125 (N_19125,N_13124,N_13080);
xnor U19126 (N_19126,N_14545,N_12952);
and U19127 (N_19127,N_14799,N_12579);
or U19128 (N_19128,N_16846,N_13187);
nor U19129 (N_19129,N_15018,N_13633);
or U19130 (N_19130,N_15223,N_15388);
nand U19131 (N_19131,N_18535,N_15821);
nand U19132 (N_19132,N_12624,N_13037);
nor U19133 (N_19133,N_16839,N_14915);
and U19134 (N_19134,N_17352,N_14301);
or U19135 (N_19135,N_14715,N_18096);
and U19136 (N_19136,N_16250,N_15080);
nor U19137 (N_19137,N_17383,N_14211);
and U19138 (N_19138,N_17394,N_16225);
or U19139 (N_19139,N_15960,N_17800);
nor U19140 (N_19140,N_18123,N_13994);
or U19141 (N_19141,N_15260,N_13607);
nand U19142 (N_19142,N_18067,N_17503);
and U19143 (N_19143,N_12750,N_17161);
nand U19144 (N_19144,N_15323,N_16944);
and U19145 (N_19145,N_15734,N_14069);
or U19146 (N_19146,N_18471,N_16998);
and U19147 (N_19147,N_15551,N_14346);
nand U19148 (N_19148,N_13221,N_18597);
xnor U19149 (N_19149,N_16145,N_14557);
or U19150 (N_19150,N_13944,N_16021);
and U19151 (N_19151,N_17687,N_13143);
and U19152 (N_19152,N_17284,N_12603);
nand U19153 (N_19153,N_16353,N_16087);
xor U19154 (N_19154,N_15415,N_13593);
or U19155 (N_19155,N_17257,N_16397);
nor U19156 (N_19156,N_12866,N_17066);
nand U19157 (N_19157,N_16750,N_14896);
and U19158 (N_19158,N_16382,N_16224);
nor U19159 (N_19159,N_15246,N_18239);
and U19160 (N_19160,N_14445,N_14037);
and U19161 (N_19161,N_14662,N_14932);
nor U19162 (N_19162,N_14582,N_17852);
xor U19163 (N_19163,N_12569,N_13272);
and U19164 (N_19164,N_16173,N_13516);
or U19165 (N_19165,N_18043,N_13194);
or U19166 (N_19166,N_17375,N_18677);
or U19167 (N_19167,N_16700,N_17803);
and U19168 (N_19168,N_16726,N_18649);
nor U19169 (N_19169,N_16182,N_16672);
and U19170 (N_19170,N_14714,N_14001);
or U19171 (N_19171,N_14623,N_13203);
nor U19172 (N_19172,N_14820,N_18202);
nor U19173 (N_19173,N_18674,N_14160);
nor U19174 (N_19174,N_17740,N_13376);
nor U19175 (N_19175,N_17057,N_14140);
or U19176 (N_19176,N_14024,N_13744);
nor U19177 (N_19177,N_12749,N_16870);
nor U19178 (N_19178,N_13732,N_15820);
and U19179 (N_19179,N_16960,N_14260);
and U19180 (N_19180,N_14635,N_15801);
nand U19181 (N_19181,N_17568,N_14434);
or U19182 (N_19182,N_14919,N_15125);
and U19183 (N_19183,N_12774,N_12753);
nand U19184 (N_19184,N_12864,N_17050);
or U19185 (N_19185,N_13181,N_12784);
nand U19186 (N_19186,N_12960,N_17405);
and U19187 (N_19187,N_15467,N_18534);
or U19188 (N_19188,N_13809,N_12574);
nor U19189 (N_19189,N_15508,N_17718);
and U19190 (N_19190,N_14765,N_18475);
nor U19191 (N_19191,N_18099,N_17840);
and U19192 (N_19192,N_15736,N_16467);
or U19193 (N_19193,N_12503,N_14220);
nand U19194 (N_19194,N_13797,N_14194);
nand U19195 (N_19195,N_16482,N_14047);
xor U19196 (N_19196,N_13369,N_16856);
or U19197 (N_19197,N_17897,N_14040);
xnor U19198 (N_19198,N_13847,N_13610);
or U19199 (N_19199,N_18291,N_13751);
or U19200 (N_19200,N_17992,N_15615);
nand U19201 (N_19201,N_13305,N_15305);
or U19202 (N_19202,N_14508,N_17214);
and U19203 (N_19203,N_15037,N_13843);
nand U19204 (N_19204,N_15845,N_13908);
xnor U19205 (N_19205,N_14898,N_16806);
nor U19206 (N_19206,N_13836,N_14030);
nor U19207 (N_19207,N_15377,N_16056);
xnor U19208 (N_19208,N_18418,N_15204);
or U19209 (N_19209,N_17207,N_17918);
nor U19210 (N_19210,N_14275,N_18747);
or U19211 (N_19211,N_12615,N_14561);
nor U19212 (N_19212,N_16383,N_18643);
or U19213 (N_19213,N_18214,N_13148);
xnor U19214 (N_19214,N_17063,N_13668);
and U19215 (N_19215,N_14288,N_16133);
nand U19216 (N_19216,N_17456,N_13161);
and U19217 (N_19217,N_14648,N_17686);
and U19218 (N_19218,N_12521,N_14899);
nor U19219 (N_19219,N_17961,N_14034);
nor U19220 (N_19220,N_13256,N_15436);
nor U19221 (N_19221,N_14812,N_18684);
nor U19222 (N_19222,N_15170,N_17583);
nor U19223 (N_19223,N_13898,N_14629);
and U19224 (N_19224,N_12795,N_14416);
nand U19225 (N_19225,N_13813,N_15273);
or U19226 (N_19226,N_18729,N_16817);
or U19227 (N_19227,N_13964,N_18577);
or U19228 (N_19228,N_17730,N_18517);
or U19229 (N_19229,N_17737,N_14050);
xnor U19230 (N_19230,N_15883,N_18655);
or U19231 (N_19231,N_14705,N_12806);
nand U19232 (N_19232,N_12672,N_13504);
and U19233 (N_19233,N_15106,N_17201);
and U19234 (N_19234,N_15144,N_14636);
or U19235 (N_19235,N_12518,N_15525);
xor U19236 (N_19236,N_12600,N_14697);
or U19237 (N_19237,N_17424,N_14519);
or U19238 (N_19238,N_15331,N_18065);
or U19239 (N_19239,N_13499,N_17580);
and U19240 (N_19240,N_17612,N_17230);
nor U19241 (N_19241,N_15944,N_14783);
and U19242 (N_19242,N_16187,N_16269);
nand U19243 (N_19243,N_13228,N_13901);
xnor U19244 (N_19244,N_12862,N_18311);
or U19245 (N_19245,N_18319,N_15713);
and U19246 (N_19246,N_12760,N_13069);
nand U19247 (N_19247,N_14930,N_17373);
nor U19248 (N_19248,N_13515,N_13676);
nor U19249 (N_19249,N_15912,N_17039);
and U19250 (N_19250,N_18739,N_16600);
nand U19251 (N_19251,N_13864,N_13168);
or U19252 (N_19252,N_12638,N_17573);
and U19253 (N_19253,N_13793,N_12770);
xor U19254 (N_19254,N_17353,N_17912);
or U19255 (N_19255,N_17941,N_13823);
nor U19256 (N_19256,N_17262,N_15962);
nand U19257 (N_19257,N_18001,N_16943);
nor U19258 (N_19258,N_14720,N_14789);
nor U19259 (N_19259,N_17738,N_15963);
nand U19260 (N_19260,N_16566,N_18283);
xor U19261 (N_19261,N_15056,N_13429);
or U19262 (N_19262,N_18546,N_16996);
xor U19263 (N_19263,N_18250,N_16799);
or U19264 (N_19264,N_14532,N_15595);
nor U19265 (N_19265,N_16956,N_13414);
or U19266 (N_19266,N_17826,N_17308);
nor U19267 (N_19267,N_13252,N_16458);
or U19268 (N_19268,N_13582,N_15329);
and U19269 (N_19269,N_16696,N_14860);
and U19270 (N_19270,N_13881,N_13658);
xnor U19271 (N_19271,N_16675,N_14481);
or U19272 (N_19272,N_18690,N_18669);
and U19273 (N_19273,N_14118,N_15955);
nand U19274 (N_19274,N_17863,N_16140);
and U19275 (N_19275,N_13631,N_17111);
or U19276 (N_19276,N_15318,N_14926);
xor U19277 (N_19277,N_18092,N_17810);
or U19278 (N_19278,N_15268,N_13359);
nand U19279 (N_19279,N_17540,N_16935);
nor U19280 (N_19280,N_16110,N_13636);
or U19281 (N_19281,N_12520,N_16013);
nor U19282 (N_19282,N_14217,N_13723);
and U19283 (N_19283,N_18222,N_13402);
and U19284 (N_19284,N_17652,N_14493);
and U19285 (N_19285,N_14684,N_13132);
nand U19286 (N_19286,N_12705,N_15126);
nor U19287 (N_19287,N_12568,N_15243);
xnor U19288 (N_19288,N_13893,N_16814);
or U19289 (N_19289,N_13192,N_17126);
or U19290 (N_19290,N_17250,N_15477);
and U19291 (N_19291,N_16737,N_18432);
and U19292 (N_19292,N_13463,N_15614);
or U19293 (N_19293,N_13053,N_12531);
or U19294 (N_19294,N_17648,N_14384);
xor U19295 (N_19295,N_18733,N_18197);
xor U19296 (N_19296,N_17981,N_16387);
and U19297 (N_19297,N_17881,N_14270);
or U19298 (N_19298,N_18343,N_17120);
or U19299 (N_19299,N_12613,N_16275);
or U19300 (N_19300,N_17229,N_18696);
or U19301 (N_19301,N_17119,N_15599);
and U19302 (N_19302,N_17898,N_14403);
nor U19303 (N_19303,N_15873,N_14660);
nand U19304 (N_19304,N_18424,N_16957);
nor U19305 (N_19305,N_13498,N_17462);
nand U19306 (N_19306,N_18497,N_12676);
nand U19307 (N_19307,N_15441,N_17631);
and U19308 (N_19308,N_15874,N_14150);
nor U19309 (N_19309,N_12827,N_13206);
nand U19310 (N_19310,N_14548,N_14023);
and U19311 (N_19311,N_13946,N_18500);
nand U19312 (N_19312,N_16311,N_15102);
xor U19313 (N_19313,N_15973,N_14039);
nor U19314 (N_19314,N_17069,N_14967);
nand U19315 (N_19315,N_17085,N_17427);
and U19316 (N_19316,N_14183,N_14805);
nand U19317 (N_19317,N_17216,N_16130);
nor U19318 (N_19318,N_16999,N_14421);
or U19319 (N_19319,N_17885,N_13986);
and U19320 (N_19320,N_18213,N_18504);
or U19321 (N_19321,N_14394,N_14020);
and U19322 (N_19322,N_16838,N_16554);
or U19323 (N_19323,N_14296,N_14337);
and U19324 (N_19324,N_15096,N_13887);
or U19325 (N_19325,N_15989,N_12607);
or U19326 (N_19326,N_15888,N_16717);
nand U19327 (N_19327,N_15811,N_17932);
and U19328 (N_19328,N_13454,N_15290);
or U19329 (N_19329,N_17679,N_15731);
and U19330 (N_19330,N_16898,N_14165);
or U19331 (N_19331,N_15741,N_12636);
and U19332 (N_19332,N_17339,N_13083);
nand U19333 (N_19333,N_17564,N_18245);
xor U19334 (N_19334,N_18467,N_17246);
nor U19335 (N_19335,N_16568,N_14506);
nor U19336 (N_19336,N_16280,N_15864);
nor U19337 (N_19337,N_14910,N_14960);
nand U19338 (N_19338,N_12831,N_18592);
nand U19339 (N_19339,N_13496,N_12930);
nor U19340 (N_19340,N_18523,N_14524);
nor U19341 (N_19341,N_12654,N_16851);
and U19342 (N_19342,N_12646,N_13654);
nor U19343 (N_19343,N_14036,N_12602);
and U19344 (N_19344,N_12819,N_18128);
nor U19345 (N_19345,N_14311,N_17887);
and U19346 (N_19346,N_15700,N_14656);
or U19347 (N_19347,N_16435,N_17286);
or U19348 (N_19348,N_13895,N_15407);
xor U19349 (N_19349,N_14488,N_13630);
nor U19350 (N_19350,N_18292,N_14567);
and U19351 (N_19351,N_14252,N_16012);
nand U19352 (N_19352,N_18720,N_13472);
nand U19353 (N_19353,N_15740,N_14502);
nor U19354 (N_19354,N_14515,N_15294);
nor U19355 (N_19355,N_16432,N_12648);
nor U19356 (N_19356,N_12659,N_17672);
and U19357 (N_19357,N_12519,N_17166);
nand U19358 (N_19358,N_18035,N_18687);
nor U19359 (N_19359,N_14829,N_14573);
nand U19360 (N_19360,N_12582,N_15770);
nand U19361 (N_19361,N_18585,N_18376);
nand U19362 (N_19362,N_15891,N_16112);
xnor U19363 (N_19363,N_13233,N_14111);
nand U19364 (N_19364,N_15123,N_13012);
and U19365 (N_19365,N_13344,N_15113);
and U19366 (N_19366,N_17049,N_15031);
xor U19367 (N_19367,N_17504,N_14376);
or U19368 (N_19368,N_15751,N_17096);
nor U19369 (N_19369,N_17688,N_18505);
or U19370 (N_19370,N_12814,N_14465);
and U19371 (N_19371,N_17408,N_13277);
xor U19372 (N_19372,N_16230,N_12740);
xnor U19373 (N_19373,N_15342,N_14227);
or U19374 (N_19374,N_18070,N_13777);
nor U19375 (N_19375,N_12619,N_16175);
nor U19376 (N_19376,N_12861,N_13858);
or U19377 (N_19377,N_15369,N_14633);
xor U19378 (N_19378,N_18647,N_12908);
and U19379 (N_19379,N_14203,N_16354);
or U19380 (N_19380,N_13989,N_18403);
or U19381 (N_19381,N_15471,N_17582);
nand U19382 (N_19382,N_15292,N_15371);
and U19383 (N_19383,N_13442,N_13099);
nor U19384 (N_19384,N_16135,N_18396);
and U19385 (N_19385,N_17235,N_15593);
nor U19386 (N_19386,N_13200,N_14531);
nand U19387 (N_19387,N_15698,N_12957);
nand U19388 (N_19388,N_13304,N_16739);
or U19389 (N_19389,N_14338,N_12911);
and U19390 (N_19390,N_17756,N_13664);
or U19391 (N_19391,N_18653,N_18435);
nor U19392 (N_19392,N_14969,N_16653);
or U19393 (N_19393,N_13320,N_12982);
or U19394 (N_19394,N_18678,N_14102);
nor U19395 (N_19395,N_12946,N_18727);
nand U19396 (N_19396,N_15908,N_17683);
or U19397 (N_19397,N_13583,N_17989);
nor U19398 (N_19398,N_14343,N_14297);
and U19399 (N_19399,N_13212,N_17575);
xor U19400 (N_19400,N_13348,N_14599);
nand U19401 (N_19401,N_18086,N_16229);
nand U19402 (N_19402,N_17919,N_17194);
or U19403 (N_19403,N_18390,N_16614);
nand U19404 (N_19404,N_13990,N_13837);
nand U19405 (N_19405,N_13670,N_12560);
or U19406 (N_19406,N_16549,N_17761);
or U19407 (N_19407,N_16000,N_17592);
or U19408 (N_19408,N_16732,N_18509);
nor U19409 (N_19409,N_16363,N_14830);
xor U19410 (N_19410,N_14486,N_13537);
nor U19411 (N_19411,N_14166,N_14827);
nor U19412 (N_19412,N_16002,N_18131);
and U19413 (N_19413,N_14494,N_12651);
nor U19414 (N_19414,N_12748,N_16901);
nor U19415 (N_19415,N_12859,N_15732);
nand U19416 (N_19416,N_14565,N_17259);
or U19417 (N_19417,N_13931,N_12544);
and U19418 (N_19418,N_12756,N_16470);
and U19419 (N_19419,N_17929,N_17939);
nand U19420 (N_19420,N_17179,N_16001);
nor U19421 (N_19421,N_17107,N_17620);
and U19422 (N_19422,N_16613,N_18541);
nand U19423 (N_19423,N_15915,N_18529);
nor U19424 (N_19424,N_15494,N_16678);
or U19425 (N_19425,N_17028,N_14157);
and U19426 (N_19426,N_14627,N_16810);
nor U19427 (N_19427,N_14836,N_15703);
nand U19428 (N_19428,N_15299,N_18410);
or U19429 (N_19429,N_17864,N_16924);
and U19430 (N_19430,N_14612,N_14630);
or U19431 (N_19431,N_14756,N_16243);
nor U19432 (N_19432,N_18062,N_17947);
nor U19433 (N_19433,N_16667,N_18562);
and U19434 (N_19434,N_15604,N_16350);
nor U19435 (N_19435,N_13642,N_17397);
nor U19436 (N_19436,N_12673,N_16584);
nor U19437 (N_19437,N_14269,N_17358);
nor U19438 (N_19438,N_18635,N_16647);
and U19439 (N_19439,N_18146,N_15300);
or U19440 (N_19440,N_13166,N_16859);
or U19441 (N_19441,N_17530,N_14852);
nor U19442 (N_19442,N_16892,N_17835);
xnor U19443 (N_19443,N_12789,N_16265);
and U19444 (N_19444,N_18459,N_17117);
and U19445 (N_19445,N_15868,N_15520);
and U19446 (N_19446,N_15169,N_15195);
nand U19447 (N_19447,N_12951,N_18153);
and U19448 (N_19448,N_17956,N_18281);
and U19449 (N_19449,N_18411,N_14226);
nor U19450 (N_19450,N_17790,N_16058);
and U19451 (N_19451,N_15493,N_14702);
nor U19452 (N_19452,N_18434,N_15328);
and U19453 (N_19453,N_16037,N_16020);
xor U19454 (N_19454,N_14174,N_14334);
nor U19455 (N_19455,N_16791,N_13919);
nand U19456 (N_19456,N_18371,N_18265);
nand U19457 (N_19457,N_17859,N_16188);
nand U19458 (N_19458,N_16946,N_12849);
nor U19459 (N_19459,N_18014,N_16171);
nor U19460 (N_19460,N_17949,N_15245);
and U19461 (N_19461,N_14008,N_15310);
xor U19462 (N_19462,N_12885,N_17153);
xnor U19463 (N_19463,N_16590,N_16226);
nand U19464 (N_19464,N_14315,N_18470);
or U19465 (N_19465,N_13488,N_17704);
or U19466 (N_19466,N_18700,N_16940);
nor U19467 (N_19467,N_17432,N_13478);
and U19468 (N_19468,N_14539,N_17567);
and U19469 (N_19469,N_13175,N_13408);
or U19470 (N_19470,N_18667,N_16864);
nor U19471 (N_19471,N_16821,N_16503);
nand U19472 (N_19472,N_13721,N_13546);
and U19473 (N_19473,N_16612,N_13955);
nand U19474 (N_19474,N_15913,N_14396);
xor U19475 (N_19475,N_12830,N_12797);
nor U19476 (N_19476,N_15898,N_14098);
nor U19477 (N_19477,N_13671,N_12668);
and U19478 (N_19478,N_16564,N_16830);
nor U19479 (N_19479,N_13090,N_17382);
nand U19480 (N_19480,N_16463,N_12853);
or U19481 (N_19481,N_16074,N_17491);
or U19482 (N_19482,N_13198,N_16661);
xnor U19483 (N_19483,N_16579,N_18416);
xor U19484 (N_19484,N_15259,N_18712);
or U19485 (N_19485,N_14634,N_15188);
nand U19486 (N_19486,N_13960,N_18383);
and U19487 (N_19487,N_13441,N_18083);
nand U19488 (N_19488,N_15336,N_14904);
nand U19489 (N_19489,N_14119,N_16891);
or U19490 (N_19490,N_13363,N_13071);
and U19491 (N_19491,N_17073,N_12649);
nand U19492 (N_19492,N_13860,N_13918);
xnor U19493 (N_19493,N_16276,N_18478);
nor U19494 (N_19494,N_14834,N_16580);
and U19495 (N_19495,N_17041,N_13355);
or U19496 (N_19496,N_17974,N_15724);
nand U19497 (N_19497,N_17130,N_18032);
or U19498 (N_19498,N_18661,N_17935);
nand U19499 (N_19499,N_17199,N_16518);
or U19500 (N_19500,N_16493,N_16158);
and U19501 (N_19501,N_12639,N_18135);
nand U19502 (N_19502,N_17651,N_13468);
or U19503 (N_19503,N_18149,N_13406);
nand U19504 (N_19504,N_13398,N_14867);
nand U19505 (N_19505,N_14122,N_13137);
nor U19506 (N_19506,N_15399,N_15889);
and U19507 (N_19507,N_17831,N_14868);
nor U19508 (N_19508,N_15910,N_16362);
nand U19509 (N_19509,N_16778,N_15951);
or U19510 (N_19510,N_15696,N_14761);
nand U19511 (N_19511,N_15117,N_13209);
nand U19512 (N_19512,N_14062,N_12792);
or U19513 (N_19513,N_14431,N_12576);
nor U19514 (N_19514,N_17888,N_12884);
nor U19515 (N_19515,N_14233,N_18602);
xnor U19516 (N_19516,N_16308,N_13033);
nor U19517 (N_19517,N_16958,N_14439);
xnor U19518 (N_19518,N_16050,N_15150);
and U19519 (N_19519,N_18732,N_14741);
nor U19520 (N_19520,N_16156,N_17816);
nor U19521 (N_19521,N_17600,N_18482);
or U19522 (N_19522,N_12936,N_13993);
or U19523 (N_19523,N_13412,N_13810);
and U19524 (N_19524,N_12691,N_12675);
xnor U19525 (N_19525,N_14428,N_15390);
and U19526 (N_19526,N_18439,N_16460);
xor U19527 (N_19527,N_15076,N_18218);
nor U19528 (N_19528,N_16023,N_16234);
or U19529 (N_19529,N_17355,N_14198);
or U19530 (N_19530,N_13952,N_13643);
xor U19531 (N_19531,N_17396,N_13530);
nand U19532 (N_19532,N_15681,N_18261);
xor U19533 (N_19533,N_16095,N_14264);
nand U19534 (N_19534,N_12899,N_17765);
or U19535 (N_19535,N_15417,N_16302);
nand U19536 (N_19536,N_16742,N_17055);
xor U19537 (N_19537,N_15357,N_16858);
nor U19538 (N_19538,N_18468,N_16962);
or U19539 (N_19539,N_12664,N_16333);
or U19540 (N_19540,N_15119,N_15976);
or U19541 (N_19541,N_13329,N_15549);
or U19542 (N_19542,N_12935,N_16202);
nand U19543 (N_19543,N_13002,N_18172);
or U19544 (N_19544,N_14282,N_14213);
or U19545 (N_19545,N_17589,N_16809);
and U19546 (N_19546,N_18412,N_16212);
or U19547 (N_19547,N_15376,N_18594);
or U19548 (N_19548,N_17186,N_18249);
nor U19549 (N_19549,N_16866,N_15836);
nor U19550 (N_19550,N_16862,N_15443);
nand U19551 (N_19551,N_14951,N_15013);
nand U19552 (N_19552,N_17030,N_15695);
or U19553 (N_19553,N_18129,N_15532);
and U19554 (N_19554,N_16118,N_12837);
or U19555 (N_19555,N_15291,N_13015);
nor U19556 (N_19556,N_14616,N_17502);
and U19557 (N_19557,N_16649,N_15680);
nor U19558 (N_19558,N_16978,N_14327);
nand U19559 (N_19559,N_14792,N_13559);
or U19560 (N_19560,N_15629,N_16753);
nor U19561 (N_19561,N_17520,N_13360);
or U19562 (N_19562,N_17832,N_13681);
nor U19563 (N_19563,N_12847,N_12637);
or U19564 (N_19564,N_14075,N_17998);
and U19565 (N_19565,N_18422,N_16168);
and U19566 (N_19566,N_16920,N_14496);
xnor U19567 (N_19567,N_15237,N_15000);
or U19568 (N_19568,N_13086,N_13700);
and U19569 (N_19569,N_18484,N_14128);
or U19570 (N_19570,N_14840,N_18104);
or U19571 (N_19571,N_12800,N_16701);
and U19572 (N_19572,N_12726,N_17033);
nor U19573 (N_19573,N_15226,N_15842);
nand U19574 (N_19574,N_12852,N_14551);
or U19575 (N_19575,N_17678,N_13817);
nor U19576 (N_19576,N_16075,N_16401);
and U19577 (N_19577,N_16239,N_18317);
nand U19578 (N_19578,N_16900,N_16835);
and U19579 (N_19579,N_13174,N_16261);
nor U19580 (N_19580,N_17276,N_16066);
nor U19581 (N_19581,N_13426,N_14619);
or U19582 (N_19582,N_17302,N_13746);
or U19583 (N_19583,N_16668,N_18454);
nor U19584 (N_19584,N_15200,N_12895);
and U19585 (N_19585,N_15312,N_14755);
nor U19586 (N_19586,N_12702,N_15781);
nor U19587 (N_19587,N_14887,N_17127);
and U19588 (N_19588,N_15430,N_14713);
nor U19589 (N_19589,N_13465,N_18028);
nand U19590 (N_19590,N_14212,N_16637);
or U19591 (N_19591,N_13353,N_17846);
nor U19592 (N_19592,N_14683,N_15896);
nand U19593 (N_19593,N_13970,N_13669);
nand U19594 (N_19594,N_13997,N_16088);
nand U19595 (N_19595,N_15737,N_15216);
nand U19596 (N_19596,N_18564,N_14240);
or U19597 (N_19597,N_18109,N_17708);
or U19598 (N_19598,N_18474,N_18324);
nor U19599 (N_19599,N_13509,N_15401);
and U19600 (N_19600,N_14536,N_16046);
or U19601 (N_19601,N_18621,N_18107);
nor U19602 (N_19602,N_17591,N_15049);
nand U19603 (N_19603,N_15902,N_12657);
xnor U19604 (N_19604,N_17087,N_12515);
xor U19605 (N_19605,N_16301,N_15872);
and U19606 (N_19606,N_16104,N_13122);
or U19607 (N_19607,N_16405,N_14793);
and U19608 (N_19608,N_15182,N_15991);
nor U19609 (N_19609,N_15067,N_17008);
nand U19610 (N_19610,N_13767,N_13757);
nand U19611 (N_19611,N_17484,N_18262);
nand U19612 (N_19612,N_15573,N_15887);
nand U19613 (N_19613,N_13151,N_13794);
nand U19614 (N_19614,N_14382,N_12977);
or U19615 (N_19615,N_16258,N_14664);
and U19616 (N_19616,N_13638,N_15324);
nor U19617 (N_19617,N_13566,N_14610);
or U19618 (N_19618,N_17658,N_14205);
nor U19619 (N_19619,N_17979,N_14722);
nand U19620 (N_19620,N_13113,N_17112);
and U19621 (N_19621,N_14358,N_13597);
nor U19622 (N_19622,N_15363,N_14833);
or U19623 (N_19623,N_14955,N_16407);
and U19624 (N_19624,N_18464,N_17335);
nor U19625 (N_19625,N_14942,N_12721);
or U19626 (N_19626,N_14738,N_15322);
nor U19627 (N_19627,N_17412,N_16936);
and U19628 (N_19628,N_16436,N_13024);
and U19629 (N_19629,N_17926,N_17438);
xor U19630 (N_19630,N_12561,N_17879);
or U19631 (N_19631,N_17793,N_16219);
or U19632 (N_19632,N_13666,N_15319);
and U19633 (N_19633,N_16323,N_14339);
xnor U19634 (N_19634,N_18047,N_18743);
nor U19635 (N_19635,N_16062,N_14920);
and U19636 (N_19636,N_16697,N_18040);
and U19637 (N_19637,N_14608,N_13387);
xor U19638 (N_19638,N_15621,N_14499);
or U19639 (N_19639,N_13786,N_13127);
nor U19640 (N_19640,N_12658,N_17071);
or U19641 (N_19641,N_17758,N_18734);
nand U19642 (N_19642,N_14590,N_18611);
nand U19643 (N_19643,N_14647,N_15772);
xor U19644 (N_19644,N_17392,N_16921);
and U19645 (N_19645,N_18537,N_15679);
nor U19646 (N_19646,N_15211,N_16380);
nor U19647 (N_19647,N_18589,N_12967);
nand U19648 (N_19648,N_14751,N_17917);
and U19649 (N_19649,N_16752,N_13357);
nand U19650 (N_19650,N_17518,N_17723);
nor U19651 (N_19651,N_17411,N_14440);
nor U19652 (N_19652,N_14734,N_13706);
nand U19653 (N_19653,N_17588,N_15884);
nand U19654 (N_19654,N_13243,N_12924);
nand U19655 (N_19655,N_17091,N_17054);
or U19656 (N_19656,N_12845,N_12807);
nand U19657 (N_19657,N_17043,N_17548);
and U19658 (N_19658,N_18741,N_18366);
nand U19659 (N_19659,N_17210,N_13147);
nand U19660 (N_19660,N_15277,N_13924);
and U19661 (N_19661,N_16628,N_15610);
and U19662 (N_19662,N_16536,N_18614);
or U19663 (N_19663,N_18305,N_13743);
nor U19664 (N_19664,N_18607,N_14710);
or U19665 (N_19665,N_14719,N_12501);
nor U19666 (N_19666,N_18193,N_15950);
and U19667 (N_19667,N_18034,N_17381);
nand U19668 (N_19668,N_18391,N_17170);
and U19669 (N_19669,N_16242,N_16833);
or U19670 (N_19670,N_15057,N_13226);
or U19671 (N_19671,N_18736,N_14175);
and U19672 (N_19672,N_17819,N_16671);
nor U19673 (N_19673,N_15225,N_17850);
and U19674 (N_19674,N_16636,N_13384);
nor U19675 (N_19675,N_12542,N_16552);
and U19676 (N_19676,N_12666,N_16933);
or U19677 (N_19677,N_12707,N_15032);
or U19678 (N_19678,N_14426,N_13423);
nand U19679 (N_19679,N_14709,N_12509);
or U19680 (N_19680,N_16530,N_12736);
or U19681 (N_19681,N_16896,N_13066);
xnor U19682 (N_19682,N_18356,N_13156);
nor U19683 (N_19683,N_17597,N_14556);
nor U19684 (N_19684,N_13018,N_17643);
nand U19685 (N_19685,N_18636,N_16873);
xnor U19686 (N_19686,N_13808,N_14293);
or U19687 (N_19687,N_15009,N_17025);
nor U19688 (N_19688,N_16259,N_13892);
nand U19689 (N_19689,N_15209,N_16581);
nor U19690 (N_19690,N_17663,N_17559);
nand U19691 (N_19691,N_15488,N_18691);
nor U19692 (N_19692,N_17856,N_16277);
and U19693 (N_19693,N_12988,N_17042);
nor U19694 (N_19694,N_18155,N_17627);
nor U19695 (N_19695,N_16228,N_17245);
nor U19696 (N_19696,N_15254,N_13351);
and U19697 (N_19697,N_17366,N_17806);
or U19698 (N_19698,N_13199,N_18746);
nand U19699 (N_19699,N_18519,N_14822);
nand U19700 (N_19700,N_14858,N_13840);
nand U19701 (N_19701,N_16131,N_13133);
nand U19702 (N_19702,N_12516,N_14247);
and U19703 (N_19703,N_18157,N_17351);
nor U19704 (N_19704,N_17895,N_15244);
nor U19705 (N_19705,N_18730,N_12902);
nand U19706 (N_19706,N_17247,N_18133);
or U19707 (N_19707,N_14448,N_13685);
and U19708 (N_19708,N_15507,N_14229);
nand U19709 (N_19709,N_13755,N_18413);
nor U19710 (N_19710,N_17637,N_16378);
nor U19711 (N_19711,N_16715,N_13974);
nand U19712 (N_19712,N_16599,N_13812);
nor U19713 (N_19713,N_16914,N_13819);
and U19714 (N_19714,N_14864,N_15256);
or U19715 (N_19715,N_15373,N_13068);
xor U19716 (N_19716,N_12912,N_16142);
nor U19717 (N_19717,N_17930,N_14094);
xnor U19718 (N_19718,N_15397,N_15414);
and U19719 (N_19719,N_15952,N_16278);
nor U19720 (N_19720,N_13640,N_15085);
nand U19721 (N_19721,N_17626,N_17717);
or U19722 (N_19722,N_16744,N_15082);
nor U19723 (N_19723,N_18340,N_17691);
nand U19724 (N_19724,N_17249,N_14678);
nand U19725 (N_19725,N_14894,N_17855);
or U19726 (N_19726,N_15235,N_12905);
or U19727 (N_19727,N_15124,N_12886);
nand U19728 (N_19728,N_18326,N_15575);
and U19729 (N_19729,N_15337,N_14609);
or U19730 (N_19730,N_16808,N_13238);
and U19731 (N_19731,N_14380,N_13644);
xor U19732 (N_19732,N_13857,N_14744);
xnor U19733 (N_19733,N_14430,N_13169);
nand U19734 (N_19734,N_17797,N_17434);
nor U19735 (N_19735,N_14335,N_13328);
or U19736 (N_19736,N_14255,N_17490);
nor U19737 (N_19737,N_14588,N_18055);
or U19738 (N_19738,N_17270,N_16231);
or U19739 (N_19739,N_13848,N_17051);
nand U19740 (N_19740,N_18363,N_16251);
nand U19741 (N_19741,N_16026,N_17880);
or U19742 (N_19742,N_12712,N_17177);
nor U19743 (N_19743,N_18278,N_13190);
or U19744 (N_19744,N_18540,N_14404);
xor U19745 (N_19745,N_16949,N_16334);
nor U19746 (N_19746,N_18042,N_16850);
or U19747 (N_19747,N_15227,N_13310);
or U19748 (N_19748,N_17313,N_18255);
or U19749 (N_19749,N_15596,N_13279);
nor U19750 (N_19750,N_14958,N_16880);
nor U19751 (N_19751,N_16139,N_14594);
xnor U19752 (N_19752,N_15925,N_17759);
nand U19753 (N_19753,N_17791,N_12923);
nand U19754 (N_19754,N_12662,N_13822);
nand U19755 (N_19755,N_18241,N_13788);
xor U19756 (N_19756,N_18584,N_17613);
or U19757 (N_19757,N_16151,N_16108);
or U19758 (N_19758,N_15878,N_16049);
or U19759 (N_19759,N_17618,N_13250);
and U19760 (N_19760,N_12713,N_15047);
nor U19761 (N_19761,N_16420,N_15608);
or U19762 (N_19762,N_12949,N_15034);
or U19763 (N_19763,N_16326,N_15784);
nand U19764 (N_19764,N_13569,N_16123);
or U19765 (N_19765,N_14791,N_13626);
and U19766 (N_19766,N_14015,N_16674);
nor U19767 (N_19767,N_16419,N_12865);
or U19768 (N_19768,N_17047,N_16938);
xnor U19769 (N_19769,N_14658,N_13052);
xor U19770 (N_19770,N_13326,N_14862);
nand U19771 (N_19771,N_14031,N_15191);
nand U19772 (N_19772,N_15626,N_17391);
or U19773 (N_19773,N_17384,N_17016);
or U19774 (N_19774,N_13467,N_13409);
nor U19775 (N_19775,N_15974,N_13267);
and U19776 (N_19776,N_12548,N_15546);
or U19777 (N_19777,N_12892,N_12536);
nand U19778 (N_19778,N_15624,N_17338);
or U19779 (N_19779,N_17328,N_14103);
or U19780 (N_19780,N_14313,N_16680);
nor U19781 (N_19781,N_13183,N_18685);
nor U19782 (N_19782,N_13098,N_15073);
and U19783 (N_19783,N_16592,N_15086);
nor U19784 (N_19784,N_18276,N_15675);
and U19785 (N_19785,N_17124,N_12644);
or U19786 (N_19786,N_12985,N_17004);
nand U19787 (N_19787,N_16486,N_12627);
xnor U19788 (N_19788,N_18722,N_14088);
nor U19789 (N_19789,N_16792,N_13832);
and U19790 (N_19790,N_17928,N_12818);
nand U19791 (N_19791,N_12510,N_17332);
xor U19792 (N_19792,N_14724,N_15416);
and U19793 (N_19793,N_17345,N_18210);
nand U19794 (N_19794,N_15899,N_13807);
nor U19795 (N_19795,N_13367,N_13158);
and U19796 (N_19796,N_12863,N_13999);
or U19797 (N_19797,N_16059,N_15958);
nand U19798 (N_19798,N_17632,N_17489);
nor U19799 (N_19799,N_14818,N_13694);
xnor U19800 (N_19800,N_12926,N_17842);
nand U19801 (N_19801,N_17181,N_16515);
xor U19802 (N_19802,N_12717,N_13780);
and U19803 (N_19803,N_14129,N_15646);
and U19804 (N_19804,N_17886,N_17779);
nand U19805 (N_19805,N_12771,N_18694);
and U19806 (N_19806,N_13049,N_13430);
and U19807 (N_19807,N_14676,N_17533);
nand U19808 (N_19808,N_18103,N_18665);
and U19809 (N_19809,N_14613,N_17144);
nand U19810 (N_19810,N_16665,N_14984);
xnor U19811 (N_19811,N_16106,N_17553);
and U19812 (N_19812,N_15431,N_16588);
or U19813 (N_19813,N_16626,N_13007);
nand U19814 (N_19814,N_14018,N_14273);
nor U19815 (N_19815,N_15411,N_16450);
and U19816 (N_19816,N_14491,N_13332);
nor U19817 (N_19817,N_16452,N_12987);
and U19818 (N_19818,N_18302,N_14801);
nand U19819 (N_19819,N_13259,N_15987);
or U19820 (N_19820,N_17344,N_14891);
nand U19821 (N_19821,N_13146,N_15714);
or U19822 (N_19822,N_15387,N_15025);
nand U19823 (N_19823,N_16312,N_17607);
nor U19824 (N_19824,N_17221,N_14929);
and U19825 (N_19825,N_18518,N_13884);
or U19826 (N_19826,N_13536,N_16611);
nand U19827 (N_19827,N_12931,N_16617);
and U19828 (N_19828,N_17138,N_15535);
and U19829 (N_19829,N_18634,N_12759);
nand U19830 (N_19830,N_15293,N_16517);
nor U19831 (N_19831,N_16124,N_14522);
nor U19832 (N_19832,N_12526,N_15617);
and U19833 (N_19833,N_13600,N_15006);
and U19834 (N_19834,N_12720,N_15749);
and U19835 (N_19835,N_18524,N_13701);
or U19836 (N_19836,N_17727,N_12858);
or U19837 (N_19837,N_15903,N_16400);
nand U19838 (N_19838,N_15867,N_12874);
and U19839 (N_19839,N_14503,N_17496);
nor U19840 (N_19840,N_17224,N_17773);
and U19841 (N_19841,N_14135,N_16698);
or U19842 (N_19842,N_14068,N_15540);
or U19843 (N_19843,N_17668,N_13801);
nor U19844 (N_19844,N_15070,N_16472);
xnor U19845 (N_19845,N_14529,N_14562);
nor U19846 (N_19846,N_17515,N_16874);
nor U19847 (N_19847,N_15093,N_18009);
xnor U19848 (N_19848,N_12642,N_17958);
nor U19849 (N_19849,N_17056,N_13244);
nand U19850 (N_19850,N_15909,N_17955);
and U19851 (N_19851,N_18152,N_16349);
and U19852 (N_19852,N_16966,N_12690);
nand U19853 (N_19853,N_13234,N_16961);
nor U19854 (N_19854,N_15658,N_16129);
nor U19855 (N_19855,N_14237,N_15861);
xor U19856 (N_19856,N_17367,N_16240);
and U19857 (N_19857,N_15107,N_16320);
xor U19858 (N_19858,N_14976,N_16338);
nand U19859 (N_19859,N_16381,N_15601);
and U19860 (N_19860,N_17029,N_17682);
nand U19861 (N_19861,N_15652,N_16783);
nor U19862 (N_19862,N_16114,N_18718);
nor U19863 (N_19863,N_17093,N_16428);
and U19864 (N_19864,N_14438,N_18121);
nor U19865 (N_19865,N_14033,N_14201);
or U19866 (N_19866,N_15327,N_15816);
nand U19867 (N_19867,N_12963,N_13781);
xor U19868 (N_19868,N_13916,N_14994);
nand U19869 (N_19869,N_13686,N_16080);
nand U19870 (N_19870,N_18393,N_14152);
or U19871 (N_19871,N_15270,N_13769);
and U19872 (N_19872,N_14185,N_17892);
and U19873 (N_19873,N_15452,N_18496);
and U19874 (N_19874,N_12975,N_18745);
and U19875 (N_19875,N_15876,N_18171);
or U19876 (N_19876,N_13561,N_13521);
or U19877 (N_19877,N_13620,N_18731);
nand U19878 (N_19878,N_12878,N_14726);
and U19879 (N_19879,N_12981,N_14089);
nor U19880 (N_19880,N_14195,N_12781);
nand U19881 (N_19881,N_18078,N_15653);
and U19882 (N_19882,N_17699,N_16684);
and U19883 (N_19883,N_15386,N_16221);
or U19884 (N_19884,N_17629,N_14704);
nand U19885 (N_19885,N_17468,N_16213);
nor U19886 (N_19886,N_12998,N_18060);
xnor U19887 (N_19887,N_16994,N_14196);
or U19888 (N_19888,N_13982,N_12527);
and U19889 (N_19889,N_14184,N_13040);
and U19890 (N_19890,N_17363,N_12743);
nand U19891 (N_19891,N_17536,N_13759);
nor U19892 (N_19892,N_15185,N_14618);
or U19893 (N_19893,N_14952,N_12643);
nor U19894 (N_19894,N_15359,N_15656);
nand U19895 (N_19895,N_17298,N_18349);
or U19896 (N_19896,N_18705,N_18138);
nand U19897 (N_19897,N_15449,N_15236);
nor U19898 (N_19898,N_14222,N_15099);
xnor U19899 (N_19899,N_13301,N_16306);
or U19900 (N_19900,N_16556,N_18480);
nor U19901 (N_19901,N_16502,N_16073);
and U19902 (N_19902,N_14280,N_18348);
nor U19903 (N_19903,N_16069,N_17675);
nand U19904 (N_19904,N_17755,N_16141);
nand U19905 (N_19905,N_14093,N_13863);
and U19906 (N_19906,N_18384,N_13574);
nor U19907 (N_19907,N_18120,N_14693);
nor U19908 (N_19908,N_14407,N_13422);
nand U19909 (N_19909,N_17354,N_16784);
and U19910 (N_19910,N_14090,N_16036);
nand U19911 (N_19911,N_17499,N_17007);
nand U19912 (N_19912,N_13347,N_14302);
or U19913 (N_19913,N_18728,N_15159);
nand U19914 (N_19914,N_17614,N_16487);
nor U19915 (N_19915,N_16722,N_17125);
nor U19916 (N_19916,N_14853,N_16262);
nor U19917 (N_19917,N_14372,N_16341);
nand U19918 (N_19918,N_16218,N_17398);
nand U19919 (N_19919,N_15691,N_14585);
and U19920 (N_19920,N_15611,N_16386);
and U19921 (N_19921,N_16909,N_16053);
and U19922 (N_19922,N_16760,N_14243);
nand U19923 (N_19923,N_14516,N_13361);
xor U19924 (N_19924,N_17774,N_13874);
xnor U19925 (N_19925,N_15859,N_14624);
or U19926 (N_19926,N_17839,N_12922);
or U19927 (N_19927,N_14168,N_17197);
xor U19928 (N_19928,N_13573,N_12572);
nor U19929 (N_19929,N_17822,N_14182);
or U19930 (N_19930,N_15483,N_14146);
nor U19931 (N_19931,N_13032,N_16247);
and U19932 (N_19932,N_16915,N_16842);
xor U19933 (N_19933,N_13586,N_15269);
or U19934 (N_19934,N_13641,N_13920);
xor U19935 (N_19935,N_14193,N_17967);
or U19936 (N_19936,N_12699,N_17265);
or U19937 (N_19937,N_14048,N_13967);
and U19938 (N_19938,N_13439,N_12671);
or U19939 (N_19939,N_14079,N_17190);
nand U19940 (N_19940,N_18227,N_14289);
nor U19941 (N_19941,N_17454,N_18441);
nand U19942 (N_19942,N_17322,N_16937);
and U19943 (N_19943,N_15907,N_13101);
nor U19944 (N_19944,N_18414,N_14559);
nor U19945 (N_19945,N_13108,N_13987);
nand U19946 (N_19946,N_14995,N_14785);
or U19947 (N_19947,N_16090,N_18050);
xor U19948 (N_19948,N_15664,N_13214);
nand U19949 (N_19949,N_17198,N_18186);
and U19950 (N_19950,N_18641,N_18100);
or U19951 (N_19951,N_16208,N_16899);
nand U19952 (N_19952,N_13268,N_14272);
nor U19953 (N_19953,N_14393,N_15383);
nand U19954 (N_19954,N_14148,N_15935);
or U19955 (N_19955,N_14305,N_18220);
nor U19956 (N_19956,N_17379,N_15400);
or U19957 (N_19957,N_15828,N_14758);
and U19958 (N_19958,N_15311,N_18080);
nor U19959 (N_19959,N_18098,N_12934);
nand U19960 (N_19960,N_17472,N_16010);
and U19961 (N_19961,N_13281,N_15919);
and U19962 (N_19962,N_14100,N_13382);
and U19963 (N_19963,N_16254,N_16689);
xor U19964 (N_19964,N_13707,N_17452);
or U19965 (N_19965,N_15385,N_15710);
xor U19966 (N_19966,N_14866,N_15473);
nand U19967 (N_19967,N_17426,N_13514);
or U19968 (N_19968,N_18402,N_13865);
nand U19969 (N_19969,N_14236,N_16651);
nor U19970 (N_19970,N_12788,N_12995);
and U19971 (N_19971,N_13867,N_18401);
or U19972 (N_19972,N_16465,N_15995);
or U19973 (N_19973,N_18225,N_17493);
nand U19974 (N_19974,N_17187,N_15602);
and U19975 (N_19975,N_13070,N_14605);
nand U19976 (N_19976,N_14939,N_13996);
xor U19977 (N_19977,N_18290,N_14642);
or U19978 (N_19978,N_16992,N_17634);
nand U19979 (N_19979,N_13737,N_13258);
or U19980 (N_19980,N_13882,N_14363);
xor U19981 (N_19981,N_18230,N_17933);
and U19982 (N_19982,N_14189,N_13399);
or U19983 (N_19983,N_17022,N_18270);
nand U19984 (N_19984,N_13754,N_12616);
nand U19985 (N_19985,N_15522,N_16894);
nand U19986 (N_19986,N_15894,N_13403);
nor U19987 (N_19987,N_17849,N_12550);
and U19988 (N_19988,N_13616,N_18106);
nor U19989 (N_19989,N_12850,N_15425);
or U19990 (N_19990,N_15735,N_17306);
nand U19991 (N_19991,N_16526,N_14477);
or U19992 (N_19992,N_14921,N_13231);
nand U19993 (N_19993,N_17485,N_15759);
nor U19994 (N_19994,N_13833,N_16456);
nor U19995 (N_19995,N_12523,N_16802);
nand U19996 (N_19996,N_14464,N_16416);
nand U19997 (N_19997,N_14651,N_15139);
or U19998 (N_19998,N_12826,N_16396);
nand U19999 (N_19999,N_15118,N_18183);
and U20000 (N_20000,N_16563,N_18456);
or U20001 (N_20001,N_14071,N_13764);
nand U20002 (N_20002,N_17232,N_12641);
or U20003 (N_20003,N_18610,N_14579);
and U20004 (N_20004,N_17188,N_15799);
nor U20005 (N_20005,N_18625,N_17292);
or U20006 (N_20006,N_13710,N_15157);
and U20007 (N_20007,N_16927,N_17638);
nor U20008 (N_20008,N_15715,N_16569);
nor U20009 (N_20009,N_18657,N_17403);
nor U20010 (N_20010,N_14364,N_13038);
nand U20011 (N_20011,N_13790,N_15959);
and U20012 (N_20012,N_14547,N_16598);
nand U20013 (N_20013,N_13095,N_18522);
nor U20014 (N_20014,N_17681,N_14472);
nand U20015 (N_20015,N_14084,N_13966);
and U20016 (N_20016,N_13331,N_15860);
nor U20017 (N_20017,N_14857,N_12972);
and U20018 (N_20018,N_16738,N_14208);
nor U20019 (N_20019,N_16030,N_16983);
xor U20020 (N_20020,N_15221,N_15040);
nor U20021 (N_20021,N_18601,N_12652);
xor U20022 (N_20022,N_16319,N_16430);
nand U20023 (N_20023,N_14996,N_18603);
and U20024 (N_20024,N_15364,N_17646);
or U20025 (N_20025,N_16492,N_13060);
xnor U20026 (N_20026,N_16521,N_16902);
nor U20027 (N_20027,N_18473,N_17053);
nand U20028 (N_20028,N_13447,N_15167);
and U20029 (N_20029,N_12552,N_16964);
nand U20030 (N_20030,N_14989,N_17316);
nand U20031 (N_20031,N_18169,N_18442);
nand U20032 (N_20032,N_14672,N_13612);
nor U20033 (N_20033,N_13528,N_15110);
nand U20034 (N_20034,N_18264,N_16886);
nand U20035 (N_20035,N_15075,N_15882);
xor U20036 (N_20036,N_16217,N_14359);
or U20037 (N_20037,N_12533,N_14971);
nor U20038 (N_20038,N_16305,N_18415);
and U20039 (N_20039,N_18143,N_17973);
or U20040 (N_20040,N_13141,N_16844);
nor U20041 (N_20041,N_16422,N_15026);
or U20042 (N_20042,N_16150,N_13473);
and U20043 (N_20043,N_17319,N_17463);
nor U20044 (N_20044,N_13783,N_18125);
or U20045 (N_20045,N_18037,N_16704);
and U20046 (N_20046,N_15819,N_18288);
nor U20047 (N_20047,N_16538,N_18557);
nand U20048 (N_20048,N_17495,N_13327);
nor U20049 (N_20049,N_17633,N_18555);
nand U20050 (N_20050,N_16627,N_17757);
or U20051 (N_20051,N_15403,N_16377);
xnor U20052 (N_20052,N_15651,N_17128);
nor U20053 (N_20053,N_18216,N_16361);
nor U20054 (N_20054,N_16403,N_17134);
or U20055 (N_20055,N_18140,N_15854);
xnor U20056 (N_20056,N_16468,N_15637);
or U20057 (N_20057,N_16965,N_17724);
or U20058 (N_20058,N_12604,N_13977);
and U20059 (N_20059,N_17753,N_15479);
and U20060 (N_20060,N_12896,N_16524);
nor U20061 (N_20061,N_18352,N_15355);
or U20062 (N_20062,N_12916,N_17995);
nor U20063 (N_20063,N_15138,N_18633);
or U20064 (N_20064,N_16604,N_18629);
nor U20065 (N_20065,N_14574,N_13307);
or U20066 (N_20066,N_13747,N_15519);
or U20067 (N_20067,N_18706,N_15598);
nor U20068 (N_20068,N_13645,N_13016);
nand U20069 (N_20069,N_17417,N_13951);
or U20070 (N_20070,N_15630,N_14759);
nand U20071 (N_20071,N_18102,N_13036);
nand U20072 (N_20072,N_16702,N_16501);
or U20073 (N_20073,N_15061,N_15378);
or U20074 (N_20074,N_17476,N_15156);
and U20075 (N_20075,N_17577,N_16709);
and U20076 (N_20076,N_14987,N_17726);
nand U20077 (N_20077,N_16664,N_12513);
nor U20078 (N_20078,N_18630,N_15584);
xor U20079 (N_20079,N_13745,N_18660);
nand U20080 (N_20080,N_16745,N_13897);
or U20081 (N_20081,N_17309,N_12782);
nand U20082 (N_20082,N_18294,N_14114);
and U20083 (N_20083,N_13534,N_15979);
nand U20084 (N_20084,N_16631,N_13672);
nand U20085 (N_20085,N_18066,N_16054);
or U20086 (N_20086,N_17714,N_16822);
or U20087 (N_20087,N_15142,N_14365);
nor U20088 (N_20088,N_17694,N_15296);
xor U20089 (N_20089,N_13163,N_18449);
and U20090 (N_20090,N_17168,N_14729);
nor U20091 (N_20091,N_17893,N_17136);
and U20092 (N_20092,N_16011,N_17494);
nor U20093 (N_20093,N_16039,N_13350);
nand U20094 (N_20094,N_17751,N_13513);
nand U20095 (N_20095,N_15810,N_17003);
nor U20096 (N_20096,N_17104,N_14366);
xnor U20097 (N_20097,N_18485,N_15513);
or U20098 (N_20098,N_13431,N_14560);
or U20099 (N_20099,N_16207,N_13309);
nor U20100 (N_20100,N_17020,N_13738);
and U20101 (N_20101,N_15730,N_17133);
or U20102 (N_20102,N_14961,N_18443);
nand U20103 (N_20103,N_12694,N_18501);
and U20104 (N_20104,N_17122,N_17571);
and U20105 (N_20105,N_16137,N_13164);
nor U20106 (N_20106,N_17925,N_13297);
nand U20107 (N_20107,N_14070,N_13735);
xor U20108 (N_20108,N_15181,N_14569);
nand U20109 (N_20109,N_12747,N_17789);
xnor U20110 (N_20110,N_15458,N_18679);
nor U20111 (N_20111,N_18735,N_18613);
nand U20112 (N_20112,N_17666,N_13845);
nor U20113 (N_20113,N_14104,N_13435);
nand U20114 (N_20114,N_15184,N_13606);
and U20115 (N_20115,N_15489,N_13784);
and U20116 (N_20116,N_12758,N_14265);
and U20117 (N_20117,N_17241,N_13802);
nor U20118 (N_20118,N_15203,N_16506);
and U20119 (N_20119,N_15706,N_14318);
or U20120 (N_20120,N_17715,N_15012);
xnor U20121 (N_20121,N_15499,N_15474);
nand U20122 (N_20122,N_17449,N_17084);
nand U20123 (N_20123,N_16679,N_17148);
or U20124 (N_20124,N_14770,N_12798);
xor U20125 (N_20125,N_16406,N_16818);
nor U20126 (N_20126,N_14471,N_15515);
or U20127 (N_20127,N_16177,N_12948);
xnor U20128 (N_20128,N_14400,N_18740);
xor U20129 (N_20129,N_14640,N_17459);
nand U20130 (N_20130,N_13680,N_13879);
nor U20131 (N_20131,N_18374,N_14347);
xnor U20132 (N_20132,N_15953,N_14615);
nand U20133 (N_20133,N_13207,N_16115);
or U20134 (N_20134,N_16852,N_17749);
and U20135 (N_20135,N_12678,N_14730);
nor U20136 (N_20136,N_14534,N_15545);
nand U20137 (N_20137,N_13126,N_16249);
nand U20138 (N_20138,N_15003,N_14941);
and U20139 (N_20139,N_18327,N_15028);
xor U20140 (N_20140,N_18408,N_18531);
or U20141 (N_20141,N_13579,N_18605);
nor U20142 (N_20142,N_14082,N_18273);
and U20143 (N_20143,N_16455,N_15585);
nor U20144 (N_20144,N_13538,N_16621);
and U20145 (N_20145,N_17871,N_12623);
or U20146 (N_20146,N_17706,N_14223);
xnor U20147 (N_20147,N_15528,N_12571);
and U20148 (N_20148,N_17480,N_16209);
or U20149 (N_20149,N_13527,N_18377);
nor U20150 (N_20150,N_12733,N_18275);
and U20151 (N_20151,N_17300,N_17546);
nor U20152 (N_20152,N_15557,N_13321);
and U20153 (N_20153,N_12893,N_18702);
xor U20154 (N_20154,N_12706,N_15877);
xor U20155 (N_20155,N_16236,N_12983);
and U20156 (N_20156,N_17100,N_15394);
or U20157 (N_20157,N_13697,N_18516);
nor U20158 (N_20158,N_15622,N_12868);
nor U20159 (N_20159,N_13503,N_17671);
xnor U20160 (N_20160,N_18373,N_12808);
nand U20161 (N_20161,N_16854,N_17421);
xnor U20162 (N_20162,N_18670,N_16948);
nand U20163 (N_20163,N_17524,N_16205);
and U20164 (N_20164,N_15800,N_14408);
or U20165 (N_20165,N_15863,N_14753);
or U20166 (N_20166,N_13922,N_13448);
xor U20167 (N_20167,N_17662,N_14544);
or U20168 (N_20168,N_15495,N_16884);
nand U20169 (N_20169,N_17811,N_15263);
and U20170 (N_20170,N_15429,N_16185);
or U20171 (N_20171,N_17560,N_14277);
nor U20172 (N_20172,N_17552,N_16379);
or U20173 (N_20173,N_18554,N_13010);
nor U20174 (N_20174,N_12752,N_16085);
xnor U20175 (N_20175,N_15504,N_12685);
nand U20176 (N_20176,N_13484,N_17390);
nand U20177 (N_20177,N_13912,N_17537);
nor U20178 (N_20178,N_15433,N_17601);
or U20179 (N_20179,N_14267,N_14974);
nand U20180 (N_20180,N_16619,N_13110);
nor U20181 (N_20181,N_14626,N_15175);
nand U20182 (N_20182,N_13693,N_16860);
and U20183 (N_20183,N_17878,N_16939);
nor U20184 (N_20184,N_18019,N_15267);
nand U20185 (N_20185,N_15600,N_14595);
nand U20186 (N_20186,N_14284,N_18224);
xnor U20187 (N_20187,N_16358,N_13914);
or U20188 (N_20188,N_17670,N_17215);
and U20189 (N_20189,N_16751,N_15472);
and U20190 (N_20190,N_18207,N_15490);
nor U20191 (N_20191,N_16454,N_17060);
and U20192 (N_20192,N_17870,N_17813);
and U20193 (N_20193,N_17883,N_13333);
or U20194 (N_20194,N_15655,N_13678);
nand U20195 (N_20195,N_15210,N_14779);
nor U20196 (N_20196,N_17693,N_17225);
and U20197 (N_20197,N_14950,N_14120);
xor U20198 (N_20198,N_18307,N_13102);
nand U20199 (N_20199,N_15780,N_14788);
and U20200 (N_20200,N_16826,N_16711);
nor U20201 (N_20201,N_17985,N_12966);
nand U20202 (N_20202,N_15627,N_17777);
nor U20203 (N_20203,N_15148,N_18624);
nor U20204 (N_20204,N_12990,N_16912);
xnor U20205 (N_20205,N_13911,N_18378);
nor U20206 (N_20206,N_12714,N_14370);
nand U20207 (N_20207,N_18682,N_17393);
xnor U20208 (N_20208,N_13112,N_16029);
xor U20209 (N_20209,N_15971,N_15581);
and U20210 (N_20210,N_13150,N_14422);
nor U20211 (N_20211,N_16633,N_14149);
or U20212 (N_20212,N_18488,N_12614);
nand U20213 (N_20213,N_16099,N_15565);
or U20214 (N_20214,N_17746,N_14513);
or U20215 (N_20215,N_13362,N_13025);
nor U20216 (N_20216,N_18695,N_12545);
nand U20217 (N_20217,N_15160,N_13709);
or U20218 (N_20218,N_15798,N_18453);
nand U20219 (N_20219,N_12581,N_16654);
nand U20220 (N_20220,N_16474,N_14180);
and U20221 (N_20221,N_18606,N_16767);
and U20222 (N_20222,N_14922,N_17700);
and U20223 (N_20223,N_15444,N_13608);
nor U20224 (N_20224,N_18033,N_15380);
and U20225 (N_20225,N_13533,N_14074);
nor U20226 (N_20226,N_14650,N_16271);
and U20227 (N_20227,N_15590,N_15326);
or U20228 (N_20228,N_13054,N_13532);
nand U20229 (N_20229,N_15348,N_15555);
and U20230 (N_20230,N_13375,N_15636);
nand U20231 (N_20231,N_14748,N_16144);
nand U20232 (N_20232,N_14991,N_17423);
and U20233 (N_20233,N_15222,N_18428);
xnor U20234 (N_20234,N_16421,N_17152);
nand U20235 (N_20235,N_12698,N_16801);
nor U20236 (N_20236,N_15663,N_13695);
and U20237 (N_20237,N_14696,N_12716);
and U20238 (N_20238,N_15372,N_15112);
xor U20239 (N_20239,N_13120,N_12904);
or U20240 (N_20240,N_16441,N_16479);
nand U20241 (N_20241,N_15011,N_13505);
or U20242 (N_20242,N_16573,N_17346);
nand U20243 (N_20243,N_13696,N_17078);
nor U20244 (N_20244,N_16245,N_15534);
nor U20245 (N_20245,N_13936,N_14000);
and U20246 (N_20246,N_13179,N_18163);
xor U20247 (N_20247,N_17021,N_14235);
or U20248 (N_20248,N_16542,N_17009);
xnor U20249 (N_20249,N_13019,N_13609);
nand U20250 (N_20250,N_15088,N_16562);
nand U20251 (N_20251,N_15709,N_14495);
nand U20252 (N_20252,N_14086,N_16583);
nor U20253 (N_20253,N_15793,N_15634);
nand U20254 (N_20254,N_16666,N_13749);
and U20255 (N_20255,N_13076,N_12838);
xor U20256 (N_20256,N_13825,N_14762);
xnor U20257 (N_20257,N_17038,N_15432);
nand U20258 (N_20258,N_13806,N_12549);
or U20259 (N_20259,N_17113,N_14892);
nor U20260 (N_20260,N_17966,N_16082);
or U20261 (N_20261,N_14242,N_18567);
and U20262 (N_20262,N_17767,N_16366);
nand U20263 (N_20263,N_13639,N_16143);
nand U20264 (N_20264,N_17848,N_16237);
nand U20265 (N_20265,N_17101,N_17551);
nor U20266 (N_20266,N_16196,N_13824);
nand U20267 (N_20267,N_17014,N_16330);
and U20268 (N_20268,N_18646,N_18251);
nand U20269 (N_20269,N_13663,N_17545);
and U20270 (N_20270,N_18419,N_13660);
and U20271 (N_20271,N_15427,N_12500);
or U20272 (N_20272,N_17896,N_17606);
and U20273 (N_20273,N_14740,N_13283);
nand U20274 (N_20274,N_15408,N_12575);
nor U20275 (N_20275,N_16495,N_13853);
or U20276 (N_20276,N_15325,N_13500);
or U20277 (N_20277,N_12953,N_13877);
or U20278 (N_20278,N_17771,N_15866);
nand U20279 (N_20279,N_14256,N_14266);
nand U20280 (N_20280,N_13720,N_18005);
nand U20281 (N_20281,N_16464,N_12746);
nor U20282 (N_20282,N_18301,N_13100);
or U20283 (N_20283,N_15999,N_18553);
nor U20284 (N_20284,N_17649,N_13318);
nand U20285 (N_20285,N_14649,N_15164);
nand U20286 (N_20286,N_17728,N_14711);
xor U20287 (N_20287,N_14807,N_15146);
or U20288 (N_20288,N_16057,N_12647);
and U20289 (N_20289,N_14291,N_15809);
and U20290 (N_20290,N_12900,N_13650);
nand U20291 (N_20291,N_13205,N_14172);
or U20292 (N_20292,N_17266,N_16461);
or U20293 (N_20293,N_16827,N_15446);
nor U20294 (N_20294,N_12799,N_15699);
nor U20295 (N_20295,N_14883,N_13300);
and U20296 (N_20296,N_17445,N_13888);
nand U20297 (N_20297,N_14249,N_13219);
or U20298 (N_20298,N_13804,N_15775);
or U20299 (N_20299,N_13971,N_17641);
or U20300 (N_20300,N_15512,N_18570);
nor U20301 (N_20301,N_15345,N_16060);
nand U20302 (N_20302,N_13915,N_15065);
nand U20303 (N_20303,N_13489,N_13418);
or U20304 (N_20304,N_13094,N_15990);
nor U20305 (N_20305,N_15729,N_15834);
nor U20306 (N_20306,N_16616,N_16981);
and U20307 (N_20307,N_18469,N_15687);
nor U20308 (N_20308,N_14286,N_14381);
nor U20309 (N_20309,N_18341,N_17044);
or U20310 (N_20310,N_15491,N_17844);
or U20311 (N_20311,N_14681,N_13123);
nand U20312 (N_20312,N_17889,N_15539);
or U20313 (N_20313,N_14437,N_14924);
nor U20314 (N_20314,N_17431,N_15783);
or U20315 (N_20315,N_13913,N_18566);
nor U20316 (N_20316,N_17326,N_17707);
nor U20317 (N_20317,N_16769,N_12994);
nor U20318 (N_20318,N_14700,N_17299);
xnor U20319 (N_20319,N_13852,N_16101);
nand U20320 (N_20320,N_14908,N_18681);
or U20321 (N_20321,N_15837,N_13020);
and U20322 (N_20322,N_15635,N_16105);
and U20323 (N_20323,N_15108,N_14533);
nand U20324 (N_20324,N_17576,N_18508);
xnor U20325 (N_20325,N_15771,N_13427);
nor U20326 (N_20326,N_14333,N_13753);
or U20327 (N_20327,N_13787,N_17720);
nand U20328 (N_20328,N_14954,N_13886);
nor U20329 (N_20329,N_17061,N_17027);
xnor U20330 (N_20330,N_16079,N_16510);
nand U20331 (N_20331,N_15349,N_14331);
and U20332 (N_20332,N_14482,N_14371);
and U20333 (N_20333,N_18639,N_14492);
or U20334 (N_20334,N_15288,N_15395);
nand U20335 (N_20335,N_18463,N_16841);
or U20336 (N_20336,N_16096,N_18711);
and U20337 (N_20337,N_18591,N_16471);
nor U20338 (N_20338,N_15858,N_14354);
xnor U20339 (N_20339,N_17067,N_14250);
nor U20340 (N_20340,N_14767,N_17220);
and U20341 (N_20341,N_16988,N_16356);
nand U20342 (N_20342,N_15402,N_17040);
nor U20343 (N_20343,N_17217,N_17587);
nor U20344 (N_20344,N_18503,N_15994);
and U20345 (N_20345,N_18683,N_18692);
nand U20346 (N_20346,N_17970,N_16575);
xnor U20347 (N_20347,N_17990,N_15343);
nand U20348 (N_20348,N_18184,N_16166);
and U20349 (N_20349,N_16201,N_13248);
nor U20350 (N_20350,N_13771,N_13834);
or U20351 (N_20351,N_13159,N_15258);
and U20352 (N_20352,N_18672,N_16688);
and U20353 (N_20353,N_13980,N_15632);
and U20354 (N_20354,N_15129,N_13477);
or U20355 (N_20355,N_14452,N_18315);
or U20356 (N_20356,N_12589,N_17903);
nor U20357 (N_20357,N_12943,N_17836);
nor U20358 (N_20358,N_15825,N_13021);
nor U20359 (N_20359,N_12860,N_13394);
nor U20360 (N_20360,N_14081,N_14737);
or U20361 (N_20361,N_16438,N_17522);
and U20362 (N_20362,N_15033,N_17162);
nand U20363 (N_20363,N_17297,N_14768);
xor U20364 (N_20364,N_15468,N_13013);
nor U20365 (N_20365,N_17320,N_13855);
or U20366 (N_20366,N_14234,N_14716);
or U20367 (N_20367,N_15212,N_16375);
xnor U20368 (N_20368,N_14509,N_16078);
nand U20369 (N_20369,N_17064,N_13073);
or U20370 (N_20370,N_16883,N_13873);
nand U20371 (N_20371,N_15036,N_14570);
and U20372 (N_20372,N_14527,N_17340);
nand U20373 (N_20373,N_16687,N_16959);
or U20374 (N_20374,N_14179,N_14011);
xnor U20375 (N_20375,N_15007,N_15917);
or U20376 (N_20376,N_16084,N_17106);
nand U20377 (N_20377,N_17163,N_15645);
or U20378 (N_20378,N_16872,N_14468);
or U20379 (N_20379,N_14295,N_13998);
nor U20380 (N_20380,N_18201,N_15966);
nand U20381 (N_20381,N_15886,N_12512);
and U20382 (N_20382,N_13287,N_15673);
and U20383 (N_20383,N_18280,N_18437);
and U20384 (N_20384,N_13507,N_16910);
xor U20385 (N_20385,N_16695,N_17555);
or U20386 (N_20386,N_18200,N_15957);
and U20387 (N_20387,N_12588,N_17705);
and U20388 (N_20388,N_16706,N_16623);
and U20389 (N_20389,N_12907,N_17867);
and U20390 (N_20390,N_15303,N_13292);
or U20391 (N_20391,N_13973,N_16197);
nor U20392 (N_20392,N_14283,N_12722);
nor U20393 (N_20393,N_16534,N_12701);
or U20394 (N_20394,N_15650,N_15218);
nor U20395 (N_20395,N_15705,N_17317);
nor U20396 (N_20396,N_15728,N_15986);
nor U20397 (N_20397,N_15098,N_12538);
xor U20398 (N_20398,N_14794,N_12880);
nand U20399 (N_20399,N_17563,N_17556);
and U20400 (N_20400,N_15231,N_17795);
and U20401 (N_20401,N_18587,N_14806);
xor U20402 (N_20402,N_14889,N_13789);
or U20403 (N_20403,N_15339,N_17654);
or U20404 (N_20404,N_18056,N_13718);
or U20405 (N_20405,N_16596,N_13953);
nand U20406 (N_20406,N_12703,N_14735);
or U20407 (N_20407,N_15321,N_16985);
nand U20408 (N_20408,N_16359,N_13798);
nand U20409 (N_20409,N_13941,N_15824);
xnor U20410 (N_20410,N_15089,N_17701);
nand U20411 (N_20411,N_18030,N_17184);
nor U20412 (N_20412,N_16708,N_16304);
or U20413 (N_20413,N_13714,N_17983);
or U20414 (N_20414,N_13763,N_13368);
or U20415 (N_20415,N_13091,N_16837);
and U20416 (N_20416,N_14776,N_16655);
and U20417 (N_20417,N_17969,N_17922);
nand U20418 (N_20418,N_16153,N_18344);
nand U20419 (N_20419,N_13590,N_15747);
or U20420 (N_20420,N_13379,N_16723);
nor U20421 (N_20421,N_16567,N_14723);
nand U20422 (N_20422,N_18132,N_17854);
and U20423 (N_20423,N_13555,N_16508);
or U20424 (N_20424,N_14959,N_13927);
nand U20425 (N_20425,N_15438,N_16392);
and U20426 (N_20426,N_14054,N_14835);
or U20427 (N_20427,N_13662,N_18027);
or U20428 (N_20428,N_15640,N_18013);
nor U20429 (N_20429,N_14418,N_17406);
nor U20430 (N_20430,N_16582,N_15350);
or U20431 (N_20431,N_17920,N_14467);
and U20432 (N_20432,N_17451,N_14760);
nand U20433 (N_20433,N_16351,N_14749);
nor U20434 (N_20434,N_14800,N_17894);
xnor U20435 (N_20435,N_17278,N_16307);
or U20436 (N_20436,N_17488,N_17838);
nor U20437 (N_20437,N_14934,N_15044);
and U20438 (N_20438,N_15787,N_18565);
nand U20439 (N_20439,N_18355,N_18084);
or U20440 (N_20440,N_13280,N_16796);
nand U20441 (N_20441,N_14577,N_14057);
or U20442 (N_20442,N_17388,N_15370);
and U20443 (N_20443,N_13482,N_18487);
or U20444 (N_20444,N_17272,N_13805);
or U20445 (N_20445,N_16775,N_12580);
xnor U20446 (N_20446,N_12653,N_17581);
and U20447 (N_20447,N_17160,N_17121);
nor U20448 (N_20448,N_14424,N_14170);
and U20449 (N_20449,N_14687,N_18698);
or U20450 (N_20450,N_15766,N_17858);
or U20451 (N_20451,N_14538,N_17080);
or U20452 (N_20452,N_15048,N_14526);
xor U20453 (N_20453,N_13818,N_16210);
nor U20454 (N_20454,N_15746,N_15274);
and U20455 (N_20455,N_17279,N_12681);
nor U20456 (N_20456,N_15931,N_14652);
nand U20457 (N_20457,N_15333,N_14055);
or U20458 (N_20458,N_12813,N_13134);
and U20459 (N_20459,N_16434,N_16565);
and U20460 (N_20460,N_16289,N_14423);
nor U20461 (N_20461,N_17982,N_17072);
nor U20462 (N_20462,N_14837,N_14085);
nand U20463 (N_20463,N_17174,N_16718);
nor U20464 (N_20464,N_17371,N_17882);
nand U20465 (N_20465,N_12577,N_12794);
xor U20466 (N_20466,N_17077,N_15911);
nor U20467 (N_20467,N_15852,N_14310);
nand U20468 (N_20468,N_17547,N_18189);
nor U20469 (N_20469,N_13299,N_17105);
nand U20470 (N_20470,N_12991,N_17812);
nor U20471 (N_20471,N_16373,N_14530);
nand U20472 (N_20472,N_18175,N_13338);
nand U20473 (N_20473,N_15521,N_16310);
nand U20474 (N_20474,N_16489,N_16656);
xnor U20475 (N_20475,N_16446,N_16170);
and U20476 (N_20476,N_16771,N_17293);
or U20477 (N_20477,N_16324,N_18721);
nor U20478 (N_20478,N_16785,N_15276);
nor U20479 (N_20479,N_18714,N_13985);
nand U20480 (N_20480,N_15697,N_16905);
or U20481 (N_20481,N_12772,N_17905);
nor U20482 (N_20482,N_17837,N_13517);
or U20483 (N_20483,N_15659,N_12598);
nand U20484 (N_20484,N_16682,N_14449);
nand U20485 (N_20485,N_14931,N_17763);
xor U20486 (N_20486,N_17255,N_13880);
or U20487 (N_20487,N_16740,N_13719);
nor U20488 (N_20488,N_13525,N_16926);
nand U20489 (N_20489,N_12971,N_12901);
and U20490 (N_20490,N_15052,N_17731);
nand U20491 (N_20491,N_17514,N_15173);
nor U20492 (N_20492,N_15208,N_15983);
nor U20493 (N_20493,N_15496,N_17192);
nand U20494 (N_20494,N_15711,N_14917);
xnor U20495 (N_20495,N_14688,N_13541);
nor U20496 (N_20496,N_14925,N_14628);
and U20497 (N_20497,N_14940,N_15554);
or U20498 (N_20498,N_16052,N_17604);
or U20499 (N_20499,N_15850,N_15485);
or U20500 (N_20500,N_17674,N_13264);
xor U20501 (N_20501,N_12932,N_15283);
and U20502 (N_20502,N_14555,N_13795);
nand U20503 (N_20503,N_18431,N_13948);
or U20504 (N_20504,N_17289,N_17528);
or U20505 (N_20505,N_15506,N_13629);
xnor U20506 (N_20506,N_16643,N_18166);
or U20507 (N_20507,N_18583,N_16490);
nor U20508 (N_20508,N_13495,N_17378);
xnor U20509 (N_20509,N_15761,N_16061);
nand U20510 (N_20510,N_14983,N_18217);
nor U20511 (N_20511,N_17833,N_14518);
and U20512 (N_20512,N_14123,N_17145);
and U20513 (N_20513,N_13899,N_16431);
xnor U20514 (N_20514,N_16868,N_12941);
nand U20515 (N_20515,N_14457,N_13023);
nand U20516 (N_20516,N_17554,N_13291);
or U20517 (N_20517,N_14202,N_13677);
nand U20518 (N_20518,N_15923,N_12867);
and U20519 (N_20519,N_13449,N_18726);
nor U20520 (N_20520,N_13263,N_14373);
nand U20521 (N_20521,N_13182,N_18093);
or U20522 (N_20522,N_17585,N_13520);
nand U20523 (N_20523,N_15039,N_15638);
nand U20524 (N_20524,N_14080,N_13762);
nor U20525 (N_20525,N_15140,N_12856);
and U20526 (N_20526,N_14436,N_16255);
or U20527 (N_20527,N_16683,N_17739);
nand U20528 (N_20528,N_13542,N_15704);
nand U20529 (N_20529,N_14355,N_17448);
nor U20530 (N_20530,N_12633,N_15949);
or U20531 (N_20531,N_13675,N_13862);
nand U20532 (N_20532,N_17685,N_16765);
nor U20533 (N_20533,N_14144,N_12999);
xnor U20534 (N_20534,N_18527,N_13896);
or U20535 (N_20535,N_12976,N_14133);
or U20536 (N_20536,N_12719,N_13518);
nor U20537 (N_20537,N_18578,N_17570);
and U20538 (N_20538,N_18156,N_13136);
nand U20539 (N_20539,N_15914,N_14173);
xnor U20540 (N_20540,N_13400,N_13006);
nor U20541 (N_20541,N_14869,N_16522);
nor U20542 (N_20542,N_18076,N_13651);
and U20543 (N_20543,N_14389,N_18164);
or U20544 (N_20544,N_15791,N_18274);
and U20545 (N_20545,N_13929,N_12634);
nand U20546 (N_20546,N_13679,N_13632);
nor U20547 (N_20547,N_18483,N_12897);
nor U20548 (N_20548,N_16220,N_12834);
nand U20549 (N_20549,N_18600,N_18612);
nand U20550 (N_20550,N_13646,N_17473);
or U20551 (N_20551,N_16466,N_15667);
xnor U20552 (N_20552,N_12945,N_12870);
nor U20553 (N_20553,N_17471,N_15450);
or U20554 (N_20554,N_15230,N_15284);
nand U20555 (N_20555,N_14895,N_14473);
nand U20556 (N_20556,N_15776,N_16586);
nor U20557 (N_20557,N_15648,N_13232);
or U20558 (N_20558,N_16483,N_18209);
nand U20559 (N_20559,N_17642,N_15068);
nand U20560 (N_20560,N_14314,N_13841);
and U20561 (N_20561,N_14028,N_15171);
nand U20562 (N_20562,N_15384,N_14916);
xor U20563 (N_20563,N_13039,N_14281);
and U20564 (N_20564,N_16537,N_14204);
nor U20565 (N_20565,N_17146,N_16459);
nor U20566 (N_20566,N_12514,N_18036);
nor U20567 (N_20567,N_16227,N_14968);
nand U20568 (N_20568,N_12817,N_18512);
nand U20569 (N_20569,N_14537,N_14977);
nor U20570 (N_20570,N_18313,N_17010);
nand U20571 (N_20571,N_12950,N_14965);
nor U20572 (N_20572,N_18176,N_17923);
or U20573 (N_20573,N_17622,N_14107);
xnor U20574 (N_20574,N_17904,N_13096);
nand U20575 (N_20575,N_13731,N_14601);
or U20576 (N_20576,N_14038,N_13846);
nor U20577 (N_20577,N_14147,N_17483);
nand U20578 (N_20578,N_18015,N_18749);
nand U20579 (N_20579,N_13346,N_14731);
nand U20580 (N_20580,N_12663,N_15484);
xor U20581 (N_20581,N_18192,N_18110);
nand U20582 (N_20582,N_13286,N_15266);
and U20583 (N_20583,N_15572,N_14845);
nand U20584 (N_20584,N_12783,N_17191);
or U20585 (N_20585,N_15022,N_13925);
and U20586 (N_20586,N_13171,N_14369);
or U20587 (N_20587,N_13432,N_17211);
or U20588 (N_20588,N_17407,N_17526);
or U20589 (N_20589,N_15078,N_18595);
nand U20590 (N_20590,N_13027,N_17115);
nand U20591 (N_20591,N_14668,N_14699);
nor U20592 (N_20592,N_17951,N_16780);
nor U20593 (N_20593,N_15189,N_18328);
nor U20594 (N_20594,N_14153,N_17676);
and U20595 (N_20595,N_15665,N_14743);
xnor U20596 (N_20596,N_18279,N_16439);
and U20597 (N_20597,N_17841,N_14435);
or U20598 (N_20598,N_18137,N_17098);
or U20599 (N_20599,N_13599,N_13595);
nor U20600 (N_20600,N_14497,N_15229);
nor U20601 (N_20601,N_12805,N_13407);
nand U20602 (N_20602,N_16244,N_15133);
or U20603 (N_20603,N_17909,N_13851);
and U20604 (N_20604,N_17946,N_13172);
nor U20605 (N_20605,N_12993,N_16008);
and U20606 (N_20606,N_13125,N_16429);
or U20607 (N_20607,N_16009,N_14646);
or U20608 (N_20608,N_14210,N_14004);
nor U20609 (N_20609,N_13373,N_16395);
or U20610 (N_20610,N_17828,N_14072);
nor U20611 (N_20611,N_17847,N_17277);
or U20612 (N_20612,N_15045,N_15404);
or U20613 (N_20613,N_13144,N_14781);
or U20614 (N_20614,N_15168,N_14817);
nor U20615 (N_20615,N_13436,N_15718);
xor U20616 (N_20616,N_16882,N_18671);
or U20617 (N_20617,N_18604,N_13294);
xor U20618 (N_20618,N_17349,N_16120);
xor U20619 (N_20619,N_18394,N_17157);
and U20620 (N_20620,N_14654,N_14849);
or U20621 (N_20621,N_13909,N_17295);
nor U20622 (N_20622,N_18167,N_18666);
nor U20623 (N_20623,N_16272,N_16528);
nand U20624 (N_20624,N_17243,N_14276);
nand U20625 (N_20625,N_14865,N_18472);
nand U20626 (N_20626,N_15301,N_15224);
or U20627 (N_20627,N_17659,N_13416);
nor U20628 (N_20628,N_13155,N_14159);
or U20629 (N_20629,N_13511,N_18515);
nand U20630 (N_20630,N_16644,N_16795);
xnor U20631 (N_20631,N_16829,N_12851);
or U20632 (N_20632,N_13471,N_12543);
and U20633 (N_20633,N_15154,N_16372);
or U20634 (N_20634,N_13050,N_13341);
xnor U20635 (N_20635,N_13092,N_15559);
nand U20636 (N_20636,N_16152,N_13424);
and U20637 (N_20637,N_18136,N_18077);
nand U20638 (N_20638,N_17082,N_18026);
or U20639 (N_20639,N_13588,N_13365);
nor U20640 (N_20640,N_13048,N_13553);
and U20641 (N_20641,N_13704,N_12980);
nor U20642 (N_20642,N_17860,N_16863);
or U20643 (N_20643,N_15250,N_15469);
and U20644 (N_20644,N_13869,N_15219);
xnor U20645 (N_20645,N_16650,N_17801);
or U20646 (N_20646,N_17696,N_17108);
nor U20647 (N_20647,N_13883,N_16594);
nand U20648 (N_20648,N_13900,N_18054);
nor U20649 (N_20649,N_15563,N_13683);
nor U20650 (N_20650,N_14558,N_14803);
nand U20651 (N_20651,N_16560,N_15965);
nand U20652 (N_20652,N_17742,N_17209);
or U20653 (N_20653,N_12843,N_16336);
nor U20654 (N_20654,N_16523,N_15725);
xor U20655 (N_20655,N_13562,N_14914);
and U20656 (N_20656,N_12556,N_16615);
or U20657 (N_20657,N_13388,N_16888);
and U20658 (N_20658,N_14938,N_13856);
nand U20659 (N_20659,N_16747,N_17329);
or U20660 (N_20660,N_15764,N_16146);
and U20661 (N_20661,N_17650,N_14427);
nand U20662 (N_20662,N_17062,N_14990);
nor U20663 (N_20663,N_14466,N_18622);
nor U20664 (N_20664,N_13866,N_15063);
and U20665 (N_20665,N_14707,N_18148);
and U20666 (N_20666,N_15024,N_16204);
or U20667 (N_20667,N_15892,N_15434);
xor U20668 (N_20668,N_12608,N_13551);
xnor U20669 (N_20669,N_15091,N_13395);
and U20670 (N_20670,N_13592,N_18609);
xor U20671 (N_20671,N_14097,N_17725);
nand U20672 (N_20672,N_14248,N_13195);
and U20673 (N_20673,N_14176,N_15518);
or U20674 (N_20674,N_14096,N_18389);
nor U20675 (N_20675,N_12883,N_18072);
nand U20676 (N_20676,N_17754,N_17015);
nor U20677 (N_20677,N_18240,N_12992);
and U20678 (N_20678,N_16559,N_18318);
or U20679 (N_20679,N_17193,N_18533);
xnor U20680 (N_20680,N_14620,N_14798);
nor U20681 (N_20681,N_17877,N_15676);
or U20682 (N_20682,N_17348,N_16798);
nand U20683 (N_20683,N_18204,N_14641);
xnor U20684 (N_20684,N_15642,N_16281);
nor U20685 (N_20685,N_16512,N_17089);
nand U20686 (N_20686,N_12689,N_14982);
xnor U20687 (N_20687,N_15660,N_18369);
or U20688 (N_20688,N_16691,N_17829);
nand U20689 (N_20689,N_17314,N_14813);
or U20690 (N_20690,N_18704,N_12833);
nor U20691 (N_20691,N_17090,N_14754);
nand U20692 (N_20692,N_13711,N_14884);
nor U20693 (N_20693,N_15143,N_18085);
nor U20694 (N_20694,N_16178,N_14067);
xor U20695 (N_20695,N_16413,N_13479);
and U20696 (N_20696,N_14199,N_14859);
or U20697 (N_20697,N_13601,N_15478);
nor U20698 (N_20698,N_14105,N_14207);
and U20699 (N_20699,N_18039,N_16119);
or U20700 (N_20700,N_15092,N_16222);
or U20701 (N_20701,N_15314,N_14125);
nor U20702 (N_20702,N_18003,N_16198);
or U20703 (N_20703,N_16005,N_16155);
or U20704 (N_20704,N_15162,N_16357);
or U20705 (N_20705,N_17024,N_18693);
nor U20706 (N_20706,N_17768,N_15503);
nand U20707 (N_20707,N_16762,N_15262);
or U20708 (N_20708,N_17347,N_16063);
or U20709 (N_20709,N_15589,N_17158);
nand U20710 (N_20710,N_12584,N_13149);
or U20711 (N_20711,N_17376,N_14854);
or U20712 (N_20712,N_17733,N_12553);
nand U20713 (N_20713,N_14130,N_17874);
nor U20714 (N_20714,N_16834,N_15334);
nand U20715 (N_20715,N_16597,N_17511);
xnor U20716 (N_20716,N_15906,N_17374);
or U20717 (N_20717,N_18499,N_16283);
or U20718 (N_20718,N_16547,N_17938);
and U20719 (N_20719,N_17213,N_13105);
or U20720 (N_20720,N_13703,N_13584);
or U20721 (N_20721,N_16348,N_12780);
xor U20722 (N_20722,N_12541,N_18011);
xnor U20723 (N_20723,N_18429,N_16183);
or U20724 (N_20724,N_13494,N_18451);
nor U20725 (N_20725,N_15451,N_13552);
nor U20726 (N_20726,N_16485,N_13044);
nor U20727 (N_20727,N_12824,N_16578);
nor U20728 (N_20728,N_18082,N_17872);
nand U20729 (N_20729,N_16743,N_15594);
nand U20730 (N_20730,N_15812,N_17914);
nand U20731 (N_20731,N_13460,N_17251);
nand U20732 (N_20732,N_15847,N_16260);
or U20733 (N_20733,N_16514,N_15338);
nor U20734 (N_20734,N_13572,N_12955);
xor U20735 (N_20735,N_17513,N_13991);
or U20736 (N_20736,N_14101,N_17954);
or U20737 (N_20737,N_17019,N_13717);
and U20738 (N_20738,N_18440,N_12650);
nor U20739 (N_20739,N_17980,N_13306);
nor U20740 (N_20740,N_18659,N_14876);
and U20741 (N_20741,N_15765,N_15613);
nor U20742 (N_20742,N_18421,N_12609);
and U20743 (N_20743,N_16919,N_14661);
or U20744 (N_20744,N_17900,N_14553);
nand U20745 (N_20745,N_15576,N_14027);
or U20746 (N_20746,N_16803,N_16890);
and U20747 (N_20747,N_17242,N_13543);
or U20748 (N_20748,N_14367,N_16516);
and U20749 (N_20749,N_14025,N_12692);
xor U20750 (N_20750,N_16979,N_18267);
and U20751 (N_20751,N_18365,N_12875);
and U20752 (N_20752,N_12910,N_18057);
nand U20753 (N_20753,N_17283,N_12879);
nand U20754 (N_20754,N_17422,N_16734);
nor U20755 (N_20755,N_18479,N_18248);
xnor U20756 (N_20756,N_17248,N_14901);
or U20757 (N_20757,N_15569,N_17735);
and U20758 (N_20758,N_16042,N_18017);
xor U20759 (N_20759,N_15008,N_16360);
or U20760 (N_20760,N_13273,N_18177);
xnor U20761 (N_20761,N_13201,N_17290);
and U20762 (N_20762,N_14572,N_18493);
xor U20763 (N_20763,N_16161,N_14294);
and U20764 (N_20764,N_15918,N_13868);
and U20765 (N_20765,N_13603,N_12903);
nand U20766 (N_20766,N_18257,N_14993);
and U20767 (N_20767,N_17712,N_13724);
nor U20768 (N_20768,N_17942,N_15105);
nor U20769 (N_20769,N_16539,N_16558);
nand U20770 (N_20770,N_17173,N_14110);
or U20771 (N_20771,N_12825,N_16761);
nand U20772 (N_20772,N_18016,N_16931);
or U20773 (N_20773,N_17058,N_13293);
nor U20774 (N_20774,N_16181,N_17965);
nor U20775 (N_20775,N_12640,N_13456);
nand U20776 (N_20776,N_18012,N_17045);
and U20777 (N_20777,N_16404,N_16963);
or U20778 (N_20778,N_16274,N_17498);
and U20779 (N_20779,N_17337,N_17324);
nor U20780 (N_20780,N_15570,N_14675);
or U20781 (N_20781,N_17361,N_17218);
nand U20782 (N_20782,N_13928,N_13547);
or U20783 (N_20783,N_14736,N_13800);
and U20784 (N_20784,N_16448,N_16004);
and U20785 (N_20785,N_16986,N_16134);
or U20786 (N_20786,N_13602,N_14774);
and U20787 (N_20787,N_13975,N_18526);
or U20788 (N_20788,N_14053,N_14029);
nor U20789 (N_20789,N_12929,N_16065);
nor U20790 (N_20790,N_12583,N_13366);
and U20791 (N_20791,N_14718,N_17079);
or U20792 (N_20792,N_15272,N_15769);
or U20793 (N_20793,N_16083,N_16815);
or U20794 (N_20794,N_12775,N_18304);
nor U20795 (N_20795,N_13965,N_14353);
or U20796 (N_20796,N_13876,N_18089);
or U20797 (N_20797,N_14003,N_14602);
nand U20798 (N_20798,N_16315,N_17523);
nor U20799 (N_20799,N_13653,N_17566);
nand U20800 (N_20800,N_13438,N_13452);
nand U20801 (N_20801,N_13910,N_17444);
xor U20802 (N_20802,N_16876,N_14811);
nor U20803 (N_20803,N_17636,N_18579);
and U20804 (N_20804,N_18162,N_17307);
nor U20805 (N_20805,N_15002,N_17509);
or U20806 (N_20806,N_14190,N_13428);
nand U20807 (N_20807,N_14433,N_13930);
or U20808 (N_20808,N_13213,N_14386);
nand U20809 (N_20809,N_16427,N_13988);
nor U20810 (N_20810,N_14566,N_13878);
and U20811 (N_20811,N_13313,N_17334);
or U20812 (N_20812,N_16779,N_18723);
or U20813 (N_20813,N_14549,N_16190);
or U20814 (N_20814,N_17331,N_18310);
or U20815 (N_20815,N_18379,N_17387);
xnor U20816 (N_20816,N_18237,N_18329);
and U20817 (N_20817,N_14117,N_13485);
nand U20818 (N_20818,N_14943,N_17446);
nor U20819 (N_20819,N_17436,N_15871);
and U20820 (N_20820,N_13739,N_17258);
and U20821 (N_20821,N_13637,N_17233);
nor U20822 (N_20822,N_15072,N_16100);
nand U20823 (N_20823,N_14625,N_15587);
or U20824 (N_20824,N_15064,N_17711);
and U20825 (N_20825,N_13497,N_12530);
and U20826 (N_20826,N_13045,N_18215);
xor U20827 (N_20827,N_15831,N_13983);
nand U20828 (N_20828,N_12683,N_13404);
nand U20829 (N_20829,N_15807,N_16571);
nand U20830 (N_20830,N_17238,N_13257);
nor U20831 (N_20831,N_16676,N_13227);
and U20832 (N_20832,N_15207,N_16125);
xnor U20833 (N_20833,N_18061,N_14300);
and U20834 (N_20834,N_14224,N_16828);
nand U20835 (N_20835,N_15662,N_17851);
and U20836 (N_20836,N_17492,N_15978);
nor U20837 (N_20837,N_17418,N_17544);
or U20838 (N_20838,N_18333,N_16993);
nor U20839 (N_20839,N_16179,N_14846);
nor U20840 (N_20840,N_18598,N_14329);
and U20841 (N_20841,N_15639,N_14850);
nor U20842 (N_20842,N_16847,N_17151);
nor U20843 (N_20843,N_14320,N_17952);
or U20844 (N_20844,N_13186,N_17621);
or U20845 (N_20845,N_12846,N_16215);
nand U20846 (N_20846,N_17095,N_13022);
nand U20847 (N_20847,N_18444,N_15813);
nor U20848 (N_20848,N_18466,N_13295);
nor U20849 (N_20849,N_15351,N_15398);
or U20850 (N_20850,N_15116,N_16172);
and U20851 (N_20851,N_17639,N_13557);
nor U20852 (N_20852,N_18596,N_16951);
nor U20853 (N_20853,N_18145,N_14893);
and U20854 (N_20854,N_15982,N_15579);
and U20855 (N_20855,N_14906,N_18111);
xnor U20856 (N_20856,N_14843,N_17615);
nor U20857 (N_20857,N_14832,N_17487);
or U20858 (N_20858,N_12551,N_16098);
or U20859 (N_20859,N_14007,N_15560);
nor U20860 (N_20860,N_16971,N_16913);
or U20861 (N_20861,N_17960,N_12511);
nand U20862 (N_20862,N_15465,N_14504);
nand U20863 (N_20863,N_18360,N_13563);
and U20864 (N_20864,N_16634,N_13162);
nor U20865 (N_20865,N_15020,N_13578);
nor U20866 (N_20866,N_18689,N_17769);
nand U20867 (N_20867,N_17395,N_13371);
nand U20868 (N_20868,N_14568,N_14692);
and U20869 (N_20869,N_18150,N_14563);
nor U20870 (N_20870,N_15234,N_12718);
nor U20871 (N_20871,N_17906,N_13451);
xnor U20872 (N_20872,N_17595,N_17261);
or U20873 (N_20873,N_16955,N_18409);
or U20874 (N_20874,N_14017,N_18399);
nand U20875 (N_20875,N_15671,N_18628);
nor U20876 (N_20876,N_18115,N_16727);
nor U20877 (N_20877,N_17931,N_16398);
nor U20878 (N_20878,N_14772,N_16805);
nand U20879 (N_20879,N_14542,N_15567);
xor U20880 (N_20880,N_16878,N_18335);
nor U20881 (N_20881,N_16040,N_12928);
nor U20882 (N_20882,N_12599,N_15564);
and U20883 (N_20883,N_16484,N_17603);
nand U20884 (N_20884,N_13282,N_16165);
xor U20885 (N_20885,N_13510,N_14432);
nor U20886 (N_20886,N_13968,N_13450);
nand U20887 (N_20887,N_17088,N_17630);
xor U20888 (N_20888,N_14614,N_16622);
and U20889 (N_20889,N_14773,N_12667);
nand U20890 (N_20890,N_13796,N_15279);
or U20891 (N_20891,N_14126,N_13440);
nor U20892 (N_20892,N_13861,N_14292);
nand U20893 (N_20893,N_13336,N_13712);
nand U20894 (N_20894,N_14809,N_15217);
nand U20895 (N_20895,N_16967,N_15439);
and U20896 (N_20896,N_17212,N_14963);
and U20897 (N_20897,N_18632,N_14352);
xor U20898 (N_20898,N_13475,N_18002);
or U20899 (N_20899,N_12562,N_18543);
nand U20900 (N_20900,N_16531,N_14665);
nor U20901 (N_20901,N_13178,N_12815);
or U20902 (N_20902,N_15808,N_15505);
or U20903 (N_20903,N_15249,N_18362);
or U20904 (N_20904,N_13523,N_17656);
nor U20905 (N_20905,N_14511,N_14988);
nor U20906 (N_20906,N_15029,N_14981);
or U20907 (N_20907,N_15308,N_17017);
nor U20908 (N_20908,N_18568,N_14151);
or U20909 (N_20909,N_15289,N_15586);
nand U20910 (N_20910,N_14045,N_16149);
and U20911 (N_20911,N_12894,N_16629);
nand U20912 (N_20912,N_16051,N_18323);
or U20913 (N_20913,N_13726,N_16365);
and U20914 (N_20914,N_17076,N_18364);
nor U20915 (N_20915,N_13389,N_17118);
xnor U20916 (N_20916,N_15242,N_14673);
nand U20917 (N_20917,N_16692,N_15993);
nor U20918 (N_20918,N_13345,N_12655);
nand U20919 (N_20919,N_14230,N_18530);
nor U20920 (N_20920,N_15790,N_14470);
and U20921 (N_20921,N_16836,N_16480);
nor U20922 (N_20922,N_14746,N_17195);
xor U20923 (N_20923,N_14708,N_17748);
nand U20924 (N_20924,N_14690,N_17853);
nor U20925 (N_20925,N_12785,N_18023);
nor U20926 (N_20926,N_18244,N_15541);
nor U20927 (N_20927,N_16608,N_17150);
or U20928 (N_20928,N_18266,N_15060);
and U20929 (N_20929,N_15202,N_14059);
nand U20930 (N_20930,N_16977,N_15754);
nand U20931 (N_20931,N_15141,N_17228);
and U20932 (N_20932,N_17206,N_17734);
or U20933 (N_20933,N_16897,N_15768);
and U20934 (N_20934,N_14253,N_17784);
or U20935 (N_20935,N_17372,N_15413);
nor U20936 (N_20936,N_14685,N_16442);
nor U20937 (N_20937,N_17760,N_14739);
nor U20938 (N_20938,N_18719,N_18004);
or U20939 (N_20939,N_13816,N_18097);
nand U20940 (N_20940,N_13215,N_14456);
nand U20941 (N_20941,N_17628,N_14964);
and U20942 (N_20942,N_13827,N_14945);
and U20943 (N_20943,N_15961,N_13142);
or U20944 (N_20944,N_12823,N_13296);
xnor U20945 (N_20945,N_18498,N_18170);
nand U20946 (N_20946,N_13337,N_17037);
and U20947 (N_20947,N_17501,N_18707);
nor U20948 (N_20948,N_16758,N_17068);
nand U20949 (N_20949,N_16264,N_14108);
nand U20950 (N_20950,N_12539,N_12629);
nand U20951 (N_20951,N_13057,N_15922);
and U20952 (N_20952,N_17865,N_14238);
nor U20953 (N_20953,N_15481,N_14540);
and U20954 (N_20954,N_15970,N_15523);
or U20955 (N_20955,N_18331,N_15738);
nand U20956 (N_20956,N_15238,N_13001);
and U20957 (N_20957,N_12763,N_13549);
nor U20958 (N_20958,N_14374,N_13298);
nor U20959 (N_20959,N_13995,N_16527);
or U20960 (N_20960,N_14263,N_14980);
nand U20961 (N_20961,N_12835,N_18284);
nand U20962 (N_20962,N_17419,N_15447);
nor U20963 (N_20963,N_16132,N_15004);
nand U20964 (N_20964,N_18506,N_16507);
nor U20965 (N_20965,N_15716,N_14598);
and U20966 (N_20966,N_15010,N_16895);
nand U20967 (N_20967,N_18154,N_15134);
or U20968 (N_20968,N_12535,N_13106);
xnor U20969 (N_20969,N_17780,N_14733);
xor U20970 (N_20970,N_14786,N_17611);
nor U20971 (N_20971,N_13814,N_17464);
nand U20972 (N_20972,N_14099,N_14228);
nor U20973 (N_20973,N_17593,N_13173);
nand U20974 (N_20974,N_14399,N_18461);
nor U20975 (N_20975,N_18144,N_12927);
nor U20976 (N_20976,N_16690,N_14728);
nand U20977 (N_20977,N_16529,N_14888);
and U20978 (N_20978,N_15201,N_16092);
nor U20979 (N_20979,N_13443,N_12565);
or U20980 (N_20980,N_15619,N_16681);
or U20981 (N_20981,N_17825,N_13831);
or U20982 (N_20982,N_16462,N_17762);
xnor U20983 (N_20983,N_17143,N_13828);
and U20984 (N_20984,N_14345,N_14274);
xor U20985 (N_20985,N_14966,N_14063);
or U20986 (N_20986,N_13103,N_14543);
nand U20987 (N_20987,N_17478,N_15094);
and U20988 (N_20988,N_18116,N_17584);
and U20989 (N_20989,N_16759,N_13434);
or U20990 (N_20990,N_13605,N_12732);
nand U20991 (N_20991,N_14725,N_16550);
and U20992 (N_20992,N_12882,N_18673);
nand U20993 (N_20993,N_12592,N_13727);
and U20994 (N_20994,N_14918,N_17370);
nand U20995 (N_20995,N_17497,N_14049);
nor U20996 (N_20996,N_12554,N_18593);
and U20997 (N_20997,N_12755,N_18481);
or U20998 (N_20998,N_17616,N_16014);
nor U20999 (N_20999,N_15053,N_18126);
xnor U21000 (N_21000,N_13733,N_18134);
nor U21001 (N_21001,N_13905,N_16355);
nor U21002 (N_21002,N_16017,N_17741);
nor U21003 (N_21003,N_12940,N_13891);
nor U21004 (N_21004,N_15393,N_15829);
nor U21005 (N_21005,N_16409,N_16917);
nand U21006 (N_21006,N_12965,N_17183);
nand U21007 (N_21007,N_17655,N_16418);
nor U21008 (N_21008,N_13531,N_13026);
or U21009 (N_21009,N_16159,N_14667);
nand U21010 (N_21010,N_15282,N_13698);
and U21011 (N_21011,N_13820,N_18370);
and U21012 (N_21012,N_18465,N_12606);
and U21013 (N_21013,N_13330,N_16433);
nand U21014 (N_21014,N_17924,N_13687);
nand U21015 (N_21015,N_16055,N_14219);
nor U21016 (N_21016,N_17817,N_17048);
or U21017 (N_21017,N_15354,N_13580);
nor U21018 (N_21018,N_13778,N_14946);
and U21019 (N_21019,N_13702,N_13635);
or U21020 (N_21020,N_15453,N_16391);
nor U21021 (N_21021,N_14903,N_17065);
nor U21022 (N_21022,N_14332,N_18031);
and U21023 (N_21023,N_15362,N_13480);
nor U21024 (N_21024,N_13943,N_18388);
nor U21025 (N_21025,N_14453,N_16763);
or U21026 (N_21026,N_16113,N_16184);
and U21027 (N_21027,N_15153,N_15135);
nand U21028 (N_21028,N_13084,N_17046);
or U21029 (N_21029,N_17624,N_15275);
and U21030 (N_21030,N_16022,N_12871);
and U21031 (N_21031,N_18561,N_13239);
nor U21032 (N_21032,N_17875,N_12765);
or U21033 (N_21033,N_14454,N_17598);
nand U21034 (N_21034,N_14517,N_14948);
or U21035 (N_21035,N_18151,N_12961);
nor U21036 (N_21036,N_15486,N_15750);
xor U21037 (N_21037,N_13444,N_13870);
and U21038 (N_21038,N_16800,N_17945);
xnor U21039 (N_21039,N_16995,N_13947);
nand U21040 (N_21040,N_13581,N_18590);
xnor U21041 (N_21041,N_14663,N_16370);
and U21042 (N_21042,N_17052,N_17815);
or U21043 (N_21043,N_12697,N_16746);
nor U21044 (N_21044,N_18436,N_17635);
and U21045 (N_21045,N_16535,N_13288);
nor U21046 (N_21046,N_15111,N_13014);
and U21047 (N_21047,N_13976,N_13352);
nor U21048 (N_21048,N_16545,N_17318);
or U21049 (N_21049,N_17169,N_13446);
nand U21050 (N_21050,N_15550,N_13390);
and U21051 (N_21051,N_16646,N_15017);
and U21052 (N_21052,N_17185,N_15767);
nor U21053 (N_21053,N_14821,N_13088);
or U21054 (N_21054,N_18372,N_18219);
and U21055 (N_21055,N_18618,N_15087);
xor U21056 (N_21056,N_14703,N_18688);
or U21057 (N_21057,N_15643,N_17116);
nor U21058 (N_21058,N_13959,N_13176);
or U21059 (N_21059,N_17469,N_13004);
and U21060 (N_21060,N_16393,N_15542);
or U21061 (N_21061,N_18006,N_14375);
and U21062 (N_21062,N_14447,N_15046);
nor U21063 (N_21063,N_13752,N_13850);
nand U21064 (N_21064,N_13185,N_13358);
nor U21065 (N_21065,N_14350,N_14241);
xnor U21066 (N_21066,N_12529,N_16703);
and U21067 (N_21067,N_18450,N_17059);
or U21068 (N_21068,N_14639,N_18314);
or U21069 (N_21069,N_17957,N_16954);
nand U21070 (N_21070,N_15368,N_18490);
and U21071 (N_21071,N_17399,N_17132);
nor U21072 (N_21072,N_12767,N_12686);
nand U21073 (N_21073,N_14875,N_15511);
or U21074 (N_21074,N_15536,N_16728);
nand U21075 (N_21075,N_15166,N_18122);
or U21076 (N_21076,N_14356,N_14584);
xnor U21077 (N_21077,N_16223,N_17486);
and U21078 (N_21078,N_18638,N_14606);
nand U21079 (N_21079,N_12591,N_14804);
xor U21080 (N_21080,N_15577,N_14136);
nand U21081 (N_21081,N_17470,N_15240);
and U21082 (N_21082,N_15137,N_16714);
nor U21083 (N_21083,N_17535,N_13902);
and U21084 (N_21084,N_16577,N_14689);
xnor U21085 (N_21085,N_17359,N_16199);
or U21086 (N_21086,N_18087,N_17416);
or U21087 (N_21087,N_17783,N_13324);
or U21088 (N_21088,N_16906,N_16804);
nand U21089 (N_21089,N_14655,N_14361);
and U21090 (N_21090,N_18058,N_12933);
or U21091 (N_21091,N_13392,N_18073);
and U21092 (N_21092,N_15745,N_18271);
and U21093 (N_21093,N_13118,N_14581);
or U21094 (N_21094,N_17285,N_17282);
nand U21095 (N_21095,N_17343,N_16138);
nor U21096 (N_21096,N_14162,N_14451);
and U21097 (N_21097,N_13589,N_14073);
nand U21098 (N_21098,N_17657,N_16544);
or U21099 (N_21099,N_14200,N_12811);
xnor U21100 (N_21100,N_15748,N_14324);
nand U21101 (N_21101,N_13958,N_17465);
and U21102 (N_21102,N_16041,N_12645);
or U21103 (N_21103,N_17665,N_14771);
and U21104 (N_21104,N_16632,N_18644);
nand U21105 (N_21105,N_13241,N_16659);
and U21106 (N_21106,N_14321,N_13210);
nand U21107 (N_21107,N_12913,N_16773);
nand U21108 (N_21108,N_17461,N_17987);
or U21109 (N_21109,N_15943,N_13312);
nor U21110 (N_21110,N_14035,N_14847);
nand U21111 (N_21111,N_13128,N_14611);
nor U21112 (N_21112,N_14137,N_17223);
or U21113 (N_21113,N_13245,N_13242);
and U21114 (N_21114,N_15702,N_14528);
and U21115 (N_21115,N_18258,N_13325);
nor U21116 (N_21116,N_13459,N_17099);
or U21117 (N_21117,N_17531,N_13736);
and U21118 (N_21118,N_12687,N_15756);
nor U21119 (N_21119,N_14419,N_17172);
nor U21120 (N_21120,N_16546,N_17692);
and U21121 (N_21121,N_13170,N_15295);
nor U21122 (N_21122,N_12508,N_17664);
and U21123 (N_21123,N_15956,N_13811);
and U21124 (N_21124,N_16111,N_12622);
nor U21125 (N_21125,N_18090,N_14796);
and U21126 (N_21126,N_14116,N_17433);
nor U21127 (N_21127,N_13844,N_15083);
nand U21128 (N_21128,N_18268,N_16016);
and U21129 (N_21129,N_13692,N_12962);
nor U21130 (N_21130,N_18569,N_13772);
xnor U21131 (N_21131,N_18652,N_15418);
xor U21132 (N_21132,N_15454,N_17171);
nor U21133 (N_21133,N_17310,N_18141);
nor U21134 (N_21134,N_13932,N_12996);
nand U21135 (N_21135,N_17968,N_17288);
nand U21136 (N_21136,N_13725,N_12984);
xor U21137 (N_21137,N_13748,N_13815);
or U21138 (N_21138,N_15176,N_18231);
and U21139 (N_21139,N_18173,N_16072);
nor U21140 (N_21140,N_18617,N_16478);
and U21141 (N_21141,N_17368,N_17669);
and U21142 (N_21142,N_14576,N_17362);
and U21143 (N_21143,N_17823,N_14268);
nand U21144 (N_21144,N_15527,N_16855);
or U21145 (N_21145,N_17677,N_16607);
or U21146 (N_21146,N_12848,N_18395);
nor U21147 (N_21147,N_15744,N_15531);
or U21148 (N_21148,N_15937,N_15927);
and U21149 (N_21149,N_17695,N_13926);
nor U21150 (N_21150,N_15071,N_16314);
nor U21151 (N_21151,N_12920,N_18676);
nand U21152 (N_21152,N_18185,N_13411);
nand U21153 (N_21153,N_14115,N_15375);
or U21154 (N_21154,N_18375,N_17075);
nor U21155 (N_21155,N_17527,N_18382);
or U21156 (N_21156,N_14890,N_15392);
xor U21157 (N_21157,N_17026,N_15287);
nand U21158 (N_21158,N_18697,N_14215);
or U21159 (N_21159,N_17680,N_13204);
or U21160 (N_21160,N_13135,N_17747);
or U21161 (N_21161,N_13587,N_17155);
nand U21162 (N_21162,N_12537,N_18022);
and U21163 (N_21163,N_12796,N_12873);
xnor U21164 (N_21164,N_16342,N_17507);
nand U21165 (N_21165,N_18044,N_13939);
or U21166 (N_21166,N_15620,N_16932);
nand U21167 (N_21167,N_17959,N_15578);
nand U21168 (N_21168,N_15517,N_12986);
nand U21169 (N_21169,N_14956,N_15670);
and U21170 (N_21170,N_12937,N_14479);
nor U21171 (N_21171,N_17156,N_13303);
or U21172 (N_21172,N_14405,N_13343);
nor U21173 (N_21173,N_17750,N_16974);
and U21174 (N_21174,N_17667,N_16670);
nor U21175 (N_21175,N_16077,N_15853);
and U21176 (N_21176,N_16603,N_15926);
nor U21177 (N_21177,N_14712,N_18178);
nand U21178 (N_21178,N_13138,N_17729);
xor U21179 (N_21179,N_13089,N_12596);
nand U21180 (N_21180,N_15900,N_17400);
or U21181 (N_21181,N_16117,N_15992);
nor U21182 (N_21182,N_13756,N_18299);
or U21183 (N_21183,N_18190,N_16831);
nor U21184 (N_21184,N_12506,N_17590);
nor U21185 (N_21185,N_14414,N_14750);
nand U21186 (N_21186,N_15558,N_14344);
xnor U21187 (N_21187,N_13673,N_13904);
or U21188 (N_21188,N_14043,N_18502);
and U21189 (N_21189,N_17219,N_15367);
nand U21190 (N_21190,N_17529,N_16494);
or U21191 (N_21191,N_14962,N_15265);
nor U21192 (N_21192,N_13364,N_14392);
nor U21193 (N_21193,N_16777,N_13104);
and U21194 (N_21194,N_17256,N_16019);
and U21195 (N_21195,N_16109,N_17703);
nor U21196 (N_21196,N_17268,N_12709);
nand U21197 (N_21197,N_17843,N_14475);
or U21198 (N_21198,N_17830,N_16861);
or U21199 (N_21199,N_17562,N_14012);
and U21200 (N_21200,N_14745,N_13129);
and U21201 (N_21201,N_17713,N_16766);
and U21202 (N_21202,N_17653,N_15786);
xor U21203 (N_21203,N_14578,N_17415);
or U21204 (N_21204,N_14886,N_17962);
nand U21205 (N_21205,N_13615,N_15967);
nor U21206 (N_21206,N_15178,N_16290);
nor U21207 (N_21207,N_15280,N_16374);
or U21208 (N_21208,N_13611,N_16385);
and U21209 (N_21209,N_17176,N_13140);
or U21210 (N_21210,N_16853,N_16496);
xnor U21211 (N_21211,N_17341,N_18118);
nand U21212 (N_21212,N_18306,N_15815);
or U21213 (N_21213,N_13506,N_15743);
nand U21214 (N_21214,N_14342,N_18226);
and U21215 (N_21215,N_16018,N_15932);
nand U21216 (N_21216,N_16755,N_14717);
nand U21217 (N_21217,N_14221,N_14550);
or U21218 (N_21218,N_15497,N_14541);
nand U21219 (N_21219,N_17164,N_17435);
nand U21220 (N_21220,N_13591,N_14258);
nand U21221 (N_21221,N_14259,N_18664);
xnor U21222 (N_21222,N_13690,N_18285);
or U21223 (N_21223,N_17321,N_18386);
nand U21224 (N_21224,N_12656,N_15712);
or U21225 (N_21225,N_13415,N_15366);
or U21226 (N_21226,N_16543,N_13061);
nor U21227 (N_21227,N_14795,N_15843);
and U21228 (N_21228,N_14056,N_15121);
or U21229 (N_21229,N_17330,N_13829);
nor U21230 (N_21230,N_18608,N_14299);
nor U21231 (N_21231,N_15833,N_14757);
nand U21232 (N_21232,N_17744,N_15016);
or U21233 (N_21233,N_13576,N_13618);
nor U21234 (N_21234,N_16318,N_13254);
nand U21235 (N_21235,N_13311,N_15684);
nor U21236 (N_21236,N_17673,N_15880);
nor U21237 (N_21237,N_16719,N_16908);
nor U21238 (N_21238,N_18074,N_17521);
nor U21239 (N_21239,N_16595,N_15264);
nor U21240 (N_21240,N_16721,N_16713);
xnor U21241 (N_21241,N_15271,N_17722);
nand U21242 (N_21242,N_17743,N_16825);
or U21243 (N_21243,N_18101,N_17006);
xor U21244 (N_21244,N_17709,N_17561);
nor U21245 (N_21245,N_18243,N_18460);
or U21246 (N_21246,N_17512,N_14442);
or U21247 (N_21247,N_16352,N_14218);
nor U21248 (N_21248,N_13011,N_16930);
xor U21249 (N_21249,N_15090,N_12857);
nor U21250 (N_21250,N_12939,N_16511);
and U21251 (N_21251,N_17409,N_14232);
and U21252 (N_21252,N_18321,N_16394);
xor U21253 (N_21253,N_14450,N_17994);
and U21254 (N_21254,N_15723,N_15682);
xnor U21255 (N_21255,N_15069,N_18381);
xnor U21256 (N_21256,N_16848,N_13225);
nand U21257 (N_21257,N_15805,N_15382);
nand U21258 (N_21258,N_15537,N_18552);
or U21259 (N_21259,N_18620,N_13474);
xor U21260 (N_21260,N_14145,N_15839);
or U21261 (N_21261,N_16976,N_14231);
and U21262 (N_21262,N_15683,N_14325);
nand U21263 (N_21263,N_15618,N_13107);
and U21264 (N_21264,N_18254,N_14653);
nor U21265 (N_21265,N_15561,N_16641);
or U21266 (N_21266,N_17716,N_12738);
nor U21267 (N_21267,N_17778,N_17380);
and U21268 (N_21268,N_18571,N_13236);
and U21269 (N_21269,N_15548,N_16662);
or U21270 (N_21270,N_15426,N_12809);
nand U21271 (N_21271,N_16328,N_16481);
nor U21272 (N_21272,N_17481,N_13502);
or U21273 (N_21273,N_18079,N_16238);
and U21274 (N_21274,N_15492,N_18000);
xnor U21275 (N_21275,N_15524,N_13380);
nor U21276 (N_21276,N_16444,N_16555);
and U21277 (N_21277,N_13625,N_18112);
nand U21278 (N_21278,N_13087,N_17357);
nand U21279 (N_21279,N_18486,N_17807);
nor U21280 (N_21280,N_12832,N_15717);
nor U21281 (N_21281,N_16941,N_14245);
or U21282 (N_21282,N_17506,N_15846);
nor U21283 (N_21283,N_15616,N_12597);
nand U21284 (N_21284,N_18572,N_18259);
nor U21285 (N_21285,N_15252,N_14022);
nor U21286 (N_21286,N_15924,N_16813);
xor U21287 (N_21287,N_15726,N_12700);
nor U21288 (N_21288,N_18658,N_13055);
nor U21289 (N_21289,N_12812,N_13560);
nor U21290 (N_21290,N_13758,N_15975);
nor U21291 (N_21291,N_13223,N_18160);
nand U21292 (N_21292,N_15131,N_16299);
xnor U21293 (N_21293,N_14698,N_16033);
nor U21294 (N_21294,N_15198,N_17690);
nor U21295 (N_21295,N_14186,N_16015);
nor U21296 (N_21296,N_15341,N_16731);
nand U21297 (N_21297,N_15997,N_14617);
and U21298 (N_21298,N_14484,N_16044);
nor U21299 (N_21299,N_17350,N_18358);
xnor U21300 (N_21300,N_14844,N_14357);
and U21301 (N_21301,N_16038,N_18417);
and U21302 (N_21302,N_17972,N_15612);
or U21303 (N_21303,N_17594,N_17517);
or U21304 (N_21304,N_13628,N_13792);
or U21305 (N_21305,N_15361,N_16180);
and U21306 (N_21306,N_18582,N_14643);
nand U21307 (N_21307,N_17915,N_13871);
xnor U21308 (N_21308,N_16189,N_18532);
and U21309 (N_21309,N_16499,N_12917);
nor U21310 (N_21310,N_16309,N_17074);
nor U21311 (N_21311,N_17647,N_16970);
and U21312 (N_21312,N_17869,N_18513);
nor U21313 (N_21313,N_15607,N_16241);
nand U21314 (N_21314,N_18575,N_12869);
nor U21315 (N_21315,N_16279,N_18357);
xnor U21316 (N_21316,N_16648,N_17254);
nor U21317 (N_21317,N_16881,N_17031);
or U21318 (N_21318,N_13271,N_17356);
nand U21319 (N_21319,N_14066,N_17018);
and U21320 (N_21320,N_15261,N_14425);
nor U21321 (N_21321,N_13826,N_16288);
or U21322 (N_21322,N_13570,N_13062);
or U21323 (N_21323,N_17890,N_18339);
or U21324 (N_21324,N_13202,N_14064);
nor U21325 (N_21325,N_14317,N_18293);
nand U21326 (N_21326,N_14564,N_16186);
nand U21327 (N_21327,N_13278,N_14485);
nand U21328 (N_21328,N_15929,N_14290);
or U21329 (N_21329,N_14383,N_18400);
xnor U21330 (N_21330,N_13340,N_14351);
and U21331 (N_21331,N_18452,N_14206);
nor U21332 (N_21332,N_17141,N_17137);
or U21333 (N_21333,N_14686,N_14429);
and U21334 (N_21334,N_13246,N_15320);
and U21335 (N_21335,N_17482,N_13119);
and U21336 (N_21336,N_15115,N_15042);
and U21337 (N_21337,N_12504,N_16045);
nor U21338 (N_21338,N_17315,N_16426);
and U21339 (N_21339,N_17602,N_16849);
or U21340 (N_21340,N_14178,N_13529);
nand U21341 (N_21341,N_15685,N_14209);
or U21342 (N_21342,N_15795,N_16570);
or U21343 (N_21343,N_16233,N_14298);
xnor U21344 (N_21344,N_18246,N_14443);
or U21345 (N_21345,N_16346,N_17304);
nand U21346 (N_21346,N_12769,N_18560);
nor U21347 (N_21347,N_16211,N_16440);
and U21348 (N_21348,N_14873,N_16705);
and U21349 (N_21349,N_15038,N_18574);
or U21350 (N_21350,N_15147,N_13854);
and U21351 (N_21351,N_15985,N_17508);
or U21352 (N_21352,N_12828,N_17269);
nor U21353 (N_21353,N_12661,N_12947);
and U21354 (N_21354,N_16160,N_13349);
nor U21355 (N_21355,N_13230,N_13661);
or U21356 (N_21356,N_18380,N_15315);
nand U21357 (N_21357,N_12776,N_17948);
and U21358 (N_21358,N_15197,N_18174);
nand U21359 (N_21359,N_18105,N_14897);
or U21360 (N_21360,N_13481,N_12974);
and U21361 (N_21361,N_16399,N_15437);
nor U21362 (N_21362,N_17291,N_15803);
and U21363 (N_21363,N_17782,N_12891);
and U21364 (N_21364,N_17149,N_15605);
nand U21365 (N_21365,N_18124,N_18332);
nor U21366 (N_21366,N_16174,N_14402);
and U21367 (N_21367,N_14076,N_17976);
or U21368 (N_21368,N_16154,N_13417);
nor U21369 (N_21369,N_12674,N_15688);
or U21370 (N_21370,N_17963,N_13617);
nor U21371 (N_21371,N_13265,N_13191);
or U21372 (N_21372,N_17550,N_17572);
nand U21373 (N_21373,N_18367,N_15623);
nand U21374 (N_21374,N_16553,N_18316);
or U21375 (N_21375,N_17140,N_14535);
or U21376 (N_21376,N_18713,N_12854);
nor U21377 (N_21377,N_14121,N_13260);
or U21378 (N_21378,N_14680,N_13017);
xor U21379 (N_21379,N_12938,N_15412);
nand U21380 (N_21380,N_15869,N_13779);
and U21381 (N_21381,N_15251,N_17899);
nor U21382 (N_21382,N_18338,N_13317);
and U21383 (N_21383,N_14784,N_14778);
and U21384 (N_21384,N_14460,N_16781);
nand U21385 (N_21385,N_18662,N_15130);
nand U21386 (N_21386,N_12547,N_17661);
or U21387 (N_21387,N_12626,N_14622);
xor U21388 (N_21388,N_18046,N_17182);
nand U21389 (N_21389,N_15633,N_14156);
nand U21390 (N_21390,N_16774,N_12532);
xor U21391 (N_21391,N_17414,N_17175);
and U21392 (N_21392,N_15628,N_17796);
nor U21393 (N_21393,N_14254,N_12737);
nand U21394 (N_21394,N_15544,N_16871);
nand U21395 (N_21395,N_12735,N_14187);
nor U21396 (N_21396,N_16609,N_14348);
nand U21397 (N_21397,N_13237,N_16443);
nand U21398 (N_21398,N_14782,N_18615);
nor U21399 (N_21399,N_15841,N_18088);
and U21400 (N_21400,N_13656,N_16437);
or U21401 (N_21401,N_14669,N_18637);
or U21402 (N_21402,N_15194,N_12517);
nand U21403 (N_21403,N_17410,N_14671);
and U21404 (N_21404,N_16782,N_13550);
nand U21405 (N_21405,N_14797,N_13803);
xnor U21406 (N_21406,N_14164,N_14169);
nor U21407 (N_21407,N_18330,N_14112);
nand U21408 (N_21408,N_13117,N_13065);
and U21409 (N_21409,N_15760,N_13240);
nand U21410 (N_21410,N_12829,N_13624);
nor U21411 (N_21411,N_18312,N_17231);
nand U21412 (N_21412,N_14046,N_16469);
xor U21413 (N_21413,N_14309,N_16316);
nand U21414 (N_21414,N_15177,N_17964);
or U21415 (N_21415,N_13490,N_14953);
nor U21416 (N_21416,N_16720,N_12979);
and U21417 (N_21417,N_15930,N_15347);
or U21418 (N_21418,N_15938,N_13220);
nand U21419 (N_21419,N_18353,N_17579);
nor U21420 (N_21420,N_17460,N_12801);
nor U21421 (N_21421,N_18325,N_13842);
nand U21422 (N_21422,N_16903,N_14078);
xor U21423 (N_21423,N_17036,N_16068);
nor U21424 (N_21424,N_15114,N_17327);
xor U21425 (N_21425,N_14597,N_15817);
nor U21426 (N_21426,N_18542,N_17977);
xnor U21427 (N_21427,N_16412,N_17519);
nor U21428 (N_21428,N_13526,N_15552);
nand U21429 (N_21429,N_17913,N_16500);
nand U21430 (N_21430,N_14225,N_15666);
or U21431 (N_21431,N_16163,N_18619);
nor U21432 (N_21432,N_13894,N_13522);
nand U21433 (N_21433,N_16024,N_18095);
nand U21434 (N_21434,N_14999,N_12898);
and U21435 (N_21435,N_14131,N_14998);
and U21436 (N_21436,N_13114,N_13875);
xor U21437 (N_21437,N_12704,N_15568);
and U21438 (N_21438,N_18556,N_16194);
and U21439 (N_21439,N_16047,N_13613);
nand U21440 (N_21440,N_18737,N_18548);
nand U21441 (N_21441,N_14124,N_13316);
or U21442 (N_21442,N_16645,N_15196);
or U21443 (N_21443,N_13319,N_15674);
and U21444 (N_21444,N_18703,N_18686);
nor U21445 (N_21445,N_15553,N_16787);
and U21446 (N_21446,N_15777,N_18581);
nor U21447 (N_21447,N_18738,N_12590);
nor U21448 (N_21448,N_16811,N_14583);
and U21449 (N_21449,N_18492,N_18476);
nand U21450 (N_21450,N_15547,N_16329);
or U21451 (N_21451,N_12730,N_15344);
xnor U21452 (N_21452,N_18551,N_14489);
nor U21453 (N_21453,N_13266,N_14839);
and U21454 (N_21454,N_16754,N_14161);
nor U21455 (N_21455,N_16975,N_17200);
or U21456 (N_21456,N_17404,N_15720);
or U21457 (N_21457,N_17244,N_16733);
and U21458 (N_21458,N_18117,N_17305);
or U21459 (N_21459,N_17114,N_14824);
nand U21460 (N_21460,N_16498,N_13131);
nor U21461 (N_21461,N_18021,N_13003);
and U21462 (N_21462,N_16757,N_13849);
nor U21463 (N_21463,N_18495,N_15678);
nand U21464 (N_21464,N_15172,N_12505);
nor U21465 (N_21465,N_17645,N_15588);
xor U21466 (N_21466,N_12595,N_14607);
nor U21467 (N_21467,N_15583,N_15298);
and U21468 (N_21468,N_18188,N_17660);
nand U21469 (N_21469,N_14520,N_18347);
and U21470 (N_21470,N_17385,N_14666);
xor U21471 (N_21471,N_12778,N_13034);
nor U21472 (N_21472,N_17154,N_17764);
and U21473 (N_21473,N_18521,N_13835);
nor U21474 (N_21474,N_14972,N_16953);
or U21475 (N_21475,N_16337,N_13699);
or U21476 (N_21476,N_15936,N_12762);
and U21477 (N_21477,N_18322,N_13575);
nor U21478 (N_21478,N_15794,N_13249);
xor U21479 (N_21479,N_15233,N_13041);
xnor U21480 (N_21480,N_18191,N_15802);
and U21481 (N_21481,N_12909,N_18195);
or U21482 (N_21482,N_13269,N_12660);
nor U21483 (N_21483,N_16952,N_14285);
or U21484 (N_21484,N_18430,N_14949);
or U21485 (N_21485,N_18680,N_15476);
nand U21486 (N_21486,N_17698,N_16606);
and U21487 (N_21487,N_16451,N_13981);
or U21488 (N_21488,N_12786,N_17227);
or U21489 (N_21489,N_17596,N_13622);
nor U21490 (N_21490,N_15050,N_18405);
nor U21491 (N_21491,N_15742,N_15435);
nand U21492 (N_21492,N_15631,N_18309);
nor U21493 (N_21493,N_15423,N_12791);
nor U21494 (N_21494,N_16408,N_14691);
nand U21495 (N_21495,N_14138,N_16989);
nand U21496 (N_21496,N_17455,N_15220);
nand U21497 (N_21497,N_17477,N_15719);
or U21498 (N_21498,N_12889,N_13469);
xnor U21499 (N_21499,N_16027,N_17386);
nand U21500 (N_21500,N_16845,N_15826);
nor U21501 (N_21501,N_18295,N_17430);
or U21502 (N_21502,N_18108,N_16071);
nor U21503 (N_21503,N_14937,N_17608);
nand U21504 (N_21504,N_16591,N_15998);
and U21505 (N_21505,N_17911,N_13284);
and U21506 (N_21506,N_16192,N_15895);
nor U21507 (N_21507,N_16043,N_12711);
nor U21508 (N_21508,N_16411,N_17792);
and U21509 (N_21509,N_13322,N_16102);
xnor U21510 (N_21510,N_15248,N_17458);
nand U21511 (N_21511,N_14415,N_12630);
or U21512 (N_21512,N_16295,N_18228);
or U21513 (N_21513,N_15074,N_17453);
and U21514 (N_21514,N_16253,N_12969);
nor U21515 (N_21515,N_13962,N_14330);
nor U21516 (N_21516,N_17908,N_16673);
and U21517 (N_21517,N_17222,N_18724);
nor U21518 (N_21518,N_14970,N_15255);
or U21519 (N_21519,N_18438,N_16322);
xor U21520 (N_21520,N_18538,N_13571);
nor U21521 (N_21521,N_13335,N_13342);
nand U21522 (N_21522,N_12919,N_18494);
or U21523 (N_21523,N_18663,N_14882);
nand U21524 (N_21524,N_17827,N_17196);
nor U21525 (N_21525,N_14016,N_13761);
nor U21526 (N_21526,N_13799,N_17937);
xnor U21527 (N_21527,N_14142,N_14512);
nand U21528 (N_21528,N_13290,N_15405);
nand U21529 (N_21529,N_16164,N_17425);
nor U21530 (N_21530,N_18573,N_18041);
or U21531 (N_21531,N_16048,N_17377);
or U21532 (N_21532,N_15353,N_12754);
and U21533 (N_21533,N_16875,N_17440);
nand U21534 (N_21534,N_14455,N_14825);
nor U21535 (N_21535,N_12958,N_18049);
nand U21536 (N_21536,N_16929,N_16193);
or U21537 (N_21537,N_12693,N_15100);
nor U21538 (N_21538,N_15192,N_14659);
nor U21539 (N_21539,N_16525,N_14900);
or U21540 (N_21540,N_18068,N_17910);
or U21541 (N_21541,N_14701,N_13274);
nand U21542 (N_21542,N_12688,N_13556);
xnor U21543 (N_21543,N_15309,N_15727);
nand U21544 (N_21544,N_16325,N_12888);
nand U21545 (N_21545,N_15969,N_13229);
or U21546 (N_21546,N_15445,N_15785);
nor U21547 (N_21547,N_17035,N_15814);
xor U21548 (N_21548,N_17619,N_16587);
and U21549 (N_21549,N_12836,N_15904);
nor U21550 (N_21550,N_17605,N_18287);
nor U21551 (N_21551,N_16824,N_17094);
nand U21552 (N_21552,N_18640,N_16294);
nand U21553 (N_21553,N_14412,N_14851);
nand U21554 (N_21554,N_18094,N_13453);
nand U21555 (N_21555,N_16167,N_17032);
and U21556 (N_21556,N_14401,N_13385);
xor U21557 (N_21557,N_17721,N_16820);
nand U21558 (N_21558,N_17439,N_15420);
or U21559 (N_21559,N_18645,N_15059);
or U21560 (N_21560,N_14947,N_14490);
and U21561 (N_21561,N_15103,N_14802);
nor U21562 (N_21562,N_16176,N_14474);
or U21563 (N_21563,N_13458,N_14032);
nor U21564 (N_21564,N_15330,N_12558);
or U21565 (N_21565,N_17102,N_14861);
xor U21566 (N_21566,N_14586,N_16298);
nand U21567 (N_21567,N_18233,N_14417);
nand U21568 (N_21568,N_15005,N_17274);
and U21569 (N_21569,N_13047,N_16367);
nand U21570 (N_21570,N_12768,N_16195);
and U21571 (N_21571,N_13218,N_12540);
nand U21572 (N_21572,N_13461,N_14368);
and U21573 (N_21573,N_15190,N_16589);
nor U21574 (N_21574,N_15199,N_15934);
xor U21575 (N_21575,N_16246,N_18272);
xor U21576 (N_21576,N_13005,N_12989);
xor U21577 (N_21577,N_18300,N_15307);
and U21578 (N_21578,N_12751,N_13917);
nand U21579 (N_21579,N_17097,N_16081);
or U21580 (N_21580,N_12766,N_13152);
or U21581 (N_21581,N_15571,N_13649);
nand U21582 (N_21582,N_17159,N_14306);
or U21583 (N_21583,N_14278,N_13413);
or U21584 (N_21584,N_17273,N_13420);
nand U21585 (N_21585,N_14819,N_13839);
and U21586 (N_21586,N_14143,N_15582);
nand U21587 (N_21587,N_18350,N_17772);
or U21588 (N_21588,N_14239,N_18447);
nor U21589 (N_21589,N_17834,N_15954);
xnor U21590 (N_21590,N_18368,N_12839);
nor U21591 (N_21591,N_16097,N_15897);
nand U21592 (N_21592,N_13859,N_17944);
nor U21593 (N_21593,N_13085,N_15501);
and U21594 (N_21594,N_16473,N_15487);
nor U21595 (N_21595,N_15529,N_16214);
nor U21596 (N_21596,N_12739,N_15055);
or U21597 (N_21597,N_14944,N_15945);
nor U21598 (N_21598,N_16447,N_13508);
or U21599 (N_21599,N_15509,N_15856);
and U21600 (N_21600,N_17123,N_17719);
or U21601 (N_21601,N_16263,N_14262);
nor U21602 (N_21602,N_14603,N_14077);
nand U21603 (N_21603,N_17180,N_17770);
or U21604 (N_21604,N_14478,N_15365);
and U21605 (N_21605,N_12842,N_16148);
nor U21606 (N_21606,N_15316,N_14158);
or U21607 (N_21607,N_15409,N_15136);
nor U21608 (N_21608,N_13180,N_15302);
and U21609 (N_21609,N_13196,N_16339);
or U21610 (N_21610,N_17927,N_15180);
nor U21611 (N_21611,N_13074,N_16660);
nand U21612 (N_21612,N_16321,N_16136);
or U21613 (N_21613,N_18297,N_13889);
nor U21614 (N_21614,N_12890,N_13059);
nor U21615 (N_21615,N_16990,N_14501);
nor U21616 (N_21616,N_18247,N_15461);
nand U21617 (N_21617,N_18159,N_14816);
xnor U21618 (N_21618,N_14155,N_17205);
or U21619 (N_21619,N_13097,N_18699);
and U21620 (N_21620,N_16519,N_17281);
nor U21621 (N_21621,N_12710,N_15066);
nand U21622 (N_21622,N_17135,N_14763);
and U21623 (N_21623,N_14091,N_17623);
nor U21624 (N_21624,N_15097,N_13619);
or U21625 (N_21625,N_12620,N_14828);
nor U21626 (N_21626,N_16928,N_17884);
nor U21627 (N_21627,N_17240,N_13652);
or U21628 (N_21628,N_16086,N_16576);
or U21629 (N_21629,N_12745,N_16268);
or U21630 (N_21630,N_18420,N_15081);
and U21631 (N_21631,N_16270,N_18263);
nand U21632 (N_21632,N_14885,N_17787);
nor U21633 (N_21633,N_18334,N_13742);
nor U21634 (N_21634,N_16064,N_15422);
or U21635 (N_21635,N_12973,N_18392);
or U21636 (N_21636,N_17253,N_14362);
nand U21637 (N_21637,N_15456,N_18675);
and U21638 (N_21638,N_18650,N_14095);
nor U21639 (N_21639,N_14874,N_14487);
and U21640 (N_21640,N_13067,N_12534);
and U21641 (N_21641,N_13109,N_18286);
nor U21642 (N_21642,N_17092,N_13370);
nand U21643 (N_21643,N_18588,N_16797);
or U21644 (N_21644,N_16287,N_16076);
nand U21645 (N_21645,N_18563,N_16984);
and U21646 (N_21646,N_13029,N_15379);
and U21647 (N_21647,N_13969,N_15132);
and U21648 (N_21648,N_17809,N_14377);
nor U21649 (N_21649,N_13539,N_14766);
or U21650 (N_21650,N_17684,N_16488);
nand U21651 (N_21651,N_16987,N_14985);
or U21652 (N_21652,N_15835,N_15693);
nand U21653 (N_21653,N_14154,N_15391);
nand U21654 (N_21654,N_12956,N_13558);
nand U21655 (N_21655,N_15689,N_15893);
nand U21656 (N_21656,N_17083,N_13554);
xor U21657 (N_21657,N_18397,N_17993);
and U21658 (N_21658,N_14902,N_14848);
nor U21659 (N_21659,N_18024,N_12557);
nand U21660 (N_21660,N_14141,N_13940);
or U21661 (N_21661,N_18626,N_18407);
or U21662 (N_21662,N_18510,N_15881);
and U21663 (N_21663,N_14326,N_13487);
or U21664 (N_21664,N_18223,N_16639);
and U21665 (N_21665,N_16548,N_17991);
nor U21666 (N_21666,N_15206,N_15947);
nor U21667 (N_21667,N_13393,N_16918);
nor U21668 (N_21668,N_14021,N_16772);
and U21669 (N_21669,N_16794,N_14042);
or U21670 (N_21670,N_14907,N_13157);
nand U21671 (N_21671,N_13145,N_17820);
nand U21672 (N_21672,N_18260,N_16889);
nand U21673 (N_21673,N_12695,N_14927);
or U21674 (N_21674,N_15849,N_16216);
nand U21675 (N_21675,N_16032,N_14409);
or U21676 (N_21676,N_14604,N_17294);
and U21677 (N_21677,N_13437,N_12567);
nor U21678 (N_21678,N_12761,N_17599);
or U21679 (N_21679,N_13308,N_15179);
and U21680 (N_21680,N_15239,N_15120);
and U21681 (N_21681,N_18580,N_13978);
nor U21682 (N_21682,N_16832,N_18139);
or U21683 (N_21683,N_15186,N_18147);
or U21684 (N_21684,N_13261,N_18168);
and U21685 (N_21685,N_14349,N_16127);
and U21686 (N_21686,N_14670,N_16300);
or U21687 (N_21687,N_14790,N_16950);
nand U21688 (N_21688,N_15460,N_16685);
and U21689 (N_21689,N_14139,N_13667);
nand U21690 (N_21690,N_13785,N_12559);
or U21691 (N_21691,N_16934,N_14510);
or U21692 (N_21692,N_18477,N_13077);
and U21693 (N_21693,N_16869,N_17237);
nor U21694 (N_21694,N_15538,N_12715);
and U21695 (N_21695,N_17543,N_15228);
nor U21696 (N_21696,N_17081,N_15708);
or U21697 (N_21697,N_18238,N_14589);
and U21698 (N_21698,N_13197,N_14923);
and U21699 (N_21699,N_15885,N_16541);
nor U21700 (N_21700,N_17360,N_13160);
nand U21701 (N_21701,N_13315,N_14523);
nand U21702 (N_21702,N_13383,N_14706);
and U21703 (N_21703,N_14308,N_16716);
and U21704 (N_21704,N_15030,N_14462);
and U21705 (N_21705,N_18113,N_18387);
and U21706 (N_21706,N_13177,N_16388);
xnor U21707 (N_21707,N_14880,N_13167);
nor U21708 (N_21708,N_18511,N_15988);
nor U21709 (N_21709,N_14051,N_16327);
xor U21710 (N_21710,N_17988,N_13512);
nand U21711 (N_21711,N_17775,N_16982);
nor U21712 (N_21712,N_17978,N_17479);
and U21713 (N_21713,N_14171,N_13954);
nand U21714 (N_21714,N_16658,N_17861);
nand U21715 (N_21715,N_18549,N_18433);
xnor U21716 (N_21716,N_13081,N_15442);
nor U21717 (N_21717,N_14682,N_15838);
or U21718 (N_21718,N_14732,N_16504);
nor U21719 (N_21719,N_18212,N_15701);
and U21720 (N_21720,N_16736,N_15592);
nand U21721 (N_21721,N_16945,N_14826);
and U21722 (N_21722,N_12635,N_14113);
nand U21723 (N_21723,N_12684,N_18361);
nand U21724 (N_21724,N_16273,N_15077);
nor U21725 (N_21725,N_14463,N_15021);
xor U21726 (N_21726,N_15574,N_15556);
xnor U21727 (N_21727,N_17467,N_18059);
and U21728 (N_21728,N_15035,N_13397);
or U21729 (N_21729,N_18406,N_15079);
xnor U21730 (N_21730,N_16369,N_18179);
nor U21731 (N_21731,N_14881,N_17516);
and U21732 (N_21732,N_14871,N_15043);
and U21733 (N_21733,N_17369,N_13648);
xor U21734 (N_21734,N_15984,N_13765);
or U21735 (N_21735,N_18038,N_13009);
and U21736 (N_21736,N_13405,N_17129);
or U21737 (N_21737,N_13491,N_13285);
or U21738 (N_21738,N_16157,N_17798);
and U21739 (N_21739,N_16980,N_16034);
and U21740 (N_21740,N_18320,N_13596);
or U21741 (N_21741,N_16973,N_18165);
nand U21742 (N_21742,N_13247,N_17876);
nand U21743 (N_21743,N_14679,N_15690);
nand U21744 (N_21744,N_14391,N_14092);
xor U21745 (N_21745,N_13830,N_17234);
nand U21746 (N_21746,N_12741,N_14645);
or U21747 (N_21747,N_17510,N_12585);
or U21748 (N_21748,N_15149,N_15374);
nand U21749 (N_21749,N_12724,N_13903);
nor U21750 (N_21750,N_14177,N_15609);
or U21751 (N_21751,N_16191,N_13933);
nand U21752 (N_21752,N_15001,N_16364);
nand U21753 (N_21753,N_12777,N_15480);
and U21754 (N_21754,N_14216,N_15580);
or U21755 (N_21755,N_13760,N_16505);
or U21756 (N_21756,N_17902,N_17131);
or U21757 (N_21757,N_12804,N_15694);
xnor U21758 (N_21758,N_15774,N_18181);
nand U21759 (N_21759,N_16070,N_16235);
nor U21760 (N_21760,N_15686,N_15533);
or U21761 (N_21761,N_13064,N_14006);
nand U21762 (N_21762,N_16823,N_16169);
or U21763 (N_21763,N_16147,N_16390);
and U21764 (N_21764,N_16819,N_18547);
nand U21765 (N_21765,N_17402,N_16907);
nor U21766 (N_21766,N_13035,N_14398);
xor U21767 (N_21767,N_15792,N_16593);
or U21768 (N_21768,N_15205,N_15865);
nor U21769 (N_21769,N_12959,N_16812);
or U21770 (N_21770,N_12524,N_15941);
or U21771 (N_21771,N_14973,N_13774);
and U21772 (N_21772,N_14480,N_14657);
nor U21773 (N_21773,N_18404,N_16625);
and U21774 (N_21774,N_14387,N_17475);
and U21775 (N_21775,N_18631,N_15733);
nand U21776 (N_21776,N_17901,N_14855);
xnor U21777 (N_21777,N_18075,N_16345);
xor U21778 (N_21778,N_17252,N_16857);
or U21779 (N_21779,N_16297,N_13262);
or U21780 (N_21780,N_16904,N_16602);
and U21781 (N_21781,N_17574,N_12968);
and U21782 (N_21782,N_18045,N_15155);
xor U21783 (N_21783,N_13253,N_15641);
nor U21784 (N_21784,N_12816,N_15763);
nand U21785 (N_21785,N_15778,N_18354);
xnor U21786 (N_21786,N_18427,N_18010);
nor U21787 (N_21787,N_17264,N_15788);
or U21788 (N_21788,N_15241,N_12822);
nor U21789 (N_21789,N_14638,N_17766);
xor U21790 (N_21790,N_13255,N_12970);
nand U21791 (N_21791,N_18018,N_15165);
and U21792 (N_21792,N_14134,N_14013);
or U21793 (N_21793,N_14044,N_12810);
or U21794 (N_21794,N_17804,N_16285);
nor U21795 (N_21795,N_12921,N_16618);
nand U21796 (N_21796,N_12563,N_16561);
and U21797 (N_21797,N_16248,N_14694);
or U21798 (N_21798,N_15332,N_17204);
or U21799 (N_21799,N_17781,N_16877);
nor U21800 (N_21800,N_12669,N_18520);
nand U21801 (N_21801,N_18385,N_18586);
nor U21802 (N_21802,N_15054,N_16741);
or U21803 (N_21803,N_16089,N_16756);
nand U21804 (N_21804,N_15122,N_14312);
nand U21805 (N_21805,N_17808,N_16638);
nor U21806 (N_21806,N_15773,N_17441);
nand U21807 (N_21807,N_13115,N_13130);
and U21808 (N_21808,N_16340,N_12586);
nand U21809 (N_21809,N_17296,N_14188);
nand U21810 (N_21810,N_13741,N_15964);
or U21811 (N_21811,N_13462,N_16669);
nor U21812 (N_21812,N_18654,N_13906);
xnor U21813 (N_21813,N_15285,N_15463);
nand U21814 (N_21814,N_14323,N_14109);
or U21815 (N_21815,N_13657,N_17002);
or U21816 (N_21816,N_12914,N_13251);
nand U21817 (N_21817,N_13768,N_14575);
xor U21818 (N_21818,N_14010,N_16410);
nor U21819 (N_21819,N_13072,N_15440);
nor U21820 (N_21820,N_17984,N_16865);
nor U21821 (N_21821,N_17802,N_17857);
nand U21822 (N_21822,N_15381,N_15470);
nand U21823 (N_21823,N_13945,N_14005);
or U21824 (N_21824,N_18709,N_17086);
nor U21825 (N_21825,N_17907,N_14870);
or U21826 (N_21826,N_16257,N_17999);
and U21827 (N_21827,N_13689,N_15161);
or U21828 (N_21828,N_15752,N_13682);
and U21829 (N_21829,N_17034,N_15356);
and U21830 (N_21830,N_13713,N_17457);
nor U21831 (N_21831,N_16686,N_18717);
and U21832 (N_21832,N_14061,N_15806);
and U21833 (N_21833,N_15051,N_13674);
xor U21834 (N_21834,N_15779,N_12764);
xor U21835 (N_21835,N_14287,N_16572);
xnor U21836 (N_21836,N_13655,N_15193);
nor U21837 (N_21837,N_17450,N_16663);
nor U21838 (N_21838,N_18336,N_15654);
nand U21839 (N_21839,N_18716,N_14192);
nand U21840 (N_21840,N_17413,N_15933);
or U21841 (N_21841,N_12617,N_15818);
nand U21842 (N_21842,N_17365,N_17500);
and U21843 (N_21843,N_13614,N_17542);
and U21844 (N_21844,N_13154,N_17541);
xor U21845 (N_21845,N_17301,N_14814);
and U21846 (N_21846,N_15905,N_12612);
nand U21847 (N_21847,N_13208,N_12593);
and U21848 (N_21848,N_17139,N_15782);
or U21849 (N_21849,N_14476,N_13222);
or U21850 (N_21850,N_12708,N_15862);
nor U21851 (N_21851,N_17578,N_17442);
nor U21852 (N_21852,N_16067,N_15827);
or U21853 (N_21853,N_18206,N_17776);
nor U21854 (N_21854,N_18203,N_15462);
nor U21855 (N_21855,N_18668,N_13564);
and U21856 (N_21856,N_17558,N_16640);
nor U21857 (N_21857,N_13378,N_15707);
nand U21858 (N_21858,N_18069,N_16793);
or U21859 (N_21859,N_18536,N_15543);
and U21860 (N_21860,N_14580,N_17539);
xnor U21861 (N_21861,N_16031,N_13921);
xnor U21862 (N_21862,N_17752,N_18081);
and U21863 (N_21863,N_14552,N_15482);
xor U21864 (N_21864,N_14340,N_14052);
and U21865 (N_21865,N_17971,N_13421);
or U21866 (N_21866,N_13963,N_14191);
and U21867 (N_21867,N_13082,N_13775);
nand U21868 (N_21868,N_16477,N_17103);
and U21869 (N_21869,N_12872,N_14483);
or U21870 (N_21870,N_15830,N_17940);
nand U21871 (N_21871,N_18161,N_13524);
or U21872 (N_21872,N_14058,N_16128);
xor U21873 (N_21873,N_17785,N_12679);
nand U21874 (N_21874,N_18020,N_16126);
xnor U21875 (N_21875,N_15545,N_13008);
or U21876 (N_21876,N_18544,N_16666);
xor U21877 (N_21877,N_14936,N_18138);
nand U21878 (N_21878,N_15786,N_13352);
nand U21879 (N_21879,N_15642,N_16609);
and U21880 (N_21880,N_16061,N_15322);
nand U21881 (N_21881,N_15612,N_14659);
or U21882 (N_21882,N_12610,N_16112);
nand U21883 (N_21883,N_18478,N_14403);
and U21884 (N_21884,N_13118,N_14900);
and U21885 (N_21885,N_13487,N_15668);
or U21886 (N_21886,N_18111,N_17977);
and U21887 (N_21887,N_14554,N_13080);
nand U21888 (N_21888,N_17197,N_18085);
and U21889 (N_21889,N_15918,N_13089);
nand U21890 (N_21890,N_14763,N_17289);
nor U21891 (N_21891,N_15591,N_18063);
and U21892 (N_21892,N_12816,N_16356);
nand U21893 (N_21893,N_17225,N_16700);
or U21894 (N_21894,N_13666,N_16565);
xor U21895 (N_21895,N_14283,N_16588);
and U21896 (N_21896,N_16518,N_13073);
nor U21897 (N_21897,N_16542,N_13658);
nor U21898 (N_21898,N_16387,N_13936);
and U21899 (N_21899,N_18373,N_16189);
xnor U21900 (N_21900,N_16947,N_13912);
or U21901 (N_21901,N_16465,N_13423);
and U21902 (N_21902,N_16887,N_14021);
nand U21903 (N_21903,N_17142,N_17110);
nor U21904 (N_21904,N_17942,N_12621);
and U21905 (N_21905,N_16562,N_17587);
and U21906 (N_21906,N_17034,N_14336);
and U21907 (N_21907,N_16057,N_13551);
xnor U21908 (N_21908,N_18254,N_12626);
nand U21909 (N_21909,N_14723,N_17343);
nor U21910 (N_21910,N_13373,N_16967);
or U21911 (N_21911,N_13086,N_13169);
or U21912 (N_21912,N_15658,N_15277);
nand U21913 (N_21913,N_18146,N_15242);
nor U21914 (N_21914,N_16816,N_17284);
nand U21915 (N_21915,N_16995,N_14685);
nand U21916 (N_21916,N_13697,N_12737);
nand U21917 (N_21917,N_14750,N_14725);
nor U21918 (N_21918,N_16505,N_15998);
nand U21919 (N_21919,N_16115,N_17997);
or U21920 (N_21920,N_13702,N_17968);
nor U21921 (N_21921,N_17397,N_12775);
and U21922 (N_21922,N_14082,N_13603);
and U21923 (N_21923,N_13945,N_13151);
or U21924 (N_21924,N_18415,N_16693);
nand U21925 (N_21925,N_17822,N_15212);
or U21926 (N_21926,N_13868,N_12985);
or U21927 (N_21927,N_14328,N_13533);
and U21928 (N_21928,N_15488,N_13982);
nand U21929 (N_21929,N_13243,N_17316);
and U21930 (N_21930,N_17769,N_15523);
and U21931 (N_21931,N_15216,N_17989);
or U21932 (N_21932,N_15515,N_16079);
nand U21933 (N_21933,N_13164,N_15715);
nor U21934 (N_21934,N_15177,N_15879);
and U21935 (N_21935,N_16120,N_14642);
and U21936 (N_21936,N_16034,N_16834);
nand U21937 (N_21937,N_16760,N_12756);
nor U21938 (N_21938,N_18161,N_14083);
xnor U21939 (N_21939,N_16984,N_16702);
nand U21940 (N_21940,N_15891,N_12736);
and U21941 (N_21941,N_17918,N_16775);
nor U21942 (N_21942,N_13680,N_15579);
or U21943 (N_21943,N_16512,N_14517);
nand U21944 (N_21944,N_15128,N_13209);
xor U21945 (N_21945,N_16644,N_15263);
nor U21946 (N_21946,N_17661,N_12987);
nor U21947 (N_21947,N_14247,N_16461);
and U21948 (N_21948,N_13809,N_15484);
nor U21949 (N_21949,N_17985,N_16612);
or U21950 (N_21950,N_15545,N_15408);
or U21951 (N_21951,N_14477,N_15563);
and U21952 (N_21952,N_14086,N_15383);
nor U21953 (N_21953,N_16748,N_14811);
nand U21954 (N_21954,N_15723,N_13092);
and U21955 (N_21955,N_14345,N_15841);
nor U21956 (N_21956,N_18106,N_17127);
xnor U21957 (N_21957,N_16248,N_14921);
or U21958 (N_21958,N_18329,N_17658);
or U21959 (N_21959,N_12904,N_15769);
nand U21960 (N_21960,N_13991,N_14646);
nand U21961 (N_21961,N_17564,N_12825);
nor U21962 (N_21962,N_16343,N_13049);
nand U21963 (N_21963,N_15133,N_17121);
nand U21964 (N_21964,N_18533,N_14431);
or U21965 (N_21965,N_13975,N_15301);
and U21966 (N_21966,N_17294,N_15297);
and U21967 (N_21967,N_16851,N_17500);
and U21968 (N_21968,N_16888,N_14219);
and U21969 (N_21969,N_13797,N_12893);
nand U21970 (N_21970,N_16592,N_17695);
and U21971 (N_21971,N_14465,N_15421);
xor U21972 (N_21972,N_14901,N_16942);
nand U21973 (N_21973,N_13617,N_16427);
or U21974 (N_21974,N_16885,N_16458);
nor U21975 (N_21975,N_15051,N_18694);
nand U21976 (N_21976,N_13128,N_14973);
nand U21977 (N_21977,N_15876,N_13610);
xor U21978 (N_21978,N_16345,N_17731);
and U21979 (N_21979,N_13230,N_17926);
nand U21980 (N_21980,N_14827,N_13125);
nor U21981 (N_21981,N_18180,N_12880);
xnor U21982 (N_21982,N_18225,N_13548);
nor U21983 (N_21983,N_16574,N_17833);
or U21984 (N_21984,N_15510,N_14944);
and U21985 (N_21985,N_18572,N_13855);
or U21986 (N_21986,N_13830,N_13270);
or U21987 (N_21987,N_13733,N_12770);
nand U21988 (N_21988,N_18406,N_18692);
and U21989 (N_21989,N_16365,N_13266);
nor U21990 (N_21990,N_14346,N_13401);
xor U21991 (N_21991,N_16262,N_17222);
nand U21992 (N_21992,N_15390,N_16494);
nor U21993 (N_21993,N_14924,N_14820);
or U21994 (N_21994,N_13610,N_17849);
nand U21995 (N_21995,N_14261,N_14014);
nor U21996 (N_21996,N_17615,N_13461);
and U21997 (N_21997,N_12822,N_14947);
xor U21998 (N_21998,N_14592,N_14155);
and U21999 (N_21999,N_17364,N_16890);
or U22000 (N_22000,N_17586,N_12884);
nand U22001 (N_22001,N_13329,N_13326);
or U22002 (N_22002,N_17868,N_13609);
and U22003 (N_22003,N_17042,N_17935);
nor U22004 (N_22004,N_16493,N_16189);
nor U22005 (N_22005,N_15173,N_18628);
nor U22006 (N_22006,N_18183,N_13281);
or U22007 (N_22007,N_13162,N_16504);
nor U22008 (N_22008,N_17399,N_16657);
and U22009 (N_22009,N_17202,N_18488);
nor U22010 (N_22010,N_13774,N_15706);
nand U22011 (N_22011,N_17814,N_17670);
or U22012 (N_22012,N_14468,N_16734);
xor U22013 (N_22013,N_14473,N_16430);
and U22014 (N_22014,N_18511,N_17253);
or U22015 (N_22015,N_15472,N_15477);
nand U22016 (N_22016,N_16635,N_13461);
nor U22017 (N_22017,N_16716,N_14819);
or U22018 (N_22018,N_15481,N_12864);
and U22019 (N_22019,N_14384,N_17683);
and U22020 (N_22020,N_14699,N_18276);
and U22021 (N_22021,N_12663,N_15074);
nor U22022 (N_22022,N_13138,N_14498);
nor U22023 (N_22023,N_16615,N_12885);
or U22024 (N_22024,N_14566,N_17177);
nor U22025 (N_22025,N_16380,N_14338);
xor U22026 (N_22026,N_13320,N_17413);
or U22027 (N_22027,N_17630,N_17199);
or U22028 (N_22028,N_16305,N_18179);
nand U22029 (N_22029,N_13780,N_12591);
and U22030 (N_22030,N_15288,N_18397);
nor U22031 (N_22031,N_17842,N_18271);
nor U22032 (N_22032,N_15103,N_15714);
or U22033 (N_22033,N_18265,N_14005);
or U22034 (N_22034,N_13729,N_15777);
and U22035 (N_22035,N_18389,N_16914);
or U22036 (N_22036,N_13060,N_16561);
nor U22037 (N_22037,N_14566,N_12608);
or U22038 (N_22038,N_12978,N_17494);
and U22039 (N_22039,N_18692,N_13235);
xor U22040 (N_22040,N_14046,N_16647);
nor U22041 (N_22041,N_17620,N_15287);
nor U22042 (N_22042,N_16625,N_12692);
xnor U22043 (N_22043,N_16077,N_15488);
nand U22044 (N_22044,N_15708,N_17808);
or U22045 (N_22045,N_13359,N_15370);
xor U22046 (N_22046,N_15058,N_17593);
nand U22047 (N_22047,N_18663,N_14038);
and U22048 (N_22048,N_18202,N_16717);
or U22049 (N_22049,N_16055,N_13252);
nor U22050 (N_22050,N_14176,N_17742);
nand U22051 (N_22051,N_15445,N_16733);
nand U22052 (N_22052,N_13447,N_13323);
nor U22053 (N_22053,N_15123,N_14248);
or U22054 (N_22054,N_12522,N_17535);
nand U22055 (N_22055,N_15117,N_16454);
nor U22056 (N_22056,N_18442,N_15843);
nand U22057 (N_22057,N_14857,N_12940);
nor U22058 (N_22058,N_14531,N_18134);
or U22059 (N_22059,N_13763,N_18184);
nor U22060 (N_22060,N_17377,N_13001);
or U22061 (N_22061,N_18635,N_17065);
and U22062 (N_22062,N_15465,N_17106);
nor U22063 (N_22063,N_14001,N_17560);
nor U22064 (N_22064,N_18090,N_17645);
nand U22065 (N_22065,N_14935,N_13609);
or U22066 (N_22066,N_18255,N_13647);
nand U22067 (N_22067,N_16364,N_18604);
nand U22068 (N_22068,N_18131,N_15063);
nand U22069 (N_22069,N_17744,N_13817);
or U22070 (N_22070,N_17677,N_14233);
or U22071 (N_22071,N_14304,N_13560);
nor U22072 (N_22072,N_14439,N_13335);
nand U22073 (N_22073,N_17982,N_13764);
or U22074 (N_22074,N_16175,N_13410);
and U22075 (N_22075,N_14357,N_14158);
nor U22076 (N_22076,N_14535,N_17497);
nor U22077 (N_22077,N_16402,N_16934);
or U22078 (N_22078,N_18178,N_14073);
xnor U22079 (N_22079,N_17629,N_13098);
or U22080 (N_22080,N_14094,N_15273);
xnor U22081 (N_22081,N_13285,N_17905);
or U22082 (N_22082,N_18170,N_16996);
nand U22083 (N_22083,N_16489,N_18377);
and U22084 (N_22084,N_14917,N_17169);
nor U22085 (N_22085,N_18356,N_13927);
nand U22086 (N_22086,N_18118,N_14552);
and U22087 (N_22087,N_14417,N_14384);
or U22088 (N_22088,N_17060,N_15570);
and U22089 (N_22089,N_15267,N_15412);
and U22090 (N_22090,N_17365,N_18581);
and U22091 (N_22091,N_17078,N_16475);
and U22092 (N_22092,N_14712,N_13958);
xor U22093 (N_22093,N_13727,N_14100);
xor U22094 (N_22094,N_14648,N_15859);
or U22095 (N_22095,N_15366,N_17743);
nand U22096 (N_22096,N_15523,N_18368);
nand U22097 (N_22097,N_13145,N_14087);
and U22098 (N_22098,N_15603,N_14487);
nand U22099 (N_22099,N_16997,N_17262);
nand U22100 (N_22100,N_13874,N_14113);
or U22101 (N_22101,N_17467,N_12529);
and U22102 (N_22102,N_15210,N_16263);
nand U22103 (N_22103,N_15051,N_18105);
and U22104 (N_22104,N_18372,N_12832);
nor U22105 (N_22105,N_17875,N_18326);
or U22106 (N_22106,N_17007,N_12536);
and U22107 (N_22107,N_15185,N_16930);
nand U22108 (N_22108,N_13611,N_17434);
nor U22109 (N_22109,N_15783,N_13930);
nand U22110 (N_22110,N_18466,N_17107);
nor U22111 (N_22111,N_16217,N_16667);
nand U22112 (N_22112,N_16743,N_13038);
and U22113 (N_22113,N_15580,N_13053);
nand U22114 (N_22114,N_14735,N_17340);
or U22115 (N_22115,N_13132,N_17374);
or U22116 (N_22116,N_18322,N_18535);
or U22117 (N_22117,N_18345,N_13100);
nor U22118 (N_22118,N_17907,N_16003);
nor U22119 (N_22119,N_14918,N_12861);
or U22120 (N_22120,N_14411,N_13391);
xor U22121 (N_22121,N_12516,N_17192);
nand U22122 (N_22122,N_18068,N_15149);
nand U22123 (N_22123,N_14150,N_15169);
and U22124 (N_22124,N_14375,N_13444);
or U22125 (N_22125,N_14347,N_13631);
nor U22126 (N_22126,N_14390,N_13259);
and U22127 (N_22127,N_17001,N_12610);
nand U22128 (N_22128,N_16828,N_15428);
nand U22129 (N_22129,N_18207,N_13538);
nand U22130 (N_22130,N_15881,N_16575);
or U22131 (N_22131,N_14867,N_13555);
or U22132 (N_22132,N_18193,N_14990);
nor U22133 (N_22133,N_17002,N_13236);
nor U22134 (N_22134,N_17915,N_13551);
and U22135 (N_22135,N_15343,N_13355);
xnor U22136 (N_22136,N_13747,N_15252);
nor U22137 (N_22137,N_12627,N_15798);
nor U22138 (N_22138,N_15258,N_16550);
or U22139 (N_22139,N_14029,N_15488);
xor U22140 (N_22140,N_13295,N_13238);
nand U22141 (N_22141,N_13290,N_16604);
nand U22142 (N_22142,N_17887,N_15546);
and U22143 (N_22143,N_16604,N_13026);
or U22144 (N_22144,N_13119,N_15926);
nor U22145 (N_22145,N_18397,N_17183);
and U22146 (N_22146,N_12500,N_17202);
or U22147 (N_22147,N_15750,N_18596);
and U22148 (N_22148,N_17435,N_13598);
or U22149 (N_22149,N_16833,N_13210);
nor U22150 (N_22150,N_15906,N_15958);
nand U22151 (N_22151,N_18162,N_17753);
and U22152 (N_22152,N_18217,N_12644);
or U22153 (N_22153,N_16132,N_13076);
nand U22154 (N_22154,N_13503,N_16699);
and U22155 (N_22155,N_18392,N_15118);
or U22156 (N_22156,N_14388,N_13677);
and U22157 (N_22157,N_18646,N_12621);
nand U22158 (N_22158,N_13670,N_18166);
and U22159 (N_22159,N_17576,N_14582);
nand U22160 (N_22160,N_15533,N_17428);
or U22161 (N_22161,N_16969,N_15747);
nand U22162 (N_22162,N_13351,N_18042);
and U22163 (N_22163,N_16263,N_13307);
or U22164 (N_22164,N_13017,N_13901);
nand U22165 (N_22165,N_13304,N_16510);
and U22166 (N_22166,N_16904,N_16577);
nand U22167 (N_22167,N_12834,N_15213);
nor U22168 (N_22168,N_17833,N_14220);
nand U22169 (N_22169,N_16826,N_14637);
xor U22170 (N_22170,N_17548,N_16152);
or U22171 (N_22171,N_15010,N_15629);
and U22172 (N_22172,N_12601,N_13346);
and U22173 (N_22173,N_14641,N_14363);
and U22174 (N_22174,N_14089,N_18479);
or U22175 (N_22175,N_16721,N_16154);
or U22176 (N_22176,N_14147,N_15617);
or U22177 (N_22177,N_15779,N_14356);
or U22178 (N_22178,N_14021,N_18229);
and U22179 (N_22179,N_18091,N_14491);
or U22180 (N_22180,N_17577,N_14116);
nand U22181 (N_22181,N_16862,N_14861);
nand U22182 (N_22182,N_17801,N_13014);
nand U22183 (N_22183,N_17028,N_18047);
nor U22184 (N_22184,N_14633,N_15816);
nor U22185 (N_22185,N_16203,N_18287);
and U22186 (N_22186,N_17245,N_16646);
nor U22187 (N_22187,N_13106,N_12911);
nand U22188 (N_22188,N_17363,N_14553);
and U22189 (N_22189,N_14439,N_14761);
and U22190 (N_22190,N_13880,N_14560);
nand U22191 (N_22191,N_15481,N_18307);
xnor U22192 (N_22192,N_13458,N_12813);
and U22193 (N_22193,N_18495,N_13455);
and U22194 (N_22194,N_17862,N_14329);
and U22195 (N_22195,N_13439,N_14967);
nor U22196 (N_22196,N_12802,N_14964);
nand U22197 (N_22197,N_14816,N_14044);
and U22198 (N_22198,N_15543,N_16043);
nand U22199 (N_22199,N_14437,N_16906);
and U22200 (N_22200,N_17712,N_15007);
nor U22201 (N_22201,N_16730,N_18089);
xnor U22202 (N_22202,N_17201,N_13649);
and U22203 (N_22203,N_13504,N_16511);
and U22204 (N_22204,N_14550,N_15413);
nand U22205 (N_22205,N_14373,N_17181);
nor U22206 (N_22206,N_17782,N_13379);
nand U22207 (N_22207,N_15412,N_13032);
and U22208 (N_22208,N_14274,N_15915);
or U22209 (N_22209,N_16439,N_17187);
nor U22210 (N_22210,N_13158,N_13436);
or U22211 (N_22211,N_14708,N_14768);
nand U22212 (N_22212,N_12600,N_12757);
nor U22213 (N_22213,N_16580,N_14234);
nor U22214 (N_22214,N_13966,N_14107);
and U22215 (N_22215,N_15849,N_13744);
nor U22216 (N_22216,N_12744,N_17106);
nand U22217 (N_22217,N_14679,N_13922);
nor U22218 (N_22218,N_17920,N_12578);
xnor U22219 (N_22219,N_18220,N_12542);
nor U22220 (N_22220,N_14746,N_17735);
xnor U22221 (N_22221,N_12811,N_16395);
nor U22222 (N_22222,N_15863,N_13732);
and U22223 (N_22223,N_14526,N_16639);
nand U22224 (N_22224,N_14441,N_13770);
xnor U22225 (N_22225,N_15169,N_13645);
nand U22226 (N_22226,N_15326,N_17031);
and U22227 (N_22227,N_13699,N_14220);
and U22228 (N_22228,N_16928,N_16515);
xor U22229 (N_22229,N_14591,N_15230);
nor U22230 (N_22230,N_17115,N_17487);
nand U22231 (N_22231,N_16740,N_18686);
nand U22232 (N_22232,N_17813,N_15610);
nand U22233 (N_22233,N_15730,N_15725);
or U22234 (N_22234,N_14577,N_15035);
or U22235 (N_22235,N_14071,N_17059);
nand U22236 (N_22236,N_17331,N_16391);
nor U22237 (N_22237,N_17914,N_16161);
or U22238 (N_22238,N_15872,N_17356);
and U22239 (N_22239,N_17982,N_15942);
nand U22240 (N_22240,N_17105,N_15696);
or U22241 (N_22241,N_17126,N_16507);
nor U22242 (N_22242,N_16956,N_14793);
nand U22243 (N_22243,N_16630,N_15751);
nand U22244 (N_22244,N_15632,N_13110);
or U22245 (N_22245,N_14407,N_17332);
and U22246 (N_22246,N_17660,N_12914);
nand U22247 (N_22247,N_15239,N_18178);
or U22248 (N_22248,N_12766,N_13646);
or U22249 (N_22249,N_17765,N_15120);
xnor U22250 (N_22250,N_16450,N_14872);
xnor U22251 (N_22251,N_15060,N_14470);
nor U22252 (N_22252,N_13515,N_16188);
nand U22253 (N_22253,N_16477,N_15852);
and U22254 (N_22254,N_16250,N_15165);
nor U22255 (N_22255,N_12767,N_15677);
xor U22256 (N_22256,N_17493,N_15554);
or U22257 (N_22257,N_15050,N_15366);
nand U22258 (N_22258,N_17818,N_18154);
nand U22259 (N_22259,N_15622,N_12947);
nor U22260 (N_22260,N_13992,N_14740);
nand U22261 (N_22261,N_12905,N_14281);
and U22262 (N_22262,N_13814,N_13514);
and U22263 (N_22263,N_17460,N_13581);
xor U22264 (N_22264,N_14351,N_14138);
or U22265 (N_22265,N_18363,N_17256);
nand U22266 (N_22266,N_14787,N_15859);
nor U22267 (N_22267,N_16288,N_14719);
or U22268 (N_22268,N_16018,N_14158);
and U22269 (N_22269,N_17968,N_13817);
nor U22270 (N_22270,N_15038,N_13337);
and U22271 (N_22271,N_18472,N_15660);
and U22272 (N_22272,N_17359,N_18131);
or U22273 (N_22273,N_17299,N_12858);
nor U22274 (N_22274,N_16255,N_14263);
nor U22275 (N_22275,N_17872,N_15240);
nand U22276 (N_22276,N_15388,N_13872);
nor U22277 (N_22277,N_16767,N_17316);
and U22278 (N_22278,N_17371,N_18285);
nor U22279 (N_22279,N_12826,N_15407);
nor U22280 (N_22280,N_14778,N_16383);
nor U22281 (N_22281,N_17372,N_16530);
nor U22282 (N_22282,N_17175,N_17826);
and U22283 (N_22283,N_18679,N_16477);
nand U22284 (N_22284,N_15486,N_14287);
nand U22285 (N_22285,N_17954,N_15013);
or U22286 (N_22286,N_15742,N_17362);
nor U22287 (N_22287,N_18084,N_17481);
or U22288 (N_22288,N_15296,N_16351);
nor U22289 (N_22289,N_17104,N_18504);
or U22290 (N_22290,N_17580,N_17712);
nand U22291 (N_22291,N_17951,N_13318);
xnor U22292 (N_22292,N_16648,N_13362);
and U22293 (N_22293,N_15149,N_17489);
nor U22294 (N_22294,N_18369,N_13816);
nand U22295 (N_22295,N_14251,N_16190);
or U22296 (N_22296,N_16612,N_18705);
and U22297 (N_22297,N_13336,N_12892);
or U22298 (N_22298,N_17345,N_16596);
xor U22299 (N_22299,N_15657,N_13454);
nor U22300 (N_22300,N_17157,N_16253);
or U22301 (N_22301,N_13787,N_14977);
or U22302 (N_22302,N_17104,N_15763);
or U22303 (N_22303,N_13445,N_14475);
or U22304 (N_22304,N_17478,N_16547);
nor U22305 (N_22305,N_12995,N_12879);
and U22306 (N_22306,N_18149,N_14060);
and U22307 (N_22307,N_15878,N_12548);
nand U22308 (N_22308,N_12714,N_13072);
and U22309 (N_22309,N_18556,N_13430);
xor U22310 (N_22310,N_14174,N_15472);
or U22311 (N_22311,N_16583,N_15409);
nand U22312 (N_22312,N_15523,N_13839);
xor U22313 (N_22313,N_15814,N_14024);
and U22314 (N_22314,N_12931,N_15093);
nor U22315 (N_22315,N_14151,N_16696);
or U22316 (N_22316,N_18516,N_16492);
nor U22317 (N_22317,N_13317,N_12962);
and U22318 (N_22318,N_15459,N_13928);
nand U22319 (N_22319,N_16851,N_16404);
nand U22320 (N_22320,N_12562,N_16649);
nor U22321 (N_22321,N_18514,N_12929);
nor U22322 (N_22322,N_17554,N_15774);
nor U22323 (N_22323,N_13518,N_12964);
or U22324 (N_22324,N_16761,N_13780);
xnor U22325 (N_22325,N_14902,N_13721);
and U22326 (N_22326,N_17232,N_17480);
or U22327 (N_22327,N_14703,N_17717);
nor U22328 (N_22328,N_18346,N_15086);
and U22329 (N_22329,N_13590,N_12706);
nand U22330 (N_22330,N_14127,N_13627);
nor U22331 (N_22331,N_13541,N_16982);
nor U22332 (N_22332,N_13634,N_17418);
nor U22333 (N_22333,N_14099,N_15449);
nor U22334 (N_22334,N_15497,N_16368);
xnor U22335 (N_22335,N_15418,N_12885);
and U22336 (N_22336,N_14818,N_18673);
nor U22337 (N_22337,N_17010,N_14896);
nand U22338 (N_22338,N_15999,N_15373);
nor U22339 (N_22339,N_16646,N_15793);
and U22340 (N_22340,N_13493,N_15646);
nand U22341 (N_22341,N_14355,N_13070);
nand U22342 (N_22342,N_16102,N_15853);
and U22343 (N_22343,N_13338,N_16447);
or U22344 (N_22344,N_15819,N_13561);
or U22345 (N_22345,N_13518,N_13012);
and U22346 (N_22346,N_16117,N_16665);
nor U22347 (N_22347,N_15808,N_18649);
xnor U22348 (N_22348,N_16849,N_17100);
or U22349 (N_22349,N_16581,N_13659);
nand U22350 (N_22350,N_13202,N_15542);
nand U22351 (N_22351,N_17083,N_15865);
nor U22352 (N_22352,N_17308,N_18278);
nor U22353 (N_22353,N_16674,N_18475);
nor U22354 (N_22354,N_17285,N_13339);
xnor U22355 (N_22355,N_15146,N_12574);
and U22356 (N_22356,N_13297,N_16192);
nor U22357 (N_22357,N_17709,N_13801);
and U22358 (N_22358,N_14517,N_13156);
nand U22359 (N_22359,N_15725,N_12963);
nor U22360 (N_22360,N_13397,N_17724);
nand U22361 (N_22361,N_17239,N_14241);
nor U22362 (N_22362,N_14906,N_13701);
or U22363 (N_22363,N_15827,N_15628);
and U22364 (N_22364,N_15054,N_14010);
or U22365 (N_22365,N_14838,N_17715);
nand U22366 (N_22366,N_16536,N_13426);
and U22367 (N_22367,N_16745,N_15874);
nor U22368 (N_22368,N_12759,N_16942);
and U22369 (N_22369,N_18479,N_15786);
xnor U22370 (N_22370,N_15509,N_15922);
nand U22371 (N_22371,N_17346,N_17140);
xor U22372 (N_22372,N_14936,N_18602);
nor U22373 (N_22373,N_18045,N_18675);
or U22374 (N_22374,N_12589,N_13752);
or U22375 (N_22375,N_13124,N_15268);
and U22376 (N_22376,N_15559,N_13631);
nor U22377 (N_22377,N_16784,N_13289);
nor U22378 (N_22378,N_18588,N_17564);
and U22379 (N_22379,N_16342,N_15132);
nand U22380 (N_22380,N_13287,N_14636);
or U22381 (N_22381,N_17704,N_13108);
nand U22382 (N_22382,N_13131,N_14388);
xor U22383 (N_22383,N_13284,N_18240);
nand U22384 (N_22384,N_13585,N_17655);
or U22385 (N_22385,N_18376,N_15889);
nand U22386 (N_22386,N_18647,N_18308);
and U22387 (N_22387,N_17739,N_13865);
and U22388 (N_22388,N_13299,N_13119);
xor U22389 (N_22389,N_14711,N_17330);
and U22390 (N_22390,N_14554,N_14257);
nand U22391 (N_22391,N_16892,N_14782);
nand U22392 (N_22392,N_16325,N_14180);
and U22393 (N_22393,N_14300,N_14810);
xor U22394 (N_22394,N_18592,N_13964);
nand U22395 (N_22395,N_17462,N_16665);
xnor U22396 (N_22396,N_16671,N_18418);
nand U22397 (N_22397,N_14140,N_16420);
and U22398 (N_22398,N_12955,N_16936);
nand U22399 (N_22399,N_18492,N_14293);
and U22400 (N_22400,N_17396,N_17205);
nand U22401 (N_22401,N_14384,N_15265);
nor U22402 (N_22402,N_14462,N_15558);
and U22403 (N_22403,N_12564,N_13592);
nand U22404 (N_22404,N_18414,N_13712);
nand U22405 (N_22405,N_18697,N_18297);
nor U22406 (N_22406,N_13307,N_14363);
and U22407 (N_22407,N_16602,N_13499);
or U22408 (N_22408,N_15687,N_12855);
or U22409 (N_22409,N_17600,N_13584);
nand U22410 (N_22410,N_15231,N_18376);
or U22411 (N_22411,N_15281,N_16899);
xnor U22412 (N_22412,N_17793,N_14375);
or U22413 (N_22413,N_13266,N_17700);
xnor U22414 (N_22414,N_13136,N_14390);
nor U22415 (N_22415,N_16225,N_17933);
nand U22416 (N_22416,N_13675,N_14673);
xnor U22417 (N_22417,N_18471,N_14224);
or U22418 (N_22418,N_18716,N_13660);
or U22419 (N_22419,N_17222,N_18108);
nand U22420 (N_22420,N_13604,N_14803);
xor U22421 (N_22421,N_13840,N_16559);
xor U22422 (N_22422,N_12715,N_14066);
or U22423 (N_22423,N_13746,N_16436);
nor U22424 (N_22424,N_18456,N_17632);
nor U22425 (N_22425,N_16020,N_13973);
nor U22426 (N_22426,N_13138,N_13852);
or U22427 (N_22427,N_16543,N_18535);
or U22428 (N_22428,N_16395,N_16439);
or U22429 (N_22429,N_17086,N_15635);
nand U22430 (N_22430,N_14806,N_14721);
nand U22431 (N_22431,N_17611,N_17140);
nand U22432 (N_22432,N_14900,N_12953);
or U22433 (N_22433,N_14685,N_18288);
nand U22434 (N_22434,N_16439,N_12585);
and U22435 (N_22435,N_18378,N_13067);
xor U22436 (N_22436,N_14663,N_15877);
nor U22437 (N_22437,N_18089,N_17384);
and U22438 (N_22438,N_18048,N_14964);
nand U22439 (N_22439,N_18552,N_17655);
and U22440 (N_22440,N_17679,N_13376);
and U22441 (N_22441,N_15166,N_14013);
nand U22442 (N_22442,N_14558,N_15705);
or U22443 (N_22443,N_15675,N_17601);
nor U22444 (N_22444,N_12915,N_17125);
xnor U22445 (N_22445,N_14538,N_13528);
xor U22446 (N_22446,N_13266,N_18388);
xor U22447 (N_22447,N_17876,N_18676);
and U22448 (N_22448,N_15245,N_14624);
nand U22449 (N_22449,N_13751,N_17093);
xnor U22450 (N_22450,N_15343,N_14381);
or U22451 (N_22451,N_12790,N_18105);
nand U22452 (N_22452,N_16033,N_15848);
and U22453 (N_22453,N_17226,N_16182);
xor U22454 (N_22454,N_13698,N_13818);
or U22455 (N_22455,N_15457,N_15517);
and U22456 (N_22456,N_13355,N_14148);
or U22457 (N_22457,N_17656,N_16639);
or U22458 (N_22458,N_12641,N_12727);
xor U22459 (N_22459,N_16115,N_15718);
and U22460 (N_22460,N_16779,N_15737);
and U22461 (N_22461,N_15343,N_17931);
or U22462 (N_22462,N_13423,N_14544);
nand U22463 (N_22463,N_14102,N_13924);
and U22464 (N_22464,N_13222,N_15458);
or U22465 (N_22465,N_14947,N_16583);
nor U22466 (N_22466,N_16162,N_14867);
or U22467 (N_22467,N_13838,N_15081);
nand U22468 (N_22468,N_16127,N_16399);
nor U22469 (N_22469,N_18593,N_16488);
or U22470 (N_22470,N_14252,N_18732);
nor U22471 (N_22471,N_18737,N_13264);
or U22472 (N_22472,N_18619,N_17880);
and U22473 (N_22473,N_15136,N_17404);
xnor U22474 (N_22474,N_18525,N_13852);
and U22475 (N_22475,N_16981,N_18635);
and U22476 (N_22476,N_17531,N_12534);
or U22477 (N_22477,N_18313,N_12944);
or U22478 (N_22478,N_14219,N_17799);
nand U22479 (N_22479,N_12957,N_14507);
and U22480 (N_22480,N_13565,N_16479);
nor U22481 (N_22481,N_14200,N_14570);
nand U22482 (N_22482,N_15518,N_12694);
xnor U22483 (N_22483,N_18609,N_15546);
nor U22484 (N_22484,N_17958,N_14489);
and U22485 (N_22485,N_16710,N_17455);
nand U22486 (N_22486,N_15700,N_13723);
xor U22487 (N_22487,N_13342,N_16012);
or U22488 (N_22488,N_15515,N_15768);
nor U22489 (N_22489,N_18369,N_16530);
and U22490 (N_22490,N_14014,N_18046);
nand U22491 (N_22491,N_13623,N_15899);
or U22492 (N_22492,N_17031,N_14938);
nor U22493 (N_22493,N_12586,N_13680);
nand U22494 (N_22494,N_17733,N_13808);
or U22495 (N_22495,N_15964,N_17055);
nor U22496 (N_22496,N_14515,N_14890);
nand U22497 (N_22497,N_18315,N_15459);
and U22498 (N_22498,N_15442,N_18245);
nand U22499 (N_22499,N_17507,N_17233);
nand U22500 (N_22500,N_12805,N_18398);
nand U22501 (N_22501,N_13894,N_16863);
nor U22502 (N_22502,N_14042,N_17573);
or U22503 (N_22503,N_13967,N_18364);
nand U22504 (N_22504,N_13728,N_13883);
and U22505 (N_22505,N_12990,N_18413);
nor U22506 (N_22506,N_18738,N_12672);
and U22507 (N_22507,N_17270,N_13489);
and U22508 (N_22508,N_18511,N_17409);
nor U22509 (N_22509,N_14113,N_16827);
or U22510 (N_22510,N_18537,N_18095);
nand U22511 (N_22511,N_18042,N_14893);
or U22512 (N_22512,N_16534,N_16141);
or U22513 (N_22513,N_17014,N_17170);
nand U22514 (N_22514,N_18371,N_15217);
or U22515 (N_22515,N_16269,N_14246);
nor U22516 (N_22516,N_17925,N_15542);
xor U22517 (N_22517,N_13440,N_15463);
and U22518 (N_22518,N_16881,N_15847);
or U22519 (N_22519,N_18175,N_17820);
nand U22520 (N_22520,N_12912,N_13291);
nand U22521 (N_22521,N_15002,N_13196);
nor U22522 (N_22522,N_16141,N_17997);
and U22523 (N_22523,N_13322,N_12829);
or U22524 (N_22524,N_13901,N_12650);
nand U22525 (N_22525,N_15544,N_13337);
xor U22526 (N_22526,N_17905,N_15679);
nor U22527 (N_22527,N_15386,N_18042);
xor U22528 (N_22528,N_12811,N_17212);
or U22529 (N_22529,N_15447,N_13964);
nand U22530 (N_22530,N_15820,N_14209);
and U22531 (N_22531,N_17547,N_16553);
or U22532 (N_22532,N_13178,N_16196);
nor U22533 (N_22533,N_15813,N_16632);
or U22534 (N_22534,N_12532,N_13527);
xor U22535 (N_22535,N_12569,N_15415);
nor U22536 (N_22536,N_15658,N_12888);
nand U22537 (N_22537,N_16233,N_15741);
or U22538 (N_22538,N_17645,N_18107);
nand U22539 (N_22539,N_16822,N_16249);
or U22540 (N_22540,N_14297,N_18088);
or U22541 (N_22541,N_15394,N_13229);
or U22542 (N_22542,N_15667,N_16400);
xnor U22543 (N_22543,N_14571,N_12509);
and U22544 (N_22544,N_16392,N_18051);
xnor U22545 (N_22545,N_18629,N_16161);
xor U22546 (N_22546,N_12604,N_13516);
nor U22547 (N_22547,N_14974,N_17105);
nand U22548 (N_22548,N_17375,N_13188);
nand U22549 (N_22549,N_14038,N_16219);
nand U22550 (N_22550,N_14669,N_16498);
nor U22551 (N_22551,N_14518,N_18548);
nor U22552 (N_22552,N_18049,N_16394);
and U22553 (N_22553,N_13735,N_12882);
or U22554 (N_22554,N_17799,N_17303);
nor U22555 (N_22555,N_17037,N_16181);
nor U22556 (N_22556,N_17546,N_16665);
xnor U22557 (N_22557,N_17619,N_17171);
nand U22558 (N_22558,N_17603,N_15129);
nand U22559 (N_22559,N_15011,N_15607);
or U22560 (N_22560,N_17165,N_16332);
nand U22561 (N_22561,N_17549,N_13021);
xnor U22562 (N_22562,N_18093,N_18356);
nor U22563 (N_22563,N_12944,N_17846);
xnor U22564 (N_22564,N_15551,N_13058);
and U22565 (N_22565,N_16091,N_14056);
or U22566 (N_22566,N_17476,N_18255);
and U22567 (N_22567,N_14135,N_16788);
xnor U22568 (N_22568,N_13089,N_12664);
and U22569 (N_22569,N_17838,N_15731);
or U22570 (N_22570,N_17202,N_12592);
xnor U22571 (N_22571,N_15864,N_18087);
or U22572 (N_22572,N_16845,N_16244);
nand U22573 (N_22573,N_17417,N_17325);
nor U22574 (N_22574,N_14836,N_13966);
nand U22575 (N_22575,N_18040,N_15207);
nor U22576 (N_22576,N_15020,N_15921);
or U22577 (N_22577,N_14963,N_16616);
or U22578 (N_22578,N_17213,N_17849);
or U22579 (N_22579,N_15789,N_15262);
nand U22580 (N_22580,N_14801,N_14047);
and U22581 (N_22581,N_14501,N_12622);
or U22582 (N_22582,N_18523,N_18246);
nand U22583 (N_22583,N_16230,N_13447);
and U22584 (N_22584,N_16834,N_17755);
and U22585 (N_22585,N_16628,N_14483);
or U22586 (N_22586,N_13301,N_14670);
or U22587 (N_22587,N_16498,N_16945);
and U22588 (N_22588,N_14804,N_18553);
or U22589 (N_22589,N_12664,N_13468);
nand U22590 (N_22590,N_13264,N_14910);
nor U22591 (N_22591,N_15693,N_18745);
nand U22592 (N_22592,N_15343,N_12566);
or U22593 (N_22593,N_14081,N_18146);
nor U22594 (N_22594,N_13148,N_12808);
or U22595 (N_22595,N_16570,N_14069);
or U22596 (N_22596,N_18704,N_16112);
nor U22597 (N_22597,N_16634,N_16532);
and U22598 (N_22598,N_18413,N_14017);
nand U22599 (N_22599,N_16096,N_14818);
or U22600 (N_22600,N_15183,N_13027);
nand U22601 (N_22601,N_13445,N_17448);
nor U22602 (N_22602,N_17978,N_12564);
xnor U22603 (N_22603,N_17765,N_13484);
nor U22604 (N_22604,N_12629,N_17910);
nor U22605 (N_22605,N_12895,N_15786);
xor U22606 (N_22606,N_13086,N_18703);
and U22607 (N_22607,N_13657,N_13016);
and U22608 (N_22608,N_14036,N_17239);
xnor U22609 (N_22609,N_17282,N_18372);
and U22610 (N_22610,N_13356,N_18452);
and U22611 (N_22611,N_18548,N_16786);
nor U22612 (N_22612,N_17049,N_12702);
nand U22613 (N_22613,N_12844,N_14395);
nand U22614 (N_22614,N_18557,N_12836);
xor U22615 (N_22615,N_14962,N_15202);
and U22616 (N_22616,N_14613,N_12722);
nor U22617 (N_22617,N_18601,N_17663);
nand U22618 (N_22618,N_12524,N_16694);
nand U22619 (N_22619,N_13209,N_17632);
nand U22620 (N_22620,N_15130,N_17234);
and U22621 (N_22621,N_13007,N_15451);
nand U22622 (N_22622,N_18032,N_13985);
nor U22623 (N_22623,N_17006,N_14868);
and U22624 (N_22624,N_14482,N_13170);
and U22625 (N_22625,N_14604,N_14329);
nor U22626 (N_22626,N_18747,N_12554);
or U22627 (N_22627,N_16910,N_13041);
or U22628 (N_22628,N_14973,N_14693);
or U22629 (N_22629,N_18347,N_18656);
and U22630 (N_22630,N_17173,N_17772);
nand U22631 (N_22631,N_16237,N_16235);
nor U22632 (N_22632,N_12886,N_15331);
nor U22633 (N_22633,N_14380,N_15868);
or U22634 (N_22634,N_12677,N_18141);
or U22635 (N_22635,N_17085,N_17081);
and U22636 (N_22636,N_17659,N_15944);
or U22637 (N_22637,N_13847,N_17382);
or U22638 (N_22638,N_15584,N_17279);
or U22639 (N_22639,N_16372,N_16352);
or U22640 (N_22640,N_17753,N_14856);
nor U22641 (N_22641,N_17875,N_14826);
or U22642 (N_22642,N_16642,N_13072);
and U22643 (N_22643,N_15773,N_12540);
nor U22644 (N_22644,N_18629,N_14373);
and U22645 (N_22645,N_18283,N_16274);
nor U22646 (N_22646,N_15003,N_18048);
and U22647 (N_22647,N_13699,N_12959);
and U22648 (N_22648,N_16773,N_15072);
nand U22649 (N_22649,N_16106,N_17982);
and U22650 (N_22650,N_13579,N_16913);
nor U22651 (N_22651,N_15533,N_13075);
nand U22652 (N_22652,N_16122,N_12734);
nand U22653 (N_22653,N_17552,N_16773);
nand U22654 (N_22654,N_17934,N_13186);
nand U22655 (N_22655,N_13962,N_18126);
nand U22656 (N_22656,N_18679,N_18693);
nor U22657 (N_22657,N_15053,N_15725);
and U22658 (N_22658,N_15092,N_14821);
or U22659 (N_22659,N_17784,N_12815);
or U22660 (N_22660,N_13103,N_15314);
nor U22661 (N_22661,N_13746,N_15642);
or U22662 (N_22662,N_14519,N_18046);
xor U22663 (N_22663,N_17978,N_17476);
xor U22664 (N_22664,N_13981,N_13523);
and U22665 (N_22665,N_13016,N_14083);
and U22666 (N_22666,N_15707,N_18028);
nand U22667 (N_22667,N_12699,N_17367);
or U22668 (N_22668,N_14270,N_14056);
and U22669 (N_22669,N_18637,N_17651);
and U22670 (N_22670,N_14907,N_18437);
xor U22671 (N_22671,N_16098,N_13845);
or U22672 (N_22672,N_13167,N_14919);
or U22673 (N_22673,N_13932,N_18425);
nor U22674 (N_22674,N_17459,N_15210);
and U22675 (N_22675,N_17252,N_17405);
and U22676 (N_22676,N_15807,N_13473);
nand U22677 (N_22677,N_17009,N_16770);
xnor U22678 (N_22678,N_13209,N_15465);
and U22679 (N_22679,N_15466,N_18005);
and U22680 (N_22680,N_18363,N_12525);
and U22681 (N_22681,N_16146,N_15569);
nor U22682 (N_22682,N_14003,N_13159);
and U22683 (N_22683,N_15912,N_15603);
nand U22684 (N_22684,N_18558,N_14428);
or U22685 (N_22685,N_16215,N_13975);
or U22686 (N_22686,N_18513,N_13563);
nor U22687 (N_22687,N_18356,N_17642);
nor U22688 (N_22688,N_17712,N_17024);
or U22689 (N_22689,N_14708,N_13368);
and U22690 (N_22690,N_14645,N_14453);
nand U22691 (N_22691,N_16801,N_14917);
nand U22692 (N_22692,N_13471,N_18620);
or U22693 (N_22693,N_17379,N_18520);
or U22694 (N_22694,N_16093,N_13019);
or U22695 (N_22695,N_14814,N_13315);
nor U22696 (N_22696,N_14517,N_17421);
nand U22697 (N_22697,N_17839,N_13319);
nand U22698 (N_22698,N_15382,N_14003);
nor U22699 (N_22699,N_14382,N_17399);
nor U22700 (N_22700,N_16145,N_16879);
and U22701 (N_22701,N_15177,N_16013);
and U22702 (N_22702,N_17195,N_15309);
or U22703 (N_22703,N_14081,N_16148);
and U22704 (N_22704,N_16505,N_18056);
and U22705 (N_22705,N_17022,N_13616);
nor U22706 (N_22706,N_14914,N_18670);
nand U22707 (N_22707,N_16035,N_15404);
and U22708 (N_22708,N_16990,N_16829);
or U22709 (N_22709,N_16545,N_12560);
or U22710 (N_22710,N_15873,N_15661);
and U22711 (N_22711,N_14847,N_15649);
or U22712 (N_22712,N_17402,N_18247);
xor U22713 (N_22713,N_17776,N_12542);
nor U22714 (N_22714,N_13546,N_15712);
and U22715 (N_22715,N_14063,N_16863);
nand U22716 (N_22716,N_15733,N_13920);
or U22717 (N_22717,N_14892,N_16945);
and U22718 (N_22718,N_12831,N_14686);
nand U22719 (N_22719,N_13110,N_18072);
nand U22720 (N_22720,N_13293,N_17883);
and U22721 (N_22721,N_13095,N_12594);
nor U22722 (N_22722,N_15536,N_16826);
xor U22723 (N_22723,N_16638,N_12588);
nand U22724 (N_22724,N_17964,N_17399);
nand U22725 (N_22725,N_16140,N_18140);
nor U22726 (N_22726,N_18093,N_14559);
xnor U22727 (N_22727,N_16547,N_16606);
nor U22728 (N_22728,N_13759,N_15911);
or U22729 (N_22729,N_17404,N_17263);
and U22730 (N_22730,N_13332,N_15113);
nand U22731 (N_22731,N_16666,N_16300);
nor U22732 (N_22732,N_17271,N_16307);
and U22733 (N_22733,N_15044,N_18599);
nor U22734 (N_22734,N_15275,N_18333);
and U22735 (N_22735,N_16144,N_16790);
and U22736 (N_22736,N_17162,N_15465);
nor U22737 (N_22737,N_18113,N_13531);
xor U22738 (N_22738,N_15667,N_14308);
nor U22739 (N_22739,N_18429,N_16003);
nor U22740 (N_22740,N_13640,N_13823);
and U22741 (N_22741,N_16479,N_16418);
nor U22742 (N_22742,N_17812,N_17533);
or U22743 (N_22743,N_16901,N_13473);
and U22744 (N_22744,N_17151,N_13268);
and U22745 (N_22745,N_14815,N_18555);
nor U22746 (N_22746,N_13066,N_18460);
or U22747 (N_22747,N_16950,N_17668);
nor U22748 (N_22748,N_13996,N_17897);
nand U22749 (N_22749,N_15807,N_15738);
nor U22750 (N_22750,N_12625,N_12566);
or U22751 (N_22751,N_12742,N_17800);
and U22752 (N_22752,N_15749,N_15563);
nand U22753 (N_22753,N_14780,N_13884);
nand U22754 (N_22754,N_13527,N_14877);
or U22755 (N_22755,N_17557,N_15095);
xor U22756 (N_22756,N_16384,N_14759);
or U22757 (N_22757,N_16364,N_13551);
nor U22758 (N_22758,N_16051,N_13405);
nand U22759 (N_22759,N_16930,N_15960);
and U22760 (N_22760,N_15339,N_13315);
nand U22761 (N_22761,N_13284,N_14124);
nor U22762 (N_22762,N_16396,N_18040);
and U22763 (N_22763,N_17231,N_15856);
nor U22764 (N_22764,N_14499,N_16310);
nor U22765 (N_22765,N_18189,N_12578);
nand U22766 (N_22766,N_13099,N_14704);
nand U22767 (N_22767,N_17984,N_18322);
nand U22768 (N_22768,N_14091,N_17926);
and U22769 (N_22769,N_17642,N_14052);
nor U22770 (N_22770,N_16938,N_17273);
nor U22771 (N_22771,N_14119,N_17916);
xor U22772 (N_22772,N_15037,N_16181);
or U22773 (N_22773,N_17789,N_15992);
or U22774 (N_22774,N_13667,N_16267);
nand U22775 (N_22775,N_15603,N_17629);
nor U22776 (N_22776,N_16555,N_15310);
and U22777 (N_22777,N_17425,N_17357);
nand U22778 (N_22778,N_16225,N_18046);
xor U22779 (N_22779,N_17061,N_18205);
nand U22780 (N_22780,N_17965,N_15314);
or U22781 (N_22781,N_17538,N_17401);
nor U22782 (N_22782,N_18132,N_17070);
nor U22783 (N_22783,N_18328,N_15060);
nand U22784 (N_22784,N_15295,N_18589);
and U22785 (N_22785,N_14832,N_15783);
and U22786 (N_22786,N_17119,N_15414);
nand U22787 (N_22787,N_12816,N_15703);
nor U22788 (N_22788,N_18246,N_13344);
xnor U22789 (N_22789,N_15579,N_16142);
nor U22790 (N_22790,N_16379,N_12558);
nand U22791 (N_22791,N_14432,N_17488);
xor U22792 (N_22792,N_14949,N_13909);
nor U22793 (N_22793,N_15705,N_14103);
nor U22794 (N_22794,N_16981,N_17762);
or U22795 (N_22795,N_13439,N_13270);
and U22796 (N_22796,N_18074,N_16287);
nor U22797 (N_22797,N_13813,N_18147);
nand U22798 (N_22798,N_18741,N_16872);
and U22799 (N_22799,N_18187,N_15988);
nand U22800 (N_22800,N_14267,N_14844);
nor U22801 (N_22801,N_15019,N_13686);
xor U22802 (N_22802,N_13977,N_15666);
nor U22803 (N_22803,N_14437,N_18476);
nor U22804 (N_22804,N_13214,N_13507);
nand U22805 (N_22805,N_12621,N_15421);
nor U22806 (N_22806,N_12884,N_16413);
nor U22807 (N_22807,N_17158,N_14107);
nor U22808 (N_22808,N_15654,N_14004);
and U22809 (N_22809,N_16112,N_18615);
and U22810 (N_22810,N_15261,N_16977);
nor U22811 (N_22811,N_17862,N_18558);
xor U22812 (N_22812,N_12587,N_13236);
xnor U22813 (N_22813,N_17309,N_18549);
xnor U22814 (N_22814,N_13512,N_13570);
nand U22815 (N_22815,N_16168,N_12942);
nand U22816 (N_22816,N_17791,N_15680);
xnor U22817 (N_22817,N_17615,N_13140);
or U22818 (N_22818,N_18662,N_17107);
nor U22819 (N_22819,N_15558,N_16629);
nand U22820 (N_22820,N_17334,N_17580);
nor U22821 (N_22821,N_13905,N_16620);
or U22822 (N_22822,N_17639,N_16938);
or U22823 (N_22823,N_18506,N_13141);
and U22824 (N_22824,N_15633,N_13389);
nor U22825 (N_22825,N_18327,N_14259);
or U22826 (N_22826,N_17048,N_14208);
and U22827 (N_22827,N_14558,N_12620);
or U22828 (N_22828,N_16756,N_13472);
nand U22829 (N_22829,N_15244,N_12838);
nor U22830 (N_22830,N_16703,N_13209);
xor U22831 (N_22831,N_18644,N_18575);
and U22832 (N_22832,N_18072,N_12895);
nand U22833 (N_22833,N_13251,N_16381);
nor U22834 (N_22834,N_15090,N_14339);
nor U22835 (N_22835,N_14946,N_17352);
or U22836 (N_22836,N_16433,N_16789);
nand U22837 (N_22837,N_16435,N_14475);
nor U22838 (N_22838,N_14376,N_13030);
or U22839 (N_22839,N_16841,N_16018);
and U22840 (N_22840,N_14065,N_16915);
or U22841 (N_22841,N_15158,N_16561);
nor U22842 (N_22842,N_17716,N_16921);
and U22843 (N_22843,N_17079,N_18120);
xnor U22844 (N_22844,N_18062,N_13230);
and U22845 (N_22845,N_12539,N_14035);
nand U22846 (N_22846,N_17729,N_14708);
or U22847 (N_22847,N_15512,N_15231);
nand U22848 (N_22848,N_13117,N_12761);
xor U22849 (N_22849,N_15781,N_16058);
and U22850 (N_22850,N_14595,N_17917);
nor U22851 (N_22851,N_16237,N_18013);
or U22852 (N_22852,N_16408,N_14169);
nand U22853 (N_22853,N_16017,N_16966);
and U22854 (N_22854,N_18637,N_16480);
or U22855 (N_22855,N_15052,N_17257);
and U22856 (N_22856,N_16273,N_13325);
nor U22857 (N_22857,N_15446,N_18555);
or U22858 (N_22858,N_17619,N_18523);
or U22859 (N_22859,N_13979,N_16084);
or U22860 (N_22860,N_13253,N_15428);
nor U22861 (N_22861,N_17521,N_14356);
or U22862 (N_22862,N_17023,N_15397);
or U22863 (N_22863,N_13892,N_18266);
xnor U22864 (N_22864,N_18735,N_12631);
or U22865 (N_22865,N_18587,N_14867);
and U22866 (N_22866,N_16386,N_16744);
and U22867 (N_22867,N_14339,N_15033);
and U22868 (N_22868,N_15718,N_15407);
nand U22869 (N_22869,N_17159,N_16169);
and U22870 (N_22870,N_14166,N_13198);
nor U22871 (N_22871,N_18277,N_16228);
and U22872 (N_22872,N_18179,N_14276);
nor U22873 (N_22873,N_18558,N_14117);
nor U22874 (N_22874,N_18601,N_12668);
nand U22875 (N_22875,N_14063,N_17717);
nor U22876 (N_22876,N_15264,N_15036);
nand U22877 (N_22877,N_13633,N_14240);
nor U22878 (N_22878,N_13278,N_15478);
nor U22879 (N_22879,N_16406,N_14208);
and U22880 (N_22880,N_12523,N_12686);
and U22881 (N_22881,N_17495,N_16466);
nand U22882 (N_22882,N_14059,N_13500);
and U22883 (N_22883,N_15716,N_17789);
xor U22884 (N_22884,N_13531,N_15321);
nor U22885 (N_22885,N_12698,N_15515);
or U22886 (N_22886,N_17665,N_14456);
or U22887 (N_22887,N_13237,N_17435);
or U22888 (N_22888,N_18067,N_17959);
nand U22889 (N_22889,N_15838,N_16745);
nand U22890 (N_22890,N_14267,N_12652);
or U22891 (N_22891,N_12506,N_12919);
nor U22892 (N_22892,N_17824,N_13309);
nor U22893 (N_22893,N_17953,N_16087);
and U22894 (N_22894,N_14529,N_16393);
nor U22895 (N_22895,N_16670,N_13482);
or U22896 (N_22896,N_16653,N_15032);
nor U22897 (N_22897,N_17158,N_16216);
nor U22898 (N_22898,N_17847,N_17347);
and U22899 (N_22899,N_14228,N_12659);
nand U22900 (N_22900,N_15043,N_12703);
and U22901 (N_22901,N_15771,N_15792);
nand U22902 (N_22902,N_14114,N_13831);
nor U22903 (N_22903,N_17055,N_16815);
or U22904 (N_22904,N_13115,N_17032);
or U22905 (N_22905,N_14833,N_15410);
or U22906 (N_22906,N_16311,N_14301);
and U22907 (N_22907,N_14131,N_14153);
and U22908 (N_22908,N_16105,N_14927);
and U22909 (N_22909,N_16023,N_17596);
or U22910 (N_22910,N_12793,N_15438);
nand U22911 (N_22911,N_16439,N_15669);
nor U22912 (N_22912,N_17521,N_17750);
and U22913 (N_22913,N_12615,N_16083);
or U22914 (N_22914,N_14065,N_15409);
and U22915 (N_22915,N_17827,N_13873);
or U22916 (N_22916,N_16423,N_18743);
nand U22917 (N_22917,N_15514,N_15810);
nor U22918 (N_22918,N_14046,N_15191);
and U22919 (N_22919,N_17258,N_13459);
or U22920 (N_22920,N_13265,N_12918);
nor U22921 (N_22921,N_16541,N_14154);
or U22922 (N_22922,N_17124,N_14890);
nand U22923 (N_22923,N_17572,N_14778);
nand U22924 (N_22924,N_14157,N_14894);
and U22925 (N_22925,N_13894,N_18596);
nor U22926 (N_22926,N_13423,N_16002);
or U22927 (N_22927,N_17703,N_13653);
nand U22928 (N_22928,N_16541,N_18744);
nor U22929 (N_22929,N_16886,N_18278);
xnor U22930 (N_22930,N_15470,N_14686);
nor U22931 (N_22931,N_13213,N_15818);
nor U22932 (N_22932,N_14742,N_17219);
or U22933 (N_22933,N_15600,N_18362);
nor U22934 (N_22934,N_17480,N_13541);
nor U22935 (N_22935,N_17956,N_15859);
and U22936 (N_22936,N_13067,N_18333);
nand U22937 (N_22937,N_13417,N_14969);
or U22938 (N_22938,N_16503,N_12535);
and U22939 (N_22939,N_18221,N_15247);
nand U22940 (N_22940,N_13187,N_15089);
and U22941 (N_22941,N_16592,N_12723);
nor U22942 (N_22942,N_18665,N_18402);
nor U22943 (N_22943,N_17301,N_14582);
and U22944 (N_22944,N_15829,N_17075);
or U22945 (N_22945,N_12596,N_14892);
nor U22946 (N_22946,N_15030,N_16649);
nor U22947 (N_22947,N_13565,N_13388);
or U22948 (N_22948,N_14782,N_14172);
and U22949 (N_22949,N_16535,N_15130);
or U22950 (N_22950,N_15628,N_14234);
nor U22951 (N_22951,N_15750,N_12790);
nand U22952 (N_22952,N_18169,N_18643);
nor U22953 (N_22953,N_16536,N_16801);
xor U22954 (N_22954,N_13583,N_15797);
xnor U22955 (N_22955,N_14531,N_14682);
or U22956 (N_22956,N_13072,N_15780);
nor U22957 (N_22957,N_16677,N_18697);
nand U22958 (N_22958,N_12936,N_16769);
and U22959 (N_22959,N_13084,N_15822);
and U22960 (N_22960,N_15734,N_17050);
nand U22961 (N_22961,N_15689,N_17319);
nor U22962 (N_22962,N_14032,N_15192);
or U22963 (N_22963,N_14269,N_16841);
or U22964 (N_22964,N_14857,N_16886);
or U22965 (N_22965,N_17394,N_15715);
xor U22966 (N_22966,N_16638,N_14066);
and U22967 (N_22967,N_16717,N_17188);
nor U22968 (N_22968,N_14937,N_13630);
or U22969 (N_22969,N_12743,N_18140);
nor U22970 (N_22970,N_12667,N_17365);
and U22971 (N_22971,N_15743,N_15448);
and U22972 (N_22972,N_14806,N_17626);
nor U22973 (N_22973,N_13729,N_13428);
and U22974 (N_22974,N_14243,N_17408);
xnor U22975 (N_22975,N_18274,N_18346);
nor U22976 (N_22976,N_16114,N_13051);
nand U22977 (N_22977,N_17784,N_13541);
xnor U22978 (N_22978,N_17096,N_12964);
or U22979 (N_22979,N_13656,N_15421);
or U22980 (N_22980,N_17610,N_14279);
nand U22981 (N_22981,N_15832,N_15096);
and U22982 (N_22982,N_18572,N_15431);
nor U22983 (N_22983,N_16287,N_12712);
nand U22984 (N_22984,N_15491,N_15874);
nand U22985 (N_22985,N_16218,N_16845);
or U22986 (N_22986,N_16540,N_17363);
nand U22987 (N_22987,N_12875,N_17205);
nand U22988 (N_22988,N_13934,N_12729);
or U22989 (N_22989,N_14846,N_12815);
nand U22990 (N_22990,N_16100,N_17722);
nand U22991 (N_22991,N_15870,N_13103);
xor U22992 (N_22992,N_14437,N_13879);
xnor U22993 (N_22993,N_15141,N_18202);
nor U22994 (N_22994,N_13164,N_13187);
and U22995 (N_22995,N_14842,N_14010);
and U22996 (N_22996,N_18133,N_18200);
nand U22997 (N_22997,N_15062,N_18069);
nand U22998 (N_22998,N_12982,N_18491);
nand U22999 (N_22999,N_14336,N_14081);
nor U23000 (N_23000,N_14822,N_17900);
nand U23001 (N_23001,N_12940,N_13188);
and U23002 (N_23002,N_12669,N_14882);
nand U23003 (N_23003,N_13246,N_14259);
nor U23004 (N_23004,N_14251,N_16024);
nor U23005 (N_23005,N_16013,N_17103);
nand U23006 (N_23006,N_13388,N_15808);
and U23007 (N_23007,N_16907,N_13227);
nor U23008 (N_23008,N_15744,N_17295);
or U23009 (N_23009,N_16630,N_14392);
nor U23010 (N_23010,N_13739,N_15347);
nand U23011 (N_23011,N_17776,N_15770);
xor U23012 (N_23012,N_12763,N_13963);
or U23013 (N_23013,N_17615,N_18550);
xor U23014 (N_23014,N_17920,N_18578);
or U23015 (N_23015,N_15177,N_17966);
nor U23016 (N_23016,N_16890,N_18395);
nor U23017 (N_23017,N_15168,N_17284);
and U23018 (N_23018,N_14958,N_13651);
and U23019 (N_23019,N_14043,N_15076);
nor U23020 (N_23020,N_15200,N_16031);
nor U23021 (N_23021,N_13623,N_14072);
or U23022 (N_23022,N_15708,N_13809);
nor U23023 (N_23023,N_17910,N_14138);
and U23024 (N_23024,N_14264,N_13045);
nand U23025 (N_23025,N_17049,N_16486);
or U23026 (N_23026,N_18043,N_17324);
and U23027 (N_23027,N_17941,N_18353);
xor U23028 (N_23028,N_17233,N_18348);
and U23029 (N_23029,N_17337,N_13989);
xnor U23030 (N_23030,N_14271,N_17978);
and U23031 (N_23031,N_15846,N_14577);
nand U23032 (N_23032,N_14069,N_13431);
nor U23033 (N_23033,N_16796,N_18613);
xnor U23034 (N_23034,N_14280,N_17702);
nand U23035 (N_23035,N_17949,N_15248);
and U23036 (N_23036,N_14439,N_14688);
or U23037 (N_23037,N_12833,N_15518);
nor U23038 (N_23038,N_14261,N_14755);
nor U23039 (N_23039,N_15137,N_15234);
nand U23040 (N_23040,N_15590,N_13110);
or U23041 (N_23041,N_13939,N_12541);
and U23042 (N_23042,N_18346,N_12545);
or U23043 (N_23043,N_17921,N_17318);
nand U23044 (N_23044,N_14520,N_16094);
xnor U23045 (N_23045,N_17425,N_17982);
nor U23046 (N_23046,N_14478,N_13259);
and U23047 (N_23047,N_13518,N_15297);
and U23048 (N_23048,N_13794,N_16204);
and U23049 (N_23049,N_18717,N_13380);
and U23050 (N_23050,N_13270,N_18727);
or U23051 (N_23051,N_17943,N_14843);
nand U23052 (N_23052,N_16671,N_15388);
nand U23053 (N_23053,N_16248,N_17684);
or U23054 (N_23054,N_15234,N_15477);
nor U23055 (N_23055,N_15617,N_13610);
nand U23056 (N_23056,N_17085,N_17747);
nand U23057 (N_23057,N_15720,N_13944);
nand U23058 (N_23058,N_13192,N_17453);
or U23059 (N_23059,N_17142,N_13529);
xor U23060 (N_23060,N_16886,N_13350);
xor U23061 (N_23061,N_18455,N_13536);
and U23062 (N_23062,N_14739,N_16471);
or U23063 (N_23063,N_14379,N_16803);
nand U23064 (N_23064,N_16981,N_15989);
or U23065 (N_23065,N_18399,N_15208);
or U23066 (N_23066,N_14403,N_14866);
nand U23067 (N_23067,N_14221,N_13504);
and U23068 (N_23068,N_15232,N_14470);
xor U23069 (N_23069,N_14348,N_16299);
and U23070 (N_23070,N_14250,N_14006);
nand U23071 (N_23071,N_17489,N_17629);
and U23072 (N_23072,N_13846,N_17947);
and U23073 (N_23073,N_14993,N_15051);
and U23074 (N_23074,N_12776,N_13730);
and U23075 (N_23075,N_12864,N_12866);
xnor U23076 (N_23076,N_18410,N_16791);
nand U23077 (N_23077,N_16742,N_18029);
nand U23078 (N_23078,N_17837,N_16376);
nand U23079 (N_23079,N_13993,N_13957);
nor U23080 (N_23080,N_15222,N_14949);
or U23081 (N_23081,N_13535,N_14951);
xor U23082 (N_23082,N_15064,N_16589);
nor U23083 (N_23083,N_15244,N_18339);
and U23084 (N_23084,N_17273,N_15885);
and U23085 (N_23085,N_13329,N_18458);
xnor U23086 (N_23086,N_17142,N_15308);
or U23087 (N_23087,N_13745,N_18049);
nand U23088 (N_23088,N_13649,N_18692);
nor U23089 (N_23089,N_18734,N_17317);
nor U23090 (N_23090,N_13514,N_16801);
or U23091 (N_23091,N_16413,N_14007);
nor U23092 (N_23092,N_17739,N_17959);
nand U23093 (N_23093,N_18149,N_12592);
nor U23094 (N_23094,N_18104,N_16090);
or U23095 (N_23095,N_12717,N_17011);
nand U23096 (N_23096,N_17875,N_18735);
nor U23097 (N_23097,N_14969,N_15191);
or U23098 (N_23098,N_15804,N_17871);
xor U23099 (N_23099,N_13190,N_13978);
or U23100 (N_23100,N_17350,N_14932);
nor U23101 (N_23101,N_14294,N_18434);
or U23102 (N_23102,N_17084,N_12721);
or U23103 (N_23103,N_17548,N_15124);
or U23104 (N_23104,N_15383,N_13085);
nand U23105 (N_23105,N_13485,N_15984);
nand U23106 (N_23106,N_14364,N_12615);
or U23107 (N_23107,N_13361,N_17350);
nand U23108 (N_23108,N_15312,N_16820);
or U23109 (N_23109,N_13944,N_14725);
or U23110 (N_23110,N_16870,N_16530);
nand U23111 (N_23111,N_13919,N_12834);
nand U23112 (N_23112,N_14823,N_14746);
and U23113 (N_23113,N_16639,N_15114);
and U23114 (N_23114,N_18572,N_14917);
nand U23115 (N_23115,N_15395,N_14156);
and U23116 (N_23116,N_12598,N_13882);
nor U23117 (N_23117,N_14477,N_17183);
nor U23118 (N_23118,N_14270,N_18017);
nor U23119 (N_23119,N_13746,N_13742);
xnor U23120 (N_23120,N_16223,N_16374);
and U23121 (N_23121,N_17319,N_17494);
or U23122 (N_23122,N_17239,N_17573);
nor U23123 (N_23123,N_15799,N_14542);
nor U23124 (N_23124,N_18414,N_12589);
or U23125 (N_23125,N_18461,N_17307);
or U23126 (N_23126,N_16595,N_15790);
nand U23127 (N_23127,N_12732,N_13870);
xnor U23128 (N_23128,N_13755,N_15454);
nand U23129 (N_23129,N_15342,N_13745);
and U23130 (N_23130,N_17088,N_17022);
nand U23131 (N_23131,N_16493,N_16964);
nor U23132 (N_23132,N_15783,N_15858);
nor U23133 (N_23133,N_15206,N_14157);
and U23134 (N_23134,N_13353,N_12850);
and U23135 (N_23135,N_17735,N_16931);
and U23136 (N_23136,N_14980,N_16960);
xnor U23137 (N_23137,N_14589,N_18097);
nand U23138 (N_23138,N_16309,N_17999);
xor U23139 (N_23139,N_14518,N_17520);
nor U23140 (N_23140,N_12764,N_15635);
and U23141 (N_23141,N_17578,N_15163);
and U23142 (N_23142,N_18050,N_16942);
and U23143 (N_23143,N_12552,N_13296);
and U23144 (N_23144,N_14597,N_15006);
or U23145 (N_23145,N_13787,N_16600);
and U23146 (N_23146,N_15139,N_17474);
nor U23147 (N_23147,N_16727,N_18688);
nand U23148 (N_23148,N_13554,N_15789);
xor U23149 (N_23149,N_17905,N_16587);
nand U23150 (N_23150,N_17608,N_14415);
nand U23151 (N_23151,N_12691,N_15273);
and U23152 (N_23152,N_18532,N_12650);
nor U23153 (N_23153,N_16502,N_17728);
nand U23154 (N_23154,N_15913,N_13381);
nand U23155 (N_23155,N_15365,N_16429);
nand U23156 (N_23156,N_15534,N_14169);
xnor U23157 (N_23157,N_15808,N_17396);
and U23158 (N_23158,N_16542,N_12626);
nand U23159 (N_23159,N_17894,N_15695);
nor U23160 (N_23160,N_13134,N_17377);
or U23161 (N_23161,N_17929,N_13478);
and U23162 (N_23162,N_15571,N_17062);
xor U23163 (N_23163,N_13913,N_15055);
nand U23164 (N_23164,N_15905,N_12647);
and U23165 (N_23165,N_17309,N_14423);
nor U23166 (N_23166,N_18402,N_15580);
and U23167 (N_23167,N_12623,N_14947);
nand U23168 (N_23168,N_16754,N_13138);
nor U23169 (N_23169,N_17847,N_13228);
and U23170 (N_23170,N_14531,N_15013);
and U23171 (N_23171,N_15976,N_16256);
nand U23172 (N_23172,N_18624,N_14150);
nor U23173 (N_23173,N_17780,N_16345);
or U23174 (N_23174,N_14726,N_14283);
nor U23175 (N_23175,N_13239,N_17117);
nor U23176 (N_23176,N_14030,N_18025);
nor U23177 (N_23177,N_12693,N_12833);
nand U23178 (N_23178,N_14507,N_15199);
or U23179 (N_23179,N_14905,N_15726);
and U23180 (N_23180,N_16968,N_13371);
xor U23181 (N_23181,N_14664,N_14620);
nand U23182 (N_23182,N_18722,N_12682);
nor U23183 (N_23183,N_14125,N_16536);
and U23184 (N_23184,N_16734,N_16807);
and U23185 (N_23185,N_14310,N_16445);
or U23186 (N_23186,N_18632,N_12706);
xor U23187 (N_23187,N_16893,N_15906);
and U23188 (N_23188,N_18253,N_14513);
or U23189 (N_23189,N_16391,N_16230);
nand U23190 (N_23190,N_13955,N_13625);
or U23191 (N_23191,N_17057,N_17627);
nand U23192 (N_23192,N_14516,N_14517);
or U23193 (N_23193,N_17035,N_18225);
and U23194 (N_23194,N_18270,N_14805);
nor U23195 (N_23195,N_17187,N_15568);
nor U23196 (N_23196,N_17130,N_13490);
nor U23197 (N_23197,N_18126,N_17344);
nor U23198 (N_23198,N_16924,N_16551);
xnor U23199 (N_23199,N_15700,N_16228);
xnor U23200 (N_23200,N_18315,N_15483);
and U23201 (N_23201,N_14634,N_17990);
and U23202 (N_23202,N_16330,N_13222);
xor U23203 (N_23203,N_12521,N_15853);
xor U23204 (N_23204,N_18542,N_12959);
and U23205 (N_23205,N_15346,N_16960);
nand U23206 (N_23206,N_14593,N_15204);
nand U23207 (N_23207,N_15445,N_13195);
nor U23208 (N_23208,N_14615,N_17695);
nand U23209 (N_23209,N_12842,N_13692);
or U23210 (N_23210,N_16279,N_18039);
or U23211 (N_23211,N_15493,N_18363);
and U23212 (N_23212,N_15416,N_15617);
and U23213 (N_23213,N_12892,N_16215);
nand U23214 (N_23214,N_13412,N_12659);
nor U23215 (N_23215,N_16392,N_17235);
nand U23216 (N_23216,N_15013,N_13925);
nor U23217 (N_23217,N_16546,N_14036);
nand U23218 (N_23218,N_15310,N_12916);
nor U23219 (N_23219,N_13133,N_15541);
nor U23220 (N_23220,N_16366,N_13322);
nand U23221 (N_23221,N_13002,N_15807);
nor U23222 (N_23222,N_14363,N_17073);
nand U23223 (N_23223,N_17474,N_13687);
nand U23224 (N_23224,N_14235,N_17729);
and U23225 (N_23225,N_15235,N_13000);
or U23226 (N_23226,N_16193,N_16118);
nor U23227 (N_23227,N_17179,N_14411);
and U23228 (N_23228,N_12720,N_13007);
nand U23229 (N_23229,N_15586,N_13236);
nor U23230 (N_23230,N_14590,N_16873);
xnor U23231 (N_23231,N_16672,N_13089);
nand U23232 (N_23232,N_13946,N_13457);
nor U23233 (N_23233,N_13739,N_18012);
and U23234 (N_23234,N_17742,N_15441);
nand U23235 (N_23235,N_14912,N_17881);
and U23236 (N_23236,N_15815,N_15768);
nand U23237 (N_23237,N_13981,N_18336);
nand U23238 (N_23238,N_16720,N_15695);
or U23239 (N_23239,N_12754,N_13714);
and U23240 (N_23240,N_12908,N_12829);
and U23241 (N_23241,N_13652,N_14823);
nor U23242 (N_23242,N_16235,N_17509);
or U23243 (N_23243,N_17495,N_17309);
nor U23244 (N_23244,N_13425,N_18299);
nand U23245 (N_23245,N_16003,N_17908);
or U23246 (N_23246,N_13059,N_15378);
nor U23247 (N_23247,N_13779,N_14107);
nor U23248 (N_23248,N_18083,N_16067);
nand U23249 (N_23249,N_13972,N_12631);
and U23250 (N_23250,N_13958,N_16978);
nor U23251 (N_23251,N_12741,N_15079);
or U23252 (N_23252,N_13273,N_15594);
and U23253 (N_23253,N_17640,N_15633);
nand U23254 (N_23254,N_13120,N_17470);
or U23255 (N_23255,N_18291,N_15522);
nand U23256 (N_23256,N_16766,N_17639);
nor U23257 (N_23257,N_18324,N_16471);
nor U23258 (N_23258,N_16397,N_16374);
nor U23259 (N_23259,N_18121,N_18184);
and U23260 (N_23260,N_18680,N_18233);
nand U23261 (N_23261,N_14512,N_15320);
nor U23262 (N_23262,N_18120,N_13480);
nand U23263 (N_23263,N_16344,N_13576);
xor U23264 (N_23264,N_17367,N_17495);
nand U23265 (N_23265,N_14668,N_15078);
nor U23266 (N_23266,N_15449,N_14864);
nor U23267 (N_23267,N_17485,N_12843);
xor U23268 (N_23268,N_14973,N_18162);
nand U23269 (N_23269,N_13250,N_17662);
nor U23270 (N_23270,N_15257,N_13991);
or U23271 (N_23271,N_14396,N_18278);
nand U23272 (N_23272,N_13381,N_18300);
nand U23273 (N_23273,N_18470,N_15672);
xnor U23274 (N_23274,N_12621,N_18477);
and U23275 (N_23275,N_14866,N_15775);
nor U23276 (N_23276,N_15889,N_16278);
nor U23277 (N_23277,N_17419,N_12944);
and U23278 (N_23278,N_14884,N_16256);
and U23279 (N_23279,N_14401,N_13989);
and U23280 (N_23280,N_17275,N_17399);
nor U23281 (N_23281,N_17175,N_16591);
and U23282 (N_23282,N_16082,N_17853);
nand U23283 (N_23283,N_14492,N_14995);
nand U23284 (N_23284,N_17475,N_15314);
xnor U23285 (N_23285,N_17219,N_12579);
nand U23286 (N_23286,N_18523,N_12644);
and U23287 (N_23287,N_14890,N_16732);
nand U23288 (N_23288,N_17560,N_14648);
and U23289 (N_23289,N_17654,N_16036);
or U23290 (N_23290,N_12931,N_17180);
and U23291 (N_23291,N_12656,N_14337);
nor U23292 (N_23292,N_13461,N_18533);
nand U23293 (N_23293,N_14767,N_15667);
nand U23294 (N_23294,N_13459,N_14614);
and U23295 (N_23295,N_14088,N_17173);
or U23296 (N_23296,N_16751,N_16988);
nor U23297 (N_23297,N_17000,N_14568);
xnor U23298 (N_23298,N_17889,N_15867);
or U23299 (N_23299,N_14313,N_17985);
and U23300 (N_23300,N_14230,N_15493);
or U23301 (N_23301,N_15767,N_17523);
nor U23302 (N_23302,N_18416,N_16878);
nor U23303 (N_23303,N_13363,N_14129);
nand U23304 (N_23304,N_15034,N_12617);
and U23305 (N_23305,N_14080,N_16120);
nor U23306 (N_23306,N_16089,N_12806);
xnor U23307 (N_23307,N_14138,N_15672);
xnor U23308 (N_23308,N_18191,N_16537);
nand U23309 (N_23309,N_14214,N_13738);
or U23310 (N_23310,N_17179,N_13403);
or U23311 (N_23311,N_14164,N_18459);
nor U23312 (N_23312,N_12507,N_17357);
and U23313 (N_23313,N_13470,N_13028);
nor U23314 (N_23314,N_16209,N_12764);
nand U23315 (N_23315,N_17409,N_18597);
and U23316 (N_23316,N_15698,N_17341);
nor U23317 (N_23317,N_14132,N_14025);
or U23318 (N_23318,N_14800,N_17981);
nor U23319 (N_23319,N_16936,N_13095);
or U23320 (N_23320,N_14245,N_15238);
xnor U23321 (N_23321,N_12845,N_12821);
nand U23322 (N_23322,N_12631,N_15730);
nand U23323 (N_23323,N_15903,N_18597);
nor U23324 (N_23324,N_16039,N_14763);
or U23325 (N_23325,N_17373,N_14467);
or U23326 (N_23326,N_13080,N_16184);
nand U23327 (N_23327,N_17254,N_15263);
nand U23328 (N_23328,N_16602,N_18329);
nor U23329 (N_23329,N_17275,N_16325);
or U23330 (N_23330,N_18024,N_16326);
nand U23331 (N_23331,N_14669,N_18563);
nand U23332 (N_23332,N_16086,N_17082);
or U23333 (N_23333,N_17303,N_17657);
nand U23334 (N_23334,N_14196,N_15328);
or U23335 (N_23335,N_16957,N_16584);
nand U23336 (N_23336,N_17070,N_16562);
nor U23337 (N_23337,N_13654,N_12965);
nor U23338 (N_23338,N_13889,N_12677);
nor U23339 (N_23339,N_13650,N_15873);
nor U23340 (N_23340,N_18667,N_12975);
nand U23341 (N_23341,N_12743,N_17757);
nand U23342 (N_23342,N_18191,N_15635);
nor U23343 (N_23343,N_18729,N_14451);
and U23344 (N_23344,N_16449,N_13370);
and U23345 (N_23345,N_16833,N_18654);
nand U23346 (N_23346,N_13938,N_18375);
nor U23347 (N_23347,N_12762,N_14692);
and U23348 (N_23348,N_13646,N_17807);
and U23349 (N_23349,N_13348,N_17581);
nand U23350 (N_23350,N_12524,N_14105);
and U23351 (N_23351,N_18036,N_14734);
nor U23352 (N_23352,N_15705,N_14987);
nor U23353 (N_23353,N_15755,N_16871);
or U23354 (N_23354,N_12634,N_17765);
nand U23355 (N_23355,N_13215,N_16223);
and U23356 (N_23356,N_12968,N_15775);
nand U23357 (N_23357,N_12962,N_14872);
nor U23358 (N_23358,N_18522,N_16431);
nor U23359 (N_23359,N_15984,N_16833);
and U23360 (N_23360,N_16565,N_16769);
and U23361 (N_23361,N_17455,N_12750);
nand U23362 (N_23362,N_14222,N_15258);
and U23363 (N_23363,N_13899,N_17933);
xnor U23364 (N_23364,N_13513,N_14488);
and U23365 (N_23365,N_13925,N_16062);
or U23366 (N_23366,N_15385,N_16751);
and U23367 (N_23367,N_14326,N_12952);
and U23368 (N_23368,N_17848,N_13624);
nor U23369 (N_23369,N_16843,N_13552);
xor U23370 (N_23370,N_16031,N_16063);
nand U23371 (N_23371,N_18069,N_18021);
and U23372 (N_23372,N_17844,N_13476);
nor U23373 (N_23373,N_14092,N_14977);
nor U23374 (N_23374,N_13129,N_15528);
xnor U23375 (N_23375,N_18367,N_13770);
or U23376 (N_23376,N_14024,N_15135);
and U23377 (N_23377,N_17941,N_18195);
or U23378 (N_23378,N_18487,N_12547);
and U23379 (N_23379,N_15613,N_15800);
nor U23380 (N_23380,N_18579,N_18609);
and U23381 (N_23381,N_17368,N_12520);
nor U23382 (N_23382,N_17645,N_14526);
or U23383 (N_23383,N_16323,N_15000);
or U23384 (N_23384,N_14336,N_17072);
nor U23385 (N_23385,N_14170,N_15435);
and U23386 (N_23386,N_14245,N_18134);
nor U23387 (N_23387,N_16045,N_17070);
nor U23388 (N_23388,N_15778,N_12862);
or U23389 (N_23389,N_13353,N_16350);
and U23390 (N_23390,N_16816,N_16131);
or U23391 (N_23391,N_12725,N_13787);
nor U23392 (N_23392,N_16220,N_18713);
xnor U23393 (N_23393,N_12626,N_14875);
and U23394 (N_23394,N_12758,N_15129);
nand U23395 (N_23395,N_13952,N_14477);
or U23396 (N_23396,N_16024,N_13019);
nand U23397 (N_23397,N_16627,N_12906);
nand U23398 (N_23398,N_13759,N_18745);
nor U23399 (N_23399,N_13653,N_13173);
nor U23400 (N_23400,N_18142,N_14632);
xnor U23401 (N_23401,N_13676,N_16335);
nor U23402 (N_23402,N_14453,N_16134);
nand U23403 (N_23403,N_14576,N_14447);
nor U23404 (N_23404,N_15440,N_17607);
nor U23405 (N_23405,N_12556,N_15797);
xnor U23406 (N_23406,N_17403,N_13341);
or U23407 (N_23407,N_15327,N_18266);
nand U23408 (N_23408,N_18420,N_14508);
xnor U23409 (N_23409,N_14229,N_18671);
and U23410 (N_23410,N_13333,N_17079);
xor U23411 (N_23411,N_18531,N_18035);
nor U23412 (N_23412,N_15314,N_16561);
nand U23413 (N_23413,N_16731,N_14529);
nor U23414 (N_23414,N_16262,N_18173);
nand U23415 (N_23415,N_14862,N_12974);
or U23416 (N_23416,N_17023,N_18158);
and U23417 (N_23417,N_17833,N_15958);
nand U23418 (N_23418,N_12886,N_17648);
or U23419 (N_23419,N_12680,N_18114);
nand U23420 (N_23420,N_13189,N_16543);
or U23421 (N_23421,N_14346,N_15561);
nand U23422 (N_23422,N_13861,N_12692);
and U23423 (N_23423,N_17884,N_16333);
nand U23424 (N_23424,N_15754,N_16482);
or U23425 (N_23425,N_14154,N_18569);
nand U23426 (N_23426,N_18516,N_13202);
and U23427 (N_23427,N_15923,N_17814);
nor U23428 (N_23428,N_14257,N_14908);
and U23429 (N_23429,N_14871,N_12743);
nor U23430 (N_23430,N_16733,N_18245);
and U23431 (N_23431,N_17341,N_14149);
nand U23432 (N_23432,N_14390,N_16204);
xor U23433 (N_23433,N_14878,N_18020);
nand U23434 (N_23434,N_14726,N_16417);
nand U23435 (N_23435,N_18446,N_15306);
or U23436 (N_23436,N_14008,N_14302);
and U23437 (N_23437,N_15863,N_17900);
and U23438 (N_23438,N_16692,N_15171);
nand U23439 (N_23439,N_12625,N_17497);
and U23440 (N_23440,N_15325,N_14420);
or U23441 (N_23441,N_18573,N_15151);
nor U23442 (N_23442,N_17037,N_17855);
or U23443 (N_23443,N_15479,N_14800);
nor U23444 (N_23444,N_13452,N_18123);
nor U23445 (N_23445,N_16219,N_18286);
nand U23446 (N_23446,N_13526,N_16729);
nand U23447 (N_23447,N_13067,N_16846);
or U23448 (N_23448,N_16005,N_14131);
and U23449 (N_23449,N_17124,N_14297);
and U23450 (N_23450,N_16155,N_15620);
and U23451 (N_23451,N_17526,N_14507);
xor U23452 (N_23452,N_16123,N_13540);
and U23453 (N_23453,N_14416,N_16197);
nor U23454 (N_23454,N_14212,N_15686);
and U23455 (N_23455,N_12849,N_14782);
and U23456 (N_23456,N_14155,N_15769);
or U23457 (N_23457,N_15175,N_15961);
nor U23458 (N_23458,N_17413,N_14780);
nor U23459 (N_23459,N_12778,N_14539);
and U23460 (N_23460,N_18245,N_15542);
nand U23461 (N_23461,N_12534,N_15855);
nand U23462 (N_23462,N_18414,N_18639);
nor U23463 (N_23463,N_14289,N_18236);
or U23464 (N_23464,N_14809,N_18317);
nor U23465 (N_23465,N_16094,N_14237);
and U23466 (N_23466,N_16275,N_18150);
or U23467 (N_23467,N_14616,N_17508);
nor U23468 (N_23468,N_17689,N_15476);
nor U23469 (N_23469,N_15734,N_15033);
or U23470 (N_23470,N_18737,N_16394);
or U23471 (N_23471,N_14806,N_12578);
and U23472 (N_23472,N_12905,N_17961);
nand U23473 (N_23473,N_13008,N_13411);
nand U23474 (N_23474,N_15499,N_15952);
nand U23475 (N_23475,N_13655,N_17371);
or U23476 (N_23476,N_18219,N_14179);
xnor U23477 (N_23477,N_16550,N_13324);
and U23478 (N_23478,N_18197,N_14789);
and U23479 (N_23479,N_15060,N_15485);
nor U23480 (N_23480,N_12505,N_16722);
xnor U23481 (N_23481,N_15793,N_17600);
nand U23482 (N_23482,N_13087,N_18614);
or U23483 (N_23483,N_15230,N_15167);
or U23484 (N_23484,N_13747,N_15381);
nor U23485 (N_23485,N_16436,N_16616);
nor U23486 (N_23486,N_17808,N_12690);
nor U23487 (N_23487,N_18393,N_16175);
and U23488 (N_23488,N_15148,N_13528);
nor U23489 (N_23489,N_15853,N_14537);
or U23490 (N_23490,N_17458,N_17018);
or U23491 (N_23491,N_14852,N_14558);
or U23492 (N_23492,N_18078,N_14564);
nand U23493 (N_23493,N_14210,N_14022);
xor U23494 (N_23494,N_14997,N_18121);
nor U23495 (N_23495,N_12915,N_17607);
xor U23496 (N_23496,N_18195,N_12827);
nand U23497 (N_23497,N_13975,N_14465);
xnor U23498 (N_23498,N_13015,N_17733);
and U23499 (N_23499,N_15835,N_15701);
nor U23500 (N_23500,N_17830,N_15752);
nand U23501 (N_23501,N_17440,N_18523);
or U23502 (N_23502,N_18046,N_18234);
or U23503 (N_23503,N_13797,N_13242);
and U23504 (N_23504,N_13938,N_18160);
nor U23505 (N_23505,N_12877,N_12730);
or U23506 (N_23506,N_13718,N_15293);
nand U23507 (N_23507,N_13741,N_14913);
nor U23508 (N_23508,N_15639,N_18582);
nor U23509 (N_23509,N_18674,N_15447);
nor U23510 (N_23510,N_14338,N_14742);
and U23511 (N_23511,N_14642,N_17775);
and U23512 (N_23512,N_12606,N_15485);
or U23513 (N_23513,N_13429,N_13885);
nor U23514 (N_23514,N_12775,N_14453);
or U23515 (N_23515,N_17203,N_15830);
nand U23516 (N_23516,N_13781,N_15573);
nor U23517 (N_23517,N_16034,N_15505);
nor U23518 (N_23518,N_16413,N_17915);
nor U23519 (N_23519,N_17435,N_16831);
or U23520 (N_23520,N_16230,N_15611);
and U23521 (N_23521,N_16309,N_13697);
and U23522 (N_23522,N_17036,N_13515);
or U23523 (N_23523,N_13182,N_16089);
nand U23524 (N_23524,N_16497,N_13195);
nand U23525 (N_23525,N_15510,N_17238);
nand U23526 (N_23526,N_12876,N_18736);
nor U23527 (N_23527,N_16316,N_16398);
or U23528 (N_23528,N_13671,N_17115);
or U23529 (N_23529,N_18087,N_13331);
or U23530 (N_23530,N_14811,N_17255);
xor U23531 (N_23531,N_15480,N_13531);
xnor U23532 (N_23532,N_17878,N_13433);
or U23533 (N_23533,N_15663,N_15768);
or U23534 (N_23534,N_17987,N_18419);
or U23535 (N_23535,N_17761,N_12577);
nand U23536 (N_23536,N_15348,N_17488);
nor U23537 (N_23537,N_16881,N_13821);
and U23538 (N_23538,N_18136,N_14910);
nor U23539 (N_23539,N_12843,N_14692);
nand U23540 (N_23540,N_17886,N_12691);
and U23541 (N_23541,N_14026,N_14047);
or U23542 (N_23542,N_13697,N_16339);
nor U23543 (N_23543,N_16790,N_18587);
nor U23544 (N_23544,N_14822,N_13589);
or U23545 (N_23545,N_18403,N_12819);
or U23546 (N_23546,N_17576,N_16990);
nand U23547 (N_23547,N_18607,N_15157);
nand U23548 (N_23548,N_17897,N_15711);
nor U23549 (N_23549,N_13445,N_14809);
nand U23550 (N_23550,N_17765,N_17077);
nor U23551 (N_23551,N_14485,N_16265);
nor U23552 (N_23552,N_15552,N_13814);
nor U23553 (N_23553,N_16155,N_17099);
and U23554 (N_23554,N_16303,N_15776);
and U23555 (N_23555,N_14590,N_13735);
nor U23556 (N_23556,N_12931,N_18092);
nor U23557 (N_23557,N_13779,N_14987);
and U23558 (N_23558,N_15292,N_17050);
or U23559 (N_23559,N_17822,N_16855);
nand U23560 (N_23560,N_13074,N_15710);
nor U23561 (N_23561,N_13104,N_13541);
and U23562 (N_23562,N_14384,N_15219);
and U23563 (N_23563,N_15258,N_13245);
and U23564 (N_23564,N_18457,N_14194);
nand U23565 (N_23565,N_16372,N_17562);
and U23566 (N_23566,N_15450,N_13268);
nor U23567 (N_23567,N_18525,N_14104);
or U23568 (N_23568,N_14856,N_12902);
nor U23569 (N_23569,N_14954,N_17857);
or U23570 (N_23570,N_12730,N_16254);
xnor U23571 (N_23571,N_15378,N_15872);
or U23572 (N_23572,N_13830,N_17355);
or U23573 (N_23573,N_14976,N_15408);
and U23574 (N_23574,N_15394,N_17187);
or U23575 (N_23575,N_12581,N_15479);
nor U23576 (N_23576,N_18672,N_15106);
xnor U23577 (N_23577,N_12809,N_12738);
and U23578 (N_23578,N_15478,N_18207);
or U23579 (N_23579,N_16584,N_17300);
and U23580 (N_23580,N_18720,N_14949);
nor U23581 (N_23581,N_17176,N_14776);
nand U23582 (N_23582,N_16996,N_18745);
nand U23583 (N_23583,N_17604,N_17445);
nand U23584 (N_23584,N_17106,N_14089);
or U23585 (N_23585,N_18083,N_16720);
or U23586 (N_23586,N_17127,N_17617);
and U23587 (N_23587,N_17648,N_17612);
nor U23588 (N_23588,N_18671,N_13578);
xor U23589 (N_23589,N_18472,N_13973);
or U23590 (N_23590,N_15986,N_16737);
xor U23591 (N_23591,N_18301,N_17431);
nor U23592 (N_23592,N_16678,N_13739);
and U23593 (N_23593,N_16483,N_13626);
or U23594 (N_23594,N_14499,N_15732);
nor U23595 (N_23595,N_15365,N_17973);
nor U23596 (N_23596,N_16494,N_12840);
or U23597 (N_23597,N_14358,N_13603);
or U23598 (N_23598,N_15766,N_14074);
or U23599 (N_23599,N_18606,N_17767);
xnor U23600 (N_23600,N_14355,N_18608);
nor U23601 (N_23601,N_15106,N_14836);
and U23602 (N_23602,N_13558,N_15920);
nor U23603 (N_23603,N_15821,N_14195);
nand U23604 (N_23604,N_12996,N_15961);
or U23605 (N_23605,N_12555,N_14000);
and U23606 (N_23606,N_13504,N_14092);
or U23607 (N_23607,N_17773,N_12842);
and U23608 (N_23608,N_15718,N_17026);
and U23609 (N_23609,N_18246,N_17474);
or U23610 (N_23610,N_18371,N_18195);
nor U23611 (N_23611,N_13671,N_17420);
nor U23612 (N_23612,N_12574,N_14774);
or U23613 (N_23613,N_17925,N_14835);
or U23614 (N_23614,N_14881,N_13726);
xor U23615 (N_23615,N_15153,N_17310);
nand U23616 (N_23616,N_17125,N_15554);
nor U23617 (N_23617,N_15909,N_17872);
and U23618 (N_23618,N_18262,N_13308);
or U23619 (N_23619,N_18463,N_18191);
nor U23620 (N_23620,N_15641,N_14501);
nor U23621 (N_23621,N_17233,N_16406);
nand U23622 (N_23622,N_18116,N_15922);
or U23623 (N_23623,N_13169,N_18296);
nand U23624 (N_23624,N_14433,N_13598);
nor U23625 (N_23625,N_15714,N_14568);
and U23626 (N_23626,N_13365,N_14411);
nand U23627 (N_23627,N_15454,N_18183);
nor U23628 (N_23628,N_15238,N_14219);
or U23629 (N_23629,N_18073,N_17831);
or U23630 (N_23630,N_14348,N_14094);
or U23631 (N_23631,N_12897,N_18548);
nand U23632 (N_23632,N_16210,N_12935);
and U23633 (N_23633,N_13583,N_15491);
or U23634 (N_23634,N_18498,N_18226);
and U23635 (N_23635,N_12951,N_13904);
or U23636 (N_23636,N_17882,N_16986);
and U23637 (N_23637,N_15790,N_16376);
or U23638 (N_23638,N_16016,N_18535);
and U23639 (N_23639,N_13164,N_14472);
and U23640 (N_23640,N_16451,N_14849);
nor U23641 (N_23641,N_16124,N_16466);
xor U23642 (N_23642,N_16084,N_16426);
and U23643 (N_23643,N_16789,N_15843);
and U23644 (N_23644,N_14377,N_14055);
and U23645 (N_23645,N_16584,N_12571);
nand U23646 (N_23646,N_18346,N_15450);
nand U23647 (N_23647,N_12739,N_15823);
xor U23648 (N_23648,N_16946,N_13420);
and U23649 (N_23649,N_17928,N_18063);
nor U23650 (N_23650,N_16606,N_13988);
nand U23651 (N_23651,N_16909,N_14006);
nor U23652 (N_23652,N_14038,N_13322);
nand U23653 (N_23653,N_14711,N_17398);
nand U23654 (N_23654,N_14789,N_13897);
and U23655 (N_23655,N_14410,N_18728);
nand U23656 (N_23656,N_12678,N_17487);
nor U23657 (N_23657,N_12523,N_15362);
or U23658 (N_23658,N_15641,N_12908);
xor U23659 (N_23659,N_12577,N_18165);
nand U23660 (N_23660,N_15460,N_17900);
nand U23661 (N_23661,N_13803,N_17386);
xor U23662 (N_23662,N_13785,N_16247);
nor U23663 (N_23663,N_18609,N_13667);
nand U23664 (N_23664,N_17879,N_18637);
and U23665 (N_23665,N_17221,N_15746);
xor U23666 (N_23666,N_17042,N_14668);
or U23667 (N_23667,N_15479,N_13325);
nand U23668 (N_23668,N_13501,N_17224);
or U23669 (N_23669,N_18297,N_12831);
nand U23670 (N_23670,N_18251,N_14905);
nor U23671 (N_23671,N_12720,N_18176);
nor U23672 (N_23672,N_14874,N_18474);
nand U23673 (N_23673,N_13676,N_17443);
nor U23674 (N_23674,N_17717,N_17097);
nor U23675 (N_23675,N_12639,N_18125);
and U23676 (N_23676,N_15082,N_13927);
xnor U23677 (N_23677,N_16630,N_14051);
nand U23678 (N_23678,N_17398,N_14079);
xor U23679 (N_23679,N_17486,N_17522);
and U23680 (N_23680,N_15467,N_14691);
and U23681 (N_23681,N_13240,N_12776);
and U23682 (N_23682,N_18059,N_16869);
xor U23683 (N_23683,N_17029,N_16443);
xor U23684 (N_23684,N_15363,N_12816);
nor U23685 (N_23685,N_14300,N_15105);
and U23686 (N_23686,N_15638,N_12865);
or U23687 (N_23687,N_15935,N_14900);
or U23688 (N_23688,N_13257,N_16188);
nor U23689 (N_23689,N_15278,N_14181);
nand U23690 (N_23690,N_18431,N_14022);
nor U23691 (N_23691,N_18635,N_13190);
and U23692 (N_23692,N_18257,N_18430);
and U23693 (N_23693,N_15499,N_17495);
or U23694 (N_23694,N_14661,N_17702);
and U23695 (N_23695,N_15959,N_16910);
nor U23696 (N_23696,N_12956,N_13696);
or U23697 (N_23697,N_13413,N_12674);
nor U23698 (N_23698,N_14573,N_17097);
or U23699 (N_23699,N_15976,N_13541);
nor U23700 (N_23700,N_15451,N_18079);
or U23701 (N_23701,N_15895,N_16505);
nor U23702 (N_23702,N_12925,N_15062);
and U23703 (N_23703,N_14716,N_17165);
nor U23704 (N_23704,N_16131,N_15383);
and U23705 (N_23705,N_16139,N_16197);
xor U23706 (N_23706,N_12714,N_18223);
and U23707 (N_23707,N_12708,N_14245);
or U23708 (N_23708,N_18655,N_17221);
or U23709 (N_23709,N_13302,N_15432);
or U23710 (N_23710,N_17235,N_18719);
nor U23711 (N_23711,N_13088,N_15666);
nand U23712 (N_23712,N_13923,N_13292);
or U23713 (N_23713,N_15386,N_18298);
nor U23714 (N_23714,N_16159,N_16485);
nor U23715 (N_23715,N_12647,N_17315);
nand U23716 (N_23716,N_17673,N_14779);
nor U23717 (N_23717,N_17386,N_16879);
or U23718 (N_23718,N_12646,N_16926);
and U23719 (N_23719,N_14067,N_16778);
xor U23720 (N_23720,N_16530,N_15007);
nand U23721 (N_23721,N_17811,N_14385);
nor U23722 (N_23722,N_15311,N_13083);
xnor U23723 (N_23723,N_14027,N_13696);
nand U23724 (N_23724,N_16492,N_18717);
nand U23725 (N_23725,N_18105,N_13155);
or U23726 (N_23726,N_15302,N_18148);
or U23727 (N_23727,N_18425,N_16995);
nor U23728 (N_23728,N_14539,N_12660);
or U23729 (N_23729,N_16243,N_14890);
nor U23730 (N_23730,N_15575,N_13817);
or U23731 (N_23731,N_13946,N_12784);
nand U23732 (N_23732,N_17763,N_13431);
nand U23733 (N_23733,N_12622,N_15626);
or U23734 (N_23734,N_17299,N_15953);
xnor U23735 (N_23735,N_16058,N_17993);
and U23736 (N_23736,N_13180,N_17524);
nor U23737 (N_23737,N_14689,N_15958);
or U23738 (N_23738,N_12597,N_17470);
or U23739 (N_23739,N_12621,N_18601);
xor U23740 (N_23740,N_12561,N_18035);
nor U23741 (N_23741,N_13089,N_16214);
and U23742 (N_23742,N_18646,N_16289);
or U23743 (N_23743,N_15513,N_18285);
and U23744 (N_23744,N_15931,N_14679);
nor U23745 (N_23745,N_16733,N_15853);
nand U23746 (N_23746,N_17476,N_18386);
and U23747 (N_23747,N_17455,N_15983);
and U23748 (N_23748,N_17041,N_13525);
xor U23749 (N_23749,N_14798,N_13689);
nor U23750 (N_23750,N_16314,N_17555);
xnor U23751 (N_23751,N_17813,N_18647);
or U23752 (N_23752,N_18628,N_13679);
nor U23753 (N_23753,N_16845,N_16022);
and U23754 (N_23754,N_17132,N_13655);
nor U23755 (N_23755,N_13913,N_16319);
and U23756 (N_23756,N_13960,N_15084);
xor U23757 (N_23757,N_16515,N_16901);
xnor U23758 (N_23758,N_17263,N_13849);
xnor U23759 (N_23759,N_16426,N_18559);
nor U23760 (N_23760,N_17994,N_13511);
nand U23761 (N_23761,N_17032,N_14066);
xnor U23762 (N_23762,N_16240,N_18602);
and U23763 (N_23763,N_13475,N_15154);
or U23764 (N_23764,N_17708,N_15716);
nand U23765 (N_23765,N_16165,N_17635);
and U23766 (N_23766,N_18630,N_12644);
nor U23767 (N_23767,N_12519,N_17993);
nand U23768 (N_23768,N_15665,N_17874);
nor U23769 (N_23769,N_15418,N_15917);
and U23770 (N_23770,N_17389,N_14967);
or U23771 (N_23771,N_15794,N_17357);
or U23772 (N_23772,N_18131,N_15206);
or U23773 (N_23773,N_15843,N_13472);
xor U23774 (N_23774,N_17254,N_15360);
and U23775 (N_23775,N_15394,N_16483);
nand U23776 (N_23776,N_12873,N_17925);
nand U23777 (N_23777,N_17153,N_17455);
or U23778 (N_23778,N_12531,N_17776);
nand U23779 (N_23779,N_14153,N_12839);
nor U23780 (N_23780,N_15926,N_16970);
or U23781 (N_23781,N_16322,N_16317);
and U23782 (N_23782,N_12533,N_18394);
nand U23783 (N_23783,N_14582,N_18103);
or U23784 (N_23784,N_16500,N_17545);
nand U23785 (N_23785,N_14905,N_17865);
and U23786 (N_23786,N_16134,N_12541);
nor U23787 (N_23787,N_13093,N_14442);
and U23788 (N_23788,N_13390,N_15508);
nand U23789 (N_23789,N_17313,N_17830);
and U23790 (N_23790,N_18119,N_13853);
xor U23791 (N_23791,N_17380,N_16767);
or U23792 (N_23792,N_17637,N_13219);
nor U23793 (N_23793,N_16572,N_13935);
nand U23794 (N_23794,N_18454,N_16021);
nor U23795 (N_23795,N_13072,N_15517);
or U23796 (N_23796,N_14514,N_18066);
nor U23797 (N_23797,N_15540,N_15826);
or U23798 (N_23798,N_15109,N_14038);
or U23799 (N_23799,N_18488,N_17384);
nor U23800 (N_23800,N_14996,N_16240);
or U23801 (N_23801,N_18547,N_15838);
or U23802 (N_23802,N_16372,N_12745);
or U23803 (N_23803,N_17890,N_16314);
or U23804 (N_23804,N_12610,N_16927);
xor U23805 (N_23805,N_15203,N_17883);
and U23806 (N_23806,N_18383,N_15266);
nor U23807 (N_23807,N_18031,N_17181);
or U23808 (N_23808,N_17318,N_15728);
nand U23809 (N_23809,N_16599,N_14576);
xnor U23810 (N_23810,N_17677,N_17177);
and U23811 (N_23811,N_14170,N_17219);
or U23812 (N_23812,N_18634,N_18065);
or U23813 (N_23813,N_14597,N_18600);
nand U23814 (N_23814,N_18595,N_16868);
and U23815 (N_23815,N_13482,N_13617);
nor U23816 (N_23816,N_17851,N_14193);
and U23817 (N_23817,N_12871,N_15181);
nand U23818 (N_23818,N_12501,N_15671);
nor U23819 (N_23819,N_15293,N_16675);
and U23820 (N_23820,N_13183,N_14868);
xor U23821 (N_23821,N_15270,N_14526);
nand U23822 (N_23822,N_16268,N_18028);
or U23823 (N_23823,N_18482,N_15833);
and U23824 (N_23824,N_13968,N_13571);
or U23825 (N_23825,N_16534,N_15258);
nor U23826 (N_23826,N_18595,N_13308);
nand U23827 (N_23827,N_14507,N_17567);
and U23828 (N_23828,N_17326,N_17215);
nand U23829 (N_23829,N_16741,N_17896);
nand U23830 (N_23830,N_16300,N_16343);
and U23831 (N_23831,N_16621,N_16528);
nand U23832 (N_23832,N_12924,N_12787);
or U23833 (N_23833,N_13713,N_13247);
nand U23834 (N_23834,N_16274,N_14991);
and U23835 (N_23835,N_17300,N_16666);
xor U23836 (N_23836,N_18200,N_14631);
nor U23837 (N_23837,N_14650,N_15486);
nor U23838 (N_23838,N_17092,N_13269);
and U23839 (N_23839,N_16701,N_13412);
and U23840 (N_23840,N_17648,N_14299);
or U23841 (N_23841,N_18712,N_17115);
xor U23842 (N_23842,N_14491,N_18371);
nor U23843 (N_23843,N_16776,N_13595);
and U23844 (N_23844,N_14281,N_18292);
nor U23845 (N_23845,N_14371,N_18615);
xor U23846 (N_23846,N_16948,N_13767);
or U23847 (N_23847,N_12867,N_13763);
nand U23848 (N_23848,N_16022,N_18168);
and U23849 (N_23849,N_18207,N_14467);
xnor U23850 (N_23850,N_14333,N_12856);
nand U23851 (N_23851,N_13030,N_13477);
nand U23852 (N_23852,N_15923,N_16786);
or U23853 (N_23853,N_15947,N_12687);
or U23854 (N_23854,N_17075,N_12537);
nand U23855 (N_23855,N_12570,N_15518);
or U23856 (N_23856,N_12539,N_16862);
and U23857 (N_23857,N_16126,N_17550);
and U23858 (N_23858,N_13334,N_15283);
nand U23859 (N_23859,N_14938,N_13872);
nand U23860 (N_23860,N_15437,N_18471);
and U23861 (N_23861,N_12618,N_16383);
nor U23862 (N_23862,N_13739,N_14331);
xnor U23863 (N_23863,N_14495,N_16950);
or U23864 (N_23864,N_17184,N_17819);
nor U23865 (N_23865,N_18254,N_13417);
or U23866 (N_23866,N_14786,N_18391);
nor U23867 (N_23867,N_18467,N_12664);
or U23868 (N_23868,N_18317,N_15002);
nand U23869 (N_23869,N_15466,N_18268);
and U23870 (N_23870,N_12672,N_17561);
or U23871 (N_23871,N_15675,N_16691);
nand U23872 (N_23872,N_14415,N_17497);
xnor U23873 (N_23873,N_16389,N_18096);
nand U23874 (N_23874,N_13972,N_18303);
nor U23875 (N_23875,N_16729,N_17650);
and U23876 (N_23876,N_15403,N_13747);
and U23877 (N_23877,N_13659,N_18045);
and U23878 (N_23878,N_12690,N_13205);
and U23879 (N_23879,N_16038,N_17224);
and U23880 (N_23880,N_14063,N_18244);
or U23881 (N_23881,N_12885,N_12777);
and U23882 (N_23882,N_14342,N_12990);
nor U23883 (N_23883,N_14508,N_18682);
nand U23884 (N_23884,N_14488,N_18126);
nor U23885 (N_23885,N_18221,N_16266);
nor U23886 (N_23886,N_18402,N_14110);
nand U23887 (N_23887,N_14878,N_16283);
nor U23888 (N_23888,N_12860,N_17140);
xor U23889 (N_23889,N_16818,N_15115);
and U23890 (N_23890,N_13820,N_17441);
nor U23891 (N_23891,N_12665,N_15924);
nand U23892 (N_23892,N_16052,N_17321);
nor U23893 (N_23893,N_17399,N_17192);
or U23894 (N_23894,N_12988,N_17958);
nand U23895 (N_23895,N_12665,N_14528);
nor U23896 (N_23896,N_16194,N_18443);
nor U23897 (N_23897,N_13762,N_12914);
or U23898 (N_23898,N_16158,N_13552);
and U23899 (N_23899,N_16515,N_13274);
and U23900 (N_23900,N_17000,N_13064);
and U23901 (N_23901,N_16151,N_15912);
xnor U23902 (N_23902,N_14598,N_17865);
nor U23903 (N_23903,N_17895,N_14731);
or U23904 (N_23904,N_12628,N_16102);
xor U23905 (N_23905,N_17682,N_13779);
nor U23906 (N_23906,N_12693,N_14074);
or U23907 (N_23907,N_16904,N_14586);
nand U23908 (N_23908,N_15682,N_17557);
nand U23909 (N_23909,N_12670,N_15615);
nand U23910 (N_23910,N_14875,N_15423);
and U23911 (N_23911,N_18267,N_13800);
nor U23912 (N_23912,N_17679,N_14190);
nor U23913 (N_23913,N_18729,N_18452);
nor U23914 (N_23914,N_14100,N_16120);
nand U23915 (N_23915,N_15885,N_12974);
nor U23916 (N_23916,N_16638,N_18717);
or U23917 (N_23917,N_15313,N_17674);
and U23918 (N_23918,N_16911,N_14131);
and U23919 (N_23919,N_13307,N_17259);
and U23920 (N_23920,N_16206,N_16241);
or U23921 (N_23921,N_15136,N_17809);
and U23922 (N_23922,N_13561,N_15124);
and U23923 (N_23923,N_15932,N_18144);
nand U23924 (N_23924,N_16706,N_15517);
and U23925 (N_23925,N_15248,N_15166);
nor U23926 (N_23926,N_17464,N_18550);
and U23927 (N_23927,N_16453,N_13118);
or U23928 (N_23928,N_12933,N_13271);
and U23929 (N_23929,N_18376,N_14233);
xnor U23930 (N_23930,N_18039,N_17496);
or U23931 (N_23931,N_12993,N_14212);
nand U23932 (N_23932,N_13948,N_12846);
nand U23933 (N_23933,N_18217,N_17382);
or U23934 (N_23934,N_17049,N_14492);
nand U23935 (N_23935,N_16982,N_17240);
nand U23936 (N_23936,N_18460,N_18155);
or U23937 (N_23937,N_16630,N_16910);
nand U23938 (N_23938,N_18722,N_17229);
and U23939 (N_23939,N_18199,N_16467);
nand U23940 (N_23940,N_17834,N_13918);
nand U23941 (N_23941,N_15413,N_14335);
nor U23942 (N_23942,N_13339,N_16520);
nor U23943 (N_23943,N_14606,N_17914);
nand U23944 (N_23944,N_12941,N_18674);
nor U23945 (N_23945,N_17308,N_13436);
or U23946 (N_23946,N_13287,N_18329);
nor U23947 (N_23947,N_16230,N_18327);
nor U23948 (N_23948,N_12875,N_13646);
nor U23949 (N_23949,N_15333,N_18359);
nand U23950 (N_23950,N_12721,N_16446);
nand U23951 (N_23951,N_14132,N_16749);
and U23952 (N_23952,N_16205,N_15123);
nand U23953 (N_23953,N_17597,N_16295);
or U23954 (N_23954,N_15546,N_15248);
and U23955 (N_23955,N_13001,N_13617);
or U23956 (N_23956,N_14392,N_18069);
xnor U23957 (N_23957,N_15908,N_15075);
nand U23958 (N_23958,N_14375,N_13008);
xnor U23959 (N_23959,N_12544,N_13806);
or U23960 (N_23960,N_18228,N_14855);
nor U23961 (N_23961,N_13341,N_15112);
nand U23962 (N_23962,N_14246,N_17855);
nor U23963 (N_23963,N_14385,N_13354);
nand U23964 (N_23964,N_15700,N_17947);
xnor U23965 (N_23965,N_15164,N_16584);
or U23966 (N_23966,N_12869,N_16174);
nor U23967 (N_23967,N_14373,N_13044);
or U23968 (N_23968,N_17430,N_13428);
nand U23969 (N_23969,N_17428,N_12735);
nand U23970 (N_23970,N_14850,N_15083);
or U23971 (N_23971,N_13948,N_12984);
xor U23972 (N_23972,N_15772,N_18404);
or U23973 (N_23973,N_18724,N_17255);
nor U23974 (N_23974,N_17192,N_13865);
nor U23975 (N_23975,N_17309,N_13783);
nand U23976 (N_23976,N_17497,N_15186);
nor U23977 (N_23977,N_18212,N_15280);
or U23978 (N_23978,N_16249,N_16535);
or U23979 (N_23979,N_17982,N_12549);
nor U23980 (N_23980,N_16476,N_17237);
nand U23981 (N_23981,N_18240,N_15152);
nor U23982 (N_23982,N_17816,N_17199);
and U23983 (N_23983,N_13629,N_16334);
nor U23984 (N_23984,N_12515,N_13313);
or U23985 (N_23985,N_12521,N_18555);
and U23986 (N_23986,N_14842,N_12883);
nor U23987 (N_23987,N_15416,N_15419);
or U23988 (N_23988,N_12869,N_15372);
and U23989 (N_23989,N_17205,N_13010);
and U23990 (N_23990,N_18710,N_13691);
and U23991 (N_23991,N_16220,N_17748);
xnor U23992 (N_23992,N_17989,N_14617);
xnor U23993 (N_23993,N_12897,N_15351);
nor U23994 (N_23994,N_14480,N_17444);
or U23995 (N_23995,N_15103,N_13628);
or U23996 (N_23996,N_18726,N_16376);
nor U23997 (N_23997,N_13011,N_13274);
nand U23998 (N_23998,N_15139,N_17217);
xor U23999 (N_23999,N_17857,N_16170);
nor U24000 (N_24000,N_15147,N_17234);
nand U24001 (N_24001,N_18005,N_15752);
nor U24002 (N_24002,N_18269,N_18133);
nand U24003 (N_24003,N_14696,N_17401);
and U24004 (N_24004,N_12560,N_13818);
and U24005 (N_24005,N_13026,N_15217);
and U24006 (N_24006,N_17209,N_14062);
nor U24007 (N_24007,N_15525,N_16007);
xor U24008 (N_24008,N_14292,N_15041);
nor U24009 (N_24009,N_16295,N_16763);
and U24010 (N_24010,N_13449,N_14964);
or U24011 (N_24011,N_15903,N_18339);
or U24012 (N_24012,N_13645,N_15292);
nand U24013 (N_24013,N_18161,N_18123);
nand U24014 (N_24014,N_16344,N_13365);
nor U24015 (N_24015,N_14181,N_13646);
nor U24016 (N_24016,N_18281,N_13965);
and U24017 (N_24017,N_14309,N_13843);
or U24018 (N_24018,N_16587,N_15281);
nor U24019 (N_24019,N_15792,N_16560);
nand U24020 (N_24020,N_16895,N_15912);
or U24021 (N_24021,N_17964,N_14304);
and U24022 (N_24022,N_16043,N_14928);
nand U24023 (N_24023,N_13421,N_17986);
xor U24024 (N_24024,N_18674,N_13932);
or U24025 (N_24025,N_13728,N_17438);
nand U24026 (N_24026,N_14530,N_14865);
or U24027 (N_24027,N_14439,N_15429);
and U24028 (N_24028,N_14450,N_12744);
nand U24029 (N_24029,N_15356,N_13650);
nand U24030 (N_24030,N_15890,N_16178);
nand U24031 (N_24031,N_12730,N_12736);
and U24032 (N_24032,N_13184,N_17577);
and U24033 (N_24033,N_13795,N_14247);
or U24034 (N_24034,N_17497,N_13889);
nand U24035 (N_24035,N_14066,N_15967);
xor U24036 (N_24036,N_17660,N_12972);
nand U24037 (N_24037,N_15824,N_13404);
nand U24038 (N_24038,N_15843,N_12677);
and U24039 (N_24039,N_17536,N_15803);
and U24040 (N_24040,N_16982,N_13950);
nand U24041 (N_24041,N_12845,N_13794);
and U24042 (N_24042,N_13788,N_14345);
or U24043 (N_24043,N_13198,N_15131);
and U24044 (N_24044,N_12837,N_16994);
nand U24045 (N_24045,N_14669,N_15789);
nand U24046 (N_24046,N_14142,N_14709);
or U24047 (N_24047,N_16173,N_12917);
nand U24048 (N_24048,N_18470,N_16093);
nor U24049 (N_24049,N_13902,N_15461);
and U24050 (N_24050,N_13848,N_17611);
xor U24051 (N_24051,N_17584,N_12838);
nand U24052 (N_24052,N_15065,N_18258);
nor U24053 (N_24053,N_16458,N_14016);
nor U24054 (N_24054,N_13888,N_14173);
and U24055 (N_24055,N_14087,N_17544);
nand U24056 (N_24056,N_13251,N_17060);
nor U24057 (N_24057,N_18270,N_16982);
or U24058 (N_24058,N_13817,N_16537);
or U24059 (N_24059,N_12829,N_17742);
nand U24060 (N_24060,N_16370,N_15136);
and U24061 (N_24061,N_18381,N_13350);
or U24062 (N_24062,N_14765,N_13344);
nand U24063 (N_24063,N_14250,N_17081);
nor U24064 (N_24064,N_14195,N_14418);
nor U24065 (N_24065,N_12541,N_13406);
or U24066 (N_24066,N_13881,N_15421);
and U24067 (N_24067,N_15240,N_14402);
nor U24068 (N_24068,N_17062,N_13025);
and U24069 (N_24069,N_12651,N_15639);
xor U24070 (N_24070,N_16692,N_13240);
and U24071 (N_24071,N_17134,N_16100);
or U24072 (N_24072,N_16895,N_15458);
xor U24073 (N_24073,N_16498,N_15990);
nor U24074 (N_24074,N_14286,N_12661);
nand U24075 (N_24075,N_15345,N_16362);
and U24076 (N_24076,N_16749,N_12539);
xnor U24077 (N_24077,N_14202,N_18115);
nand U24078 (N_24078,N_12811,N_14362);
or U24079 (N_24079,N_17627,N_12523);
or U24080 (N_24080,N_17019,N_15850);
nor U24081 (N_24081,N_14655,N_13379);
xor U24082 (N_24082,N_15583,N_15909);
xnor U24083 (N_24083,N_14407,N_17756);
nor U24084 (N_24084,N_18237,N_13727);
nor U24085 (N_24085,N_17621,N_18136);
nor U24086 (N_24086,N_15100,N_17957);
nor U24087 (N_24087,N_13200,N_17505);
xor U24088 (N_24088,N_18097,N_13958);
xnor U24089 (N_24089,N_14642,N_14236);
and U24090 (N_24090,N_13306,N_15058);
or U24091 (N_24091,N_15493,N_15602);
nor U24092 (N_24092,N_12678,N_13669);
nand U24093 (N_24093,N_17330,N_16152);
or U24094 (N_24094,N_12938,N_16972);
nor U24095 (N_24095,N_16030,N_13617);
or U24096 (N_24096,N_18516,N_17919);
nand U24097 (N_24097,N_18657,N_15622);
or U24098 (N_24098,N_16323,N_12700);
nor U24099 (N_24099,N_13373,N_15875);
nand U24100 (N_24100,N_12734,N_16034);
or U24101 (N_24101,N_16416,N_12610);
or U24102 (N_24102,N_14174,N_13725);
nor U24103 (N_24103,N_15550,N_17956);
or U24104 (N_24104,N_16875,N_14689);
nor U24105 (N_24105,N_15589,N_16811);
xnor U24106 (N_24106,N_13893,N_15424);
nor U24107 (N_24107,N_13651,N_18552);
nor U24108 (N_24108,N_14407,N_15669);
nand U24109 (N_24109,N_14189,N_17291);
xor U24110 (N_24110,N_18655,N_13909);
nand U24111 (N_24111,N_16427,N_15216);
nand U24112 (N_24112,N_12953,N_14909);
and U24113 (N_24113,N_17654,N_15852);
or U24114 (N_24114,N_15829,N_12751);
and U24115 (N_24115,N_14887,N_14562);
or U24116 (N_24116,N_16855,N_15085);
nor U24117 (N_24117,N_13887,N_15690);
nor U24118 (N_24118,N_18150,N_13940);
or U24119 (N_24119,N_16426,N_15513);
nor U24120 (N_24120,N_15396,N_13483);
nand U24121 (N_24121,N_12998,N_14461);
nor U24122 (N_24122,N_12825,N_15525);
nor U24123 (N_24123,N_13801,N_15071);
or U24124 (N_24124,N_16411,N_14563);
nor U24125 (N_24125,N_13739,N_14057);
nor U24126 (N_24126,N_12738,N_13528);
or U24127 (N_24127,N_17801,N_13437);
nor U24128 (N_24128,N_16111,N_17239);
and U24129 (N_24129,N_12580,N_18224);
or U24130 (N_24130,N_18242,N_15501);
nand U24131 (N_24131,N_14153,N_17459);
nor U24132 (N_24132,N_15010,N_16038);
and U24133 (N_24133,N_15704,N_18499);
nor U24134 (N_24134,N_15869,N_15657);
nor U24135 (N_24135,N_16256,N_15836);
xnor U24136 (N_24136,N_17418,N_16819);
nor U24137 (N_24137,N_17400,N_14715);
and U24138 (N_24138,N_15852,N_15041);
nor U24139 (N_24139,N_12781,N_13166);
nand U24140 (N_24140,N_17261,N_15694);
nand U24141 (N_24141,N_16720,N_18012);
or U24142 (N_24142,N_13249,N_13019);
or U24143 (N_24143,N_13626,N_12947);
nand U24144 (N_24144,N_12613,N_13380);
and U24145 (N_24145,N_16880,N_17054);
and U24146 (N_24146,N_12508,N_15054);
nor U24147 (N_24147,N_15158,N_14369);
nand U24148 (N_24148,N_14702,N_14110);
nor U24149 (N_24149,N_15586,N_14245);
and U24150 (N_24150,N_12792,N_13692);
xnor U24151 (N_24151,N_18410,N_17549);
or U24152 (N_24152,N_13587,N_16757);
and U24153 (N_24153,N_12873,N_18409);
nand U24154 (N_24154,N_17434,N_16451);
xor U24155 (N_24155,N_17154,N_15465);
or U24156 (N_24156,N_17841,N_16127);
nand U24157 (N_24157,N_16895,N_17700);
xor U24158 (N_24158,N_16542,N_13745);
nand U24159 (N_24159,N_14399,N_17887);
or U24160 (N_24160,N_17540,N_15313);
nor U24161 (N_24161,N_15916,N_17031);
nand U24162 (N_24162,N_12527,N_12819);
nand U24163 (N_24163,N_18691,N_12602);
nand U24164 (N_24164,N_15407,N_16799);
xnor U24165 (N_24165,N_17741,N_14161);
nor U24166 (N_24166,N_17426,N_15566);
nand U24167 (N_24167,N_14619,N_17608);
or U24168 (N_24168,N_15987,N_16423);
nor U24169 (N_24169,N_15923,N_14630);
and U24170 (N_24170,N_12719,N_16373);
nand U24171 (N_24171,N_12504,N_18425);
xor U24172 (N_24172,N_14743,N_13953);
or U24173 (N_24173,N_18600,N_15368);
nand U24174 (N_24174,N_13380,N_14852);
and U24175 (N_24175,N_14799,N_18590);
and U24176 (N_24176,N_18285,N_16866);
or U24177 (N_24177,N_16886,N_17945);
or U24178 (N_24178,N_13648,N_15102);
and U24179 (N_24179,N_14645,N_14177);
or U24180 (N_24180,N_13602,N_18688);
or U24181 (N_24181,N_16773,N_16574);
or U24182 (N_24182,N_18720,N_18729);
nor U24183 (N_24183,N_15893,N_13481);
or U24184 (N_24184,N_13560,N_15915);
nand U24185 (N_24185,N_18063,N_14940);
xor U24186 (N_24186,N_14510,N_16564);
nor U24187 (N_24187,N_17044,N_15534);
or U24188 (N_24188,N_14753,N_18482);
nor U24189 (N_24189,N_13167,N_12914);
nor U24190 (N_24190,N_15359,N_14245);
or U24191 (N_24191,N_13628,N_17299);
nor U24192 (N_24192,N_13113,N_13234);
and U24193 (N_24193,N_12845,N_12681);
nand U24194 (N_24194,N_13239,N_18162);
nor U24195 (N_24195,N_14849,N_16695);
nor U24196 (N_24196,N_13424,N_16213);
nor U24197 (N_24197,N_13636,N_14441);
nor U24198 (N_24198,N_15957,N_16307);
nor U24199 (N_24199,N_12608,N_12880);
nand U24200 (N_24200,N_16711,N_17115);
or U24201 (N_24201,N_17023,N_17425);
nor U24202 (N_24202,N_18645,N_16876);
or U24203 (N_24203,N_15781,N_17718);
and U24204 (N_24204,N_15879,N_18257);
and U24205 (N_24205,N_18136,N_15053);
nand U24206 (N_24206,N_14165,N_13381);
or U24207 (N_24207,N_16296,N_14628);
or U24208 (N_24208,N_14932,N_15420);
or U24209 (N_24209,N_16837,N_14431);
nand U24210 (N_24210,N_15993,N_15039);
and U24211 (N_24211,N_15037,N_17252);
nand U24212 (N_24212,N_15307,N_17467);
or U24213 (N_24213,N_18347,N_18088);
or U24214 (N_24214,N_17584,N_13994);
xnor U24215 (N_24215,N_15250,N_18625);
nor U24216 (N_24216,N_12967,N_12946);
nor U24217 (N_24217,N_14510,N_17030);
xnor U24218 (N_24218,N_13670,N_15394);
nor U24219 (N_24219,N_17497,N_16196);
nand U24220 (N_24220,N_18419,N_18649);
or U24221 (N_24221,N_18429,N_18515);
and U24222 (N_24222,N_14248,N_13738);
nand U24223 (N_24223,N_16633,N_15908);
nor U24224 (N_24224,N_14652,N_13674);
nor U24225 (N_24225,N_15633,N_16325);
nand U24226 (N_24226,N_15115,N_15209);
or U24227 (N_24227,N_16632,N_18616);
nand U24228 (N_24228,N_17210,N_17078);
nand U24229 (N_24229,N_14647,N_15355);
or U24230 (N_24230,N_18268,N_15324);
nor U24231 (N_24231,N_13204,N_14184);
nor U24232 (N_24232,N_13849,N_17021);
or U24233 (N_24233,N_12625,N_13696);
and U24234 (N_24234,N_17820,N_16616);
nor U24235 (N_24235,N_15240,N_17863);
nor U24236 (N_24236,N_18605,N_12543);
or U24237 (N_24237,N_15964,N_12906);
nor U24238 (N_24238,N_15625,N_15624);
xnor U24239 (N_24239,N_14818,N_13700);
nor U24240 (N_24240,N_16228,N_16062);
and U24241 (N_24241,N_15193,N_17719);
and U24242 (N_24242,N_18375,N_13193);
and U24243 (N_24243,N_13299,N_14964);
nand U24244 (N_24244,N_17528,N_18387);
nand U24245 (N_24245,N_17217,N_14431);
or U24246 (N_24246,N_13215,N_16558);
nand U24247 (N_24247,N_16265,N_12741);
nor U24248 (N_24248,N_12500,N_17027);
nor U24249 (N_24249,N_13621,N_15316);
or U24250 (N_24250,N_16582,N_18101);
nor U24251 (N_24251,N_18575,N_16284);
or U24252 (N_24252,N_15615,N_16092);
or U24253 (N_24253,N_15108,N_15315);
nor U24254 (N_24254,N_13947,N_13848);
or U24255 (N_24255,N_12866,N_15983);
and U24256 (N_24256,N_15035,N_17725);
nor U24257 (N_24257,N_14468,N_18387);
and U24258 (N_24258,N_16907,N_17676);
nand U24259 (N_24259,N_15141,N_17003);
xnor U24260 (N_24260,N_17794,N_14682);
nand U24261 (N_24261,N_15753,N_14246);
nor U24262 (N_24262,N_12686,N_13396);
nand U24263 (N_24263,N_18656,N_18366);
and U24264 (N_24264,N_12805,N_16486);
nand U24265 (N_24265,N_16987,N_16512);
and U24266 (N_24266,N_13552,N_18298);
nor U24267 (N_24267,N_18004,N_16980);
or U24268 (N_24268,N_18033,N_14688);
nand U24269 (N_24269,N_13951,N_14680);
nand U24270 (N_24270,N_18112,N_13738);
or U24271 (N_24271,N_13880,N_14428);
and U24272 (N_24272,N_13544,N_14062);
or U24273 (N_24273,N_17201,N_16565);
or U24274 (N_24274,N_14436,N_16128);
or U24275 (N_24275,N_17596,N_14567);
or U24276 (N_24276,N_14352,N_14587);
or U24277 (N_24277,N_18576,N_13951);
or U24278 (N_24278,N_17865,N_17710);
nor U24279 (N_24279,N_17439,N_16242);
and U24280 (N_24280,N_15156,N_14427);
and U24281 (N_24281,N_12757,N_15482);
or U24282 (N_24282,N_16069,N_13127);
or U24283 (N_24283,N_15051,N_17550);
and U24284 (N_24284,N_18619,N_13775);
and U24285 (N_24285,N_18435,N_17118);
nor U24286 (N_24286,N_13915,N_18397);
nand U24287 (N_24287,N_12749,N_17548);
nand U24288 (N_24288,N_14660,N_15985);
and U24289 (N_24289,N_15275,N_18026);
or U24290 (N_24290,N_16962,N_14138);
nor U24291 (N_24291,N_12677,N_12721);
nand U24292 (N_24292,N_17866,N_13962);
nand U24293 (N_24293,N_15631,N_14056);
and U24294 (N_24294,N_16083,N_13115);
nor U24295 (N_24295,N_18664,N_15863);
or U24296 (N_24296,N_16883,N_16020);
and U24297 (N_24297,N_17602,N_16842);
nor U24298 (N_24298,N_18638,N_14057);
and U24299 (N_24299,N_15095,N_17874);
nand U24300 (N_24300,N_15799,N_15180);
or U24301 (N_24301,N_18050,N_12823);
or U24302 (N_24302,N_16995,N_13139);
or U24303 (N_24303,N_16461,N_15937);
nand U24304 (N_24304,N_18628,N_17734);
nand U24305 (N_24305,N_12556,N_15694);
nand U24306 (N_24306,N_14357,N_13490);
nand U24307 (N_24307,N_14210,N_13385);
and U24308 (N_24308,N_17699,N_17656);
nand U24309 (N_24309,N_14452,N_17901);
nand U24310 (N_24310,N_17999,N_18273);
nor U24311 (N_24311,N_14540,N_18089);
nand U24312 (N_24312,N_14003,N_14162);
and U24313 (N_24313,N_16006,N_16214);
and U24314 (N_24314,N_18106,N_16506);
nor U24315 (N_24315,N_17670,N_16913);
nand U24316 (N_24316,N_15966,N_17826);
and U24317 (N_24317,N_16300,N_17648);
or U24318 (N_24318,N_16782,N_14838);
and U24319 (N_24319,N_15133,N_12784);
or U24320 (N_24320,N_17129,N_14463);
or U24321 (N_24321,N_14025,N_13639);
and U24322 (N_24322,N_14390,N_16292);
and U24323 (N_24323,N_17777,N_18625);
and U24324 (N_24324,N_18525,N_13228);
nor U24325 (N_24325,N_16020,N_14133);
and U24326 (N_24326,N_17548,N_15216);
xor U24327 (N_24327,N_17966,N_17457);
xor U24328 (N_24328,N_15443,N_17510);
or U24329 (N_24329,N_17873,N_18496);
xnor U24330 (N_24330,N_14186,N_14524);
or U24331 (N_24331,N_15851,N_18265);
or U24332 (N_24332,N_18041,N_16325);
or U24333 (N_24333,N_15513,N_16260);
or U24334 (N_24334,N_12657,N_18566);
or U24335 (N_24335,N_14725,N_14597);
nor U24336 (N_24336,N_16753,N_17890);
nand U24337 (N_24337,N_17394,N_17367);
nor U24338 (N_24338,N_17980,N_16607);
nor U24339 (N_24339,N_14103,N_16438);
nand U24340 (N_24340,N_16282,N_17080);
nand U24341 (N_24341,N_17500,N_15422);
nand U24342 (N_24342,N_17960,N_14879);
and U24343 (N_24343,N_13612,N_15906);
xnor U24344 (N_24344,N_15138,N_15872);
xor U24345 (N_24345,N_16830,N_13189);
or U24346 (N_24346,N_15691,N_16825);
and U24347 (N_24347,N_12537,N_16322);
nand U24348 (N_24348,N_16614,N_15812);
nand U24349 (N_24349,N_12832,N_13268);
and U24350 (N_24350,N_15892,N_15235);
nand U24351 (N_24351,N_16922,N_18013);
and U24352 (N_24352,N_14943,N_18503);
nand U24353 (N_24353,N_18419,N_17986);
nor U24354 (N_24354,N_18063,N_17746);
nand U24355 (N_24355,N_13507,N_17812);
or U24356 (N_24356,N_15033,N_17640);
and U24357 (N_24357,N_13362,N_16003);
or U24358 (N_24358,N_15341,N_14767);
and U24359 (N_24359,N_12504,N_12644);
nor U24360 (N_24360,N_13212,N_16724);
or U24361 (N_24361,N_14977,N_13789);
nor U24362 (N_24362,N_12566,N_17723);
nor U24363 (N_24363,N_16054,N_14981);
nor U24364 (N_24364,N_16185,N_17463);
and U24365 (N_24365,N_18000,N_14869);
nand U24366 (N_24366,N_17679,N_14096);
nor U24367 (N_24367,N_14205,N_18132);
or U24368 (N_24368,N_16920,N_13440);
or U24369 (N_24369,N_17662,N_15862);
xnor U24370 (N_24370,N_13393,N_16083);
or U24371 (N_24371,N_18231,N_17340);
and U24372 (N_24372,N_14617,N_17054);
xor U24373 (N_24373,N_14473,N_15834);
and U24374 (N_24374,N_15293,N_12742);
xnor U24375 (N_24375,N_14598,N_15913);
nand U24376 (N_24376,N_14241,N_14434);
nor U24377 (N_24377,N_13232,N_15465);
and U24378 (N_24378,N_12641,N_16904);
and U24379 (N_24379,N_15627,N_13808);
or U24380 (N_24380,N_17463,N_15232);
nor U24381 (N_24381,N_17937,N_17643);
nand U24382 (N_24382,N_14709,N_14378);
and U24383 (N_24383,N_16986,N_17181);
and U24384 (N_24384,N_14569,N_16630);
or U24385 (N_24385,N_14449,N_15919);
and U24386 (N_24386,N_16771,N_12871);
xnor U24387 (N_24387,N_17491,N_13160);
and U24388 (N_24388,N_17871,N_14506);
and U24389 (N_24389,N_16401,N_13483);
nand U24390 (N_24390,N_13422,N_17777);
and U24391 (N_24391,N_17066,N_17919);
and U24392 (N_24392,N_16532,N_15400);
and U24393 (N_24393,N_17236,N_15152);
nand U24394 (N_24394,N_14402,N_14155);
nor U24395 (N_24395,N_16113,N_12891);
nand U24396 (N_24396,N_15249,N_17506);
and U24397 (N_24397,N_16819,N_17562);
or U24398 (N_24398,N_15344,N_15905);
xor U24399 (N_24399,N_15927,N_16035);
nor U24400 (N_24400,N_12801,N_12928);
nor U24401 (N_24401,N_14916,N_18354);
and U24402 (N_24402,N_15468,N_13798);
xnor U24403 (N_24403,N_16020,N_18653);
nand U24404 (N_24404,N_17606,N_14228);
nor U24405 (N_24405,N_18402,N_13896);
nand U24406 (N_24406,N_16864,N_14181);
nand U24407 (N_24407,N_18525,N_15697);
or U24408 (N_24408,N_18107,N_18275);
and U24409 (N_24409,N_17403,N_17936);
nand U24410 (N_24410,N_16472,N_17239);
or U24411 (N_24411,N_17692,N_12738);
nor U24412 (N_24412,N_16264,N_15125);
xnor U24413 (N_24413,N_13493,N_13837);
xor U24414 (N_24414,N_15421,N_15917);
nor U24415 (N_24415,N_16904,N_12964);
and U24416 (N_24416,N_18603,N_12871);
and U24417 (N_24417,N_13265,N_18707);
nor U24418 (N_24418,N_17825,N_14440);
and U24419 (N_24419,N_15617,N_13401);
nor U24420 (N_24420,N_15599,N_14496);
and U24421 (N_24421,N_13942,N_15117);
nand U24422 (N_24422,N_15081,N_17898);
nor U24423 (N_24423,N_13899,N_16845);
and U24424 (N_24424,N_15709,N_12869);
xor U24425 (N_24425,N_13378,N_14363);
nand U24426 (N_24426,N_16684,N_15391);
nor U24427 (N_24427,N_15448,N_16641);
nor U24428 (N_24428,N_16401,N_12960);
nand U24429 (N_24429,N_12697,N_18371);
xnor U24430 (N_24430,N_16902,N_14266);
nand U24431 (N_24431,N_18563,N_15614);
or U24432 (N_24432,N_15462,N_16339);
nand U24433 (N_24433,N_15270,N_17701);
or U24434 (N_24434,N_16973,N_16780);
nand U24435 (N_24435,N_18143,N_17736);
nand U24436 (N_24436,N_16816,N_17397);
nand U24437 (N_24437,N_17562,N_18670);
nand U24438 (N_24438,N_15527,N_12629);
and U24439 (N_24439,N_13005,N_14831);
and U24440 (N_24440,N_18693,N_14993);
xor U24441 (N_24441,N_14881,N_15305);
nor U24442 (N_24442,N_15491,N_12795);
xnor U24443 (N_24443,N_15655,N_18267);
xor U24444 (N_24444,N_17759,N_17825);
or U24445 (N_24445,N_15011,N_14418);
xor U24446 (N_24446,N_13556,N_14203);
or U24447 (N_24447,N_15549,N_14474);
and U24448 (N_24448,N_15079,N_13989);
and U24449 (N_24449,N_17721,N_17724);
or U24450 (N_24450,N_17347,N_17054);
or U24451 (N_24451,N_17444,N_17698);
xnor U24452 (N_24452,N_13120,N_15791);
nor U24453 (N_24453,N_15714,N_17212);
nand U24454 (N_24454,N_16405,N_18153);
and U24455 (N_24455,N_17840,N_15667);
or U24456 (N_24456,N_15312,N_16629);
nor U24457 (N_24457,N_14490,N_13070);
nand U24458 (N_24458,N_17707,N_17053);
nor U24459 (N_24459,N_16219,N_12933);
xnor U24460 (N_24460,N_17076,N_18493);
or U24461 (N_24461,N_18715,N_12936);
xnor U24462 (N_24462,N_12642,N_18194);
or U24463 (N_24463,N_13531,N_16872);
nand U24464 (N_24464,N_14704,N_17593);
nor U24465 (N_24465,N_13188,N_17926);
or U24466 (N_24466,N_14716,N_15502);
and U24467 (N_24467,N_18636,N_15532);
or U24468 (N_24468,N_17522,N_14784);
nand U24469 (N_24469,N_14662,N_13744);
nand U24470 (N_24470,N_14380,N_16751);
nand U24471 (N_24471,N_14472,N_14090);
and U24472 (N_24472,N_15478,N_16441);
and U24473 (N_24473,N_15133,N_12826);
nand U24474 (N_24474,N_14383,N_12690);
and U24475 (N_24475,N_12821,N_14387);
nand U24476 (N_24476,N_13438,N_14065);
nor U24477 (N_24477,N_18137,N_13317);
or U24478 (N_24478,N_12592,N_14631);
nand U24479 (N_24479,N_13696,N_14794);
nor U24480 (N_24480,N_14380,N_17833);
or U24481 (N_24481,N_15239,N_13403);
nand U24482 (N_24482,N_15741,N_13614);
nor U24483 (N_24483,N_14048,N_17986);
nand U24484 (N_24484,N_16057,N_13618);
and U24485 (N_24485,N_14722,N_12583);
nor U24486 (N_24486,N_16083,N_14652);
and U24487 (N_24487,N_17172,N_13486);
and U24488 (N_24488,N_13430,N_17340);
nor U24489 (N_24489,N_16234,N_17083);
nand U24490 (N_24490,N_13412,N_13469);
nor U24491 (N_24491,N_18288,N_12847);
or U24492 (N_24492,N_13105,N_17249);
and U24493 (N_24493,N_16482,N_13040);
and U24494 (N_24494,N_17825,N_16246);
and U24495 (N_24495,N_17576,N_12804);
nor U24496 (N_24496,N_17428,N_18427);
and U24497 (N_24497,N_15015,N_15262);
or U24498 (N_24498,N_12563,N_13477);
or U24499 (N_24499,N_16234,N_15992);
nor U24500 (N_24500,N_18588,N_14409);
and U24501 (N_24501,N_12719,N_18158);
and U24502 (N_24502,N_17728,N_17725);
or U24503 (N_24503,N_17398,N_13647);
nor U24504 (N_24504,N_16411,N_12901);
nand U24505 (N_24505,N_14118,N_15238);
or U24506 (N_24506,N_18115,N_15494);
nand U24507 (N_24507,N_17422,N_15192);
and U24508 (N_24508,N_14813,N_17544);
nand U24509 (N_24509,N_16177,N_15998);
xor U24510 (N_24510,N_18640,N_15693);
and U24511 (N_24511,N_15437,N_12710);
and U24512 (N_24512,N_17562,N_14372);
nand U24513 (N_24513,N_15334,N_15439);
nor U24514 (N_24514,N_14835,N_15940);
xor U24515 (N_24515,N_17792,N_16482);
or U24516 (N_24516,N_16316,N_18352);
xnor U24517 (N_24517,N_16354,N_15941);
nor U24518 (N_24518,N_17323,N_12909);
nor U24519 (N_24519,N_16422,N_18247);
and U24520 (N_24520,N_12745,N_12975);
and U24521 (N_24521,N_17783,N_18749);
and U24522 (N_24522,N_13757,N_16894);
or U24523 (N_24523,N_12537,N_15919);
or U24524 (N_24524,N_13955,N_16921);
nor U24525 (N_24525,N_17928,N_16709);
nand U24526 (N_24526,N_15947,N_15908);
or U24527 (N_24527,N_13956,N_17470);
nor U24528 (N_24528,N_15414,N_17812);
and U24529 (N_24529,N_14217,N_12609);
or U24530 (N_24530,N_18177,N_17058);
nor U24531 (N_24531,N_15443,N_17279);
nand U24532 (N_24532,N_17257,N_14614);
nand U24533 (N_24533,N_17704,N_12739);
nor U24534 (N_24534,N_15165,N_17466);
nor U24535 (N_24535,N_16671,N_18436);
xnor U24536 (N_24536,N_14041,N_15319);
nor U24537 (N_24537,N_15756,N_14497);
or U24538 (N_24538,N_16526,N_12998);
xnor U24539 (N_24539,N_14410,N_14926);
nand U24540 (N_24540,N_14739,N_16263);
or U24541 (N_24541,N_18722,N_13876);
or U24542 (N_24542,N_15033,N_13500);
nand U24543 (N_24543,N_15786,N_16952);
and U24544 (N_24544,N_15186,N_14720);
nand U24545 (N_24545,N_17883,N_15329);
and U24546 (N_24546,N_14410,N_13355);
and U24547 (N_24547,N_14179,N_14524);
nor U24548 (N_24548,N_15447,N_16425);
nand U24549 (N_24549,N_14328,N_15492);
and U24550 (N_24550,N_12993,N_14225);
nor U24551 (N_24551,N_16638,N_14904);
and U24552 (N_24552,N_15156,N_18227);
nand U24553 (N_24553,N_18502,N_18399);
and U24554 (N_24554,N_14552,N_17339);
nand U24555 (N_24555,N_13278,N_18179);
nand U24556 (N_24556,N_13983,N_15001);
xnor U24557 (N_24557,N_16068,N_17712);
nor U24558 (N_24558,N_16680,N_17052);
xor U24559 (N_24559,N_16230,N_12679);
or U24560 (N_24560,N_14413,N_17377);
nand U24561 (N_24561,N_15120,N_17162);
and U24562 (N_24562,N_12672,N_14238);
or U24563 (N_24563,N_16850,N_15875);
xor U24564 (N_24564,N_15051,N_17461);
nor U24565 (N_24565,N_17609,N_18224);
or U24566 (N_24566,N_14863,N_15142);
or U24567 (N_24567,N_14415,N_17096);
nand U24568 (N_24568,N_13838,N_15397);
nor U24569 (N_24569,N_15458,N_15318);
and U24570 (N_24570,N_13635,N_16985);
and U24571 (N_24571,N_14322,N_17412);
nand U24572 (N_24572,N_12851,N_17031);
and U24573 (N_24573,N_17829,N_12976);
or U24574 (N_24574,N_16008,N_12510);
nor U24575 (N_24575,N_13982,N_13541);
nor U24576 (N_24576,N_18693,N_13105);
and U24577 (N_24577,N_18424,N_18051);
nor U24578 (N_24578,N_14962,N_15530);
nand U24579 (N_24579,N_15738,N_17310);
and U24580 (N_24580,N_16122,N_15607);
nor U24581 (N_24581,N_17818,N_16221);
nor U24582 (N_24582,N_16644,N_15023);
and U24583 (N_24583,N_14362,N_14905);
nand U24584 (N_24584,N_12761,N_16692);
nand U24585 (N_24585,N_15239,N_12647);
xor U24586 (N_24586,N_14018,N_16900);
nor U24587 (N_24587,N_17811,N_16927);
xor U24588 (N_24588,N_14493,N_18316);
nor U24589 (N_24589,N_15767,N_17396);
nor U24590 (N_24590,N_14359,N_17500);
and U24591 (N_24591,N_17466,N_12557);
xnor U24592 (N_24592,N_17972,N_15413);
nand U24593 (N_24593,N_17986,N_18664);
nor U24594 (N_24594,N_17479,N_14228);
or U24595 (N_24595,N_17236,N_12781);
nor U24596 (N_24596,N_12786,N_18451);
or U24597 (N_24597,N_16738,N_15893);
nor U24598 (N_24598,N_15569,N_14051);
or U24599 (N_24599,N_16153,N_18030);
nand U24600 (N_24600,N_18107,N_17663);
xor U24601 (N_24601,N_13521,N_16840);
or U24602 (N_24602,N_17788,N_17933);
nand U24603 (N_24603,N_15784,N_13893);
nor U24604 (N_24604,N_15041,N_18666);
and U24605 (N_24605,N_17007,N_16524);
or U24606 (N_24606,N_13474,N_13606);
or U24607 (N_24607,N_18476,N_18354);
nand U24608 (N_24608,N_13170,N_14739);
nor U24609 (N_24609,N_15204,N_13757);
or U24610 (N_24610,N_13261,N_13157);
and U24611 (N_24611,N_14487,N_13610);
xor U24612 (N_24612,N_13558,N_17598);
nor U24613 (N_24613,N_18454,N_17458);
nor U24614 (N_24614,N_14433,N_15360);
nor U24615 (N_24615,N_16938,N_13683);
nor U24616 (N_24616,N_13685,N_17118);
and U24617 (N_24617,N_18230,N_14211);
and U24618 (N_24618,N_16383,N_17436);
and U24619 (N_24619,N_16681,N_17080);
and U24620 (N_24620,N_14501,N_15144);
or U24621 (N_24621,N_13704,N_12952);
or U24622 (N_24622,N_16358,N_15481);
or U24623 (N_24623,N_13984,N_14500);
xnor U24624 (N_24624,N_18569,N_13462);
nor U24625 (N_24625,N_15937,N_17470);
or U24626 (N_24626,N_15088,N_12710);
and U24627 (N_24627,N_16156,N_16896);
xor U24628 (N_24628,N_14792,N_14261);
and U24629 (N_24629,N_14699,N_12735);
nand U24630 (N_24630,N_15898,N_15963);
or U24631 (N_24631,N_12601,N_14118);
xor U24632 (N_24632,N_14152,N_17569);
nor U24633 (N_24633,N_17713,N_14319);
nor U24634 (N_24634,N_16601,N_15610);
nand U24635 (N_24635,N_12818,N_13393);
and U24636 (N_24636,N_18695,N_12961);
nand U24637 (N_24637,N_13497,N_15141);
nor U24638 (N_24638,N_18100,N_13253);
nor U24639 (N_24639,N_18504,N_16078);
nor U24640 (N_24640,N_17030,N_16154);
and U24641 (N_24641,N_17878,N_16440);
or U24642 (N_24642,N_14491,N_18220);
xnor U24643 (N_24643,N_13395,N_16304);
or U24644 (N_24644,N_14677,N_13316);
and U24645 (N_24645,N_15178,N_14968);
nor U24646 (N_24646,N_12788,N_13799);
nand U24647 (N_24647,N_18697,N_16729);
nor U24648 (N_24648,N_17348,N_15041);
nor U24649 (N_24649,N_14766,N_17303);
nand U24650 (N_24650,N_13391,N_18155);
nand U24651 (N_24651,N_12857,N_13516);
and U24652 (N_24652,N_18096,N_18692);
and U24653 (N_24653,N_14747,N_14778);
and U24654 (N_24654,N_17021,N_17923);
nand U24655 (N_24655,N_17204,N_12839);
nand U24656 (N_24656,N_13280,N_13003);
and U24657 (N_24657,N_16243,N_15164);
nand U24658 (N_24658,N_17099,N_14309);
xnor U24659 (N_24659,N_14287,N_12524);
nor U24660 (N_24660,N_17685,N_16175);
nand U24661 (N_24661,N_12970,N_15456);
nor U24662 (N_24662,N_13042,N_18740);
nand U24663 (N_24663,N_18209,N_18060);
or U24664 (N_24664,N_14458,N_17575);
nor U24665 (N_24665,N_15383,N_15560);
nor U24666 (N_24666,N_18346,N_17556);
and U24667 (N_24667,N_18088,N_14915);
nor U24668 (N_24668,N_13597,N_15330);
or U24669 (N_24669,N_16611,N_15384);
nand U24670 (N_24670,N_15232,N_15490);
nand U24671 (N_24671,N_17091,N_15603);
xor U24672 (N_24672,N_13012,N_17979);
nand U24673 (N_24673,N_16399,N_12788);
xor U24674 (N_24674,N_17897,N_14890);
nand U24675 (N_24675,N_15035,N_13822);
and U24676 (N_24676,N_17214,N_14525);
and U24677 (N_24677,N_14067,N_14714);
or U24678 (N_24678,N_12512,N_15406);
and U24679 (N_24679,N_13922,N_13511);
and U24680 (N_24680,N_16887,N_16443);
nand U24681 (N_24681,N_15546,N_14535);
nor U24682 (N_24682,N_16403,N_16604);
or U24683 (N_24683,N_14832,N_14791);
nand U24684 (N_24684,N_13542,N_17751);
and U24685 (N_24685,N_17089,N_16877);
xor U24686 (N_24686,N_12949,N_18562);
and U24687 (N_24687,N_15856,N_14287);
nor U24688 (N_24688,N_16357,N_12798);
nand U24689 (N_24689,N_15293,N_14302);
and U24690 (N_24690,N_18358,N_12746);
nand U24691 (N_24691,N_15929,N_13266);
and U24692 (N_24692,N_15562,N_14981);
nor U24693 (N_24693,N_17170,N_16240);
or U24694 (N_24694,N_13144,N_15070);
or U24695 (N_24695,N_14206,N_13943);
or U24696 (N_24696,N_16812,N_16761);
or U24697 (N_24697,N_13145,N_16052);
nor U24698 (N_24698,N_15821,N_14109);
and U24699 (N_24699,N_14536,N_17999);
and U24700 (N_24700,N_16091,N_16020);
nor U24701 (N_24701,N_17762,N_17068);
nand U24702 (N_24702,N_13779,N_18479);
nand U24703 (N_24703,N_17588,N_17156);
nor U24704 (N_24704,N_16972,N_17786);
or U24705 (N_24705,N_14674,N_14775);
and U24706 (N_24706,N_17671,N_15930);
and U24707 (N_24707,N_16426,N_13895);
or U24708 (N_24708,N_18651,N_12699);
or U24709 (N_24709,N_13029,N_14964);
and U24710 (N_24710,N_17046,N_12858);
xnor U24711 (N_24711,N_13918,N_16313);
nor U24712 (N_24712,N_17637,N_18096);
or U24713 (N_24713,N_17350,N_15144);
nand U24714 (N_24714,N_14876,N_17301);
nor U24715 (N_24715,N_13218,N_16252);
nand U24716 (N_24716,N_15572,N_13310);
or U24717 (N_24717,N_13298,N_18345);
nand U24718 (N_24718,N_15286,N_14394);
or U24719 (N_24719,N_18564,N_17977);
and U24720 (N_24720,N_17880,N_15157);
or U24721 (N_24721,N_15948,N_15236);
nor U24722 (N_24722,N_16574,N_15391);
nand U24723 (N_24723,N_18094,N_17408);
nor U24724 (N_24724,N_17371,N_16623);
and U24725 (N_24725,N_16485,N_16770);
or U24726 (N_24726,N_17951,N_13048);
and U24727 (N_24727,N_16880,N_14286);
and U24728 (N_24728,N_15327,N_16652);
or U24729 (N_24729,N_17806,N_16209);
nand U24730 (N_24730,N_14420,N_15976);
nor U24731 (N_24731,N_14269,N_14516);
or U24732 (N_24732,N_14878,N_15011);
nand U24733 (N_24733,N_14341,N_17027);
and U24734 (N_24734,N_15269,N_12607);
or U24735 (N_24735,N_14519,N_14239);
or U24736 (N_24736,N_17692,N_15135);
and U24737 (N_24737,N_15080,N_16510);
and U24738 (N_24738,N_17272,N_13914);
and U24739 (N_24739,N_17777,N_18440);
nand U24740 (N_24740,N_13320,N_13240);
or U24741 (N_24741,N_16442,N_16535);
nor U24742 (N_24742,N_12848,N_14295);
nor U24743 (N_24743,N_15835,N_16264);
nand U24744 (N_24744,N_13291,N_16757);
and U24745 (N_24745,N_15980,N_14983);
or U24746 (N_24746,N_18042,N_14039);
nand U24747 (N_24747,N_15312,N_16855);
and U24748 (N_24748,N_18228,N_18653);
and U24749 (N_24749,N_18737,N_17095);
nand U24750 (N_24750,N_18000,N_16037);
nor U24751 (N_24751,N_15584,N_17669);
nand U24752 (N_24752,N_17387,N_17749);
nor U24753 (N_24753,N_13264,N_16106);
nor U24754 (N_24754,N_12766,N_17172);
nand U24755 (N_24755,N_16664,N_15289);
nor U24756 (N_24756,N_17605,N_17468);
nand U24757 (N_24757,N_14625,N_18404);
xnor U24758 (N_24758,N_13314,N_17533);
and U24759 (N_24759,N_13431,N_14370);
nand U24760 (N_24760,N_18430,N_15526);
and U24761 (N_24761,N_15102,N_13092);
nor U24762 (N_24762,N_17939,N_18426);
or U24763 (N_24763,N_17640,N_15384);
and U24764 (N_24764,N_17924,N_14116);
nor U24765 (N_24765,N_18057,N_17681);
nand U24766 (N_24766,N_14314,N_14290);
nor U24767 (N_24767,N_14074,N_16167);
nand U24768 (N_24768,N_18661,N_16738);
nor U24769 (N_24769,N_18431,N_14963);
nand U24770 (N_24770,N_14477,N_15406);
nand U24771 (N_24771,N_13750,N_15119);
and U24772 (N_24772,N_15650,N_16936);
or U24773 (N_24773,N_13099,N_14878);
nor U24774 (N_24774,N_14623,N_13287);
and U24775 (N_24775,N_15374,N_17428);
and U24776 (N_24776,N_17728,N_15830);
xnor U24777 (N_24777,N_17334,N_14593);
or U24778 (N_24778,N_15561,N_13263);
nor U24779 (N_24779,N_18738,N_17328);
nor U24780 (N_24780,N_12771,N_15172);
and U24781 (N_24781,N_16309,N_13501);
nor U24782 (N_24782,N_13430,N_13166);
and U24783 (N_24783,N_17694,N_12755);
and U24784 (N_24784,N_16691,N_15899);
nand U24785 (N_24785,N_15015,N_14885);
and U24786 (N_24786,N_13428,N_13377);
nand U24787 (N_24787,N_16918,N_16340);
nor U24788 (N_24788,N_15169,N_13615);
or U24789 (N_24789,N_15780,N_12922);
nor U24790 (N_24790,N_15709,N_17834);
xnor U24791 (N_24791,N_17418,N_18466);
and U24792 (N_24792,N_15750,N_18348);
and U24793 (N_24793,N_14259,N_14250);
nor U24794 (N_24794,N_15340,N_12659);
and U24795 (N_24795,N_12849,N_16334);
and U24796 (N_24796,N_12838,N_17132);
and U24797 (N_24797,N_12858,N_12988);
and U24798 (N_24798,N_18232,N_15026);
or U24799 (N_24799,N_17204,N_18656);
or U24800 (N_24800,N_14414,N_15197);
nand U24801 (N_24801,N_13928,N_15253);
nor U24802 (N_24802,N_15902,N_17629);
nand U24803 (N_24803,N_14416,N_14496);
nor U24804 (N_24804,N_14996,N_13043);
and U24805 (N_24805,N_18474,N_18082);
nand U24806 (N_24806,N_12765,N_14942);
nor U24807 (N_24807,N_18073,N_12702);
and U24808 (N_24808,N_14488,N_15392);
or U24809 (N_24809,N_17095,N_18685);
nor U24810 (N_24810,N_14625,N_18527);
and U24811 (N_24811,N_18133,N_15700);
xnor U24812 (N_24812,N_12587,N_14471);
nor U24813 (N_24813,N_14071,N_16682);
nand U24814 (N_24814,N_13705,N_17282);
nand U24815 (N_24815,N_16428,N_16546);
and U24816 (N_24816,N_17171,N_12740);
nor U24817 (N_24817,N_16224,N_14590);
nor U24818 (N_24818,N_12536,N_16953);
nand U24819 (N_24819,N_18304,N_15489);
and U24820 (N_24820,N_14128,N_17608);
nor U24821 (N_24821,N_17720,N_12760);
or U24822 (N_24822,N_18423,N_14622);
nor U24823 (N_24823,N_18560,N_13724);
and U24824 (N_24824,N_13075,N_14953);
nor U24825 (N_24825,N_13236,N_17423);
or U24826 (N_24826,N_16391,N_18717);
nor U24827 (N_24827,N_14077,N_15078);
nor U24828 (N_24828,N_16545,N_12594);
nor U24829 (N_24829,N_15262,N_13229);
nand U24830 (N_24830,N_16817,N_18414);
xnor U24831 (N_24831,N_12792,N_13474);
nand U24832 (N_24832,N_13143,N_15852);
xnor U24833 (N_24833,N_12585,N_16020);
xnor U24834 (N_24834,N_17884,N_15153);
nand U24835 (N_24835,N_18229,N_18423);
or U24836 (N_24836,N_14336,N_14978);
or U24837 (N_24837,N_18703,N_14453);
and U24838 (N_24838,N_13504,N_17115);
and U24839 (N_24839,N_13014,N_15692);
or U24840 (N_24840,N_14441,N_16145);
and U24841 (N_24841,N_12812,N_12717);
and U24842 (N_24842,N_17454,N_12788);
xor U24843 (N_24843,N_17378,N_17450);
nand U24844 (N_24844,N_15866,N_15307);
or U24845 (N_24845,N_15343,N_16218);
nor U24846 (N_24846,N_15652,N_16692);
nand U24847 (N_24847,N_14029,N_18732);
nand U24848 (N_24848,N_16236,N_16927);
and U24849 (N_24849,N_16172,N_17150);
nand U24850 (N_24850,N_16146,N_16377);
or U24851 (N_24851,N_14539,N_15094);
nand U24852 (N_24852,N_16710,N_13646);
and U24853 (N_24853,N_12706,N_14505);
nand U24854 (N_24854,N_18656,N_17574);
and U24855 (N_24855,N_13645,N_15311);
nor U24856 (N_24856,N_14236,N_17224);
and U24857 (N_24857,N_15305,N_16532);
nand U24858 (N_24858,N_13812,N_17837);
xnor U24859 (N_24859,N_16514,N_16573);
nor U24860 (N_24860,N_15197,N_12929);
nor U24861 (N_24861,N_17465,N_14242);
nand U24862 (N_24862,N_16284,N_18535);
nor U24863 (N_24863,N_12532,N_12817);
or U24864 (N_24864,N_18646,N_12729);
or U24865 (N_24865,N_15920,N_13495);
or U24866 (N_24866,N_14312,N_15584);
or U24867 (N_24867,N_18409,N_16880);
nor U24868 (N_24868,N_14263,N_12603);
nand U24869 (N_24869,N_15456,N_18346);
or U24870 (N_24870,N_14030,N_17144);
nand U24871 (N_24871,N_13517,N_17017);
and U24872 (N_24872,N_17093,N_13759);
nand U24873 (N_24873,N_18251,N_13893);
and U24874 (N_24874,N_15243,N_17432);
xor U24875 (N_24875,N_16087,N_15947);
nand U24876 (N_24876,N_13191,N_17986);
or U24877 (N_24877,N_17892,N_12851);
nor U24878 (N_24878,N_14615,N_13834);
and U24879 (N_24879,N_17434,N_13609);
nand U24880 (N_24880,N_17097,N_18246);
or U24881 (N_24881,N_14616,N_15442);
or U24882 (N_24882,N_15056,N_15121);
or U24883 (N_24883,N_13176,N_17330);
xor U24884 (N_24884,N_13060,N_17684);
and U24885 (N_24885,N_16047,N_14944);
nand U24886 (N_24886,N_14869,N_17010);
nor U24887 (N_24887,N_16388,N_18670);
nor U24888 (N_24888,N_13442,N_17712);
and U24889 (N_24889,N_16138,N_17838);
xor U24890 (N_24890,N_18063,N_18078);
nor U24891 (N_24891,N_13955,N_13395);
nor U24892 (N_24892,N_18566,N_15943);
and U24893 (N_24893,N_14643,N_16583);
xor U24894 (N_24894,N_17305,N_18056);
nand U24895 (N_24895,N_15687,N_18664);
nor U24896 (N_24896,N_18188,N_17983);
nand U24897 (N_24897,N_15998,N_17578);
or U24898 (N_24898,N_17736,N_14990);
and U24899 (N_24899,N_16572,N_13250);
nor U24900 (N_24900,N_16587,N_17869);
nor U24901 (N_24901,N_17285,N_16795);
or U24902 (N_24902,N_17894,N_16684);
xor U24903 (N_24903,N_14461,N_14130);
nand U24904 (N_24904,N_16670,N_14073);
or U24905 (N_24905,N_18293,N_18400);
nand U24906 (N_24906,N_15599,N_17461);
nor U24907 (N_24907,N_17592,N_14373);
xnor U24908 (N_24908,N_16589,N_14212);
and U24909 (N_24909,N_18265,N_15257);
or U24910 (N_24910,N_17767,N_18287);
and U24911 (N_24911,N_15552,N_14797);
nor U24912 (N_24912,N_15149,N_17725);
or U24913 (N_24913,N_17200,N_12557);
nor U24914 (N_24914,N_15295,N_16382);
or U24915 (N_24915,N_18096,N_17876);
xor U24916 (N_24916,N_15768,N_17660);
nand U24917 (N_24917,N_16100,N_13414);
nand U24918 (N_24918,N_15977,N_15853);
xor U24919 (N_24919,N_16146,N_16326);
or U24920 (N_24920,N_15025,N_13365);
nor U24921 (N_24921,N_12931,N_14902);
or U24922 (N_24922,N_17865,N_14121);
nor U24923 (N_24923,N_12747,N_15549);
and U24924 (N_24924,N_16635,N_15698);
and U24925 (N_24925,N_17663,N_13371);
or U24926 (N_24926,N_13357,N_14161);
and U24927 (N_24927,N_15462,N_13306);
and U24928 (N_24928,N_17157,N_14777);
and U24929 (N_24929,N_13723,N_13782);
nor U24930 (N_24930,N_13718,N_14787);
and U24931 (N_24931,N_14077,N_12533);
and U24932 (N_24932,N_17786,N_16640);
and U24933 (N_24933,N_12892,N_17843);
and U24934 (N_24934,N_12985,N_17933);
or U24935 (N_24935,N_18377,N_15680);
nor U24936 (N_24936,N_14835,N_17953);
and U24937 (N_24937,N_16169,N_14528);
or U24938 (N_24938,N_12621,N_14426);
nand U24939 (N_24939,N_15080,N_15610);
and U24940 (N_24940,N_13854,N_15967);
xor U24941 (N_24941,N_15150,N_17782);
or U24942 (N_24942,N_16094,N_15981);
xor U24943 (N_24943,N_16231,N_13768);
or U24944 (N_24944,N_18470,N_14742);
and U24945 (N_24945,N_15159,N_18074);
nand U24946 (N_24946,N_16619,N_15123);
nor U24947 (N_24947,N_15182,N_12641);
xnor U24948 (N_24948,N_14989,N_16308);
nand U24949 (N_24949,N_14034,N_17271);
and U24950 (N_24950,N_14112,N_18129);
nand U24951 (N_24951,N_17445,N_14542);
nor U24952 (N_24952,N_14261,N_18490);
xnor U24953 (N_24953,N_12609,N_15245);
and U24954 (N_24954,N_16988,N_16059);
nor U24955 (N_24955,N_14934,N_14792);
and U24956 (N_24956,N_17135,N_17643);
nand U24957 (N_24957,N_16270,N_14059);
nand U24958 (N_24958,N_16026,N_15338);
and U24959 (N_24959,N_16396,N_14200);
nor U24960 (N_24960,N_12978,N_13680);
nand U24961 (N_24961,N_17102,N_12583);
nor U24962 (N_24962,N_14466,N_16423);
nand U24963 (N_24963,N_12985,N_14275);
and U24964 (N_24964,N_18447,N_17943);
or U24965 (N_24965,N_14183,N_14644);
or U24966 (N_24966,N_17303,N_17892);
nand U24967 (N_24967,N_16396,N_13783);
or U24968 (N_24968,N_17165,N_15458);
and U24969 (N_24969,N_16100,N_17522);
and U24970 (N_24970,N_15732,N_15729);
xor U24971 (N_24971,N_13360,N_13993);
xnor U24972 (N_24972,N_14969,N_16656);
and U24973 (N_24973,N_13281,N_13216);
or U24974 (N_24974,N_16196,N_13709);
and U24975 (N_24975,N_13022,N_13066);
xnor U24976 (N_24976,N_13885,N_15000);
nor U24977 (N_24977,N_12974,N_15141);
nor U24978 (N_24978,N_14543,N_14211);
nand U24979 (N_24979,N_17788,N_13120);
nor U24980 (N_24980,N_14367,N_15190);
and U24981 (N_24981,N_14319,N_14823);
nand U24982 (N_24982,N_15578,N_16429);
xor U24983 (N_24983,N_16763,N_16422);
nor U24984 (N_24984,N_16598,N_17419);
or U24985 (N_24985,N_18026,N_15152);
nor U24986 (N_24986,N_17009,N_14731);
xnor U24987 (N_24987,N_16170,N_14860);
nor U24988 (N_24988,N_18077,N_13018);
and U24989 (N_24989,N_12802,N_15996);
nand U24990 (N_24990,N_18478,N_15157);
nor U24991 (N_24991,N_18572,N_15034);
and U24992 (N_24992,N_16890,N_12735);
xnor U24993 (N_24993,N_16963,N_13073);
nor U24994 (N_24994,N_17643,N_14656);
xor U24995 (N_24995,N_15598,N_17518);
and U24996 (N_24996,N_15876,N_12991);
xor U24997 (N_24997,N_12973,N_16696);
nand U24998 (N_24998,N_15253,N_15286);
or U24999 (N_24999,N_14255,N_16487);
nor UO_0 (O_0,N_20039,N_20624);
nand UO_1 (O_1,N_21230,N_22542);
and UO_2 (O_2,N_22281,N_22128);
nor UO_3 (O_3,N_20816,N_23880);
and UO_4 (O_4,N_20857,N_19336);
or UO_5 (O_5,N_22697,N_23043);
nor UO_6 (O_6,N_21258,N_23537);
and UO_7 (O_7,N_24628,N_24946);
nand UO_8 (O_8,N_18962,N_23538);
or UO_9 (O_9,N_21266,N_20671);
xnor UO_10 (O_10,N_20078,N_23777);
or UO_11 (O_11,N_19265,N_19206);
nor UO_12 (O_12,N_19883,N_23574);
nor UO_13 (O_13,N_19074,N_18988);
xnor UO_14 (O_14,N_23263,N_18788);
or UO_15 (O_15,N_23396,N_22563);
or UO_16 (O_16,N_21440,N_20855);
or UO_17 (O_17,N_22097,N_24937);
or UO_18 (O_18,N_24940,N_24246);
or UO_19 (O_19,N_21574,N_23959);
nor UO_20 (O_20,N_24724,N_22915);
and UO_21 (O_21,N_23367,N_19506);
and UO_22 (O_22,N_19992,N_22182);
nand UO_23 (O_23,N_24179,N_19886);
or UO_24 (O_24,N_23774,N_21813);
nor UO_25 (O_25,N_23868,N_19570);
nor UO_26 (O_26,N_22522,N_22176);
nor UO_27 (O_27,N_19953,N_24368);
or UO_28 (O_28,N_20151,N_21035);
xnor UO_29 (O_29,N_23531,N_21822);
nor UO_30 (O_30,N_18886,N_22352);
or UO_31 (O_31,N_21107,N_20248);
and UO_32 (O_32,N_21277,N_23147);
nor UO_33 (O_33,N_19306,N_19798);
and UO_34 (O_34,N_22939,N_20715);
or UO_35 (O_35,N_23495,N_21537);
or UO_36 (O_36,N_22952,N_20993);
or UO_37 (O_37,N_20174,N_24473);
and UO_38 (O_38,N_21158,N_23181);
nand UO_39 (O_39,N_22526,N_19926);
nand UO_40 (O_40,N_23055,N_23818);
nor UO_41 (O_41,N_20745,N_20055);
nor UO_42 (O_42,N_23625,N_22641);
nor UO_43 (O_43,N_20010,N_22459);
or UO_44 (O_44,N_23614,N_24359);
nor UO_45 (O_45,N_24977,N_21009);
nor UO_46 (O_46,N_20867,N_21522);
nand UO_47 (O_47,N_19865,N_20167);
and UO_48 (O_48,N_22519,N_20599);
and UO_49 (O_49,N_19572,N_21951);
xnor UO_50 (O_50,N_22359,N_24003);
or UO_51 (O_51,N_18890,N_19157);
nand UO_52 (O_52,N_22096,N_18923);
nor UO_53 (O_53,N_22370,N_20142);
and UO_54 (O_54,N_20277,N_19346);
nor UO_55 (O_55,N_24458,N_20061);
nor UO_56 (O_56,N_23566,N_22560);
nor UO_57 (O_57,N_22077,N_23720);
or UO_58 (O_58,N_23634,N_23655);
and UO_59 (O_59,N_22203,N_21501);
nand UO_60 (O_60,N_23394,N_23028);
xor UO_61 (O_61,N_20721,N_20552);
nand UO_62 (O_62,N_24611,N_24395);
nand UO_63 (O_63,N_19780,N_19793);
xnor UO_64 (O_64,N_20642,N_19555);
nand UO_65 (O_65,N_21379,N_18853);
xor UO_66 (O_66,N_20355,N_21106);
or UO_67 (O_67,N_20408,N_21469);
xor UO_68 (O_68,N_22187,N_20196);
nor UO_69 (O_69,N_24440,N_23782);
nor UO_70 (O_70,N_21183,N_24386);
or UO_71 (O_71,N_23129,N_19356);
xor UO_72 (O_72,N_19522,N_19921);
xor UO_73 (O_73,N_21449,N_20481);
or UO_74 (O_74,N_20881,N_23350);
nand UO_75 (O_75,N_22590,N_23685);
nand UO_76 (O_76,N_24963,N_22103);
and UO_77 (O_77,N_23800,N_20116);
nand UO_78 (O_78,N_24270,N_22523);
nand UO_79 (O_79,N_20237,N_22801);
and UO_80 (O_80,N_23528,N_20361);
nor UO_81 (O_81,N_22511,N_20211);
and UO_82 (O_82,N_22461,N_24064);
nor UO_83 (O_83,N_21546,N_21356);
or UO_84 (O_84,N_21204,N_20949);
xnor UO_85 (O_85,N_24139,N_22981);
and UO_86 (O_86,N_21502,N_20690);
nand UO_87 (O_87,N_20755,N_19267);
xnor UO_88 (O_88,N_20156,N_19408);
nor UO_89 (O_89,N_21066,N_24303);
and UO_90 (O_90,N_21394,N_24055);
nand UO_91 (O_91,N_21519,N_24991);
or UO_92 (O_92,N_24466,N_19456);
nand UO_93 (O_93,N_22098,N_19355);
nand UO_94 (O_94,N_21135,N_23796);
nand UO_95 (O_95,N_19095,N_19612);
nor UO_96 (O_96,N_21834,N_22914);
nor UO_97 (O_97,N_20178,N_22022);
xnor UO_98 (O_98,N_22917,N_19537);
nand UO_99 (O_99,N_18781,N_23109);
nand UO_100 (O_100,N_22372,N_19811);
and UO_101 (O_101,N_18939,N_23308);
nor UO_102 (O_102,N_24435,N_24239);
nand UO_103 (O_103,N_19937,N_22159);
and UO_104 (O_104,N_24413,N_24105);
xnor UO_105 (O_105,N_23451,N_21268);
nand UO_106 (O_106,N_22169,N_21542);
nor UO_107 (O_107,N_20127,N_23389);
nand UO_108 (O_108,N_24966,N_24643);
or UO_109 (O_109,N_20776,N_24698);
and UO_110 (O_110,N_24360,N_24416);
nand UO_111 (O_111,N_19340,N_19017);
xnor UO_112 (O_112,N_22266,N_21599);
nand UO_113 (O_113,N_21410,N_19731);
nand UO_114 (O_114,N_20475,N_23914);
nor UO_115 (O_115,N_24528,N_22823);
nand UO_116 (O_116,N_24975,N_22439);
nor UO_117 (O_117,N_19814,N_23596);
and UO_118 (O_118,N_21857,N_19762);
nand UO_119 (O_119,N_22789,N_18915);
and UO_120 (O_120,N_20807,N_21903);
or UO_121 (O_121,N_23667,N_19078);
or UO_122 (O_122,N_23524,N_22013);
and UO_123 (O_123,N_22601,N_19342);
and UO_124 (O_124,N_22113,N_19149);
nor UO_125 (O_125,N_19884,N_19256);
nor UO_126 (O_126,N_24747,N_19740);
xor UO_127 (O_127,N_19042,N_22210);
and UO_128 (O_128,N_24625,N_20732);
nor UO_129 (O_129,N_24207,N_23086);
and UO_130 (O_130,N_19171,N_22615);
and UO_131 (O_131,N_22771,N_20346);
or UO_132 (O_132,N_23038,N_22111);
or UO_133 (O_133,N_23465,N_20786);
and UO_134 (O_134,N_22313,N_20068);
and UO_135 (O_135,N_23187,N_24681);
or UO_136 (O_136,N_23155,N_19044);
nand UO_137 (O_137,N_21797,N_19386);
nand UO_138 (O_138,N_23455,N_19751);
nor UO_139 (O_139,N_22496,N_24186);
nor UO_140 (O_140,N_22390,N_21874);
nor UO_141 (O_141,N_23330,N_21417);
nor UO_142 (O_142,N_19877,N_21886);
and UO_143 (O_143,N_20468,N_19376);
or UO_144 (O_144,N_21563,N_23069);
nand UO_145 (O_145,N_19505,N_21400);
nand UO_146 (O_146,N_23602,N_20158);
and UO_147 (O_147,N_19908,N_21307);
nor UO_148 (O_148,N_21705,N_22742);
and UO_149 (O_149,N_22277,N_20222);
and UO_150 (O_150,N_23553,N_20806);
and UO_151 (O_151,N_21012,N_19410);
nor UO_152 (O_152,N_24608,N_24477);
xor UO_153 (O_153,N_20903,N_24581);
xnor UO_154 (O_154,N_22260,N_23152);
or UO_155 (O_155,N_20144,N_19518);
nor UO_156 (O_156,N_24140,N_21901);
and UO_157 (O_157,N_19727,N_24768);
nor UO_158 (O_158,N_20549,N_22451);
xor UO_159 (O_159,N_20630,N_22885);
and UO_160 (O_160,N_22125,N_24565);
nand UO_161 (O_161,N_19321,N_21128);
and UO_162 (O_162,N_24505,N_22320);
and UO_163 (O_163,N_21531,N_24956);
nand UO_164 (O_164,N_20841,N_23987);
or UO_165 (O_165,N_23754,N_21856);
nand UO_166 (O_166,N_21240,N_19175);
or UO_167 (O_167,N_23933,N_20575);
nand UO_168 (O_168,N_24805,N_19805);
and UO_169 (O_169,N_22990,N_21638);
nor UO_170 (O_170,N_23710,N_20956);
nand UO_171 (O_171,N_20843,N_24155);
nand UO_172 (O_172,N_19797,N_24892);
nor UO_173 (O_173,N_24065,N_24312);
or UO_174 (O_174,N_20305,N_24124);
nor UO_175 (O_175,N_19493,N_23965);
and UO_176 (O_176,N_19899,N_20467);
nor UO_177 (O_177,N_21124,N_24832);
and UO_178 (O_178,N_19446,N_21138);
nand UO_179 (O_179,N_22814,N_21500);
or UO_180 (O_180,N_22014,N_21166);
nand UO_181 (O_181,N_24936,N_24717);
xnor UO_182 (O_182,N_18889,N_18864);
nand UO_183 (O_183,N_19985,N_24542);
nand UO_184 (O_184,N_20938,N_23049);
xor UO_185 (O_185,N_18812,N_21585);
or UO_186 (O_186,N_23581,N_20594);
nand UO_187 (O_187,N_20496,N_18960);
nor UO_188 (O_188,N_22855,N_23841);
and UO_189 (O_189,N_20273,N_19394);
nor UO_190 (O_190,N_22513,N_22397);
nor UO_191 (O_191,N_22751,N_19070);
nor UO_192 (O_192,N_19402,N_19212);
or UO_193 (O_193,N_19671,N_20518);
nand UO_194 (O_194,N_21717,N_19794);
nor UO_195 (O_195,N_22890,N_24405);
nand UO_196 (O_196,N_21391,N_21809);
nor UO_197 (O_197,N_22265,N_24471);
nand UO_198 (O_198,N_23241,N_22919);
xor UO_199 (O_199,N_20676,N_20922);
xnor UO_200 (O_200,N_20455,N_22579);
or UO_201 (O_201,N_19893,N_21071);
nor UO_202 (O_202,N_24159,N_19289);
and UO_203 (O_203,N_22688,N_22254);
and UO_204 (O_204,N_24373,N_24476);
and UO_205 (O_205,N_21283,N_20527);
xnor UO_206 (O_206,N_18973,N_19163);
and UO_207 (O_207,N_24070,N_22105);
and UO_208 (O_208,N_21781,N_21595);
nor UO_209 (O_209,N_19576,N_20201);
and UO_210 (O_210,N_23355,N_23989);
nor UO_211 (O_211,N_24446,N_23003);
or UO_212 (O_212,N_19434,N_22351);
nand UO_213 (O_213,N_20637,N_20299);
nand UO_214 (O_214,N_21582,N_21249);
nor UO_215 (O_215,N_23768,N_22487);
nand UO_216 (O_216,N_22104,N_21475);
nand UO_217 (O_217,N_23924,N_18855);
or UO_218 (O_218,N_22668,N_24729);
nor UO_219 (O_219,N_24875,N_20413);
nor UO_220 (O_220,N_24927,N_19511);
nor UO_221 (O_221,N_19809,N_24015);
or UO_222 (O_222,N_19416,N_24109);
nor UO_223 (O_223,N_22786,N_22179);
or UO_224 (O_224,N_20685,N_21487);
nor UO_225 (O_225,N_21403,N_20325);
nand UO_226 (O_226,N_21498,N_20308);
or UO_227 (O_227,N_20450,N_22471);
or UO_228 (O_228,N_22674,N_22813);
or UO_229 (O_229,N_22494,N_22779);
and UO_230 (O_230,N_21215,N_20348);
nand UO_231 (O_231,N_21934,N_23936);
and UO_232 (O_232,N_24419,N_22854);
and UO_233 (O_233,N_23556,N_19297);
nor UO_234 (O_234,N_19427,N_24042);
nand UO_235 (O_235,N_21507,N_24853);
nand UO_236 (O_236,N_19023,N_21991);
xnor UO_237 (O_237,N_21312,N_22879);
xor UO_238 (O_238,N_23213,N_19140);
nor UO_239 (O_239,N_20820,N_20953);
nor UO_240 (O_240,N_20388,N_21444);
nor UO_241 (O_241,N_22395,N_24796);
nor UO_242 (O_242,N_22761,N_21182);
and UO_243 (O_243,N_23864,N_24095);
xor UO_244 (O_244,N_21114,N_23638);
or UO_245 (O_245,N_20684,N_24817);
nand UO_246 (O_246,N_24409,N_21656);
nand UO_247 (O_247,N_23877,N_20853);
nor UO_248 (O_248,N_20316,N_24089);
and UO_249 (O_249,N_19514,N_18909);
nor UO_250 (O_250,N_24241,N_21769);
or UO_251 (O_251,N_22754,N_22886);
nand UO_252 (O_252,N_23885,N_20957);
or UO_253 (O_253,N_20653,N_18885);
or UO_254 (O_254,N_24320,N_18769);
xnor UO_255 (O_255,N_22241,N_19106);
nor UO_256 (O_256,N_23324,N_22566);
nor UO_257 (O_257,N_23184,N_23470);
or UO_258 (O_258,N_23658,N_24700);
xnor UO_259 (O_259,N_20389,N_21662);
nor UO_260 (O_260,N_19471,N_19792);
nor UO_261 (O_261,N_22706,N_19349);
xor UO_262 (O_262,N_19222,N_20788);
or UO_263 (O_263,N_23024,N_20851);
or UO_264 (O_264,N_24561,N_23557);
and UO_265 (O_265,N_24526,N_19967);
or UO_266 (O_266,N_18869,N_21105);
and UO_267 (O_267,N_23466,N_20161);
nand UO_268 (O_268,N_19347,N_22454);
nor UO_269 (O_269,N_21959,N_24499);
and UO_270 (O_270,N_22605,N_20424);
nor UO_271 (O_271,N_19606,N_21055);
and UO_272 (O_272,N_22979,N_20138);
nand UO_273 (O_273,N_18767,N_20882);
and UO_274 (O_274,N_18773,N_20125);
and UO_275 (O_275,N_19320,N_20106);
nand UO_276 (O_276,N_18893,N_20535);
nor UO_277 (O_277,N_22377,N_21784);
and UO_278 (O_278,N_19642,N_19103);
nand UO_279 (O_279,N_19257,N_20281);
nand UO_280 (O_280,N_22108,N_21751);
and UO_281 (O_281,N_22787,N_21227);
or UO_282 (O_282,N_20283,N_18850);
or UO_283 (O_283,N_19414,N_19770);
nand UO_284 (O_284,N_20326,N_21434);
and UO_285 (O_285,N_19359,N_24890);
nand UO_286 (O_286,N_18816,N_18813);
nor UO_287 (O_287,N_24230,N_23781);
or UO_288 (O_288,N_23127,N_21146);
and UO_289 (O_289,N_24792,N_23714);
and UO_290 (O_290,N_20360,N_19463);
and UO_291 (O_291,N_21297,N_22198);
or UO_292 (O_292,N_23812,N_19835);
or UO_293 (O_293,N_20626,N_22122);
or UO_294 (O_294,N_23518,N_24712);
and UO_295 (O_295,N_24813,N_19228);
nand UO_296 (O_296,N_20708,N_20207);
nand UO_297 (O_297,N_21641,N_22725);
nand UO_298 (O_298,N_19812,N_19861);
nand UO_299 (O_299,N_22472,N_22527);
nor UO_300 (O_300,N_23401,N_20371);
nand UO_301 (O_301,N_24380,N_22410);
nand UO_302 (O_302,N_20908,N_21879);
xnor UO_303 (O_303,N_21059,N_23104);
or UO_304 (O_304,N_22201,N_22388);
nand UO_305 (O_305,N_20534,N_20625);
xor UO_306 (O_306,N_21827,N_18825);
and UO_307 (O_307,N_22246,N_22693);
and UO_308 (O_308,N_19079,N_18881);
nand UO_309 (O_309,N_24928,N_18846);
nand UO_310 (O_310,N_24461,N_19482);
and UO_311 (O_311,N_19684,N_22287);
or UO_312 (O_312,N_22790,N_23122);
or UO_313 (O_313,N_19191,N_21718);
nand UO_314 (O_314,N_24949,N_20289);
nand UO_315 (O_315,N_21042,N_24020);
xor UO_316 (O_316,N_22655,N_22047);
and UO_317 (O_317,N_22596,N_22404);
xnor UO_318 (O_318,N_18873,N_23066);
and UO_319 (O_319,N_20378,N_22799);
xnor UO_320 (O_320,N_22977,N_19341);
nand UO_321 (O_321,N_19557,N_24554);
nor UO_322 (O_322,N_24742,N_23650);
nand UO_323 (O_323,N_20069,N_19838);
nor UO_324 (O_324,N_21628,N_22131);
and UO_325 (O_325,N_22237,N_21317);
nor UO_326 (O_326,N_24512,N_23420);
nor UO_327 (O_327,N_22980,N_21908);
xnor UO_328 (O_328,N_19911,N_22962);
and UO_329 (O_329,N_22431,N_22045);
nand UO_330 (O_330,N_23772,N_20414);
nor UO_331 (O_331,N_21304,N_19343);
and UO_332 (O_332,N_22819,N_23487);
nor UO_333 (O_333,N_20543,N_22035);
or UO_334 (O_334,N_21488,N_20441);
nor UO_335 (O_335,N_24079,N_22647);
nor UO_336 (O_336,N_23858,N_19932);
and UO_337 (O_337,N_23371,N_20007);
nand UO_338 (O_338,N_21726,N_24904);
and UO_339 (O_339,N_20542,N_20996);
xor UO_340 (O_340,N_20410,N_21261);
or UO_341 (O_341,N_21402,N_20592);
or UO_342 (O_342,N_24997,N_24494);
or UO_343 (O_343,N_23364,N_20876);
xnor UO_344 (O_344,N_24663,N_24502);
or UO_345 (O_345,N_21068,N_19858);
or UO_346 (O_346,N_20253,N_22434);
nor UO_347 (O_347,N_22509,N_18984);
or UO_348 (O_348,N_18847,N_18768);
nand UO_349 (O_349,N_24986,N_21795);
xor UO_350 (O_350,N_20910,N_22611);
or UO_351 (O_351,N_19290,N_20815);
and UO_352 (O_352,N_22606,N_22099);
nor UO_353 (O_353,N_23597,N_20500);
nand UO_354 (O_354,N_24970,N_22012);
nand UO_355 (O_355,N_23787,N_22541);
nand UO_356 (O_356,N_19974,N_21333);
and UO_357 (O_357,N_22945,N_19739);
nor UO_358 (O_358,N_22669,N_21063);
and UO_359 (O_359,N_24343,N_19726);
nand UO_360 (O_360,N_20146,N_20048);
nand UO_361 (O_361,N_23173,N_22685);
xnor UO_362 (O_362,N_22091,N_23598);
nand UO_363 (O_363,N_24418,N_22336);
xor UO_364 (O_364,N_20317,N_20704);
nand UO_365 (O_365,N_21850,N_22161);
xor UO_366 (O_366,N_22084,N_18959);
or UO_367 (O_367,N_19126,N_20090);
or UO_368 (O_368,N_21573,N_22178);
and UO_369 (O_369,N_23141,N_20364);
nor UO_370 (O_370,N_22670,N_23399);
and UO_371 (O_371,N_23853,N_24745);
or UO_372 (O_372,N_20465,N_20327);
nor UO_373 (O_373,N_23376,N_18876);
nor UO_374 (O_374,N_21415,N_19357);
nor UO_375 (O_375,N_23418,N_21949);
and UO_376 (O_376,N_22763,N_20973);
nor UO_377 (O_377,N_23369,N_20803);
or UO_378 (O_378,N_22943,N_24046);
xnor UO_379 (O_379,N_22257,N_20310);
nor UO_380 (O_380,N_19277,N_21131);
nor UO_381 (O_381,N_24807,N_22735);
xnor UO_382 (O_382,N_23273,N_24880);
xor UO_383 (O_383,N_24519,N_21778);
nand UO_384 (O_384,N_23203,N_22941);
or UO_385 (O_385,N_19763,N_19657);
nor UO_386 (O_386,N_22803,N_19246);
nor UO_387 (O_387,N_22272,N_23228);
and UO_388 (O_388,N_21604,N_24921);
nor UO_389 (O_389,N_18823,N_21544);
xor UO_390 (O_390,N_23332,N_24788);
and UO_391 (O_391,N_20054,N_24075);
xnor UO_392 (O_392,N_24309,N_24690);
and UO_393 (O_393,N_23794,N_21979);
or UO_394 (O_394,N_19808,N_23652);
and UO_395 (O_395,N_22049,N_24901);
nand UO_396 (O_396,N_23622,N_23271);
or UO_397 (O_397,N_19235,N_21997);
and UO_398 (O_398,N_18833,N_20366);
nor UO_399 (O_399,N_21859,N_20674);
xor UO_400 (O_400,N_19348,N_24769);
and UO_401 (O_401,N_22074,N_23776);
xnor UO_402 (O_402,N_22329,N_23690);
nand UO_403 (O_403,N_19328,N_22518);
or UO_404 (O_404,N_21962,N_19821);
and UO_405 (O_405,N_24896,N_23629);
nor UO_406 (O_406,N_19011,N_21987);
nor UO_407 (O_407,N_23926,N_24014);
nand UO_408 (O_408,N_22645,N_18910);
and UO_409 (O_409,N_23696,N_23494);
nor UO_410 (O_410,N_19707,N_24456);
or UO_411 (O_411,N_22238,N_21301);
or UO_412 (O_412,N_22838,N_22374);
nor UO_413 (O_413,N_22559,N_19586);
nand UO_414 (O_414,N_23306,N_23039);
and UO_415 (O_415,N_22151,N_19239);
or UO_416 (O_416,N_21559,N_22398);
or UO_417 (O_417,N_24612,N_21075);
nand UO_418 (O_418,N_21933,N_20403);
xnor UO_419 (O_419,N_23456,N_22441);
and UO_420 (O_420,N_19645,N_21891);
or UO_421 (O_421,N_22212,N_21642);
nor UO_422 (O_422,N_23608,N_23969);
and UO_423 (O_423,N_23407,N_20350);
nor UO_424 (O_424,N_21939,N_20115);
or UO_425 (O_425,N_21036,N_22894);
and UO_426 (O_426,N_21973,N_21735);
nand UO_427 (O_427,N_24265,N_20062);
nor UO_428 (O_428,N_22139,N_23788);
and UO_429 (O_429,N_20379,N_18927);
or UO_430 (O_430,N_22224,N_21306);
nand UO_431 (O_431,N_21852,N_22333);
or UO_432 (O_432,N_19663,N_23115);
nand UO_433 (O_433,N_22759,N_19300);
and UO_434 (O_434,N_23105,N_19435);
and UO_435 (O_435,N_19991,N_22168);
nor UO_436 (O_436,N_21272,N_21525);
and UO_437 (O_437,N_22443,N_24961);
and UO_438 (O_438,N_19183,N_18888);
or UO_439 (O_439,N_22581,N_19715);
nand UO_440 (O_440,N_22102,N_19539);
and UO_441 (O_441,N_22913,N_22529);
xnor UO_442 (O_442,N_24423,N_20173);
and UO_443 (O_443,N_22063,N_21601);
or UO_444 (O_444,N_19528,N_23044);
and UO_445 (O_445,N_23511,N_23291);
nand UO_446 (O_446,N_20656,N_19847);
and UO_447 (O_447,N_22418,N_19851);
nand UO_448 (O_448,N_22248,N_21898);
nor UO_449 (O_449,N_21443,N_23693);
and UO_450 (O_450,N_24391,N_23870);
nand UO_451 (O_451,N_20618,N_22396);
and UO_452 (O_452,N_22192,N_24973);
nor UO_453 (O_453,N_19148,N_23680);
and UO_454 (O_454,N_19688,N_19479);
nand UO_455 (O_455,N_19081,N_18917);
nand UO_456 (O_456,N_23326,N_22259);
nand UO_457 (O_457,N_21341,N_20362);
and UO_458 (O_458,N_21149,N_23178);
nand UO_459 (O_459,N_22033,N_19029);
and UO_460 (O_460,N_23731,N_23210);
nor UO_461 (O_461,N_24190,N_18807);
xnor UO_462 (O_462,N_24527,N_18851);
or UO_463 (O_463,N_24731,N_24804);
and UO_464 (O_464,N_23911,N_19466);
xor UO_465 (O_465,N_19609,N_24669);
and UO_466 (O_466,N_21362,N_24686);
nor UO_467 (O_467,N_24059,N_19919);
nand UO_468 (O_468,N_23615,N_19056);
xnor UO_469 (O_469,N_20794,N_24259);
nand UO_470 (O_470,N_19238,N_19680);
nor UO_471 (O_471,N_24371,N_20569);
xnor UO_472 (O_472,N_22216,N_20503);
or UO_473 (O_473,N_20112,N_23252);
nor UO_474 (O_474,N_22640,N_21942);
nand UO_475 (O_475,N_19654,N_23527);
nor UO_476 (O_476,N_24291,N_23064);
nand UO_477 (O_477,N_19643,N_21494);
nor UO_478 (O_478,N_23771,N_19830);
and UO_479 (O_479,N_24776,N_18894);
nand UO_480 (O_480,N_21584,N_23994);
nand UO_481 (O_481,N_23033,N_20770);
nand UO_482 (O_482,N_20638,N_20890);
nand UO_483 (O_483,N_19020,N_20145);
or UO_484 (O_484,N_19536,N_21967);
nand UO_485 (O_485,N_23117,N_23599);
or UO_486 (O_486,N_22162,N_20886);
nand UO_487 (O_487,N_24665,N_22452);
and UO_488 (O_488,N_21422,N_20854);
nand UO_489 (O_489,N_22505,N_20221);
nand UO_490 (O_490,N_24737,N_20731);
xnor UO_491 (O_491,N_24100,N_18778);
or UO_492 (O_492,N_20714,N_23239);
and UO_493 (O_493,N_22951,N_20471);
nand UO_494 (O_494,N_23436,N_24363);
nand UO_495 (O_495,N_19634,N_19988);
nand UO_496 (O_496,N_23520,N_20064);
and UO_497 (O_497,N_21163,N_19871);
nand UO_498 (O_498,N_20336,N_24389);
nand UO_499 (O_499,N_18872,N_22691);
nand UO_500 (O_500,N_24825,N_19362);
nand UO_501 (O_501,N_22678,N_21296);
xor UO_502 (O_502,N_20148,N_23499);
nand UO_503 (O_503,N_20784,N_22833);
nand UO_504 (O_504,N_20452,N_20734);
nor UO_505 (O_505,N_19240,N_21424);
or UO_506 (O_506,N_22409,N_24680);
nand UO_507 (O_507,N_21080,N_24049);
or UO_508 (O_508,N_21041,N_21586);
nor UO_509 (O_509,N_21274,N_23095);
and UO_510 (O_510,N_19443,N_23819);
and UO_511 (O_511,N_23515,N_24097);
or UO_512 (O_512,N_24585,N_22358);
and UO_513 (O_513,N_24604,N_20801);
nor UO_514 (O_514,N_22068,N_24688);
xnor UO_515 (O_515,N_21216,N_19702);
nor UO_516 (O_516,N_23218,N_19025);
xor UO_517 (O_517,N_22317,N_24277);
and UO_518 (O_518,N_23684,N_22448);
and UO_519 (O_519,N_22969,N_23387);
nor UO_520 (O_520,N_22467,N_18845);
nand UO_521 (O_521,N_22304,N_22144);
nand UO_522 (O_522,N_22873,N_19326);
and UO_523 (O_523,N_24062,N_24287);
nand UO_524 (O_524,N_19111,N_22734);
nor UO_525 (O_525,N_20774,N_22954);
or UO_526 (O_526,N_23521,N_23755);
nand UO_527 (O_527,N_20466,N_24842);
nor UO_528 (O_528,N_24091,N_19819);
and UO_529 (O_529,N_23360,N_20216);
nor UO_530 (O_530,N_20143,N_22389);
or UO_531 (O_531,N_22984,N_19141);
nand UO_532 (O_532,N_19521,N_22090);
and UO_533 (O_533,N_22484,N_20826);
nor UO_534 (O_534,N_21129,N_19108);
nor UO_535 (O_535,N_20561,N_19488);
xor UO_536 (O_536,N_20613,N_24846);
and UO_537 (O_537,N_19364,N_24749);
xor UO_538 (O_538,N_22177,N_23861);
nor UO_539 (O_539,N_22155,N_18865);
nand UO_540 (O_540,N_19382,N_21195);
nor UO_541 (O_541,N_22570,N_18785);
nor UO_542 (O_542,N_23992,N_22861);
and UO_543 (O_543,N_24172,N_19579);
or UO_544 (O_544,N_24587,N_21019);
or UO_545 (O_545,N_18826,N_23222);
nor UO_546 (O_546,N_19824,N_21456);
or UO_547 (O_547,N_21961,N_19066);
or UO_548 (O_548,N_22637,N_18996);
xnor UO_549 (O_549,N_19407,N_24073);
nor UO_550 (O_550,N_18877,N_24603);
and UO_551 (O_551,N_22805,N_20027);
or UO_552 (O_552,N_21926,N_20384);
xor UO_553 (O_553,N_21539,N_22251);
and UO_554 (O_554,N_21536,N_21408);
nand UO_555 (O_555,N_21017,N_19255);
nor UO_556 (O_556,N_23294,N_23457);
and UO_557 (O_557,N_22375,N_22106);
and UO_558 (O_558,N_21074,N_21575);
and UO_559 (O_559,N_22293,N_20075);
nor UO_560 (O_560,N_20985,N_20703);
and UO_561 (O_561,N_22392,N_23266);
nor UO_562 (O_562,N_21855,N_24252);
nand UO_563 (O_563,N_22430,N_18815);
nor UO_564 (O_564,N_19554,N_22092);
nor UO_565 (O_565,N_18983,N_19962);
and UO_566 (O_566,N_22651,N_20066);
nand UO_567 (O_567,N_22623,N_24001);
or UO_568 (O_568,N_19465,N_21923);
nand UO_569 (O_569,N_21496,N_21712);
or UO_570 (O_570,N_21521,N_19491);
nor UO_571 (O_571,N_19777,N_23372);
nor UO_572 (O_572,N_20385,N_20935);
and UO_573 (O_573,N_24231,N_22413);
nand UO_574 (O_574,N_22256,N_19943);
or UO_575 (O_575,N_24408,N_19818);
xor UO_576 (O_576,N_23862,N_22447);
or UO_577 (O_577,N_18844,N_19698);
or UO_578 (O_578,N_22043,N_19330);
nand UO_579 (O_579,N_22261,N_21888);
nand UO_580 (O_580,N_20505,N_24488);
nand UO_581 (O_581,N_21843,N_20622);
and UO_582 (O_582,N_22944,N_20406);
and UO_583 (O_583,N_24150,N_18981);
nor UO_584 (O_584,N_23770,N_23604);
nor UO_585 (O_585,N_24546,N_23208);
and UO_586 (O_586,N_22476,N_18796);
or UO_587 (O_587,N_24232,N_24216);
xnor UO_588 (O_588,N_20271,N_19031);
nand UO_589 (O_589,N_20047,N_23888);
and UO_590 (O_590,N_23314,N_21289);
or UO_591 (O_591,N_19325,N_21904);
nand UO_592 (O_592,N_18907,N_19411);
and UO_593 (O_593,N_19128,N_20516);
nor UO_594 (O_594,N_20160,N_21695);
nand UO_595 (O_595,N_22909,N_23896);
and UO_596 (O_596,N_20028,N_21915);
and UO_597 (O_597,N_23939,N_19948);
xor UO_598 (O_598,N_21767,N_19556);
and UO_599 (O_599,N_19880,N_24344);
nand UO_600 (O_600,N_21619,N_19307);
nand UO_601 (O_601,N_21435,N_20259);
and UO_602 (O_602,N_18829,N_20825);
or UO_603 (O_603,N_21145,N_23229);
nor UO_604 (O_604,N_21322,N_21490);
and UO_605 (O_605,N_20192,N_21734);
nor UO_606 (O_606,N_20084,N_19086);
nor UO_607 (O_607,N_19405,N_21047);
and UO_608 (O_608,N_19598,N_20269);
or UO_609 (O_609,N_22094,N_24547);
xor UO_610 (O_610,N_20762,N_22580);
nor UO_611 (O_611,N_23426,N_22378);
nor UO_612 (O_612,N_23976,N_24624);
and UO_613 (O_613,N_23167,N_22639);
or UO_614 (O_614,N_20354,N_21037);
nor UO_615 (O_615,N_19100,N_21515);
nand UO_616 (O_616,N_24384,N_21889);
nor UO_617 (O_617,N_24213,N_20837);
nor UO_618 (O_618,N_22334,N_18979);
or UO_619 (O_619,N_23368,N_19501);
nand UO_620 (O_620,N_22757,N_22483);
and UO_621 (O_621,N_21064,N_19428);
or UO_622 (O_622,N_21337,N_21348);
or UO_623 (O_623,N_21686,N_24610);
or UO_624 (O_624,N_19475,N_23526);
or UO_625 (O_625,N_23078,N_18786);
nand UO_626 (O_626,N_19295,N_23806);
or UO_627 (O_627,N_18912,N_20526);
or UO_628 (O_628,N_22054,N_19032);
nand UO_629 (O_629,N_21450,N_23253);
or UO_630 (O_630,N_23445,N_20456);
or UO_631 (O_631,N_18903,N_20157);
xnor UO_632 (O_632,N_24274,N_20967);
or UO_633 (O_633,N_21351,N_21405);
nor UO_634 (O_634,N_19510,N_24630);
or UO_635 (O_635,N_22780,N_21706);
nor UO_636 (O_636,N_23142,N_20194);
and UO_637 (O_637,N_21673,N_20603);
and UO_638 (O_638,N_21893,N_22220);
and UO_639 (O_639,N_24117,N_19845);
xnor UO_640 (O_640,N_19433,N_21083);
xnor UO_641 (O_641,N_22501,N_22696);
nor UO_642 (O_642,N_22064,N_24402);
and UO_643 (O_643,N_21680,N_19773);
nand UO_644 (O_644,N_20665,N_21224);
nand UO_645 (O_645,N_19571,N_19993);
xnor UO_646 (O_646,N_19010,N_18752);
or UO_647 (O_647,N_23586,N_23380);
nand UO_648 (O_648,N_21027,N_18811);
and UO_649 (O_649,N_18852,N_23193);
nor UO_650 (O_650,N_22314,N_24228);
and UO_651 (O_651,N_23215,N_23883);
or UO_652 (O_652,N_24615,N_20647);
or UO_653 (O_653,N_21015,N_22116);
and UO_654 (O_654,N_24167,N_18814);
nand UO_655 (O_655,N_22728,N_22732);
and UO_656 (O_656,N_19977,N_18931);
and UO_657 (O_657,N_24131,N_19406);
nor UO_658 (O_658,N_19907,N_19936);
and UO_659 (O_659,N_22046,N_22868);
nor UO_660 (O_660,N_21389,N_21094);
or UO_661 (O_661,N_23627,N_20494);
or UO_662 (O_662,N_24247,N_19143);
xor UO_663 (O_663,N_22893,N_19316);
nand UO_664 (O_664,N_21110,N_19214);
and UO_665 (O_665,N_19652,N_20610);
or UO_666 (O_666,N_23508,N_20793);
nor UO_667 (O_667,N_19904,N_24008);
nor UO_668 (O_668,N_20578,N_21766);
nor UO_669 (O_669,N_18802,N_24590);
and UO_670 (O_670,N_24356,N_23639);
nor UO_671 (O_671,N_20911,N_24452);
nand UO_672 (O_672,N_22339,N_18934);
nand UO_673 (O_673,N_21504,N_20675);
nand UO_674 (O_674,N_20296,N_23458);
nand UO_675 (O_675,N_21460,N_24704);
and UO_676 (O_676,N_20290,N_20891);
nand UO_677 (O_677,N_20607,N_22185);
or UO_678 (O_678,N_24248,N_20122);
or UO_679 (O_679,N_24960,N_24040);
xor UO_680 (O_680,N_21896,N_22479);
and UO_681 (O_681,N_24026,N_22709);
and UO_682 (O_682,N_20562,N_23159);
and UO_683 (O_683,N_18782,N_21884);
nand UO_684 (O_684,N_22935,N_21560);
nand UO_685 (O_685,N_22196,N_19527);
or UO_686 (O_686,N_20641,N_24021);
and UO_687 (O_687,N_21970,N_20171);
nand UO_688 (O_688,N_19339,N_24152);
nor UO_689 (O_689,N_20530,N_19467);
nor UO_690 (O_690,N_22052,N_19636);
and UO_691 (O_691,N_22684,N_23352);
nand UO_692 (O_692,N_21730,N_23817);
nand UO_693 (O_693,N_22283,N_18902);
xor UO_694 (O_694,N_22726,N_24974);
nand UO_695 (O_695,N_20279,N_22184);
nand UO_696 (O_696,N_21438,N_20376);
nor UO_697 (O_697,N_19384,N_20363);
or UO_698 (O_698,N_21630,N_24451);
nor UO_699 (O_699,N_23320,N_23533);
or UO_700 (O_700,N_20419,N_22997);
or UO_701 (O_701,N_24330,N_19176);
nor UO_702 (O_702,N_23982,N_22995);
nor UO_703 (O_703,N_20003,N_23220);
nor UO_704 (O_704,N_21489,N_23315);
or UO_705 (O_705,N_21708,N_24234);
nand UO_706 (O_706,N_21173,N_19396);
nor UO_707 (O_707,N_24349,N_24687);
nand UO_708 (O_708,N_18980,N_20646);
or UO_709 (O_709,N_24619,N_19849);
and UO_710 (O_710,N_23763,N_23626);
xnor UO_711 (O_711,N_21980,N_19398);
xnor UO_712 (O_712,N_19146,N_20134);
and UO_713 (O_713,N_20941,N_24714);
or UO_714 (O_714,N_21860,N_22319);
nor UO_715 (O_715,N_18883,N_24829);
and UO_716 (O_716,N_21830,N_21527);
or UO_717 (O_717,N_22510,N_20687);
or UO_718 (O_718,N_22698,N_22627);
or UO_719 (O_719,N_23128,N_23889);
or UO_720 (O_720,N_21065,N_24319);
or UO_721 (O_721,N_22549,N_19594);
and UO_722 (O_722,N_24509,N_20262);
nand UO_723 (O_723,N_21029,N_19368);
nand UO_724 (O_724,N_21655,N_24910);
and UO_725 (O_725,N_22062,N_23378);
nand UO_726 (O_726,N_23961,N_19236);
nand UO_727 (O_727,N_23928,N_22872);
and UO_728 (O_728,N_22572,N_22089);
or UO_729 (O_729,N_24490,N_18783);
nand UO_730 (O_730,N_22661,N_22810);
nand UO_731 (O_731,N_19714,N_21078);
and UO_732 (O_732,N_21890,N_22081);
or UO_733 (O_733,N_22286,N_21749);
nor UO_734 (O_734,N_22856,N_24197);
or UO_735 (O_735,N_24931,N_24286);
or UO_736 (O_736,N_21344,N_21786);
nand UO_737 (O_737,N_23825,N_22847);
and UO_738 (O_738,N_19841,N_22553);
or UO_739 (O_739,N_19939,N_22804);
nor UO_740 (O_740,N_21323,N_18761);
nand UO_741 (O_741,N_18860,N_20868);
and UO_742 (O_742,N_18926,N_20792);
or UO_743 (O_743,N_24850,N_24626);
nand UO_744 (O_744,N_18754,N_23686);
nand UO_745 (O_745,N_20324,N_22986);
nor UO_746 (O_746,N_20885,N_23962);
and UO_747 (O_747,N_23042,N_24920);
nor UO_748 (O_748,N_22059,N_22007);
and UO_749 (O_749,N_20591,N_20560);
or UO_750 (O_750,N_23751,N_20711);
or UO_751 (O_751,N_19531,N_23940);
nand UO_752 (O_752,N_24969,N_24457);
and UO_753 (O_753,N_19813,N_19882);
nand UO_754 (O_754,N_19543,N_22632);
nand UO_755 (O_755,N_18946,N_20584);
nor UO_756 (O_756,N_20838,N_24218);
and UO_757 (O_757,N_20486,N_19085);
or UO_758 (O_758,N_24596,N_24563);
nand UO_759 (O_759,N_23905,N_19131);
nand UO_760 (O_760,N_19765,N_19960);
nand UO_761 (O_761,N_24169,N_18766);
or UO_762 (O_762,N_19534,N_24153);
and UO_763 (O_763,N_20136,N_23202);
and UO_764 (O_764,N_24444,N_20320);
nor UO_765 (O_765,N_22228,N_24614);
and UO_766 (O_766,N_24233,N_22444);
and UO_767 (O_767,N_22603,N_18838);
and UO_768 (O_768,N_18995,N_20013);
or UO_769 (O_769,N_24854,N_23821);
nor UO_770 (O_770,N_24534,N_19736);
or UO_771 (O_771,N_23440,N_22964);
and UO_772 (O_772,N_22862,N_24862);
nand UO_773 (O_773,N_22284,N_20532);
and UO_774 (O_774,N_24039,N_24044);
or UO_775 (O_775,N_18800,N_23492);
nor UO_776 (O_776,N_23663,N_24116);
nand UO_777 (O_777,N_23237,N_22841);
nand UO_778 (O_778,N_20254,N_20619);
nor UO_779 (O_779,N_22120,N_22921);
and UO_780 (O_780,N_20664,N_20445);
and UO_781 (O_781,N_19145,N_22453);
nor UO_782 (O_782,N_23106,N_23851);
nor UO_783 (O_783,N_24414,N_24562);
nor UO_784 (O_784,N_24771,N_18913);
nand UO_785 (O_785,N_22183,N_23304);
xor UO_786 (O_786,N_22762,N_19460);
or UO_787 (O_787,N_21353,N_19914);
nand UO_788 (O_788,N_24024,N_23644);
nand UO_789 (O_789,N_20012,N_21054);
and UO_790 (O_790,N_24013,N_22731);
xor UO_791 (O_791,N_21452,N_23477);
or UO_792 (O_792,N_19973,N_21566);
nand UO_793 (O_793,N_21924,N_21433);
nand UO_794 (O_794,N_20393,N_20228);
xor UO_795 (O_795,N_22381,N_20670);
or UO_796 (O_796,N_22361,N_24900);
nand UO_797 (O_797,N_24962,N_23668);
and UO_798 (O_798,N_23300,N_19437);
or UO_799 (O_799,N_21155,N_23886);
nand UO_800 (O_800,N_24908,N_20576);
nor UO_801 (O_801,N_21902,N_24600);
and UO_802 (O_802,N_21750,N_23747);
nor UO_803 (O_803,N_24564,N_21725);
nand UO_804 (O_804,N_21736,N_19373);
nand UO_805 (O_805,N_20274,N_19801);
or UO_806 (O_806,N_21409,N_20332);
xor UO_807 (O_807,N_24481,N_24178);
or UO_808 (O_808,N_19273,N_23699);
or UO_809 (O_809,N_19258,N_22275);
nand UO_810 (O_810,N_19743,N_23611);
and UO_811 (O_811,N_21593,N_24634);
nor UO_812 (O_812,N_24644,N_19538);
nand UO_813 (O_813,N_20088,N_23133);
and UO_814 (O_814,N_21451,N_23148);
nor UO_815 (O_815,N_22365,N_20547);
nor UO_816 (O_816,N_20866,N_19144);
and UO_817 (O_817,N_19621,N_23946);
or UO_818 (O_818,N_21388,N_20559);
or UO_819 (O_819,N_22001,N_24238);
nor UO_820 (O_820,N_19679,N_22845);
and UO_821 (O_821,N_19429,N_23761);
and UO_822 (O_822,N_24795,N_22598);
nor UO_823 (O_823,N_21298,N_21108);
nor UO_824 (O_824,N_18880,N_22621);
or UO_825 (O_825,N_21815,N_24204);
nor UO_826 (O_826,N_23941,N_21147);
and UO_827 (O_827,N_19164,N_19963);
nand UO_828 (O_828,N_20033,N_24128);
nand UO_829 (O_829,N_20582,N_22963);
xor UO_830 (O_830,N_21210,N_19984);
and UO_831 (O_831,N_24459,N_20049);
and UO_832 (O_832,N_20545,N_22053);
nor UO_833 (O_833,N_19615,N_24187);
or UO_834 (O_834,N_20773,N_24348);
nor UO_835 (O_835,N_23186,N_19895);
or UO_836 (O_836,N_19217,N_21144);
xor UO_837 (O_837,N_20688,N_20437);
and UO_838 (O_838,N_24137,N_20571);
nor UO_839 (O_839,N_20369,N_24952);
nor UO_840 (O_840,N_22978,N_20214);
and UO_841 (O_841,N_20380,N_20929);
nor UO_842 (O_842,N_24327,N_24941);
xnor UO_843 (O_843,N_21109,N_23810);
nand UO_844 (O_844,N_24308,N_18897);
and UO_845 (O_845,N_23031,N_24164);
nand UO_846 (O_846,N_23060,N_19299);
or UO_847 (O_847,N_20447,N_18993);
or UO_848 (O_848,N_18791,N_21548);
and UO_849 (O_849,N_21023,N_19752);
nor UO_850 (O_850,N_21871,N_24557);
nor UO_851 (O_851,N_24635,N_24636);
nand UO_852 (O_852,N_22385,N_24281);
nor UO_853 (O_853,N_21264,N_19596);
and UO_854 (O_854,N_20697,N_22827);
or UO_855 (O_855,N_23554,N_19523);
nand UO_856 (O_856,N_21723,N_19132);
and UO_857 (O_857,N_20415,N_22620);
and UO_858 (O_858,N_22034,N_22672);
xor UO_859 (O_859,N_20869,N_22524);
nand UO_860 (O_860,N_19755,N_24828);
xnor UO_861 (O_861,N_19490,N_21779);
or UO_862 (O_862,N_24083,N_20719);
or UO_863 (O_863,N_22557,N_20373);
nor UO_864 (O_864,N_19894,N_22264);
nor UO_865 (O_865,N_22341,N_21697);
or UO_866 (O_866,N_23348,N_20874);
nor UO_867 (O_867,N_22044,N_20709);
and UO_868 (O_868,N_19223,N_20865);
and UO_869 (O_869,N_23739,N_19492);
nor UO_870 (O_870,N_19933,N_20778);
or UO_871 (O_871,N_19387,N_24379);
nor UO_872 (O_872,N_21853,N_19450);
or UO_873 (O_873,N_24261,N_24843);
and UO_874 (O_874,N_21254,N_22546);
nor UO_875 (O_875,N_20463,N_20117);
or UO_876 (O_876,N_20528,N_21895);
or UO_877 (O_877,N_24392,N_23158);
nand UO_878 (O_878,N_24654,N_23432);
or UO_879 (O_879,N_19495,N_19431);
nor UO_880 (O_880,N_19639,N_24180);
nor UO_881 (O_881,N_23633,N_24345);
or UO_882 (O_882,N_23292,N_23180);
nor UO_883 (O_883,N_22117,N_19409);
or UO_884 (O_884,N_24280,N_22880);
or UO_885 (O_885,N_21596,N_20073);
and UO_886 (O_886,N_24236,N_24885);
and UO_887 (O_887,N_20072,N_19439);
and UO_888 (O_888,N_23734,N_20895);
and UO_889 (O_889,N_23645,N_19269);
nor UO_890 (O_890,N_24043,N_20394);
nand UO_891 (O_891,N_21651,N_20329);
nand UO_892 (O_892,N_19053,N_23802);
xor UO_893 (O_893,N_19250,N_23999);
nand UO_894 (O_894,N_24715,N_19421);
and UO_895 (O_895,N_20747,N_21270);
nor UO_896 (O_896,N_22394,N_22350);
nand UO_897 (O_897,N_20473,N_20696);
or UO_898 (O_898,N_21558,N_24183);
nor UO_899 (O_899,N_19658,N_21263);
xor UO_900 (O_900,N_24383,N_23848);
nand UO_901 (O_901,N_19477,N_21999);
nor UO_902 (O_902,N_24181,N_24831);
or UO_903 (O_903,N_21600,N_21788);
nor UO_904 (O_904,N_21554,N_21916);
nand UO_905 (O_905,N_19979,N_23729);
or UO_906 (O_906,N_22492,N_19678);
xnor UO_907 (O_907,N_22137,N_20700);
nand UO_908 (O_908,N_20978,N_23592);
nand UO_909 (O_909,N_22512,N_20404);
nor UO_910 (O_910,N_20686,N_22474);
xnor UO_911 (O_911,N_21633,N_24907);
or UO_912 (O_912,N_24911,N_21239);
and UO_913 (O_913,N_21985,N_21777);
nand UO_914 (O_914,N_19637,N_20761);
and UO_915 (O_915,N_23207,N_23165);
and UO_916 (O_916,N_24732,N_18859);
and UO_917 (O_917,N_22239,N_23157);
nand UO_918 (O_918,N_22039,N_19213);
xnor UO_919 (O_919,N_22892,N_22820);
xor UO_920 (O_920,N_22171,N_21458);
nor UO_921 (O_921,N_21010,N_24114);
nor UO_922 (O_922,N_23080,N_20052);
and UO_923 (O_923,N_21420,N_22715);
nor UO_924 (O_924,N_24720,N_23079);
nand UO_925 (O_925,N_22331,N_23678);
and UO_926 (O_926,N_22072,N_23041);
nor UO_927 (O_927,N_23061,N_20011);
nand UO_928 (O_928,N_19889,N_20218);
nor UO_929 (O_929,N_24378,N_20234);
nand UO_930 (O_930,N_21740,N_24770);
and UO_931 (O_931,N_20944,N_22811);
or UO_932 (O_932,N_20241,N_23792);
nor UO_933 (O_933,N_23475,N_20189);
nand UO_934 (O_934,N_22400,N_22673);
nor UO_935 (O_935,N_24943,N_21345);
nand UO_936 (O_936,N_20733,N_22547);
and UO_937 (O_937,N_22976,N_24271);
or UO_938 (O_938,N_23582,N_19512);
or UO_939 (O_939,N_24998,N_20266);
nand UO_940 (O_940,N_24762,N_24058);
and UO_941 (O_941,N_20431,N_18868);
nand UO_942 (O_942,N_18937,N_22029);
and UO_943 (O_943,N_23471,N_21868);
xor UO_944 (O_944,N_24733,N_18809);
and UO_945 (O_945,N_23956,N_22478);
nand UO_946 (O_946,N_20103,N_21207);
nand UO_947 (O_947,N_23415,N_19098);
nand UO_948 (O_948,N_20848,N_20872);
nor UO_949 (O_949,N_22382,N_22427);
nor UO_950 (O_950,N_19928,N_21984);
nand UO_951 (O_951,N_20730,N_20738);
and UO_952 (O_952,N_21562,N_23713);
nand UO_953 (O_953,N_19425,N_23856);
and UO_954 (O_954,N_24725,N_23280);
nand UO_955 (O_955,N_19703,N_21211);
and UO_956 (O_956,N_22617,N_23170);
or UO_957 (O_957,N_24553,N_22038);
nor UO_958 (O_958,N_22435,N_20635);
and UO_959 (O_959,N_19593,N_20386);
and UO_960 (O_960,N_22743,N_20149);
nand UO_961 (O_961,N_20175,N_19583);
nor UO_962 (O_962,N_18882,N_19562);
or UO_963 (O_963,N_23548,N_19776);
or UO_964 (O_964,N_21320,N_23444);
nor UO_965 (O_965,N_23733,N_23689);
nand UO_966 (O_966,N_23312,N_23855);
or UO_967 (O_967,N_22741,N_23666);
nor UO_968 (O_968,N_18956,N_18966);
xnor UO_969 (O_969,N_22996,N_19644);
nand UO_970 (O_970,N_24726,N_20524);
nor UO_971 (O_971,N_22475,N_21621);
or UO_972 (O_972,N_20102,N_24815);
nor UO_973 (O_973,N_20937,N_21226);
nand UO_974 (O_974,N_19084,N_21459);
nor UO_975 (O_975,N_21325,N_24810);
nand UO_976 (O_976,N_22695,N_20099);
or UO_977 (O_977,N_20692,N_24282);
or UO_978 (O_978,N_21423,N_23767);
nand UO_979 (O_979,N_24135,N_19618);
nor UO_980 (O_980,N_18887,N_24310);
xnor UO_981 (O_981,N_21334,N_23004);
nand UO_982 (O_982,N_23545,N_24255);
and UO_983 (O_983,N_22869,N_20137);
and UO_984 (O_984,N_19741,N_19048);
nand UO_985 (O_985,N_19462,N_22851);
or UO_986 (O_986,N_20553,N_20902);
nor UO_987 (O_987,N_22278,N_22408);
and UO_988 (O_988,N_23577,N_24641);
and UO_989 (O_989,N_21335,N_20442);
nor UO_990 (O_990,N_24514,N_20875);
nand UO_991 (O_991,N_22303,N_22130);
nor UO_992 (O_992,N_19831,N_21892);
or UO_993 (O_993,N_21143,N_24202);
or UO_994 (O_994,N_22701,N_21008);
nor UO_995 (O_995,N_24739,N_20831);
xor UO_996 (O_996,N_23410,N_24305);
nand UO_997 (O_997,N_20556,N_21835);
or UO_998 (O_998,N_23342,N_21371);
nor UO_999 (O_999,N_21004,N_24182);
nor UO_1000 (O_1000,N_22321,N_24082);
xor UO_1001 (O_1001,N_20766,N_24809);
nand UO_1002 (O_1002,N_19890,N_21048);
and UO_1003 (O_1003,N_23059,N_18920);
nand UO_1004 (O_1004,N_24755,N_24464);
or UO_1005 (O_1005,N_19153,N_21053);
nor UO_1006 (O_1006,N_19507,N_21689);
or UO_1007 (O_1007,N_23931,N_24283);
or UO_1008 (O_1008,N_23068,N_20758);
nor UO_1009 (O_1009,N_22421,N_21545);
and UO_1010 (O_1010,N_20971,N_21918);
nor UO_1011 (O_1011,N_22705,N_23564);
xor UO_1012 (O_1012,N_22877,N_24084);
or UO_1013 (O_1013,N_24166,N_18784);
xnor UO_1014 (O_1014,N_23704,N_19054);
or UO_1015 (O_1015,N_24814,N_19249);
and UO_1016 (O_1016,N_19254,N_22777);
and UO_1017 (O_1017,N_23595,N_19829);
nor UO_1018 (O_1018,N_23430,N_20001);
nand UO_1019 (O_1019,N_21352,N_23840);
nand UO_1020 (O_1020,N_21024,N_19710);
nor UO_1021 (O_1021,N_21447,N_24602);
nor UO_1022 (O_1022,N_23694,N_20022);
nand UO_1023 (O_1023,N_19975,N_20974);
nand UO_1024 (O_1024,N_23009,N_21281);
nand UO_1025 (O_1025,N_19582,N_23569);
nor UO_1026 (O_1026,N_19478,N_22057);
and UO_1027 (O_1027,N_24397,N_19614);
nor UO_1028 (O_1028,N_20628,N_23773);
or UO_1029 (O_1029,N_22157,N_22036);
nand UO_1030 (O_1030,N_22225,N_19935);
and UO_1031 (O_1031,N_21679,N_22906);
nor UO_1032 (O_1032,N_22573,N_24366);
nand UO_1033 (O_1033,N_19284,N_19082);
nor UO_1034 (O_1034,N_19286,N_19365);
nand UO_1035 (O_1035,N_24474,N_23010);
xnor UO_1036 (O_1036,N_22515,N_22189);
nor UO_1037 (O_1037,N_24942,N_21693);
or UO_1038 (O_1038,N_19202,N_20152);
and UO_1039 (O_1039,N_18837,N_19392);
or UO_1040 (O_1040,N_19689,N_19696);
xor UO_1041 (O_1041,N_21644,N_19862);
nand UO_1042 (O_1042,N_24697,N_24648);
nand UO_1043 (O_1043,N_23558,N_22583);
or UO_1044 (O_1044,N_24388,N_20434);
nand UO_1045 (O_1045,N_24210,N_23981);
or UO_1046 (O_1046,N_21253,N_20521);
nor UO_1047 (O_1047,N_23854,N_21603);
or UO_1048 (O_1048,N_19184,N_21526);
or UO_1049 (O_1049,N_24670,N_21060);
nand UO_1050 (O_1050,N_20889,N_19156);
nor UO_1051 (O_1051,N_23235,N_23804);
nand UO_1052 (O_1052,N_23780,N_23500);
nand UO_1053 (O_1053,N_24774,N_20219);
nand UO_1054 (O_1054,N_21005,N_20238);
and UO_1055 (O_1055,N_24276,N_20045);
or UO_1056 (O_1056,N_23205,N_23421);
and UO_1057 (O_1057,N_24351,N_21646);
nand UO_1058 (O_1058,N_19173,N_19035);
nor UO_1059 (O_1059,N_19137,N_22959);
nor UO_1060 (O_1060,N_23648,N_22006);
nand UO_1061 (O_1061,N_23409,N_23917);
or UO_1062 (O_1062,N_23512,N_23579);
and UO_1063 (O_1063,N_20554,N_21481);
nor UO_1064 (O_1064,N_19520,N_24226);
nor UO_1065 (O_1065,N_19891,N_21632);
and UO_1066 (O_1066,N_19014,N_19629);
nand UO_1067 (O_1067,N_23140,N_24574);
nand UO_1068 (O_1068,N_19113,N_20032);
nor UO_1069 (O_1069,N_19853,N_22923);
nor UO_1070 (O_1070,N_24918,N_22677);
or UO_1071 (O_1071,N_19264,N_23570);
and UO_1072 (O_1072,N_21937,N_24009);
and UO_1073 (O_1073,N_24483,N_24570);
nor UO_1074 (O_1074,N_23912,N_24863);
or UO_1075 (O_1075,N_24406,N_24989);
or UO_1076 (O_1076,N_18875,N_23084);
or UO_1077 (O_1077,N_21785,N_23984);
and UO_1078 (O_1078,N_20905,N_23784);
nor UO_1079 (O_1079,N_20095,N_24399);
or UO_1080 (O_1080,N_19481,N_18810);
nand UO_1081 (O_1081,N_24802,N_22428);
xor UO_1082 (O_1082,N_23647,N_22806);
xor UO_1083 (O_1083,N_20800,N_22965);
xnor UO_1084 (O_1084,N_23555,N_20307);
and UO_1085 (O_1085,N_19498,N_18817);
nand UO_1086 (O_1086,N_24462,N_20357);
and UO_1087 (O_1087,N_24744,N_24957);
xnor UO_1088 (O_1088,N_20041,N_22005);
nor UO_1089 (O_1089,N_22069,N_24549);
or UO_1090 (O_1090,N_22543,N_23833);
or UO_1091 (O_1091,N_24185,N_20695);
or UO_1092 (O_1092,N_20344,N_19968);
xor UO_1093 (O_1093,N_21721,N_24328);
nand UO_1094 (O_1094,N_24967,N_20495);
and UO_1095 (O_1095,N_18832,N_19225);
nand UO_1096 (O_1096,N_19220,N_19530);
nor UO_1097 (O_1097,N_20514,N_22449);
or UO_1098 (O_1098,N_21790,N_24301);
or UO_1099 (O_1099,N_20517,N_24045);
or UO_1100 (O_1100,N_21201,N_22562);
nor UO_1101 (O_1101,N_24751,N_23901);
and UO_1102 (O_1102,N_21694,N_21565);
or UO_1103 (O_1103,N_23046,N_20919);
or UO_1104 (O_1104,N_23539,N_19363);
and UO_1105 (O_1105,N_24449,N_19055);
nand UO_1106 (O_1106,N_22482,N_21972);
nor UO_1107 (O_1107,N_20920,N_19093);
nand UO_1108 (O_1108,N_19951,N_19109);
or UO_1109 (O_1109,N_23978,N_23303);
or UO_1110 (O_1110,N_22839,N_21465);
nand UO_1111 (O_1111,N_23649,N_23665);
nor UO_1112 (O_1112,N_23323,N_23587);
and UO_1113 (O_1113,N_19472,N_22739);
and UO_1114 (O_1114,N_23980,N_19909);
nand UO_1115 (O_1115,N_20432,N_20934);
or UO_1116 (O_1116,N_23514,N_19252);
nand UO_1117 (O_1117,N_19656,N_22247);
nand UO_1118 (O_1118,N_19305,N_23636);
nor UO_1119 (O_1119,N_23468,N_22292);
nor UO_1120 (O_1120,N_23227,N_22252);
and UO_1121 (O_1121,N_24662,N_19438);
or UO_1122 (O_1122,N_22858,N_22172);
nor UO_1123 (O_1123,N_19692,N_22019);
nor UO_1124 (O_1124,N_21618,N_20513);
or UO_1125 (O_1125,N_23996,N_24538);
nor UO_1126 (O_1126,N_20006,N_19377);
or UO_1127 (O_1127,N_21658,N_21622);
and UO_1128 (O_1128,N_21462,N_20531);
nor UO_1129 (O_1129,N_19417,N_23025);
and UO_1130 (O_1130,N_20682,N_19785);
and UO_1131 (O_1131,N_24417,N_20164);
xor UO_1132 (O_1132,N_24870,N_20382);
and UO_1133 (O_1133,N_21606,N_24053);
and UO_1134 (O_1134,N_21911,N_23803);
nand UO_1135 (O_1135,N_19957,N_21577);
nor UO_1136 (O_1136,N_21089,N_22604);
nand UO_1137 (O_1137,N_24317,N_22765);
and UO_1138 (O_1138,N_21355,N_19165);
nand UO_1139 (O_1139,N_23211,N_22469);
nor UO_1140 (O_1140,N_19059,N_19509);
and UO_1141 (O_1141,N_21365,N_24450);
nor UO_1142 (O_1142,N_22587,N_22023);
nand UO_1143 (O_1143,N_20683,N_20677);
or UO_1144 (O_1144,N_21838,N_24867);
nand UO_1145 (O_1145,N_21395,N_19279);
nor UO_1146 (O_1146,N_24403,N_24223);
nor UO_1147 (O_1147,N_22903,N_24205);
and UO_1148 (O_1148,N_22085,N_20147);
and UO_1149 (O_1149,N_24161,N_22692);
or UO_1150 (O_1150,N_19210,N_23899);
nand UO_1151 (O_1151,N_24659,N_24639);
nor UO_1152 (O_1152,N_23197,N_22383);
nor UO_1153 (O_1153,N_23485,N_22156);
and UO_1154 (O_1154,N_24127,N_24582);
xor UO_1155 (O_1155,N_21819,N_21457);
and UO_1156 (O_1156,N_22233,N_22618);
or UO_1157 (O_1157,N_20193,N_19121);
and UO_1158 (O_1158,N_21783,N_19069);
or UO_1159 (O_1159,N_24924,N_20409);
and UO_1160 (O_1160,N_24794,N_21994);
or UO_1161 (O_1161,N_22289,N_24995);
nand UO_1162 (O_1162,N_22355,N_24072);
or UO_1163 (O_1163,N_24198,N_23643);
nor UO_1164 (O_1164,N_24243,N_23008);
nand UO_1165 (O_1165,N_22080,N_21763);
nor UO_1166 (O_1166,N_24529,N_23549);
or UO_1167 (O_1167,N_19902,N_22616);
nor UO_1168 (O_1168,N_19848,N_24987);
and UO_1169 (O_1169,N_23224,N_24120);
xnor UO_1170 (O_1170,N_23472,N_21483);
and UO_1171 (O_1171,N_24597,N_20702);
xor UO_1172 (O_1172,N_19308,N_20187);
nor UO_1173 (O_1173,N_24660,N_24374);
nand UO_1174 (O_1174,N_20478,N_19449);
nand UO_1175 (O_1175,N_24189,N_20133);
and UO_1176 (O_1176,N_21557,N_23343);
nand UO_1177 (O_1177,N_24988,N_24782);
and UO_1178 (O_1178,N_18961,N_20295);
or UO_1179 (O_1179,N_21543,N_23160);
nor UO_1180 (O_1180,N_20574,N_19107);
and UO_1181 (O_1181,N_24981,N_21326);
and UO_1182 (O_1182,N_23013,N_23612);
or UO_1183 (O_1183,N_19000,N_20347);
or UO_1184 (O_1184,N_23260,N_19027);
nor UO_1185 (O_1185,N_20880,N_21373);
xor UO_1186 (O_1186,N_21666,N_18969);
nand UO_1187 (O_1187,N_22665,N_22132);
nand UO_1188 (O_1188,N_22714,N_23603);
and UO_1189 (O_1189,N_23530,N_22532);
nand UO_1190 (O_1190,N_20396,N_19774);
nor UO_1191 (O_1191,N_19242,N_24438);
nand UO_1192 (O_1192,N_20525,N_24682);
nand UO_1193 (O_1193,N_22752,N_24445);
and UO_1194 (O_1194,N_23561,N_21761);
or UO_1195 (O_1195,N_23030,N_19361);
nand UO_1196 (O_1196,N_21252,N_24827);
or UO_1197 (O_1197,N_19781,N_23460);
nor UO_1198 (O_1198,N_23765,N_23881);
nor UO_1199 (O_1199,N_20830,N_21250);
and UO_1200 (O_1200,N_22088,N_19870);
nor UO_1201 (O_1201,N_21636,N_21826);
and UO_1202 (O_1202,N_22686,N_23836);
nand UO_1203 (O_1203,N_19647,N_21237);
and UO_1204 (O_1204,N_19946,N_19790);
nor UO_1205 (O_1205,N_22766,N_24877);
and UO_1206 (O_1206,N_19201,N_24051);
nand UO_1207 (O_1207,N_24041,N_20444);
nand UO_1208 (O_1208,N_19903,N_22650);
xor UO_1209 (O_1209,N_19660,N_19390);
nor UO_1210 (O_1210,N_19464,N_20439);
xnor UO_1211 (O_1211,N_23448,N_22197);
and UO_1212 (O_1212,N_24029,N_24919);
nand UO_1213 (O_1213,N_22609,N_19700);
or UO_1214 (O_1214,N_19205,N_21380);
xor UO_1215 (O_1215,N_23826,N_19344);
nand UO_1216 (O_1216,N_22288,N_18857);
nor UO_1217 (O_1217,N_22550,N_23986);
nand UO_1218 (O_1218,N_20926,N_24761);
nor UO_1219 (O_1219,N_24606,N_22783);
nor UO_1220 (O_1220,N_20023,N_24699);
nor UO_1221 (O_1221,N_22369,N_18964);
nor UO_1222 (O_1222,N_18755,N_21104);
or UO_1223 (O_1223,N_24579,N_20693);
or UO_1224 (O_1224,N_19381,N_21426);
nor UO_1225 (O_1225,N_22307,N_20402);
or UO_1226 (O_1226,N_21115,N_24253);
nand UO_1227 (O_1227,N_19567,N_22831);
nor UO_1228 (O_1228,N_23876,N_21248);
and UO_1229 (O_1229,N_23110,N_18822);
or UO_1230 (O_1230,N_23798,N_21448);
nor UO_1231 (O_1231,N_19092,N_19080);
nor UO_1232 (O_1232,N_20139,N_19532);
nor UO_1233 (O_1233,N_19262,N_23908);
and UO_1234 (O_1234,N_20827,N_20339);
nand UO_1235 (O_1235,N_20727,N_21876);
xor UO_1236 (O_1236,N_19756,N_24047);
nor UO_1237 (O_1237,N_19551,N_19312);
or UO_1238 (O_1238,N_22537,N_23143);
nor UO_1239 (O_1239,N_20081,N_19566);
or UO_1240 (O_1240,N_22488,N_24906);
nand UO_1241 (O_1241,N_21431,N_24723);
nand UO_1242 (O_1242,N_21700,N_19385);
or UO_1243 (O_1243,N_24684,N_24077);
nor UO_1244 (O_1244,N_19980,N_20725);
or UO_1245 (O_1245,N_20483,N_21947);
nor UO_1246 (O_1246,N_22648,N_23726);
nand UO_1247 (O_1247,N_23226,N_21363);
nand UO_1248 (O_1248,N_23551,N_24209);
nand UO_1249 (O_1249,N_20400,N_19120);
or UO_1250 (O_1250,N_24173,N_21343);
nand UO_1251 (O_1251,N_22681,N_21513);
nand UO_1252 (O_1252,N_19820,N_19002);
nand UO_1253 (O_1253,N_20210,N_21589);
nand UO_1254 (O_1254,N_19457,N_22795);
nor UO_1255 (O_1255,N_23264,N_22181);
nor UO_1256 (O_1256,N_19959,N_19496);
xor UO_1257 (O_1257,N_22055,N_21471);
xnor UO_1258 (O_1258,N_22245,N_22594);
nor UO_1259 (O_1259,N_19207,N_23828);
nand UO_1260 (O_1260,N_23977,N_23842);
or UO_1261 (O_1261,N_20860,N_23523);
nand UO_1262 (O_1262,N_19151,N_23968);
xnor UO_1263 (O_1263,N_20541,N_22625);
xor UO_1264 (O_1264,N_21375,N_20859);
xor UO_1265 (O_1265,N_18794,N_19389);
and UO_1266 (O_1266,N_24410,N_19683);
or UO_1267 (O_1267,N_24511,N_20506);
nand UO_1268 (O_1268,N_21191,N_23321);
nand UO_1269 (O_1269,N_19666,N_24431);
xnor UO_1270 (O_1270,N_19260,N_22565);
or UO_1271 (O_1271,N_24080,N_21849);
xnor UO_1272 (O_1272,N_21752,N_20297);
and UO_1273 (O_1273,N_19130,N_24493);
nand UO_1274 (O_1274,N_19589,N_18798);
nor UO_1275 (O_1275,N_24983,N_22899);
nor UO_1276 (O_1276,N_19622,N_21152);
nand UO_1277 (O_1277,N_20252,N_22828);
nand UO_1278 (O_1278,N_22152,N_24932);
and UO_1279 (O_1279,N_22652,N_22750);
and UO_1280 (O_1280,N_19052,N_22736);
and UO_1281 (O_1281,N_21703,N_23698);
nor UO_1282 (O_1282,N_19965,N_22174);
nand UO_1283 (O_1283,N_19412,N_18862);
xnor UO_1284 (O_1284,N_19747,N_21591);
and UO_1285 (O_1285,N_20457,N_22818);
nand UO_1286 (O_1286,N_24355,N_24496);
or UO_1287 (O_1287,N_20909,N_20349);
and UO_1288 (O_1288,N_23149,N_19816);
nand UO_1289 (O_1289,N_20877,N_19005);
xor UO_1290 (O_1290,N_22009,N_23453);
and UO_1291 (O_1291,N_24023,N_21235);
or UO_1292 (O_1292,N_23146,N_23692);
nor UO_1293 (O_1293,N_19041,N_19982);
and UO_1294 (O_1294,N_23522,N_19033);
nand UO_1295 (O_1295,N_20126,N_21463);
nand UO_1296 (O_1296,N_23716,N_18941);
xnor UO_1297 (O_1297,N_21927,N_23136);
or UO_1298 (O_1298,N_18762,N_24953);
and UO_1299 (O_1299,N_20170,N_22342);
or UO_1300 (O_1300,N_23691,N_24777);
or UO_1301 (O_1301,N_18858,N_22507);
nor UO_1302 (O_1302,N_20981,N_20844);
nor UO_1303 (O_1303,N_21722,N_21672);
and UO_1304 (O_1304,N_19826,N_22755);
and UO_1305 (O_1305,N_23701,N_23150);
xor UO_1306 (O_1306,N_19859,N_23027);
xnor UO_1307 (O_1307,N_24369,N_19135);
nor UO_1308 (O_1308,N_20176,N_20735);
nor UO_1309 (O_1309,N_23384,N_23878);
and UO_1310 (O_1310,N_21214,N_22680);
nand UO_1311 (O_1311,N_19568,N_23808);
nor UO_1312 (O_1312,N_21455,N_20461);
or UO_1313 (O_1313,N_22646,N_22405);
or UO_1314 (O_1314,N_21816,N_24237);
nand UO_1315 (O_1315,N_23903,N_24818);
nor UO_1316 (O_1316,N_23474,N_23532);
xor UO_1317 (O_1317,N_19950,N_22219);
xor UO_1318 (O_1318,N_22500,N_20723);
and UO_1319 (O_1319,N_19147,N_18797);
and UO_1320 (O_1320,N_24575,N_23664);
nor UO_1321 (O_1321,N_18840,N_19110);
or UO_1322 (O_1322,N_23035,N_20340);
nor UO_1323 (O_1323,N_19424,N_18776);
and UO_1324 (O_1324,N_19221,N_21880);
and UO_1325 (O_1325,N_21547,N_24422);
or UO_1326 (O_1326,N_18830,N_18925);
or UO_1327 (O_1327,N_24394,N_24506);
nor UO_1328 (O_1328,N_22274,N_24336);
nor UO_1329 (O_1329,N_19253,N_23637);
or UO_1330 (O_1330,N_20824,N_23831);
nor UO_1331 (O_1331,N_24176,N_20557);
nor UO_1332 (O_1332,N_22363,N_21671);
or UO_1333 (O_1333,N_24147,N_20914);
nand UO_1334 (O_1334,N_19015,N_19918);
nand UO_1335 (O_1335,N_24074,N_20585);
or UO_1336 (O_1336,N_20713,N_19423);
or UO_1337 (O_1337,N_19709,N_22682);
nand UO_1338 (O_1338,N_19400,N_20718);
or UO_1339 (O_1339,N_23311,N_20572);
and UO_1340 (O_1340,N_22654,N_21025);
nand UO_1341 (O_1341,N_23048,N_21194);
nor UO_1342 (O_1342,N_22802,N_22070);
nand UO_1343 (O_1343,N_21794,N_20129);
xor UO_1344 (O_1344,N_19182,N_20226);
or UO_1345 (O_1345,N_22531,N_20659);
and UO_1346 (O_1346,N_24513,N_23081);
and UO_1347 (O_1347,N_24708,N_24269);
and UO_1348 (O_1348,N_18831,N_23900);
nor UO_1349 (O_1349,N_21206,N_23302);
nor UO_1350 (O_1350,N_23964,N_24497);
nor UO_1351 (O_1351,N_22458,N_24121);
and UO_1352 (O_1352,N_24257,N_21773);
or UO_1353 (O_1353,N_24254,N_24719);
nor UO_1354 (O_1354,N_20654,N_20230);
nor UO_1355 (O_1355,N_21607,N_20768);
or UO_1356 (O_1356,N_22535,N_23925);
xnor UO_1357 (O_1357,N_24525,N_21653);
nand UO_1358 (O_1358,N_21347,N_22300);
nor UO_1359 (O_1359,N_23756,N_19383);
nor UO_1360 (O_1360,N_20309,N_24951);
and UO_1361 (O_1361,N_22465,N_21361);
and UO_1362 (O_1362,N_24784,N_18836);
nand UO_1363 (O_1363,N_22712,N_22520);
nand UO_1364 (O_1364,N_22503,N_21414);
xnor UO_1365 (O_1365,N_19789,N_20789);
or UO_1366 (O_1366,N_20135,N_22634);
nor UO_1367 (O_1367,N_18790,N_24367);
xor UO_1368 (O_1368,N_21134,N_21594);
nand UO_1369 (O_1369,N_21170,N_23107);
or UO_1370 (O_1370,N_19766,N_22356);
or UO_1371 (O_1371,N_24661,N_24819);
xnor UO_1372 (O_1372,N_24398,N_21900);
and UO_1373 (O_1373,N_22146,N_24331);
and UO_1374 (O_1374,N_21275,N_21432);
or UO_1375 (O_1375,N_20304,N_24930);
nand UO_1376 (O_1376,N_21988,N_21076);
or UO_1377 (O_1377,N_20790,N_18763);
nand UO_1378 (O_1378,N_22998,N_21209);
nor UO_1379 (O_1379,N_24306,N_20180);
and UO_1380 (O_1380,N_19746,N_21878);
nand UO_1381 (O_1381,N_22470,N_24289);
or UO_1382 (O_1382,N_21120,N_23375);
or UO_1383 (O_1383,N_24094,N_23413);
or UO_1384 (O_1384,N_20159,N_22874);
and UO_1385 (O_1385,N_24019,N_20722);
nand UO_1386 (O_1386,N_19215,N_21225);
and UO_1387 (O_1387,N_21099,N_20529);
and UO_1388 (O_1388,N_19599,N_21177);
and UO_1389 (O_1389,N_22136,N_21556);
or UO_1390 (O_1390,N_24341,N_20987);
and UO_1391 (O_1391,N_22310,N_21992);
nor UO_1392 (O_1392,N_19924,N_23635);
or UO_1393 (O_1393,N_23656,N_23882);
nand UO_1394 (O_1394,N_24244,N_23433);
nor UO_1395 (O_1395,N_21111,N_23676);
and UO_1396 (O_1396,N_22947,N_20537);
xor UO_1397 (O_1397,N_22071,N_19758);
nand UO_1398 (O_1398,N_19846,N_21213);
nor UO_1399 (O_1399,N_19404,N_23249);
or UO_1400 (O_1400,N_22561,N_21611);
nor UO_1401 (O_1401,N_23975,N_20184);
nor UO_1402 (O_1402,N_20464,N_19319);
and UO_1403 (O_1403,N_22597,N_20426);
and UO_1404 (O_1404,N_19198,N_20583);
nand UO_1405 (O_1405,N_21506,N_24362);
and UO_1406 (O_1406,N_20989,N_24584);
nand UO_1407 (O_1407,N_24364,N_20213);
nand UO_1408 (O_1408,N_21535,N_21160);
nand UO_1409 (O_1409,N_20172,N_20512);
and UO_1410 (O_1410,N_23101,N_22269);
nand UO_1411 (O_1411,N_24212,N_21701);
nand UO_1412 (O_1412,N_23406,N_19317);
or UO_1413 (O_1413,N_22973,N_21518);
and UO_1414 (O_1414,N_19504,N_20894);
nor UO_1415 (O_1415,N_23057,N_19969);
or UO_1416 (O_1416,N_23740,N_19775);
xnor UO_1417 (O_1417,N_24650,N_20650);
and UO_1418 (O_1418,N_24859,N_22694);
or UO_1419 (O_1419,N_20453,N_24673);
nand UO_1420 (O_1420,N_20300,N_24693);
xnor UO_1421 (O_1421,N_23124,N_22041);
or UO_1422 (O_1422,N_22975,N_20429);
nand UO_1423 (O_1423,N_24758,N_21719);
or UO_1424 (O_1424,N_24353,N_21178);
and UO_1425 (O_1425,N_24093,N_23849);
or UO_1426 (O_1426,N_22315,N_24463);
nor UO_1427 (O_1427,N_20190,N_22371);
nor UO_1428 (O_1428,N_21392,N_20482);
nor UO_1429 (O_1429,N_20970,N_19301);
nor UO_1430 (O_1430,N_19971,N_24016);
nand UO_1431 (O_1431,N_19976,N_21123);
or UO_1432 (O_1432,N_21245,N_23052);
and UO_1433 (O_1433,N_21745,N_18989);
or UO_1434 (O_1434,N_20356,N_24914);
nand UO_1435 (O_1435,N_19913,N_24240);
or UO_1436 (O_1436,N_19274,N_19261);
nand UO_1437 (O_1437,N_24878,N_18895);
and UO_1438 (O_1438,N_19393,N_21461);
nor UO_1439 (O_1439,N_19995,N_20864);
nand UO_1440 (O_1440,N_21218,N_23927);
nor UO_1441 (O_1441,N_23221,N_19559);
nand UO_1442 (O_1442,N_22109,N_24500);
and UO_1443 (O_1443,N_21676,N_24132);
nand UO_1444 (O_1444,N_24743,N_21189);
nor UO_1445 (O_1445,N_23727,N_20334);
and UO_1446 (O_1446,N_24104,N_24821);
nand UO_1447 (O_1447,N_20454,N_24426);
nand UO_1448 (O_1448,N_24790,N_23750);
or UO_1449 (O_1449,N_22495,N_20182);
and UO_1450 (O_1450,N_19994,N_22027);
nor UO_1451 (O_1451,N_20294,N_18891);
or UO_1452 (O_1452,N_20558,N_19717);
or UO_1453 (O_1453,N_23584,N_18789);
nand UO_1454 (O_1454,N_24299,N_22730);
nor UO_1455 (O_1455,N_20132,N_21030);
and UO_1456 (O_1456,N_20994,N_23198);
nor UO_1457 (O_1457,N_21315,N_20243);
nor UO_1458 (O_1458,N_20536,N_21532);
xnor UO_1459 (O_1459,N_20480,N_19007);
nor UO_1460 (O_1460,N_18843,N_21180);
nand UO_1461 (O_1461,N_22165,N_23144);
and UO_1462 (O_1462,N_23988,N_18770);
nor UO_1463 (O_1463,N_22445,N_22250);
or UO_1464 (O_1464,N_23957,N_19978);
and UO_1465 (O_1465,N_20208,N_24443);
nand UO_1466 (O_1466,N_19796,N_19167);
and UO_1467 (O_1467,N_24050,N_21406);
nor UO_1468 (O_1468,N_21652,N_24599);
nand UO_1469 (O_1469,N_20915,N_19197);
or UO_1470 (O_1470,N_19170,N_21493);
and UO_1471 (O_1471,N_24469,N_24215);
nor UO_1472 (O_1472,N_20019,N_24595);
and UO_1473 (O_1473,N_22916,N_22663);
and UO_1474 (O_1474,N_21682,N_19723);
nand UO_1475 (O_1475,N_21436,N_23299);
and UO_1476 (O_1476,N_21378,N_19329);
or UO_1477 (O_1477,N_18803,N_24760);
and UO_1478 (O_1478,N_22271,N_20835);
and UO_1479 (O_1479,N_20658,N_24235);
nor UO_1480 (O_1480,N_19229,N_21257);
and UO_1481 (O_1481,N_20341,N_21905);
or UO_1482 (O_1482,N_21223,N_19783);
or UO_1483 (O_1483,N_20999,N_21588);
and UO_1484 (O_1484,N_22521,N_21840);
and UO_1485 (O_1485,N_23601,N_24005);
nand UO_1486 (O_1486,N_24467,N_22614);
or UO_1487 (O_1487,N_22291,N_21753);
or UO_1488 (O_1488,N_20303,N_20976);
nand UO_1489 (O_1489,N_22386,N_24061);
nand UO_1490 (O_1490,N_18977,N_21865);
or UO_1491 (O_1491,N_20632,N_21818);
and UO_1492 (O_1492,N_20131,N_21861);
and UO_1493 (O_1493,N_24676,N_18842);
xnor UO_1494 (O_1494,N_22540,N_21208);
nor UO_1495 (O_1495,N_24365,N_23185);
or UO_1496 (O_1496,N_24407,N_21681);
and UO_1497 (O_1497,N_21446,N_18982);
or UO_1498 (O_1498,N_18904,N_20472);
or UO_1499 (O_1499,N_22213,N_22721);
xor UO_1500 (O_1500,N_23269,N_19778);
nor UO_1501 (O_1501,N_22166,N_24934);
xor UO_1502 (O_1502,N_24048,N_21724);
nand UO_1503 (O_1503,N_21174,N_22713);
and UO_1504 (O_1504,N_23357,N_20623);
and UO_1505 (O_1505,N_24334,N_24979);
nor UO_1506 (O_1506,N_21079,N_23891);
nor UO_1507 (O_1507,N_22767,N_24954);
or UO_1508 (O_1508,N_24649,N_19833);
nand UO_1509 (O_1509,N_20050,N_24092);
nand UO_1510 (O_1510,N_18908,N_22346);
nand UO_1511 (O_1511,N_20287,N_21772);
and UO_1512 (O_1512,N_21095,N_19602);
and UO_1513 (O_1513,N_22800,N_22330);
and UO_1514 (O_1514,N_22551,N_22364);
or UO_1515 (O_1515,N_19211,N_22417);
and UO_1516 (O_1516,N_24335,N_24915);
nor UO_1517 (O_1517,N_23479,N_22745);
nand UO_1518 (O_1518,N_19724,N_20548);
or UO_1519 (O_1519,N_20961,N_23659);
nor UO_1520 (O_1520,N_20313,N_20427);
or UO_1521 (O_1521,N_21058,N_22822);
or UO_1522 (O_1522,N_19546,N_20753);
and UO_1523 (O_1523,N_18759,N_19930);
and UO_1524 (O_1524,N_22076,N_23679);
nor UO_1525 (O_1525,N_20611,N_21592);
nand UO_1526 (O_1526,N_19897,N_23449);
nor UO_1527 (O_1527,N_20487,N_21747);
nand UO_1528 (O_1528,N_20383,N_18808);
xor UO_1529 (O_1529,N_21164,N_20821);
xnor UO_1530 (O_1530,N_20546,N_22675);
nand UO_1531 (O_1531,N_20939,N_19230);
nor UO_1532 (O_1532,N_23762,N_23616);
or UO_1533 (O_1533,N_24066,N_23329);
or UO_1534 (O_1534,N_20565,N_22205);
and UO_1535 (O_1535,N_21670,N_21416);
nand UO_1536 (O_1536,N_19515,N_20352);
nor UO_1537 (O_1537,N_19718,N_18828);
or UO_1538 (O_1538,N_21051,N_19516);
nor UO_1539 (O_1539,N_20763,N_21964);
nor UO_1540 (O_1540,N_23278,N_23214);
nand UO_1541 (O_1541,N_23243,N_19868);
and UO_1542 (O_1542,N_20278,N_23578);
or UO_1543 (O_1543,N_21186,N_22222);
nor UO_1544 (O_1544,N_22934,N_20067);
or UO_1545 (O_1545,N_21176,N_20185);
or UO_1546 (O_1546,N_22414,N_18974);
xnor UO_1547 (O_1547,N_23593,N_23745);
xor UO_1548 (O_1548,N_21077,N_23053);
nand UO_1549 (O_1549,N_24938,N_23037);
nor UO_1550 (O_1550,N_20029,N_19187);
or UO_1551 (O_1551,N_20951,N_20783);
nand UO_1552 (O_1552,N_19058,N_22729);
nand UO_1553 (O_1553,N_21762,N_18879);
nand UO_1554 (O_1554,N_21683,N_19234);
or UO_1555 (O_1555,N_20589,N_21113);
xor UO_1556 (O_1556,N_19916,N_22920);
or UO_1557 (O_1557,N_19912,N_23286);
xnor UO_1558 (O_1558,N_18751,N_24017);
and UO_1559 (O_1559,N_22514,N_20017);
nand UO_1560 (O_1560,N_19061,N_19218);
nor UO_1561 (O_1561,N_23906,N_20280);
nor UO_1562 (O_1562,N_20836,N_23175);
or UO_1563 (O_1563,N_22306,N_23967);
xor UO_1564 (O_1564,N_20927,N_20249);
nand UO_1565 (O_1565,N_24482,N_20345);
or UO_1566 (O_1566,N_18834,N_24069);
nor UO_1567 (O_1567,N_23307,N_22048);
nand UO_1568 (O_1568,N_23970,N_20094);
and UO_1569 (O_1569,N_24290,N_19708);
nand UO_1570 (O_1570,N_21851,N_24057);
or UO_1571 (O_1571,N_23993,N_23135);
xnor UO_1572 (O_1572,N_22837,N_22585);
nand UO_1573 (O_1573,N_21664,N_21931);
or UO_1574 (O_1574,N_24793,N_19662);
and UO_1575 (O_1575,N_24882,N_20282);
nand UO_1576 (O_1576,N_19097,N_20962);
nor UO_1577 (O_1577,N_20405,N_19196);
or UO_1578 (O_1578,N_20651,N_21020);
and UO_1579 (O_1579,N_21293,N_20799);
nand UO_1580 (O_1580,N_20810,N_21709);
and UO_1581 (O_1581,N_19542,N_21153);
xnor UO_1582 (O_1582,N_24655,N_18841);
nor UO_1583 (O_1583,N_23757,N_21811);
nor UO_1584 (O_1584,N_24165,N_24487);
nand UO_1585 (O_1585,N_23092,N_19990);
nor UO_1586 (O_1586,N_20251,N_24766);
or UO_1587 (O_1587,N_21910,N_21119);
and UO_1588 (O_1588,N_21360,N_20051);
or UO_1589 (O_1589,N_21804,N_19625);
nor UO_1590 (O_1590,N_20673,N_20850);
or UO_1591 (O_1591,N_19732,N_23189);
nand UO_1592 (O_1592,N_22798,N_24425);
or UO_1593 (O_1593,N_20181,N_19595);
and UO_1594 (O_1594,N_24773,N_23859);
nand UO_1595 (O_1595,N_20948,N_24677);
nand UO_1596 (O_1596,N_24262,N_23382);
or UO_1597 (O_1597,N_21419,N_19966);
nor UO_1598 (O_1598,N_20917,N_19685);
nand UO_1599 (O_1599,N_23385,N_24136);
nand UO_1600 (O_1600,N_20913,N_21963);
and UO_1601 (O_1601,N_21728,N_23702);
or UO_1602 (O_1602,N_22040,N_20417);
nand UO_1603 (O_1603,N_21491,N_23543);
and UO_1604 (O_1604,N_19200,N_23476);
or UO_1605 (O_1605,N_24652,N_20813);
and UO_1606 (O_1606,N_22657,N_23339);
xnor UO_1607 (O_1607,N_23613,N_21003);
nand UO_1608 (O_1608,N_23442,N_21026);
xnor UO_1609 (O_1609,N_24781,N_19263);
nor UO_1610 (O_1610,N_20021,N_23276);
nor UO_1611 (O_1611,N_21966,N_19872);
or UO_1612 (O_1612,N_20015,N_20655);
nor UO_1613 (O_1613,N_24830,N_24468);
and UO_1614 (O_1614,N_23707,N_23623);
and UO_1615 (O_1615,N_20563,N_23071);
nand UO_1616 (O_1616,N_23866,N_24480);
or UO_1617 (O_1617,N_22857,N_19874);
and UO_1618 (O_1618,N_19524,N_19635);
nand UO_1619 (O_1619,N_23588,N_23305);
or UO_1620 (O_1620,N_23017,N_23942);
and UO_1621 (O_1621,N_22544,N_19956);
nand UO_1622 (O_1622,N_21647,N_24142);
and UO_1623 (O_1623,N_19879,N_23743);
nor UO_1624 (O_1624,N_20490,N_24982);
nand UO_1625 (O_1625,N_19166,N_23607);
and UO_1626 (O_1626,N_22622,N_22932);
and UO_1627 (O_1627,N_22145,N_22610);
xor UO_1628 (O_1628,N_24605,N_22744);
nand UO_1629 (O_1629,N_19101,N_21965);
xnor UO_1630 (O_1630,N_21484,N_24933);
nor UO_1631 (O_1631,N_19315,N_23338);
nor UO_1632 (O_1632,N_24631,N_21609);
nand UO_1633 (O_1633,N_24503,N_22270);
nor UO_1634 (O_1634,N_22556,N_22517);
xnor UO_1635 (O_1635,N_23997,N_20065);
or UO_1636 (O_1636,N_24779,N_21061);
and UO_1637 (O_1637,N_23125,N_20972);
nor UO_1638 (O_1638,N_22832,N_20476);
xor UO_1639 (O_1639,N_24889,N_24696);
nor UO_1640 (O_1640,N_23935,N_21912);
nor UO_1641 (O_1641,N_23573,N_21007);
and UO_1642 (O_1642,N_19735,N_24025);
and UO_1643 (O_1643,N_21290,N_24820);
nand UO_1644 (O_1644,N_20177,N_23463);
nor UO_1645 (O_1645,N_18998,N_20958);
nand UO_1646 (O_1646,N_23746,N_23016);
or UO_1647 (O_1647,N_23450,N_21713);
nand UO_1648 (O_1648,N_21070,N_20606);
nand UO_1649 (O_1649,N_23091,N_18978);
or UO_1650 (O_1650,N_21102,N_21704);
nor UO_1651 (O_1651,N_24321,N_18799);
nor UO_1652 (O_1652,N_22925,N_20710);
xor UO_1653 (O_1653,N_19296,N_22087);
or UO_1654 (O_1654,N_22140,N_23137);
nor UO_1655 (O_1655,N_20030,N_20097);
and UO_1656 (O_1656,N_24917,N_20318);
nand UO_1657 (O_1657,N_20840,N_24018);
and UO_1658 (O_1658,N_24537,N_19360);
or UO_1659 (O_1659,N_22423,N_23669);
and UO_1660 (O_1660,N_24199,N_22150);
nand UO_1661 (O_1661,N_19873,N_20828);
and UO_1662 (O_1662,N_23705,N_21782);
nor UO_1663 (O_1663,N_23219,N_20522);
nand UO_1664 (O_1664,N_19318,N_23973);
nor UO_1665 (O_1665,N_21288,N_20643);
xor UO_1666 (O_1666,N_20616,N_23653);
and UO_1667 (O_1667,N_19302,N_19669);
nor UO_1668 (O_1668,N_24370,N_20242);
nor UO_1669 (O_1669,N_22107,N_20873);
and UO_1670 (O_1670,N_23116,N_20008);
nand UO_1671 (O_1671,N_19415,N_19233);
nor UO_1672 (O_1672,N_19138,N_22738);
nor UO_1673 (O_1673,N_18775,N_23327);
nand UO_1674 (O_1674,N_21847,N_24835);
and UO_1675 (O_1675,N_19445,N_23164);
and UO_1676 (O_1676,N_23063,N_24454);
nor UO_1677 (O_1677,N_22253,N_22193);
and UO_1678 (O_1678,N_24645,N_20016);
nor UO_1679 (O_1679,N_22924,N_22929);
or UO_1680 (O_1680,N_23654,N_23661);
xor UO_1681 (O_1681,N_21190,N_21299);
nand UO_1682 (O_1682,N_20814,N_19270);
and UO_1683 (O_1683,N_19915,N_23022);
nand UO_1684 (O_1684,N_21665,N_22871);
xor UO_1685 (O_1685,N_24266,N_22968);
nand UO_1686 (O_1686,N_18985,N_19632);
nor UO_1687 (O_1687,N_19026,N_22619);
nand UO_1688 (O_1688,N_20140,N_19192);
or UO_1689 (O_1689,N_21014,N_23915);
or UO_1690 (O_1690,N_22628,N_20652);
xnor UO_1691 (O_1691,N_21661,N_19836);
and UO_1692 (O_1692,N_24653,N_22121);
nor UO_1693 (O_1693,N_24703,N_23290);
nand UO_1694 (O_1694,N_23119,N_20796);
nor UO_1695 (O_1695,N_24583,N_23824);
and UO_1696 (O_1696,N_24347,N_22834);
nor UO_1697 (O_1697,N_22209,N_19038);
and UO_1698 (O_1698,N_22826,N_23909);
nor UO_1699 (O_1699,N_24174,N_19021);
nor UO_1700 (O_1700,N_20823,N_23898);
nor UO_1701 (O_1701,N_21940,N_19767);
nand UO_1702 (O_1702,N_24864,N_20153);
nand UO_1703 (O_1703,N_20988,N_19800);
nor UO_1704 (O_1704,N_20155,N_22770);
or UO_1705 (O_1705,N_24849,N_20071);
xor UO_1706 (O_1706,N_21116,N_24978);
and UO_1707 (O_1707,N_24713,N_21354);
nand UO_1708 (O_1708,N_24860,N_23166);
nand UO_1709 (O_1709,N_24465,N_24706);
and UO_1710 (O_1710,N_21464,N_21188);
nor UO_1711 (O_1711,N_21056,N_19860);
or UO_1712 (O_1712,N_23505,N_24716);
nor UO_1713 (O_1713,N_20014,N_21977);
or UO_1714 (O_1714,N_24568,N_20229);
xor UO_1715 (O_1715,N_21675,N_20435);
nand UO_1716 (O_1716,N_24160,N_21445);
nor UO_1717 (O_1717,N_23179,N_22683);
nor UO_1718 (O_1718,N_20276,N_24125);
or UO_1719 (O_1719,N_19311,N_19832);
nand UO_1720 (O_1720,N_18874,N_24433);
xor UO_1721 (O_1721,N_24633,N_24442);
nor UO_1722 (O_1722,N_19670,N_20141);
nor UO_1723 (O_1723,N_22028,N_23257);
xnor UO_1724 (O_1724,N_23953,N_20154);
nor UO_1725 (O_1725,N_23381,N_21615);
and UO_1726 (O_1726,N_22717,N_23801);
and UO_1727 (O_1727,N_22863,N_21978);
xor UO_1728 (O_1728,N_19022,N_21167);
nand UO_1729 (O_1729,N_23918,N_22536);
and UO_1730 (O_1730,N_23816,N_22031);
and UO_1731 (O_1731,N_23529,N_24090);
and UO_1732 (O_1732,N_22901,N_24004);
and UO_1733 (O_1733,N_23121,N_18951);
nand UO_1734 (O_1734,N_20507,N_21421);
xnor UO_1735 (O_1735,N_19952,N_22896);
or UO_1736 (O_1736,N_18878,N_22624);
nor UO_1737 (O_1737,N_22720,N_22776);
or UO_1738 (O_1738,N_21523,N_21430);
nor UO_1739 (O_1739,N_23493,N_20120);
xnor UO_1740 (O_1740,N_22870,N_19722);
nor UO_1741 (O_1741,N_23517,N_23958);
nor UO_1742 (O_1742,N_24533,N_19802);
and UO_1743 (O_1743,N_22368,N_19454);
or UO_1744 (O_1744,N_21768,N_20811);
and UO_1745 (O_1745,N_22966,N_20351);
or UO_1746 (O_1746,N_19804,N_22399);
or UO_1747 (O_1747,N_20901,N_23349);
and UO_1748 (O_1748,N_22555,N_23217);
nand UO_1749 (O_1749,N_20694,N_21626);
or UO_1750 (O_1750,N_24171,N_22928);
or UO_1751 (O_1751,N_23846,N_22931);
xor UO_1752 (O_1752,N_21684,N_22308);
and UO_1753 (O_1753,N_21265,N_21571);
nand UO_1754 (O_1754,N_24515,N_18849);
and UO_1755 (O_1755,N_21031,N_24947);
or UO_1756 (O_1756,N_23431,N_22402);
or UO_1757 (O_1757,N_19631,N_24958);
or UO_1758 (O_1758,N_22158,N_21453);
nand UO_1759 (O_1759,N_21552,N_21597);
xnor UO_1760 (O_1760,N_21714,N_19577);
nand UO_1761 (O_1761,N_19071,N_18867);
nand UO_1762 (O_1762,N_21021,N_20119);
and UO_1763 (O_1763,N_20035,N_23002);
nand UO_1764 (O_1764,N_19118,N_23062);
or UO_1765 (O_1765,N_20186,N_21756);
nor UO_1766 (O_1766,N_24718,N_23190);
or UO_1767 (O_1767,N_20511,N_20446);
and UO_1768 (O_1768,N_23503,N_24923);
nand UO_1769 (O_1769,N_21710,N_24249);
nand UO_1770 (O_1770,N_21468,N_23461);
nand UO_1771 (O_1771,N_23504,N_23156);
nand UO_1772 (O_1772,N_21881,N_19158);
or UO_1773 (O_1773,N_19691,N_21669);
or UO_1774 (O_1774,N_22753,N_19461);
and UO_1775 (O_1775,N_20268,N_23054);
and UO_1776 (O_1776,N_20246,N_21583);
nor UO_1777 (O_1777,N_20847,N_21524);
nand UO_1778 (O_1778,N_19397,N_24823);
or UO_1779 (O_1779,N_22875,N_19706);
nor UO_1780 (O_1780,N_21136,N_20918);
nor UO_1781 (O_1781,N_21100,N_22327);
nor UO_1782 (O_1782,N_24339,N_19248);
or UO_1783 (O_1783,N_22882,N_20298);
xnor UO_1784 (O_1784,N_23949,N_22030);
nor UO_1785 (O_1785,N_22051,N_22737);
nor UO_1786 (O_1786,N_22481,N_19483);
xnor UO_1787 (O_1787,N_20198,N_23391);
or UO_1788 (O_1788,N_24390,N_23006);
nor UO_1789 (O_1789,N_22635,N_22180);
or UO_1790 (O_1790,N_23454,N_19077);
or UO_1791 (O_1791,N_22332,N_20750);
or UO_1792 (O_1792,N_24479,N_24701);
or UO_1793 (O_1793,N_21897,N_24925);
and UO_1794 (O_1794,N_19283,N_22232);
and UO_1795 (O_1795,N_20368,N_20497);
and UO_1796 (O_1796,N_21303,N_22994);
nor UO_1797 (O_1797,N_19232,N_23820);
nand UO_1798 (O_1798,N_24149,N_21259);
nor UO_1799 (O_1799,N_20225,N_21340);
nand UO_1800 (O_1800,N_22061,N_20689);
nor UO_1801 (O_1801,N_21232,N_23014);
and UO_1802 (O_1802,N_20797,N_23317);
nor UO_1803 (O_1803,N_22477,N_21598);
nor UO_1804 (O_1804,N_24916,N_22037);
nand UO_1805 (O_1805,N_22768,N_20232);
nand UO_1806 (O_1806,N_21743,N_20969);
nand UO_1807 (O_1807,N_23247,N_21631);
or UO_1808 (O_1808,N_20025,N_22455);
or UO_1809 (O_1809,N_21412,N_22173);
nor UO_1810 (O_1810,N_24168,N_19247);
nor UO_1811 (O_1811,N_23560,N_19855);
and UO_1812 (O_1812,N_22756,N_22865);
xor UO_1813 (O_1813,N_21690,N_19673);
nand UO_1814 (O_1814,N_23000,N_23488);
nor UO_1815 (O_1815,N_23963,N_23823);
and UO_1816 (O_1816,N_23363,N_20428);
nor UO_1817 (O_1817,N_20418,N_18975);
and UO_1818 (O_1818,N_22642,N_22235);
xnor UO_1819 (O_1819,N_22086,N_24727);
or UO_1820 (O_1820,N_19638,N_22296);
nor UO_1821 (O_1821,N_20742,N_24472);
or UO_1822 (O_1822,N_24656,N_24112);
or UO_1823 (O_1823,N_19375,N_22050);
nor UO_1824 (O_1824,N_23497,N_21780);
and UO_1825 (O_1825,N_21913,N_20319);
nor UO_1826 (O_1826,N_23139,N_24295);
xnor UO_1827 (O_1827,N_22956,N_22190);
nand UO_1828 (O_1828,N_23865,N_23632);
or UO_1829 (O_1829,N_21096,N_19188);
nand UO_1830 (O_1830,N_24858,N_21956);
nor UO_1831 (O_1831,N_22335,N_24640);
and UO_1832 (O_1832,N_24848,N_20705);
xnor UO_1833 (O_1833,N_23513,N_19219);
nor UO_1834 (O_1834,N_23346,N_23452);
xor UO_1835 (O_1835,N_20121,N_21486);
nor UO_1836 (O_1836,N_21287,N_23182);
nor UO_1837 (O_1837,N_18965,N_19114);
or UO_1838 (O_1838,N_23916,N_18935);
and UO_1839 (O_1839,N_22793,N_19310);
nand UO_1840 (O_1840,N_24138,N_22357);
nor UO_1841 (O_1841,N_23194,N_23483);
nand UO_1842 (O_1842,N_22633,N_24288);
nor UO_1843 (O_1843,N_24067,N_21087);
nand UO_1844 (O_1844,N_19422,N_24707);
nand UO_1845 (O_1845,N_21814,N_21952);
nand UO_1846 (O_1846,N_23675,N_23834);
and UO_1847 (O_1847,N_19540,N_21580);
and UO_1848 (O_1848,N_22056,N_22015);
and UO_1849 (O_1849,N_24736,N_24175);
and UO_1850 (O_1850,N_20089,N_23657);
nor UO_1851 (O_1851,N_23244,N_19769);
nor UO_1852 (O_1852,N_19529,N_19282);
nor UO_1853 (O_1853,N_23469,N_20086);
and UO_1854 (O_1854,N_22204,N_24358);
and UO_1855 (O_1855,N_21739,N_22649);
and UO_1856 (O_1856,N_19193,N_21715);
nand UO_1857 (O_1857,N_20451,N_22955);
nor UO_1858 (O_1858,N_22067,N_23591);
and UO_1859 (O_1859,N_22442,N_24242);
and UO_1860 (O_1860,N_22318,N_23544);
xnor UO_1861 (O_1861,N_19068,N_20587);
nand UO_1862 (O_1862,N_19142,N_21118);
nand UO_1863 (O_1863,N_22498,N_20921);
nor UO_1864 (O_1864,N_19997,N_21088);
xnor UO_1865 (O_1865,N_24214,N_22017);
nand UO_1866 (O_1866,N_19931,N_20887);
or UO_1867 (O_1867,N_24184,N_24031);
or UO_1868 (O_1868,N_24891,N_24322);
nand UO_1869 (O_1869,N_21049,N_23744);
nand UO_1870 (O_1870,N_22942,N_21649);
nor UO_1871 (O_1871,N_20263,N_19940);
or UO_1872 (O_1872,N_24948,N_23735);
nand UO_1873 (O_1873,N_19550,N_19345);
or UO_1874 (O_1874,N_21168,N_21610);
nor UO_1875 (O_1875,N_22456,N_19584);
nor UO_1876 (O_1876,N_20306,N_22486);
nand UO_1877 (O_1877,N_24569,N_21579);
nor UO_1878 (O_1878,N_20629,N_18955);
nand UO_1879 (O_1879,N_22362,N_22999);
nor UO_1880 (O_1880,N_21331,N_21383);
and UO_1881 (O_1881,N_19420,N_20060);
nand UO_1882 (O_1882,N_18861,N_24929);
and UO_1883 (O_1883,N_20863,N_20407);
nand UO_1884 (O_1884,N_22348,N_23519);
and UO_1885 (O_1885,N_21028,N_20936);
nor UO_1886 (O_1886,N_21172,N_19288);
and UO_1887 (O_1887,N_22953,N_23397);
nor UO_1888 (O_1888,N_21495,N_22387);
nand UO_1889 (O_1889,N_18901,N_19782);
or UO_1890 (O_1890,N_23879,N_19352);
or UO_1891 (O_1891,N_24787,N_24753);
and UO_1892 (O_1892,N_21311,N_24260);
nor UO_1893 (O_1893,N_21271,N_21273);
nand UO_1894 (O_1894,N_21514,N_23076);
and UO_1895 (O_1895,N_23093,N_20588);
nand UO_1896 (O_1896,N_22493,N_24412);
nand UO_1897 (O_1897,N_22792,N_22568);
nand UO_1898 (O_1898,N_22571,N_22719);
nand UO_1899 (O_1899,N_22215,N_22429);
or UO_1900 (O_1900,N_19508,N_21339);
nor UO_1901 (O_1901,N_24002,N_23791);
xnor UO_1902 (O_1902,N_19251,N_19309);
nand UO_1903 (O_1903,N_22608,N_18793);
or UO_1904 (O_1904,N_21748,N_20791);
nand UO_1905 (O_1905,N_20421,N_22480);
xor UO_1906 (O_1906,N_20716,N_20150);
nand UO_1907 (O_1907,N_23026,N_24873);
and UO_1908 (O_1908,N_20082,N_24789);
or UO_1909 (O_1909,N_24012,N_20191);
nand UO_1910 (O_1910,N_20667,N_23571);
nor UO_1911 (O_1911,N_23542,N_23919);
nor UO_1912 (O_1912,N_19367,N_18945);
xnor UO_1913 (O_1913,N_21255,N_23845);
xnor UO_1914 (O_1914,N_24340,N_22584);
nand UO_1915 (O_1915,N_21707,N_21159);
nand UO_1916 (O_1916,N_18827,N_24778);
or UO_1917 (O_1917,N_23356,N_22948);
nor UO_1918 (O_1918,N_20817,N_23873);
or UO_1919 (O_1919,N_18971,N_18818);
nor UO_1920 (O_1920,N_24361,N_21928);
nor UO_1921 (O_1921,N_23265,N_19497);
and UO_1922 (O_1922,N_20070,N_23496);
nor UO_1923 (O_1923,N_21643,N_19474);
and UO_1924 (O_1924,N_24556,N_24530);
nor UO_1925 (O_1925,N_21877,N_24078);
or UO_1926 (O_1926,N_22309,N_24841);
nor UO_1927 (O_1927,N_22126,N_22936);
and UO_1928 (O_1928,N_19303,N_23811);
xnor UO_1929 (O_1929,N_22773,N_23481);
or UO_1930 (O_1930,N_23795,N_20808);
nor UO_1931 (O_1931,N_24812,N_24689);
nor UO_1932 (O_1932,N_23340,N_23872);
and UO_1933 (O_1933,N_22200,N_21774);
nor UO_1934 (O_1934,N_23706,N_22949);
nand UO_1935 (O_1935,N_21957,N_23287);
or UO_1936 (O_1936,N_21117,N_24899);
nand UO_1937 (O_1937,N_21200,N_24421);
nand UO_1938 (O_1938,N_18948,N_21097);
nor UO_1939 (O_1939,N_22961,N_19469);
and UO_1940 (O_1940,N_24342,N_19597);
and UO_1941 (O_1941,N_24294,N_24196);
and UO_1942 (O_1942,N_22207,N_21637);
nand UO_1943 (O_1943,N_20250,N_19690);
and UO_1944 (O_1944,N_24601,N_19771);
or UO_1945 (O_1945,N_24279,N_20100);
nand UO_1946 (O_1946,N_23437,N_23223);
nor UO_1947 (O_1947,N_23403,N_24902);
nand UO_1948 (O_1948,N_21564,N_24099);
nor UO_1949 (O_1949,N_19073,N_21509);
xor UO_1950 (O_1950,N_22659,N_23805);
and UO_1951 (O_1951,N_24492,N_21038);
or UO_1952 (O_1952,N_20107,N_22895);
nand UO_1953 (O_1953,N_22154,N_22078);
or UO_1954 (O_1954,N_24872,N_19958);
xor UO_1955 (O_1955,N_20302,N_24221);
nand UO_1956 (O_1956,N_21238,N_23563);
and UO_1957 (O_1957,N_24618,N_20227);
or UO_1958 (O_1958,N_23123,N_24567);
nand UO_1959 (O_1959,N_24491,N_23887);
and UO_1960 (O_1960,N_21141,N_21279);
nor UO_1961 (O_1961,N_23473,N_24945);
or UO_1962 (O_1962,N_23283,N_23703);
nand UO_1963 (O_1963,N_19451,N_24134);
nand UO_1964 (O_1964,N_19807,N_21376);
and UO_1965 (O_1965,N_21282,N_21184);
and UO_1966 (O_1966,N_22664,N_19440);
or UO_1967 (O_1967,N_21640,N_23188);
nor UO_1968 (O_1968,N_24903,N_19060);
and UO_1969 (O_1969,N_20573,N_22280);
and UO_1970 (O_1970,N_22700,N_24263);
or UO_1971 (O_1971,N_23955,N_21986);
and UO_1972 (O_1972,N_24552,N_20166);
nor UO_1973 (O_1973,N_23902,N_18898);
nor UO_1974 (O_1974,N_19623,N_21161);
nand UO_1975 (O_1975,N_20649,N_22878);
and UO_1976 (O_1976,N_24133,N_19030);
xnor UO_1977 (O_1977,N_19613,N_23541);
and UO_1978 (O_1978,N_21624,N_20782);
or UO_1979 (O_1979,N_21657,N_21260);
or UO_1980 (O_1980,N_23417,N_22138);
nor UO_1981 (O_1981,N_23281,N_22967);
nor UO_1982 (O_1982,N_24855,N_22747);
and UO_1983 (O_1983,N_24672,N_23416);
and UO_1984 (O_1984,N_19476,N_24560);
nor UO_1985 (O_1985,N_23895,N_18870);
or UO_1986 (O_1986,N_22326,N_19513);
and UO_1987 (O_1987,N_24350,N_23267);
nand UO_1988 (O_1988,N_19278,N_19828);
nor UO_1989 (O_1989,N_19955,N_20586);
nor UO_1990 (O_1990,N_24922,N_23284);
nor UO_1991 (O_1991,N_19779,N_22807);
and UO_1992 (O_1992,N_21319,N_21650);
xnor UO_1993 (O_1993,N_24115,N_24338);
nor UO_1994 (O_1994,N_24894,N_22345);
nor UO_1995 (O_1995,N_23199,N_23344);
nor UO_1996 (O_1996,N_24088,N_20564);
or UO_1997 (O_1997,N_24037,N_22671);
or UO_1998 (O_1998,N_22312,N_23238);
or UO_1999 (O_1999,N_24141,N_23151);
or UO_2000 (O_2000,N_24730,N_20353);
xor UO_2001 (O_2001,N_24085,N_20896);
or UO_2002 (O_2002,N_22211,N_19791);
or UO_2003 (O_2003,N_23402,N_21086);
xnor UO_2004 (O_2004,N_21368,N_18854);
and UO_2005 (O_2005,N_24123,N_20460);
nor UO_2006 (O_2006,N_20264,N_21428);
and UO_2007 (O_2007,N_20662,N_24201);
and UO_2008 (O_2008,N_19687,N_24478);
xor UO_2009 (O_2009,N_22407,N_24909);
xor UO_2010 (O_2010,N_19159,N_23429);
or UO_2011 (O_2011,N_22112,N_24510);
nand UO_2012 (O_2012,N_22202,N_21805);
nand UO_2013 (O_2013,N_22491,N_21540);
nor UO_2014 (O_2014,N_21974,N_24151);
or UO_2015 (O_2015,N_23719,N_23728);
or UO_2016 (O_2016,N_19875,N_19046);
nor UO_2017 (O_2017,N_20640,N_24278);
and UO_2018 (O_2018,N_22373,N_23869);
and UO_2019 (O_2019,N_19204,N_23631);
and UO_2020 (O_2020,N_23427,N_23089);
and UO_2021 (O_2021,N_23952,N_23018);
nor UO_2022 (O_2022,N_19489,N_22338);
nand UO_2023 (O_2023,N_19259,N_24006);
and UO_2024 (O_2024,N_24592,N_24411);
xnor UO_2025 (O_2025,N_19742,N_24126);
nand UO_2026 (O_2026,N_24038,N_19954);
nand UO_2027 (O_2027,N_21867,N_23943);
and UO_2028 (O_2028,N_22337,N_20195);
and UO_2029 (O_2029,N_23126,N_20663);
and UO_2030 (O_2030,N_20018,N_24990);
and UO_2031 (O_2031,N_19699,N_19581);
or UO_2032 (O_2032,N_18976,N_21787);
or UO_2033 (O_2033,N_19039,N_19332);
and UO_2034 (O_2034,N_18928,N_21567);
or UO_2035 (O_2035,N_23335,N_20504);
or UO_2036 (O_2036,N_20245,N_24851);
nand UO_2037 (O_2037,N_21367,N_20639);
nor UO_2038 (O_2038,N_24119,N_19004);
nor UO_2039 (O_2039,N_23775,N_23671);
or UO_2040 (O_2040,N_19749,N_22115);
and UO_2041 (O_2041,N_23246,N_24504);
or UO_2042 (O_2042,N_21678,N_23738);
or UO_2043 (O_2043,N_21346,N_24071);
and UO_2044 (O_2044,N_24404,N_20197);
or UO_2045 (O_2045,N_21057,N_23328);
nand UO_2046 (O_2046,N_19293,N_21938);
xor UO_2047 (O_2047,N_20375,N_23695);
nor UO_2048 (O_2048,N_23242,N_23374);
nand UO_2049 (O_2049,N_22024,N_22191);
nand UO_2050 (O_2050,N_23145,N_22163);
nor UO_2051 (O_2051,N_19172,N_20964);
nor UO_2052 (O_2052,N_21338,N_23758);
or UO_2053 (O_2053,N_22353,N_20374);
and UO_2054 (O_2054,N_20739,N_20858);
and UO_2055 (O_2055,N_24824,N_19216);
or UO_2056 (O_2056,N_20477,N_19112);
or UO_2057 (O_2057,N_19185,N_20101);
nor UO_2058 (O_2058,N_21623,N_21220);
or UO_2059 (O_2059,N_22960,N_21198);
and UO_2060 (O_2060,N_21833,N_24297);
and UO_2061 (O_2061,N_22842,N_24573);
nor UO_2062 (O_2062,N_20600,N_24540);
or UO_2063 (O_2063,N_22528,N_24566);
or UO_2064 (O_2064,N_19867,N_22908);
nand UO_2065 (O_2065,N_23950,N_20046);
or UO_2066 (O_2066,N_23711,N_24035);
and UO_2067 (O_2067,N_20312,N_20236);
nand UO_2068 (O_2068,N_19616,N_20681);
nor UO_2069 (O_2069,N_23337,N_24800);
or UO_2070 (O_2070,N_23163,N_24439);
or UO_2071 (O_2071,N_22796,N_19815);
nand UO_2072 (O_2072,N_19243,N_18758);
nor UO_2073 (O_2073,N_21807,N_24705);
nor UO_2074 (O_2074,N_23769,N_20215);
and UO_2075 (O_2075,N_22299,N_19134);
and UO_2076 (O_2076,N_21276,N_18997);
and UO_2077 (O_2077,N_23040,N_20036);
nor UO_2078 (O_2078,N_20931,N_19761);
nor UO_2079 (O_2079,N_24337,N_24157);
or UO_2080 (O_2080,N_24470,N_19195);
nand UO_2081 (O_2081,N_23435,N_21899);
nor UO_2082 (O_2082,N_24323,N_20301);
and UO_2083 (O_2083,N_20740,N_20470);
nor UO_2084 (O_2084,N_24441,N_22403);
nand UO_2085 (O_2085,N_20728,N_22188);
xnor UO_2086 (O_2086,N_20108,N_21427);
nand UO_2087 (O_2087,N_23070,N_21733);
nor UO_2088 (O_2088,N_21084,N_20449);
nor UO_2089 (O_2089,N_21244,N_23047);
xor UO_2090 (O_2090,N_19964,N_23749);
nand UO_2091 (O_2091,N_20699,N_20110);
or UO_2092 (O_2092,N_20392,N_19628);
and UO_2093 (O_2093,N_22349,N_21308);
nor UO_2094 (O_2094,N_19525,N_21758);
nor UO_2095 (O_2095,N_23502,N_19544);
and UO_2096 (O_2096,N_21872,N_21698);
nor UO_2097 (O_2097,N_24764,N_19672);
or UO_2098 (O_2098,N_20980,N_22114);
or UO_2099 (O_2099,N_24211,N_23100);
nor UO_2100 (O_2100,N_23297,N_20787);
nor UO_2101 (O_2101,N_22746,N_20798);
nor UO_2102 (O_2102,N_22436,N_23096);
nand UO_2103 (O_2103,N_22926,N_19124);
or UO_2104 (O_2104,N_24122,N_23809);
nand UO_2105 (O_2105,N_21823,N_24741);
and UO_2106 (O_2106,N_24816,N_21983);
nand UO_2107 (O_2107,N_22457,N_19353);
or UO_2108 (O_2108,N_23827,N_19016);
and UO_2109 (O_2109,N_23099,N_19099);
or UO_2110 (O_2110,N_23525,N_24847);
nor UO_2111 (O_2111,N_23617,N_20330);
nor UO_2112 (O_2112,N_23216,N_23920);
and UO_2113 (O_2113,N_22876,N_21137);
and UO_2114 (O_2114,N_23682,N_19677);
and UO_2115 (O_2115,N_21384,N_21614);
nor UO_2116 (O_2116,N_24780,N_19105);
and UO_2117 (O_2117,N_20862,N_24797);
xor UO_2118 (O_2118,N_19294,N_22708);
nand UO_2119 (O_2119,N_22325,N_22704);
nand UO_2120 (O_2120,N_21667,N_18804);
or UO_2121 (O_2121,N_20818,N_24170);
and UO_2122 (O_2122,N_20943,N_23688);
and UO_2123 (O_2123,N_19561,N_22255);
and UO_2124 (O_2124,N_24507,N_20950);
nand UO_2125 (O_2125,N_24826,N_20680);
nand UO_2126 (O_2126,N_22489,N_19028);
xnor UO_2127 (O_2127,N_21072,N_24307);
nand UO_2128 (O_2128,N_23875,N_24783);
nand UO_2129 (O_2129,N_20781,N_21181);
nand UO_2130 (O_2130,N_19102,N_24887);
xor UO_2131 (O_2131,N_20743,N_22026);
and UO_2132 (O_2132,N_22784,N_19563);
or UO_2133 (O_2133,N_22083,N_22718);
nand UO_2134 (O_2134,N_24523,N_20849);
or UO_2135 (O_2135,N_20907,N_21817);
and UO_2136 (O_2136,N_21696,N_24869);
or UO_2137 (O_2137,N_21776,N_23752);
or UO_2138 (O_2138,N_24318,N_21332);
or UO_2139 (O_2139,N_19989,N_24267);
nor UO_2140 (O_2140,N_22273,N_19089);
xor UO_2141 (O_2141,N_20712,N_20188);
xor UO_2142 (O_2142,N_20096,N_23660);
nor UO_2143 (O_2143,N_21799,N_20759);
nor UO_2144 (O_2144,N_24415,N_22988);
xnor UO_2145 (O_2145,N_24076,N_21869);
nand UO_2146 (O_2146,N_20756,N_21062);
nand UO_2147 (O_2147,N_23510,N_20038);
nand UO_2148 (O_2148,N_24382,N_22133);
nand UO_2149 (O_2149,N_18949,N_21324);
nor UO_2150 (O_2150,N_24111,N_24545);
nor UO_2151 (O_2151,N_19961,N_23085);
xor UO_2152 (O_2152,N_23153,N_19155);
or UO_2153 (O_2153,N_20777,N_21476);
or UO_2154 (O_2154,N_20469,N_22460);
xnor UO_2155 (O_2155,N_24324,N_21801);
xnor UO_2156 (O_2156,N_19354,N_23478);
nand UO_2157 (O_2157,N_24993,N_20111);
nor UO_2158 (O_2158,N_21663,N_21846);
or UO_2159 (O_2159,N_22836,N_20878);
nor UO_2160 (O_2160,N_19585,N_21473);
or UO_2161 (O_2161,N_21466,N_19575);
and UO_2162 (O_2162,N_18987,N_22989);
nand UO_2163 (O_2163,N_22263,N_24754);
xnor UO_2164 (O_2164,N_24113,N_20566);
nor UO_2165 (O_2165,N_20780,N_21046);
xnor UO_2166 (O_2166,N_24275,N_24543);
nand UO_2167 (O_2167,N_22075,N_22234);
and UO_2168 (O_2168,N_21995,N_23272);
nor UO_2169 (O_2169,N_20771,N_24256);
and UO_2170 (O_2170,N_24548,N_19378);
xor UO_2171 (O_2171,N_23712,N_21437);
nand UO_2172 (O_2172,N_23501,N_24385);
nor UO_2173 (O_2173,N_24516,N_21792);
nand UO_2174 (O_2174,N_20621,N_20163);
nand UO_2175 (O_2175,N_24354,N_21085);
xnor UO_2176 (O_2176,N_22577,N_22095);
and UO_2177 (O_2177,N_22433,N_22687);
nor UO_2178 (O_2178,N_19499,N_19695);
and UO_2179 (O_2179,N_20200,N_24609);
nor UO_2180 (O_2180,N_21616,N_24300);
nand UO_2181 (O_2181,N_24430,N_22676);
and UO_2182 (O_2182,N_20395,N_21382);
and UO_2183 (O_2183,N_24304,N_20678);
or UO_2184 (O_2184,N_22602,N_24130);
and UO_2185 (O_2185,N_20795,N_21169);
and UO_2186 (O_2186,N_19799,N_21016);
nor UO_2187 (O_2187,N_19754,N_20765);
or UO_2188 (O_2188,N_20059,N_22631);
and UO_2189 (O_2189,N_20443,N_22900);
or UO_2190 (O_2190,N_21958,N_21764);
nand UO_2191 (O_2191,N_20724,N_23535);
xnor UO_2192 (O_2192,N_23011,N_21629);
or UO_2193 (O_2193,N_24898,N_24056);
or UO_2194 (O_2194,N_20484,N_19494);
and UO_2195 (O_2195,N_21133,N_21330);
or UO_2196 (O_2196,N_22391,N_20267);
and UO_2197 (O_2197,N_20502,N_18932);
and UO_2198 (O_2198,N_23132,N_23944);
or UO_2199 (O_2199,N_21836,N_24888);
nand UO_2200 (O_2200,N_23404,N_19281);
and UO_2201 (O_2201,N_22065,N_23923);
nor UO_2202 (O_2202,N_20042,N_19827);
nand UO_2203 (O_2203,N_24617,N_24268);
nand UO_2204 (O_2204,N_22740,N_20672);
or UO_2205 (O_2205,N_19972,N_22018);
nor UO_2206 (O_2206,N_23697,N_21467);
xnor UO_2207 (O_2207,N_20538,N_20884);
or UO_2208 (O_2208,N_24588,N_19619);
nand UO_2209 (O_2209,N_24866,N_21691);
nand UO_2210 (O_2210,N_18848,N_21292);
xor UO_2211 (O_2211,N_21090,N_24838);
or UO_2212 (O_2212,N_23874,N_19304);
or UO_2213 (O_2213,N_22902,N_23112);
xor UO_2214 (O_2214,N_22552,N_23778);
nand UO_2215 (O_2215,N_21006,N_22772);
nor UO_2216 (O_2216,N_23621,N_21385);
nand UO_2217 (O_2217,N_24000,N_20924);
or UO_2218 (O_2218,N_19942,N_22983);
and UO_2219 (O_2219,N_22393,N_20462);
xor UO_2220 (O_2220,N_19122,N_21418);
nor UO_2221 (O_2221,N_22912,N_19999);
and UO_2222 (O_2222,N_23830,N_23347);
nand UO_2223 (O_2223,N_21130,N_19419);
nor UO_2224 (O_2224,N_20769,N_20314);
or UO_2225 (O_2225,N_23405,N_23250);
or UO_2226 (O_2226,N_21635,N_24302);
nor UO_2227 (O_2227,N_24163,N_22236);
xnor UO_2228 (O_2228,N_24436,N_24559);
nor UO_2229 (O_2229,N_24657,N_21499);
nor UO_2230 (O_2230,N_21404,N_21318);
nor UO_2231 (O_2231,N_19705,N_20293);
nor UO_2232 (O_2232,N_21914,N_21771);
xnor UO_2233 (O_2233,N_24876,N_23546);
or UO_2234 (O_2234,N_19983,N_21760);
or UO_2235 (O_2235,N_24623,N_23015);
nand UO_2236 (O_2236,N_18795,N_22905);
and UO_2237 (O_2237,N_23191,N_21578);
xnor UO_2238 (O_2238,N_24803,N_21236);
nand UO_2239 (O_2239,N_20520,N_20076);
nand UO_2240 (O_2240,N_22282,N_22658);
nand UO_2241 (O_2241,N_23829,N_24518);
nand UO_2242 (O_2242,N_21907,N_20668);
nand UO_2243 (O_2243,N_23590,N_21945);
and UO_2244 (O_2244,N_23624,N_23019);
and UO_2245 (O_2245,N_23309,N_22231);
and UO_2246 (O_2246,N_21309,N_23742);
nor UO_2247 (O_2247,N_24455,N_21142);
nand UO_2248 (O_2248,N_24775,N_24593);
and UO_2249 (O_2249,N_20767,N_21291);
nor UO_2250 (O_2250,N_21866,N_22887);
and UO_2251 (O_2251,N_21551,N_22911);
xnor UO_2252 (O_2252,N_22415,N_23562);
nor UO_2253 (O_2253,N_22160,N_23559);
and UO_2254 (O_2254,N_22463,N_21825);
and UO_2255 (O_2255,N_24448,N_18866);
or UO_2256 (O_2256,N_21944,N_19920);
nor UO_2257 (O_2257,N_18821,N_19917);
nand UO_2258 (O_2258,N_20982,N_20954);
xor UO_2259 (O_2259,N_22764,N_18968);
nand UO_2260 (O_2260,N_24671,N_24292);
or UO_2261 (O_2261,N_20063,N_23797);
nand UO_2262 (O_2262,N_24200,N_20321);
and UO_2263 (O_2263,N_20220,N_23857);
nor UO_2264 (O_2264,N_24193,N_20720);
nor UO_2265 (O_2265,N_19923,N_24589);
nand UO_2266 (O_2266,N_18991,N_22376);
and UO_2267 (O_2267,N_24555,N_19665);
or UO_2268 (O_2268,N_24486,N_19667);
and UO_2269 (O_2269,N_24905,N_24194);
and UO_2270 (O_2270,N_21247,N_21793);
nand UO_2271 (O_2271,N_22569,N_21256);
nor UO_2272 (O_2272,N_23687,N_20423);
xnor UO_2273 (O_2273,N_21350,N_21602);
nand UO_2274 (O_2274,N_21538,N_23852);
nor UO_2275 (O_2275,N_20381,N_24629);
and UO_2276 (O_2276,N_23948,N_19617);
or UO_2277 (O_2277,N_20779,N_23838);
nor UO_2278 (O_2278,N_20644,N_22016);
nand UO_2279 (O_2279,N_21960,N_21505);
and UO_2280 (O_2280,N_19104,N_22897);
nor UO_2281 (O_2281,N_24401,N_20995);
and UO_2282 (O_2282,N_20261,N_20940);
nor UO_2283 (O_2283,N_20247,N_22268);
nand UO_2284 (O_2284,N_24508,N_19881);
nor UO_2285 (O_2285,N_24959,N_22785);
xor UO_2286 (O_2286,N_20130,N_20834);
or UO_2287 (O_2287,N_22124,N_20285);
nand UO_2288 (O_2288,N_22933,N_21336);
nand UO_2289 (O_2289,N_21820,N_19391);
or UO_2290 (O_2290,N_20053,N_18774);
and UO_2291 (O_2291,N_19704,N_21568);
nand UO_2292 (O_2292,N_24735,N_24188);
or UO_2293 (O_2293,N_22110,N_24258);
nor UO_2294 (O_2294,N_19413,N_21941);
and UO_2295 (O_2295,N_24868,N_20959);
or UO_2296 (O_2296,N_21812,N_19090);
and UO_2297 (O_2297,N_22644,N_23594);
or UO_2298 (O_2298,N_23484,N_21327);
or UO_2299 (O_2299,N_23606,N_21503);
and UO_2300 (O_2300,N_23718,N_23370);
or UO_2301 (O_2301,N_19701,N_22825);
xnor UO_2302 (O_2302,N_23154,N_21620);
or UO_2303 (O_2303,N_21953,N_20577);
nand UO_2304 (O_2304,N_20315,N_21796);
nor UO_2305 (O_2305,N_21982,N_24143);
nand UO_2306 (O_2306,N_19047,N_20923);
nor UO_2307 (O_2307,N_20058,N_20235);
nor UO_2308 (O_2308,N_20359,N_23641);
and UO_2309 (O_2309,N_23540,N_21757);
and UO_2310 (O_2310,N_19280,N_24666);
nor UO_2311 (O_2311,N_20691,N_18856);
or UO_2312 (O_2312,N_18958,N_21950);
nor UO_2313 (O_2313,N_20199,N_22613);
or UO_2314 (O_2314,N_24146,N_21930);
nor UO_2315 (O_2315,N_18933,N_22530);
or UO_2316 (O_2316,N_22322,N_24326);
or UO_2317 (O_2317,N_19037,N_23195);
and UO_2318 (O_2318,N_24145,N_19333);
nor UO_2319 (O_2319,N_19910,N_24377);
or UO_2320 (O_2320,N_24227,N_21674);
nand UO_2321 (O_2321,N_23334,N_19323);
xor UO_2322 (O_2322,N_22462,N_19324);
or UO_2323 (O_2323,N_22992,N_24786);
xor UO_2324 (O_2324,N_22907,N_21534);
xnor UO_2325 (O_2325,N_21358,N_21359);
xor UO_2326 (O_2326,N_20871,N_20822);
nand UO_2327 (O_2327,N_23930,N_21439);
nor UO_2328 (O_2328,N_19591,N_19327);
and UO_2329 (O_2329,N_22279,N_24811);
xor UO_2330 (O_2330,N_23609,N_21755);
nor UO_2331 (O_2331,N_23065,N_19817);
or UO_2332 (O_2332,N_21685,N_19447);
and UO_2333 (O_2333,N_22748,N_20741);
nor UO_2334 (O_2334,N_19331,N_19753);
nand UO_2335 (O_2335,N_24400,N_20493);
nand UO_2336 (O_2336,N_24837,N_23293);
or UO_2337 (O_2337,N_20540,N_22815);
xnor UO_2338 (O_2338,N_22574,N_23279);
and UO_2339 (O_2339,N_22290,N_20893);
and UO_2340 (O_2340,N_19436,N_22506);
and UO_2341 (O_2341,N_23345,N_24293);
or UO_2342 (O_2342,N_22148,N_23934);
and UO_2343 (O_2343,N_21828,N_21157);
nand UO_2344 (O_2344,N_19745,N_20204);
xnor UO_2345 (O_2345,N_21932,N_19869);
and UO_2346 (O_2346,N_21605,N_24642);
nor UO_2347 (O_2347,N_19067,N_21711);
and UO_2348 (O_2348,N_20433,N_19123);
nand UO_2349 (O_2349,N_20932,N_23168);
and UO_2350 (O_2350,N_22971,N_19854);
or UO_2351 (O_2351,N_24501,N_19825);
or UO_2352 (O_2352,N_24939,N_22630);
nor UO_2353 (O_2353,N_23736,N_23423);
or UO_2354 (O_2354,N_20079,N_22267);
and UO_2355 (O_2355,N_20501,N_21011);
or UO_2356 (O_2356,N_24632,N_23438);
nor UO_2357 (O_2357,N_22343,N_22690);
nand UO_2358 (O_2358,N_21050,N_20555);
or UO_2359 (O_2359,N_22420,N_21746);
or UO_2360 (O_2360,N_20009,N_21998);
nor UO_2361 (O_2361,N_22972,N_20291);
nor UO_2362 (O_2362,N_19901,N_22419);
or UO_2363 (O_2363,N_21175,N_20595);
nand UO_2364 (O_2364,N_20604,N_20631);
xnor UO_2365 (O_2365,N_24535,N_21996);
xnor UO_2366 (O_2366,N_21231,N_24646);
and UO_2367 (O_2367,N_23985,N_20037);
and UO_2368 (O_2368,N_20515,N_19605);
or UO_2369 (O_2369,N_22240,N_21553);
nor UO_2370 (O_2370,N_20579,N_24674);
and UO_2371 (O_2371,N_20952,N_20906);
nor UO_2372 (O_2372,N_23005,N_19075);
xor UO_2373 (O_2373,N_24313,N_23428);
or UO_2374 (O_2374,N_23177,N_22797);
or UO_2375 (O_2375,N_22846,N_21387);
or UO_2376 (O_2376,N_19180,N_23174);
nand UO_2377 (O_2377,N_20492,N_22244);
nor UO_2378 (O_2378,N_20209,N_23822);
nand UO_2379 (O_2379,N_19970,N_24429);
and UO_2380 (O_2380,N_22440,N_24785);
nand UO_2381 (O_2381,N_24968,N_21364);
nand UO_2382 (O_2382,N_24298,N_24036);
or UO_2383 (O_2383,N_20785,N_19611);
and UO_2384 (O_2384,N_22101,N_21612);
or UO_2385 (O_2385,N_19168,N_23486);
nor UO_2386 (O_2386,N_21112,N_22545);
nand UO_2387 (O_2387,N_23547,N_21316);
xor UO_2388 (O_2388,N_21328,N_22760);
or UO_2389 (O_2389,N_19944,N_24852);
nand UO_2390 (O_2390,N_24834,N_21044);
and UO_2391 (O_2391,N_19231,N_21954);
or UO_2392 (O_2392,N_19941,N_23029);
nor UO_2393 (O_2393,N_21732,N_21922);
or UO_2394 (O_2394,N_20975,N_24844);
xnor UO_2395 (O_2395,N_21882,N_20124);
nand UO_2396 (O_2396,N_24822,N_23892);
and UO_2397 (O_2397,N_18779,N_23325);
nor UO_2398 (O_2398,N_22534,N_21477);
or UO_2399 (O_2399,N_21441,N_20615);
nand UO_2400 (O_2400,N_23589,N_20648);
and UO_2401 (O_2401,N_23414,N_21280);
nor UO_2402 (O_2402,N_21154,N_24086);
nand UO_2403 (O_2403,N_19372,N_19441);
and UO_2404 (O_2404,N_21407,N_20510);
nand UO_2405 (O_2405,N_23087,N_20657);
and UO_2406 (O_2406,N_21770,N_20448);
or UO_2407 (O_2407,N_22599,N_19610);
nor UO_2408 (O_2408,N_23568,N_21754);
nor UO_2409 (O_2409,N_20539,N_19998);
xor UO_2410 (O_2410,N_21150,N_19864);
or UO_2411 (O_2411,N_21001,N_21045);
nand UO_2412 (O_2412,N_23748,N_20270);
nand UO_2413 (O_2413,N_20123,N_23083);
or UO_2414 (O_2414,N_22724,N_24245);
or UO_2415 (O_2415,N_21688,N_20485);
nand UO_2416 (O_2416,N_21196,N_18942);
nor UO_2417 (O_2417,N_22066,N_22446);
or UO_2418 (O_2418,N_24836,N_23979);
and UO_2419 (O_2419,N_22791,N_20105);
or UO_2420 (O_2420,N_23619,N_21919);
and UO_2421 (O_2421,N_24372,N_22607);
xnor UO_2422 (O_2422,N_20717,N_21887);
nor UO_2423 (O_2423,N_24622,N_18922);
and UO_2424 (O_2424,N_24667,N_20031);
nor UO_2425 (O_2425,N_18772,N_19526);
xnor UO_2426 (O_2426,N_22412,N_19686);
nor UO_2427 (O_2427,N_20370,N_23491);
nor UO_2428 (O_2428,N_19949,N_22853);
or UO_2429 (O_2429,N_23760,N_24984);
nand UO_2430 (O_2430,N_23353,N_24541);
nand UO_2431 (O_2431,N_23113,N_19006);
or UO_2432 (O_2432,N_23318,N_19119);
nand UO_2433 (O_2433,N_22548,N_22840);
nor UO_2434 (O_2434,N_22206,N_23847);
nand UO_2435 (O_2435,N_22276,N_23236);
nand UO_2436 (O_2436,N_21935,N_19981);
nand UO_2437 (O_2437,N_19878,N_18957);
or UO_2438 (O_2438,N_19468,N_19169);
or UO_2439 (O_2439,N_23672,N_23023);
nor UO_2440 (O_2440,N_22508,N_22425);
and UO_2441 (O_2441,N_23045,N_20080);
nor UO_2442 (O_2442,N_20128,N_19174);
or UO_2443 (O_2443,N_19287,N_22937);
nand UO_2444 (O_2444,N_20391,N_20567);
nor UO_2445 (O_2445,N_23012,N_24955);
or UO_2446 (O_2446,N_22958,N_21808);
or UO_2447 (O_2447,N_23576,N_19837);
or UO_2448 (O_2448,N_21193,N_19925);
or UO_2449 (O_2449,N_24427,N_23799);
or UO_2450 (O_2450,N_20679,N_23832);
or UO_2451 (O_2451,N_20272,N_19633);
and UO_2452 (O_2452,N_22829,N_22485);
or UO_2453 (O_2453,N_19573,N_24748);
and UO_2454 (O_2454,N_23201,N_21222);
and UO_2455 (O_2455,N_20113,N_24710);
or UO_2456 (O_2456,N_23516,N_19403);
and UO_2457 (O_2457,N_19927,N_22889);
xnor UO_2458 (O_2458,N_19453,N_23572);
or UO_2459 (O_2459,N_19129,N_22593);
or UO_2460 (O_2460,N_23425,N_24329);
and UO_2461 (O_2461,N_20256,N_19945);
and UO_2462 (O_2462,N_22504,N_20508);
nor UO_2463 (O_2463,N_22079,N_20963);
xor UO_2464 (O_2464,N_21069,N_21267);
nand UO_2465 (O_2465,N_19649,N_22539);
nand UO_2466 (O_2466,N_24558,N_21082);
xnor UO_2467 (O_2467,N_21179,N_23673);
and UO_2468 (O_2468,N_19374,N_22564);
nor UO_2469 (O_2469,N_20203,N_24935);
nor UO_2470 (O_2470,N_23232,N_23021);
or UO_2471 (O_2471,N_24881,N_23884);
nor UO_2472 (O_2472,N_20118,N_21366);
nor UO_2473 (O_2473,N_19127,N_20083);
nand UO_2474 (O_2474,N_20669,N_22186);
nor UO_2475 (O_2475,N_23971,N_23814);
and UO_2476 (O_2476,N_18750,N_19694);
or UO_2477 (O_2477,N_24801,N_23618);
and UO_2478 (O_2478,N_23871,N_20612);
nand UO_2479 (O_2479,N_21634,N_19136);
and UO_2480 (O_2480,N_24722,N_20829);
and UO_2481 (O_2481,N_24434,N_18972);
xor UO_2482 (O_2482,N_23813,N_21883);
and UO_2483 (O_2483,N_24217,N_23007);
or UO_2484 (O_2484,N_20104,N_19626);
or UO_2485 (O_2485,N_20288,N_21660);
nor UO_2486 (O_2486,N_22127,N_19697);
and UO_2487 (O_2487,N_24691,N_19096);
xor UO_2488 (O_2488,N_19693,N_23462);
nor UO_2489 (O_2489,N_19604,N_19648);
and UO_2490 (O_2490,N_20892,N_21052);
or UO_2491 (O_2491,N_23386,N_20390);
xnor UO_2492 (O_2492,N_23724,N_20752);
and UO_2493 (O_2493,N_24637,N_22667);
and UO_2494 (O_2494,N_22366,N_22643);
or UO_2495 (O_2495,N_23913,N_19588);
nand UO_2496 (O_2496,N_22170,N_24118);
nand UO_2497 (O_2497,N_18916,N_22666);
nor UO_2498 (O_2498,N_19045,N_22781);
nor UO_2499 (O_2499,N_23600,N_22008);
or UO_2500 (O_2500,N_21549,N_22258);
or UO_2501 (O_2501,N_19072,N_21845);
nor UO_2502 (O_2502,N_22576,N_20533);
nor UO_2503 (O_2503,N_23277,N_24522);
nor UO_2504 (O_2504,N_21478,N_22558);
nor UO_2505 (O_2505,N_19444,N_21171);
and UO_2506 (O_2506,N_20968,N_19395);
nand UO_2507 (O_2507,N_19905,N_19019);
and UO_2508 (O_2508,N_22223,N_24311);
nor UO_2509 (O_2509,N_24586,N_22295);
nand UO_2510 (O_2510,N_20992,N_19892);
and UO_2511 (O_2511,N_24833,N_20024);
or UO_2512 (O_2512,N_20365,N_18792);
nand UO_2513 (O_2513,N_19719,N_19009);
nand UO_2514 (O_2514,N_23789,N_24428);
xnor UO_2515 (O_2515,N_20257,N_21529);
nand UO_2516 (O_2516,N_21569,N_22788);
xor UO_2517 (O_2517,N_23361,N_18765);
and UO_2518 (O_2518,N_20746,N_22866);
nand UO_2519 (O_2519,N_18943,N_20205);
nand UO_2520 (O_2520,N_23620,N_21401);
and UO_2521 (O_2521,N_21205,N_19043);
and UO_2522 (O_2522,N_20706,N_20165);
nor UO_2523 (O_2523,N_24580,N_20474);
xnor UO_2524 (O_2524,N_22214,N_18936);
and UO_2525 (O_2525,N_23082,N_19051);
nand UO_2526 (O_2526,N_20499,N_23171);
nand UO_2527 (O_2527,N_22437,N_23844);
or UO_2528 (O_2528,N_20842,N_22525);
or UO_2529 (O_2529,N_21894,N_23464);
or UO_2530 (O_2530,N_23443,N_20342);
or UO_2531 (O_2531,N_22993,N_18900);
nand UO_2532 (O_2532,N_22242,N_22135);
nand UO_2533 (O_2533,N_21185,N_23575);
nand UO_2534 (O_2534,N_24759,N_24752);
nor UO_2535 (O_2535,N_21246,N_24616);
nand UO_2536 (O_2536,N_21975,N_23793);
or UO_2537 (O_2537,N_24702,N_24664);
nand UO_2538 (O_2538,N_19057,N_24325);
xnor UO_2539 (O_2539,N_20946,N_20459);
xnor UO_2540 (O_2540,N_24871,N_19810);
or UO_2541 (O_2541,N_22891,N_19459);
or UO_2542 (O_2542,N_21570,N_23907);
and UO_2543 (O_2543,N_22592,N_21731);
xnor UO_2544 (O_2544,N_21576,N_24976);
xnor UO_2545 (O_2545,N_24437,N_18819);
or UO_2546 (O_2546,N_19922,N_21397);
nand UO_2547 (O_2547,N_24222,N_20748);
or UO_2548 (O_2548,N_23998,N_23316);
nor UO_2549 (O_2549,N_23130,N_22612);
nor UO_2550 (O_2550,N_20701,N_19592);
nand UO_2551 (O_2551,N_23904,N_19713);
or UO_2552 (O_2552,N_22567,N_22149);
nor UO_2553 (O_2553,N_19448,N_23785);
nand UO_2554 (O_2554,N_21492,N_19502);
or UO_2555 (O_2555,N_19380,N_19737);
or UO_2556 (O_2556,N_19655,N_19040);
and UO_2557 (O_2557,N_21470,N_19150);
nand UO_2558 (O_2558,N_20645,N_21824);
and UO_2559 (O_2559,N_21393,N_20590);
and UO_2560 (O_2560,N_22699,N_24420);
nand UO_2561 (O_2561,N_23259,N_23937);
nand UO_2562 (O_2562,N_22311,N_19008);
xor UO_2563 (O_2563,N_20491,N_24156);
nand UO_2564 (O_2564,N_20666,N_18805);
and UO_2565 (O_2565,N_20275,N_19203);
or UO_2566 (O_2566,N_24453,N_21269);
xnor UO_2567 (O_2567,N_23192,N_21039);
and UO_2568 (O_2568,N_23628,N_22297);
nand UO_2569 (O_2569,N_24746,N_22848);
nand UO_2570 (O_2570,N_22922,N_19091);
nor UO_2571 (O_2571,N_20034,N_19906);
or UO_2572 (O_2572,N_22401,N_21374);
nand UO_2573 (O_2573,N_19569,N_18994);
nand UO_2574 (O_2574,N_20608,N_22229);
or UO_2575 (O_2575,N_20523,N_19620);
and UO_2576 (O_2576,N_19659,N_24996);
or UO_2577 (O_2577,N_19834,N_19839);
and UO_2578 (O_2578,N_22301,N_19179);
nand UO_2579 (O_2579,N_21474,N_23815);
or UO_2580 (O_2580,N_21203,N_23783);
nand UO_2581 (O_2581,N_24856,N_19885);
nand UO_2582 (O_2582,N_22727,N_20005);
nand UO_2583 (O_2583,N_22422,N_24550);
or UO_2584 (O_2584,N_19716,N_23313);
or UO_2585 (O_2585,N_23843,N_21148);
and UO_2586 (O_2586,N_19866,N_19651);
nor UO_2587 (O_2587,N_22142,N_23196);
nand UO_2588 (O_2588,N_23073,N_22578);
xor UO_2589 (O_2589,N_24273,N_24376);
and UO_2590 (O_2590,N_19947,N_24489);
nand UO_2591 (O_2591,N_19083,N_19291);
nor UO_2592 (O_2592,N_19366,N_23480);
or UO_2593 (O_2593,N_20802,N_20286);
xor UO_2594 (O_2594,N_24765,N_21485);
or UO_2595 (O_2595,N_20399,N_23274);
or UO_2596 (O_2596,N_20707,N_21741);
nand UO_2597 (O_2597,N_22042,N_19549);
nor UO_2598 (O_2598,N_23102,N_23285);
and UO_2599 (O_2599,N_24857,N_24272);
nor UO_2600 (O_2600,N_22970,N_24791);
or UO_2601 (O_2601,N_24106,N_21342);
xnor UO_2602 (O_2602,N_24203,N_21806);
nand UO_2603 (O_2603,N_24685,N_22636);
or UO_2604 (O_2604,N_24102,N_20040);
nor UO_2605 (O_2605,N_21530,N_21687);
or UO_2606 (O_2606,N_22930,N_20984);
nand UO_2607 (O_2607,N_22354,N_21192);
nand UO_2608 (O_2608,N_23725,N_23929);
and UO_2609 (O_2609,N_23094,N_21921);
nand UO_2610 (O_2610,N_24658,N_19887);
and UO_2611 (O_2611,N_24206,N_19552);
and UO_2612 (O_2612,N_19503,N_20997);
or UO_2613 (O_2613,N_20736,N_19244);
and UO_2614 (O_2614,N_19603,N_19852);
and UO_2615 (O_2615,N_21314,N_24063);
nand UO_2616 (O_2616,N_20580,N_23890);
nand UO_2617 (O_2617,N_19676,N_24346);
and UO_2618 (O_2618,N_19759,N_21482);
nor UO_2619 (O_2619,N_19733,N_24536);
xor UO_2620 (O_2620,N_23231,N_22021);
nand UO_2621 (O_2621,N_20925,N_19241);
or UO_2622 (O_2622,N_24108,N_22199);
or UO_2623 (O_2623,N_21870,N_22533);
nor UO_2624 (O_2624,N_19139,N_19470);
nor UO_2625 (O_2625,N_19088,N_18963);
nand UO_2626 (O_2626,N_22195,N_23256);
or UO_2627 (O_2627,N_20223,N_21716);
nor UO_2628 (O_2628,N_24571,N_23310);
xor UO_2629 (O_2629,N_19896,N_20331);
or UO_2630 (O_2630,N_23536,N_20550);
nand UO_2631 (O_2631,N_24387,N_24695);
nor UO_2632 (O_2632,N_22774,N_20244);
and UO_2633 (O_2633,N_20812,N_19843);
nand UO_2634 (O_2634,N_23759,N_24154);
and UO_2635 (O_2635,N_23358,N_24572);
nor UO_2636 (O_2636,N_22812,N_24022);
or UO_2637 (O_2637,N_23251,N_18757);
nand UO_2638 (O_2638,N_23245,N_22884);
and UO_2639 (O_2639,N_23482,N_23709);
or UO_2640 (O_2640,N_18905,N_22164);
nand UO_2641 (O_2641,N_24030,N_19087);
or UO_2642 (O_2642,N_23910,N_18899);
nand UO_2643 (O_2643,N_22707,N_24806);
nor UO_2644 (O_2644,N_20091,N_22143);
and UO_2645 (O_2645,N_20912,N_21369);
xnor UO_2646 (O_2646,N_21219,N_21349);
nor UO_2647 (O_2647,N_23261,N_20000);
and UO_2648 (O_2648,N_19938,N_21990);
and UO_2649 (O_2649,N_22093,N_20239);
nor UO_2650 (O_2650,N_19013,N_23051);
and UO_2651 (O_2651,N_20043,N_19601);
or UO_2652 (O_2652,N_21425,N_22473);
nor UO_2653 (O_2653,N_19768,N_23610);
and UO_2654 (O_2654,N_21413,N_22940);
xor UO_2655 (O_2655,N_19823,N_19335);
and UO_2656 (O_2656,N_21098,N_22011);
nand UO_2657 (O_2657,N_23388,N_24296);
or UO_2658 (O_2658,N_19245,N_21517);
nand UO_2659 (O_2659,N_24980,N_22384);
and UO_2660 (O_2660,N_19152,N_23422);
nor UO_2661 (O_2661,N_23206,N_23766);
and UO_2662 (O_2662,N_18992,N_20387);
nor UO_2663 (O_2663,N_24098,N_19664);
or UO_2664 (O_2664,N_21013,N_19787);
and UO_2665 (O_2665,N_19194,N_20726);
or UO_2666 (O_2666,N_23398,N_23583);
nor UO_2667 (O_2667,N_24192,N_19608);
nor UO_2668 (O_2668,N_23605,N_19519);
xor UO_2669 (O_2669,N_21429,N_20425);
xor UO_2670 (O_2670,N_22119,N_20979);
and UO_2671 (O_2671,N_19720,N_21262);
or UO_2672 (O_2672,N_24424,N_22733);
nor UO_2673 (O_2673,N_21442,N_24250);
nand UO_2674 (O_2674,N_18780,N_23395);
xor UO_2675 (O_2675,N_22025,N_23954);
or UO_2676 (O_2676,N_22946,N_19442);
and UO_2677 (O_2677,N_21132,N_19728);
and UO_2678 (O_2678,N_20775,N_19712);
nor UO_2679 (O_2679,N_23379,N_23262);
nor UO_2680 (O_2680,N_24087,N_22302);
nand UO_2681 (O_2681,N_22985,N_23322);
nand UO_2682 (O_2682,N_21873,N_24475);
nor UO_2683 (O_2683,N_22490,N_23111);
or UO_2684 (O_2684,N_21702,N_24158);
or UO_2685 (O_2685,N_20509,N_24865);
or UO_2686 (O_2686,N_19199,N_22867);
nand UO_2687 (O_2687,N_21479,N_21480);
nor UO_2688 (O_2688,N_21165,N_20087);
nand UO_2689 (O_2689,N_19117,N_20900);
nand UO_2690 (O_2690,N_21313,N_20401);
xnor UO_2691 (O_2691,N_21775,N_24485);
and UO_2692 (O_2692,N_23056,N_21411);
nor UO_2693 (O_2693,N_22950,N_22344);
or UO_2694 (O_2694,N_21906,N_20358);
and UO_2695 (O_2695,N_22147,N_19757);
or UO_2696 (O_2696,N_23732,N_21302);
xnor UO_2697 (O_2697,N_21199,N_23447);
or UO_2698 (O_2698,N_21357,N_22082);
or UO_2699 (O_2699,N_23441,N_19285);
nand UO_2700 (O_2700,N_22380,N_23034);
nand UO_2701 (O_2701,N_19987,N_19266);
or UO_2702 (O_2702,N_24484,N_20292);
or UO_2703 (O_2703,N_24110,N_20323);
or UO_2704 (O_2704,N_24950,N_24621);
xnor UO_2705 (O_2705,N_20179,N_20206);
or UO_2706 (O_2706,N_18970,N_23662);
and UO_2707 (O_2707,N_21968,N_20845);
and UO_2708 (O_2708,N_22864,N_23721);
nor UO_2709 (O_2709,N_20942,N_19545);
and UO_2710 (O_2710,N_19788,N_19600);
or UO_2711 (O_2711,N_23893,N_23134);
and UO_2712 (O_2712,N_19116,N_19565);
or UO_2713 (O_2713,N_18919,N_24799);
nor UO_2714 (O_2714,N_21862,N_19842);
nand UO_2715 (O_2715,N_22850,N_19682);
nor UO_2716 (O_2716,N_22898,N_19452);
nor UO_2717 (O_2717,N_22711,N_23359);
and UO_2718 (O_2718,N_24683,N_23103);
and UO_2719 (O_2719,N_20436,N_23067);
nor UO_2720 (O_2720,N_20990,N_23365);
nand UO_2721 (O_2721,N_19036,N_21969);
nor UO_2722 (O_2722,N_21920,N_19322);
or UO_2723 (O_2723,N_18990,N_21212);
and UO_2724 (O_2724,N_24524,N_21854);
nor UO_2725 (O_2725,N_23972,N_21516);
xor UO_2726 (O_2726,N_24060,N_23209);
xnor UO_2727 (O_2727,N_24531,N_20233);
or UO_2728 (O_2728,N_22328,N_22516);
nor UO_2729 (O_2729,N_21929,N_18764);
or UO_2730 (O_2730,N_22859,N_22134);
and UO_2731 (O_2731,N_19574,N_19844);
xor UO_2732 (O_2732,N_21550,N_19760);
xor UO_2733 (O_2733,N_21073,N_24068);
and UO_2734 (O_2734,N_22416,N_20114);
nand UO_2735 (O_2735,N_23459,N_24432);
nor UO_2736 (O_2736,N_24895,N_23282);
and UO_2737 (O_2737,N_21831,N_20231);
or UO_2738 (O_2738,N_19876,N_20839);
nor UO_2739 (O_2739,N_19012,N_21699);
nor UO_2740 (O_2740,N_23509,N_21284);
or UO_2741 (O_2741,N_21613,N_20620);
nand UO_2742 (O_2742,N_19208,N_24738);
and UO_2743 (O_2743,N_19856,N_21286);
or UO_2744 (O_2744,N_23118,N_24381);
nor UO_2745 (O_2745,N_23947,N_24578);
and UO_2746 (O_2746,N_23424,N_19640);
and UO_2747 (O_2747,N_22340,N_21765);
nor UO_2748 (O_2748,N_23295,N_20092);
nand UO_2749 (O_2749,N_23254,N_19271);
or UO_2750 (O_2750,N_21742,N_20258);
nand UO_2751 (O_2751,N_24999,N_18801);
xor UO_2752 (O_2752,N_24972,N_24208);
and UO_2753 (O_2753,N_20983,N_21234);
nand UO_2754 (O_2754,N_23534,N_19711);
or UO_2755 (O_2755,N_21803,N_24756);
and UO_2756 (O_2756,N_18892,N_20960);
nand UO_2757 (O_2757,N_21590,N_24162);
xnor UO_2758 (O_2758,N_19379,N_23289);
and UO_2759 (O_2759,N_20897,N_24638);
and UO_2760 (O_2760,N_19661,N_19560);
and UO_2761 (O_2761,N_18947,N_18863);
nand UO_2762 (O_2762,N_22497,N_19161);
nor UO_2763 (O_2763,N_21294,N_20397);
or UO_2764 (O_2764,N_22749,N_24532);
or UO_2765 (O_2765,N_22816,N_19063);
and UO_2766 (O_2766,N_18787,N_19822);
nand UO_2767 (O_2767,N_20833,N_24314);
and UO_2768 (O_2768,N_23098,N_24964);
nor UO_2769 (O_2769,N_23467,N_24396);
nor UO_2770 (O_2770,N_22860,N_19480);
nand UO_2771 (O_2771,N_22782,N_19178);
or UO_2772 (O_2772,N_23786,N_22194);
and UO_2773 (O_2773,N_24096,N_22775);
or UO_2774 (O_2774,N_23651,N_20109);
or UO_2775 (O_2775,N_20260,N_21217);
or UO_2776 (O_2776,N_21528,N_19292);
xnor UO_2777 (O_2777,N_22141,N_20057);
nor UO_2778 (O_2778,N_19486,N_20614);
or UO_2779 (O_2779,N_23585,N_22153);
and UO_2780 (O_2780,N_18938,N_23240);
nand UO_2781 (O_2781,N_20930,N_22918);
nor UO_2782 (O_2782,N_20498,N_21022);
and UO_2783 (O_2783,N_24460,N_19738);
nand UO_2784 (O_2784,N_18777,N_21300);
nand UO_2785 (O_2785,N_21242,N_24495);
and UO_2786 (O_2786,N_19772,N_21955);
nand UO_2787 (O_2787,N_21221,N_22716);
nand UO_2788 (O_2788,N_23951,N_22249);
and UO_2789 (O_2789,N_18918,N_18871);
and UO_2790 (O_2790,N_18986,N_18954);
nand UO_2791 (O_2791,N_24517,N_21229);
and UO_2792 (O_2792,N_22589,N_19517);
nor UO_2793 (O_2793,N_19587,N_24191);
nand UO_2794 (O_2794,N_21587,N_20772);
or UO_2795 (O_2795,N_20488,N_21789);
or UO_2796 (O_2796,N_19485,N_23717);
and UO_2797 (O_2797,N_24620,N_19177);
nor UO_2798 (O_2798,N_23183,N_19806);
nand UO_2799 (O_2799,N_23991,N_23921);
xnor UO_2800 (O_2800,N_23162,N_23807);
or UO_2801 (O_2801,N_22835,N_24129);
nor UO_2802 (O_2802,N_22073,N_22656);
nand UO_2803 (O_2803,N_19024,N_20898);
nor UO_2804 (O_2804,N_20879,N_21093);
and UO_2805 (O_2805,N_24839,N_19062);
and UO_2806 (O_2806,N_24539,N_21810);
xor UO_2807 (O_2807,N_21839,N_21002);
and UO_2808 (O_2808,N_20367,N_19076);
nor UO_2809 (O_2809,N_21677,N_23753);
nand UO_2810 (O_2810,N_23275,N_24694);
nor UO_2811 (O_2811,N_20183,N_18884);
and UO_2812 (O_2812,N_19418,N_23715);
nand UO_2813 (O_2813,N_20398,N_18940);
or UO_2814 (O_2814,N_21295,N_21372);
nand UO_2815 (O_2815,N_19986,N_21829);
nand UO_2816 (O_2816,N_20596,N_21122);
nand UO_2817 (O_2817,N_19154,N_21510);
nand UO_2818 (O_2818,N_21508,N_19064);
nor UO_2819 (O_2819,N_24607,N_22703);
nor UO_2820 (O_2820,N_18921,N_19888);
or UO_2821 (O_2821,N_23072,N_23077);
xor UO_2822 (O_2822,N_23683,N_24576);
nand UO_2823 (O_2823,N_20224,N_22004);
or UO_2824 (O_2824,N_23983,N_21399);
or UO_2825 (O_2825,N_21692,N_23552);
and UO_2826 (O_2826,N_20568,N_19553);
and UO_2827 (O_2827,N_20804,N_22927);
and UO_2828 (O_2828,N_22957,N_23108);
nor UO_2829 (O_2829,N_19034,N_23258);
or UO_2830 (O_2830,N_21228,N_20202);
or UO_2831 (O_2831,N_19314,N_23779);
or UO_2832 (O_2832,N_24551,N_19189);
nand UO_2833 (O_2833,N_19725,N_24316);
nor UO_2834 (O_2834,N_23730,N_19430);
nor UO_2835 (O_2835,N_24220,N_24944);
or UO_2836 (O_2836,N_24285,N_19721);
nand UO_2837 (O_2837,N_19298,N_23176);
nand UO_2838 (O_2838,N_21497,N_23506);
nand UO_2839 (O_2839,N_21472,N_20883);
and UO_2840 (O_2840,N_23074,N_22032);
or UO_2841 (O_2841,N_22426,N_23646);
nand UO_2842 (O_2842,N_20757,N_21034);
and UO_2843 (O_2843,N_18835,N_19541);
nand UO_2844 (O_2844,N_23863,N_21000);
nor UO_2845 (O_2845,N_22010,N_19226);
and UO_2846 (O_2846,N_20422,N_21233);
or UO_2847 (O_2847,N_23131,N_24032);
xnor UO_2848 (O_2848,N_22227,N_19487);
nand UO_2849 (O_2849,N_23408,N_23670);
and UO_2850 (O_2850,N_24052,N_19646);
nor UO_2851 (O_2851,N_22000,N_20861);
and UO_2852 (O_2852,N_22809,N_22679);
xor UO_2853 (O_2853,N_19748,N_23565);
or UO_2854 (O_2854,N_22710,N_20420);
or UO_2855 (O_2855,N_22653,N_20634);
nand UO_2856 (O_2856,N_22830,N_19369);
xnor UO_2857 (O_2857,N_21081,N_22294);
and UO_2858 (O_2858,N_20933,N_19564);
or UO_2859 (O_2859,N_19857,N_20479);
or UO_2860 (O_2860,N_23894,N_19898);
nor UO_2861 (O_2861,N_23172,N_23392);
xnor UO_2862 (O_2862,N_20416,N_24897);
and UO_2863 (O_2863,N_20284,N_23204);
nand UO_2864 (O_2864,N_21043,N_20255);
or UO_2865 (O_2865,N_20998,N_22629);
and UO_2866 (O_2866,N_22824,N_21202);
and UO_2867 (O_2867,N_18952,N_24375);
nor UO_2868 (O_2868,N_22638,N_24750);
nor UO_2869 (O_2869,N_21555,N_21875);
or UO_2870 (O_2870,N_23268,N_22464);
nand UO_2871 (O_2871,N_21251,N_22468);
nand UO_2872 (O_2872,N_23960,N_21654);
nand UO_2873 (O_2873,N_21759,N_23640);
and UO_2874 (O_2874,N_22849,N_24757);
and UO_2875 (O_2875,N_20372,N_19432);
nor UO_2876 (O_2876,N_19784,N_24971);
and UO_2877 (O_2877,N_18771,N_22002);
nor UO_2878 (O_2878,N_20991,N_24225);
and UO_2879 (O_2879,N_23489,N_24498);
xnor UO_2880 (O_2880,N_22058,N_21841);
nor UO_2881 (O_2881,N_19049,N_24798);
nand UO_2882 (O_2882,N_23390,N_21278);
xnor UO_2883 (O_2883,N_24893,N_23248);
nand UO_2884 (O_2884,N_24598,N_20764);
nand UO_2885 (O_2885,N_22466,N_19334);
xor UO_2886 (O_2886,N_19786,N_24675);
and UO_2887 (O_2887,N_24965,N_21101);
or UO_2888 (O_2888,N_23850,N_19227);
or UO_2889 (O_2889,N_24913,N_21842);
xor UO_2890 (O_2890,N_22285,N_22218);
and UO_2891 (O_2891,N_22591,N_21581);
nand UO_2892 (O_2892,N_21541,N_23837);
nor UO_2893 (O_2893,N_19181,N_20335);
nor UO_2894 (O_2894,N_24081,N_24332);
and UO_2895 (O_2895,N_23097,N_20928);
xor UO_2896 (O_2896,N_23580,N_23234);
and UO_2897 (O_2897,N_24679,N_19641);
or UO_2898 (O_2898,N_20098,N_22432);
or UO_2899 (O_2899,N_20819,N_19580);
or UO_2900 (O_2900,N_19160,N_22538);
and UO_2901 (O_2901,N_19535,N_21561);
and UO_2902 (O_2902,N_22582,N_22910);
nor UO_2903 (O_2903,N_21241,N_18806);
nor UO_2904 (O_2904,N_21127,N_21285);
nor UO_2905 (O_2905,N_21151,N_20846);
and UO_2906 (O_2906,N_20605,N_19313);
xor UO_2907 (O_2907,N_23867,N_22360);
nor UO_2908 (O_2908,N_22499,N_24883);
or UO_2909 (O_2909,N_23366,N_21729);
nand UO_2910 (O_2910,N_23400,N_24879);
nor UO_2911 (O_2911,N_18929,N_20333);
and UO_2912 (O_2912,N_23377,N_19558);
nand UO_2913 (O_2913,N_24594,N_23708);
nand UO_2914 (O_2914,N_21858,N_22817);
nand UO_2915 (O_2915,N_20636,N_19473);
and UO_2916 (O_2916,N_20888,N_23362);
or UO_2917 (O_2917,N_24912,N_20751);
nand UO_2918 (O_2918,N_21126,N_20337);
or UO_2919 (O_2919,N_20633,N_21844);
xnor UO_2920 (O_2920,N_21645,N_24352);
or UO_2921 (O_2921,N_18911,N_21946);
xor UO_2922 (O_2922,N_23974,N_19272);
and UO_2923 (O_2923,N_22502,N_21798);
or UO_2924 (O_2924,N_19578,N_23439);
nand UO_2925 (O_2925,N_21310,N_20729);
nand UO_2926 (O_2926,N_22888,N_20338);
nor UO_2927 (O_2927,N_22411,N_22100);
nor UO_2928 (O_2928,N_20311,N_21032);
or UO_2929 (O_2929,N_23169,N_21832);
xnor UO_2930 (O_2930,N_24393,N_21981);
and UO_2931 (O_2931,N_21821,N_21139);
xnor UO_2932 (O_2932,N_22660,N_20544);
and UO_2933 (O_2933,N_24721,N_19607);
and UO_2934 (O_2934,N_24011,N_23681);
and UO_2935 (O_2935,N_23001,N_23550);
or UO_2936 (O_2936,N_21909,N_23839);
and UO_2937 (O_2937,N_21800,N_19224);
and UO_2938 (O_2938,N_21386,N_24740);
or UO_2939 (O_2939,N_21572,N_22987);
nand UO_2940 (O_2940,N_23945,N_23897);
and UO_2941 (O_2941,N_24034,N_22689);
nor UO_2942 (O_2942,N_22208,N_20698);
or UO_2943 (O_2943,N_22167,N_24010);
and UO_2944 (O_2944,N_24767,N_22626);
xor UO_2945 (O_2945,N_18753,N_22217);
nand UO_2946 (O_2946,N_22298,N_23411);
and UO_2947 (O_2947,N_19624,N_20458);
nand UO_2948 (O_2948,N_23200,N_20977);
xnor UO_2949 (O_2949,N_19337,N_19209);
or UO_2950 (O_2950,N_24447,N_24709);
nand UO_2951 (O_2951,N_23075,N_19590);
nor UO_2952 (O_2952,N_23050,N_21993);
xor UO_2953 (O_2953,N_20899,N_19370);
nor UO_2954 (O_2954,N_24148,N_19996);
nor UO_2955 (O_2955,N_20660,N_19358);
or UO_2956 (O_2956,N_19533,N_23412);
nand UO_2957 (O_2957,N_20609,N_20093);
nor UO_2958 (O_2958,N_23288,N_18999);
xor UO_2959 (O_2959,N_19338,N_23058);
nand UO_2960 (O_2960,N_19003,N_21737);
nor UO_2961 (O_2961,N_24591,N_22904);
nand UO_2962 (O_2962,N_23419,N_24101);
or UO_2963 (O_2963,N_22175,N_23161);
and UO_2964 (O_2964,N_20212,N_23507);
and UO_2965 (O_2965,N_18953,N_23036);
nand UO_2966 (O_2966,N_22367,N_18824);
and UO_2967 (O_2967,N_24647,N_24520);
nor UO_2968 (O_2968,N_24177,N_24219);
or UO_2969 (O_2969,N_22883,N_23446);
and UO_2970 (O_2970,N_19764,N_22938);
and UO_2971 (O_2971,N_22843,N_23938);
nor UO_2972 (O_2972,N_19803,N_23498);
or UO_2973 (O_2973,N_22662,N_22324);
xor UO_2974 (O_2974,N_20412,N_21627);
xor UO_2975 (O_2975,N_22243,N_23331);
nor UO_2976 (O_2976,N_24651,N_20240);
nand UO_2977 (O_2977,N_23860,N_24763);
nand UO_2978 (O_2978,N_20074,N_20440);
and UO_2979 (O_2979,N_19681,N_21668);
and UO_2980 (O_2980,N_19401,N_24264);
or UO_2981 (O_2981,N_20162,N_21398);
xnor UO_2982 (O_2982,N_21659,N_24874);
nand UO_2983 (O_2983,N_19268,N_18967);
nand UO_2984 (O_2984,N_24613,N_23790);
nor UO_2985 (O_2985,N_20965,N_24840);
nand UO_2986 (O_2986,N_21197,N_22722);
and UO_2987 (O_2987,N_22323,N_23490);
nand UO_2988 (O_2988,N_23741,N_21390);
or UO_2989 (O_2989,N_19399,N_19929);
nor UO_2990 (O_2990,N_24033,N_24007);
nor UO_2991 (O_2991,N_22588,N_24577);
nor UO_2992 (O_2992,N_23319,N_24251);
or UO_2993 (O_2993,N_21943,N_22702);
nor UO_2994 (O_2994,N_19351,N_20805);
xnor UO_2995 (O_2995,N_20077,N_22778);
nor UO_2996 (O_2996,N_22438,N_20168);
nand UO_2997 (O_2997,N_22221,N_22262);
or UO_2998 (O_2998,N_24544,N_19484);
nand UO_2999 (O_2999,N_22844,N_20916);
endmodule