module basic_750_5000_1000_10_levels_1xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nor U0 (N_0,In_244,In_499);
xnor U1 (N_1,In_362,In_482);
or U2 (N_2,In_249,In_297);
nand U3 (N_3,In_389,In_627);
nand U4 (N_4,In_506,In_6);
or U5 (N_5,In_17,In_301);
or U6 (N_6,In_584,In_196);
nand U7 (N_7,In_293,In_708);
and U8 (N_8,In_167,In_523);
nand U9 (N_9,In_258,In_673);
and U10 (N_10,In_284,In_97);
nor U11 (N_11,In_593,In_236);
and U12 (N_12,In_158,In_594);
nor U13 (N_13,In_644,In_736);
or U14 (N_14,In_342,In_512);
and U15 (N_15,In_378,In_697);
nand U16 (N_16,In_491,In_291);
or U17 (N_17,In_374,In_615);
nand U18 (N_18,In_495,In_115);
and U19 (N_19,In_407,In_273);
nor U20 (N_20,In_398,In_292);
and U21 (N_21,In_534,In_687);
nand U22 (N_22,In_746,In_324);
and U23 (N_23,In_738,In_340);
nand U24 (N_24,In_24,In_698);
and U25 (N_25,In_371,In_353);
or U26 (N_26,In_520,In_671);
and U27 (N_27,In_35,In_426);
nand U28 (N_28,In_60,In_605);
or U29 (N_29,In_667,In_99);
or U30 (N_30,In_119,In_717);
and U31 (N_31,In_424,In_542);
nand U32 (N_32,In_150,In_30);
nor U33 (N_33,In_98,In_388);
or U34 (N_34,In_136,In_25);
or U35 (N_35,In_114,In_201);
nand U36 (N_36,In_451,In_303);
nor U37 (N_37,In_566,In_664);
or U38 (N_38,In_455,In_326);
or U39 (N_39,In_210,In_406);
or U40 (N_40,In_476,In_39);
and U41 (N_41,In_264,In_127);
nand U42 (N_42,In_529,In_51);
and U43 (N_43,In_16,In_176);
and U44 (N_44,In_704,In_442);
nor U45 (N_45,In_507,In_254);
nor U46 (N_46,In_550,In_487);
nor U47 (N_47,In_357,In_415);
or U48 (N_48,In_350,In_372);
and U49 (N_49,In_654,In_103);
or U50 (N_50,In_700,In_689);
nand U51 (N_51,In_314,In_94);
or U52 (N_52,In_530,In_272);
or U53 (N_53,In_440,In_492);
nor U54 (N_54,In_624,In_490);
nand U55 (N_55,In_547,In_445);
or U56 (N_56,In_574,In_635);
nand U57 (N_57,In_4,In_443);
nor U58 (N_58,In_515,In_125);
or U59 (N_59,In_749,In_100);
nor U60 (N_60,In_76,In_302);
and U61 (N_61,In_257,In_377);
nor U62 (N_62,In_582,In_437);
nor U63 (N_63,In_557,In_65);
and U64 (N_64,In_674,In_545);
or U65 (N_65,In_485,In_164);
and U66 (N_66,In_657,In_448);
and U67 (N_67,In_188,In_247);
nor U68 (N_68,In_603,In_113);
or U69 (N_69,In_732,In_248);
xnor U70 (N_70,In_253,In_570);
and U71 (N_71,In_500,In_628);
or U72 (N_72,In_385,In_89);
and U73 (N_73,In_536,In_466);
nor U74 (N_74,In_225,In_430);
and U75 (N_75,In_280,In_447);
nor U76 (N_76,In_590,In_524);
or U77 (N_77,In_327,In_243);
nand U78 (N_78,In_538,In_218);
nor U79 (N_79,In_222,In_427);
and U80 (N_80,In_505,In_414);
nand U81 (N_81,In_170,In_509);
nor U82 (N_82,In_211,In_259);
nand U83 (N_83,In_58,In_493);
and U84 (N_84,In_488,In_434);
or U85 (N_85,In_431,In_300);
or U86 (N_86,In_632,In_358);
nor U87 (N_87,In_501,In_686);
nor U88 (N_88,In_337,In_436);
and U89 (N_89,In_726,In_304);
and U90 (N_90,In_422,In_26);
nand U91 (N_91,In_472,In_90);
nand U92 (N_92,In_70,In_360);
nand U93 (N_93,In_359,In_595);
nand U94 (N_94,In_688,In_88);
or U95 (N_95,In_577,In_496);
nand U96 (N_96,In_335,In_600);
and U97 (N_97,In_638,In_20);
and U98 (N_98,In_33,In_567);
nor U99 (N_99,In_27,In_172);
nand U100 (N_100,In_339,In_614);
or U101 (N_101,In_652,In_152);
nor U102 (N_102,In_93,In_479);
and U103 (N_103,In_276,In_636);
nand U104 (N_104,In_647,In_260);
and U105 (N_105,In_428,In_556);
or U106 (N_106,In_625,In_117);
nand U107 (N_107,In_129,In_18);
nor U108 (N_108,In_399,In_111);
nand U109 (N_109,In_279,In_723);
or U110 (N_110,In_610,In_576);
or U111 (N_111,In_46,In_290);
nor U112 (N_112,In_444,In_658);
nand U113 (N_113,In_581,In_352);
or U114 (N_114,In_695,In_197);
and U115 (N_115,In_413,In_747);
nor U116 (N_116,In_382,In_40);
or U117 (N_117,In_468,In_561);
nand U118 (N_118,In_611,In_522);
nand U119 (N_119,In_267,In_59);
and U120 (N_120,In_151,In_165);
nand U121 (N_121,In_669,In_183);
or U122 (N_122,In_475,In_441);
nor U123 (N_123,In_195,In_517);
nor U124 (N_124,In_663,In_226);
nand U125 (N_125,In_121,In_438);
or U126 (N_126,In_580,In_602);
nand U127 (N_127,In_137,In_84);
or U128 (N_128,In_345,In_465);
or U129 (N_129,In_457,In_564);
nand U130 (N_130,In_333,In_696);
or U131 (N_131,In_516,In_618);
nor U132 (N_132,In_470,In_510);
and U133 (N_133,In_571,In_720);
or U134 (N_134,In_416,In_2);
nand U135 (N_135,In_401,In_693);
nand U136 (N_136,In_518,In_640);
nand U137 (N_137,In_138,In_91);
or U138 (N_138,In_552,In_64);
and U139 (N_139,In_660,In_462);
nand U140 (N_140,In_474,In_642);
nor U141 (N_141,In_721,In_713);
nand U142 (N_142,In_316,In_251);
nand U143 (N_143,In_684,In_289);
nor U144 (N_144,In_271,In_232);
nor U145 (N_145,In_395,In_296);
or U146 (N_146,In_57,In_87);
nor U147 (N_147,In_206,In_380);
or U148 (N_148,In_743,In_5);
or U149 (N_149,In_458,In_308);
nand U150 (N_150,In_95,In_425);
and U151 (N_151,In_347,In_692);
or U152 (N_152,In_420,In_404);
or U153 (N_153,In_393,In_126);
and U154 (N_154,In_366,In_562);
nand U155 (N_155,In_429,In_322);
nand U156 (N_156,In_541,In_268);
or U157 (N_157,In_453,In_643);
nor U158 (N_158,In_400,In_634);
nor U159 (N_159,In_539,In_67);
nor U160 (N_160,In_23,In_234);
nor U161 (N_161,In_41,In_531);
nor U162 (N_162,In_174,In_344);
nand U163 (N_163,In_80,In_473);
nor U164 (N_164,In_733,In_15);
and U165 (N_165,In_486,In_553);
nor U166 (N_166,In_265,In_239);
and U167 (N_167,In_596,In_146);
or U168 (N_168,In_159,In_219);
nor U169 (N_169,In_134,In_659);
nand U170 (N_170,In_629,In_144);
nand U171 (N_171,In_537,In_528);
nand U172 (N_172,In_107,In_682);
nor U173 (N_173,In_200,In_221);
or U174 (N_174,In_592,In_707);
nand U175 (N_175,In_139,In_554);
nor U176 (N_176,In_702,In_135);
nand U177 (N_177,In_148,In_143);
or U178 (N_178,In_587,In_348);
nor U179 (N_179,In_722,In_277);
or U180 (N_180,In_320,In_63);
or U181 (N_181,In_619,In_169);
and U182 (N_182,In_588,In_367);
nand U183 (N_183,In_675,In_50);
nand U184 (N_184,In_421,In_412);
nor U185 (N_185,In_551,In_641);
or U186 (N_186,In_665,In_275);
or U187 (N_187,In_452,In_410);
nand U188 (N_188,In_494,In_61);
xor U189 (N_189,In_52,In_356);
or U190 (N_190,In_325,In_616);
and U191 (N_191,In_282,In_12);
nor U192 (N_192,In_132,In_368);
and U193 (N_193,In_394,In_199);
or U194 (N_194,In_184,In_256);
nand U195 (N_195,In_432,In_28);
nand U196 (N_196,In_655,In_92);
nor U197 (N_197,In_163,In_423);
or U198 (N_198,In_71,In_43);
xor U199 (N_199,In_578,In_202);
nor U200 (N_200,In_730,In_307);
and U201 (N_201,In_250,In_319);
nor U202 (N_202,In_104,In_212);
nor U203 (N_203,In_569,In_503);
nor U204 (N_204,In_646,In_245);
nor U205 (N_205,In_179,In_508);
nand U206 (N_206,In_729,In_118);
nand U207 (N_207,In_31,In_14);
nor U208 (N_208,In_710,In_224);
and U209 (N_209,In_706,In_355);
or U210 (N_210,In_124,In_82);
and U211 (N_211,In_128,In_548);
and U212 (N_212,In_691,In_227);
nand U213 (N_213,In_261,In_108);
and U214 (N_214,In_213,In_73);
or U215 (N_215,In_310,In_477);
and U216 (N_216,In_328,In_598);
or U217 (N_217,In_228,In_651);
nand U218 (N_218,In_209,In_287);
or U219 (N_219,In_417,In_311);
nand U220 (N_220,In_364,In_181);
and U221 (N_221,In_678,In_719);
nand U222 (N_222,In_601,In_361);
nor U223 (N_223,In_155,In_365);
or U224 (N_224,In_392,In_712);
nand U225 (N_225,In_266,In_0);
and U226 (N_226,In_315,In_3);
nor U227 (N_227,In_583,In_504);
and U228 (N_228,In_262,In_405);
and U229 (N_229,In_75,In_563);
nand U230 (N_230,In_381,In_386);
and U231 (N_231,In_403,In_446);
nand U232 (N_232,In_252,In_724);
nor U233 (N_233,In_185,In_109);
nor U234 (N_234,In_81,In_662);
or U235 (N_235,In_630,In_645);
nor U236 (N_236,In_175,In_532);
or U237 (N_237,In_10,In_141);
nand U238 (N_238,In_317,In_391);
and U239 (N_239,In_513,In_229);
nor U240 (N_240,In_180,In_727);
and U241 (N_241,In_330,In_734);
and U242 (N_242,In_384,In_460);
nor U243 (N_243,In_55,In_572);
or U244 (N_244,In_639,In_123);
and U245 (N_245,In_408,In_68);
and U246 (N_246,In_157,In_110);
nand U247 (N_247,In_613,In_8);
and U248 (N_248,In_469,In_612);
nand U249 (N_249,In_742,In_681);
nand U250 (N_250,In_573,In_661);
nand U251 (N_251,In_685,In_205);
and U252 (N_252,In_116,In_69);
nand U253 (N_253,In_543,In_631);
or U254 (N_254,In_263,In_38);
nor U255 (N_255,In_597,In_668);
or U256 (N_256,In_306,In_411);
nand U257 (N_257,In_173,In_278);
nor U258 (N_258,In_449,In_161);
and U259 (N_259,In_255,In_79);
or U260 (N_260,In_715,In_220);
nor U261 (N_261,In_145,In_49);
or U262 (N_262,In_177,In_699);
nor U263 (N_263,In_332,In_683);
nand U264 (N_264,In_21,In_166);
and U265 (N_265,In_483,In_122);
nor U266 (N_266,In_191,In_383);
and U267 (N_267,In_521,In_725);
nor U268 (N_268,In_498,In_29);
nor U269 (N_269,In_728,In_617);
or U270 (N_270,In_608,In_242);
xnor U271 (N_271,In_526,In_656);
nand U272 (N_272,In_189,In_533);
nand U273 (N_273,In_182,In_633);
or U274 (N_274,In_419,In_471);
nand U275 (N_275,In_459,In_149);
and U276 (N_276,In_418,In_238);
or U277 (N_277,In_679,In_666);
or U278 (N_278,In_555,In_193);
nand U279 (N_279,In_489,In_606);
and U280 (N_280,In_741,In_274);
nand U281 (N_281,In_709,In_231);
and U282 (N_282,In_36,In_96);
or U283 (N_283,In_120,In_54);
xor U284 (N_284,In_599,In_74);
and U285 (N_285,In_535,In_546);
nor U286 (N_286,In_154,In_269);
nand U287 (N_287,In_215,In_13);
and U288 (N_288,In_396,In_343);
or U289 (N_289,In_650,In_497);
nand U290 (N_290,In_62,In_37);
or U291 (N_291,In_637,In_349);
or U292 (N_292,In_230,In_153);
or U293 (N_293,In_190,In_237);
nand U294 (N_294,In_680,In_66);
nand U295 (N_295,In_106,In_716);
or U296 (N_296,In_147,In_77);
and U297 (N_297,In_204,In_101);
and U298 (N_298,In_511,In_216);
nand U299 (N_299,In_171,In_207);
or U300 (N_300,In_346,In_22);
and U301 (N_301,In_288,In_214);
or U302 (N_302,In_456,In_373);
nand U303 (N_303,In_241,In_740);
nor U304 (N_304,In_439,In_478);
or U305 (N_305,In_514,In_246);
or U306 (N_306,In_329,In_622);
nor U307 (N_307,In_45,In_586);
and U308 (N_308,In_701,In_47);
nor U309 (N_309,In_379,In_744);
and U310 (N_310,In_318,In_620);
nand U311 (N_311,In_34,In_240);
and U312 (N_312,In_464,In_677);
and U313 (N_313,In_321,In_112);
or U314 (N_314,In_105,In_558);
nor U315 (N_315,In_72,In_454);
and U316 (N_316,In_203,In_560);
nand U317 (N_317,In_575,In_323);
and U318 (N_318,In_44,In_1);
and U319 (N_319,In_56,In_194);
or U320 (N_320,In_156,In_142);
nand U321 (N_321,In_649,In_375);
or U322 (N_322,In_519,In_286);
nand U323 (N_323,In_168,In_387);
or U324 (N_324,In_133,In_559);
or U325 (N_325,In_463,In_591);
and U326 (N_326,In_653,In_283);
or U327 (N_327,In_294,In_299);
and U328 (N_328,In_670,In_705);
or U329 (N_329,In_42,In_694);
or U330 (N_330,In_78,In_281);
or U331 (N_331,In_85,In_160);
or U332 (N_332,In_363,In_376);
nand U333 (N_333,In_233,In_402);
and U334 (N_334,In_186,In_481);
nor U335 (N_335,In_192,In_731);
nand U336 (N_336,In_626,In_527);
and U337 (N_337,In_198,In_48);
or U338 (N_338,In_309,In_131);
nand U339 (N_339,In_285,In_19);
nor U340 (N_340,In_390,In_270);
and U341 (N_341,In_739,In_208);
nor U342 (N_342,In_690,In_86);
and U343 (N_343,In_604,In_737);
nand U344 (N_344,In_217,In_748);
or U345 (N_345,In_648,In_9);
and U346 (N_346,In_549,In_579);
or U347 (N_347,In_369,In_480);
or U348 (N_348,In_565,In_338);
nor U349 (N_349,In_140,In_718);
or U350 (N_350,In_7,In_623);
nor U351 (N_351,In_672,In_295);
or U352 (N_352,In_313,In_370);
or U353 (N_353,In_102,In_312);
or U354 (N_354,In_502,In_162);
nand U355 (N_355,In_609,In_53);
and U356 (N_356,In_607,In_341);
nor U357 (N_357,In_676,In_450);
nor U358 (N_358,In_745,In_484);
nand U359 (N_359,In_409,In_187);
nor U360 (N_360,In_336,In_298);
nor U361 (N_361,In_223,In_83);
or U362 (N_362,In_305,In_397);
nand U363 (N_363,In_178,In_334);
or U364 (N_364,In_735,In_467);
and U365 (N_365,In_544,In_589);
or U366 (N_366,In_331,In_130);
or U367 (N_367,In_525,In_351);
and U368 (N_368,In_621,In_585);
nor U369 (N_369,In_703,In_11);
nor U370 (N_370,In_568,In_235);
nand U371 (N_371,In_711,In_433);
and U372 (N_372,In_540,In_435);
and U373 (N_373,In_32,In_354);
nand U374 (N_374,In_714,In_461);
and U375 (N_375,In_727,In_560);
nor U376 (N_376,In_430,In_569);
nor U377 (N_377,In_506,In_589);
nand U378 (N_378,In_374,In_377);
nand U379 (N_379,In_245,In_349);
nor U380 (N_380,In_36,In_427);
and U381 (N_381,In_279,In_255);
nand U382 (N_382,In_43,In_168);
nand U383 (N_383,In_37,In_583);
nand U384 (N_384,In_3,In_172);
nand U385 (N_385,In_478,In_138);
nand U386 (N_386,In_106,In_155);
and U387 (N_387,In_268,In_510);
nand U388 (N_388,In_80,In_412);
nand U389 (N_389,In_300,In_294);
and U390 (N_390,In_549,In_232);
nor U391 (N_391,In_392,In_69);
nor U392 (N_392,In_669,In_412);
nor U393 (N_393,In_531,In_186);
or U394 (N_394,In_719,In_434);
and U395 (N_395,In_139,In_303);
and U396 (N_396,In_710,In_331);
nand U397 (N_397,In_389,In_747);
or U398 (N_398,In_189,In_337);
and U399 (N_399,In_685,In_229);
nor U400 (N_400,In_593,In_202);
or U401 (N_401,In_610,In_394);
or U402 (N_402,In_177,In_720);
and U403 (N_403,In_570,In_175);
nand U404 (N_404,In_370,In_575);
nor U405 (N_405,In_642,In_418);
or U406 (N_406,In_175,In_531);
nand U407 (N_407,In_437,In_624);
and U408 (N_408,In_339,In_16);
and U409 (N_409,In_245,In_179);
nor U410 (N_410,In_156,In_325);
and U411 (N_411,In_691,In_488);
and U412 (N_412,In_690,In_22);
nor U413 (N_413,In_158,In_162);
or U414 (N_414,In_381,In_382);
nor U415 (N_415,In_269,In_271);
or U416 (N_416,In_624,In_400);
nand U417 (N_417,In_644,In_590);
nand U418 (N_418,In_362,In_41);
nor U419 (N_419,In_589,In_546);
and U420 (N_420,In_663,In_96);
nor U421 (N_421,In_21,In_674);
nand U422 (N_422,In_745,In_425);
nor U423 (N_423,In_448,In_305);
or U424 (N_424,In_616,In_570);
nor U425 (N_425,In_85,In_623);
nand U426 (N_426,In_166,In_334);
nand U427 (N_427,In_154,In_228);
nand U428 (N_428,In_565,In_420);
nand U429 (N_429,In_361,In_23);
or U430 (N_430,In_43,In_329);
nor U431 (N_431,In_282,In_594);
nand U432 (N_432,In_731,In_705);
nand U433 (N_433,In_70,In_207);
or U434 (N_434,In_511,In_623);
and U435 (N_435,In_224,In_447);
nor U436 (N_436,In_455,In_707);
or U437 (N_437,In_516,In_238);
or U438 (N_438,In_265,In_382);
nand U439 (N_439,In_396,In_246);
or U440 (N_440,In_199,In_597);
nand U441 (N_441,In_506,In_242);
nor U442 (N_442,In_550,In_392);
and U443 (N_443,In_506,In_137);
and U444 (N_444,In_745,In_677);
nor U445 (N_445,In_477,In_605);
nor U446 (N_446,In_257,In_138);
nand U447 (N_447,In_444,In_741);
and U448 (N_448,In_682,In_164);
and U449 (N_449,In_425,In_58);
and U450 (N_450,In_200,In_192);
nand U451 (N_451,In_25,In_466);
nor U452 (N_452,In_616,In_522);
nor U453 (N_453,In_735,In_101);
nand U454 (N_454,In_263,In_78);
or U455 (N_455,In_94,In_26);
or U456 (N_456,In_466,In_212);
or U457 (N_457,In_461,In_96);
nor U458 (N_458,In_101,In_350);
or U459 (N_459,In_667,In_616);
nor U460 (N_460,In_452,In_289);
or U461 (N_461,In_29,In_12);
nand U462 (N_462,In_341,In_309);
or U463 (N_463,In_8,In_221);
or U464 (N_464,In_302,In_164);
nor U465 (N_465,In_714,In_220);
or U466 (N_466,In_733,In_336);
or U467 (N_467,In_338,In_350);
or U468 (N_468,In_619,In_333);
or U469 (N_469,In_553,In_171);
nor U470 (N_470,In_561,In_330);
and U471 (N_471,In_49,In_433);
nor U472 (N_472,In_353,In_207);
and U473 (N_473,In_109,In_366);
nor U474 (N_474,In_533,In_629);
or U475 (N_475,In_611,In_137);
nor U476 (N_476,In_432,In_315);
nor U477 (N_477,In_203,In_250);
nand U478 (N_478,In_30,In_613);
and U479 (N_479,In_426,In_323);
nor U480 (N_480,In_463,In_541);
nor U481 (N_481,In_255,In_746);
nand U482 (N_482,In_343,In_109);
or U483 (N_483,In_744,In_503);
nand U484 (N_484,In_326,In_258);
or U485 (N_485,In_460,In_154);
or U486 (N_486,In_224,In_678);
nor U487 (N_487,In_5,In_120);
or U488 (N_488,In_348,In_499);
and U489 (N_489,In_176,In_688);
or U490 (N_490,In_703,In_55);
and U491 (N_491,In_696,In_123);
nand U492 (N_492,In_32,In_500);
nor U493 (N_493,In_692,In_48);
and U494 (N_494,In_155,In_709);
and U495 (N_495,In_67,In_422);
nand U496 (N_496,In_361,In_419);
nand U497 (N_497,In_427,In_202);
nand U498 (N_498,In_234,In_250);
or U499 (N_499,In_416,In_190);
or U500 (N_500,N_430,N_384);
or U501 (N_501,N_306,N_426);
nor U502 (N_502,N_470,N_70);
and U503 (N_503,N_302,N_254);
or U504 (N_504,N_461,N_399);
and U505 (N_505,N_276,N_50);
nor U506 (N_506,N_443,N_427);
nor U507 (N_507,N_487,N_498);
nor U508 (N_508,N_150,N_425);
and U509 (N_509,N_134,N_28);
or U510 (N_510,N_336,N_123);
or U511 (N_511,N_52,N_259);
nor U512 (N_512,N_92,N_135);
or U513 (N_513,N_88,N_347);
nor U514 (N_514,N_244,N_31);
nand U515 (N_515,N_251,N_233);
and U516 (N_516,N_294,N_469);
nor U517 (N_517,N_483,N_34);
nor U518 (N_518,N_220,N_475);
or U519 (N_519,N_203,N_262);
nand U520 (N_520,N_42,N_51);
nor U521 (N_521,N_112,N_129);
or U522 (N_522,N_218,N_121);
or U523 (N_523,N_444,N_143);
and U524 (N_524,N_55,N_58);
or U525 (N_525,N_73,N_125);
and U526 (N_526,N_142,N_131);
nor U527 (N_527,N_354,N_368);
nor U528 (N_528,N_192,N_414);
nor U529 (N_529,N_24,N_11);
nand U530 (N_530,N_326,N_381);
and U531 (N_531,N_473,N_261);
nand U532 (N_532,N_246,N_268);
and U533 (N_533,N_372,N_228);
and U534 (N_534,N_235,N_253);
or U535 (N_535,N_63,N_84);
and U536 (N_536,N_115,N_272);
nor U537 (N_537,N_286,N_155);
nand U538 (N_538,N_89,N_157);
nand U539 (N_539,N_35,N_97);
or U540 (N_540,N_394,N_391);
nand U541 (N_541,N_418,N_257);
and U542 (N_542,N_85,N_489);
nand U543 (N_543,N_59,N_386);
and U544 (N_544,N_434,N_17);
nand U545 (N_545,N_66,N_248);
and U546 (N_546,N_488,N_455);
nor U547 (N_547,N_232,N_119);
nand U548 (N_548,N_324,N_18);
or U549 (N_549,N_39,N_456);
or U550 (N_550,N_329,N_447);
and U551 (N_551,N_330,N_343);
nor U552 (N_552,N_3,N_169);
nor U553 (N_553,N_114,N_457);
nand U554 (N_554,N_260,N_44);
nor U555 (N_555,N_40,N_280);
or U556 (N_556,N_205,N_138);
and U557 (N_557,N_122,N_15);
nor U558 (N_558,N_188,N_486);
nand U559 (N_559,N_385,N_497);
nand U560 (N_560,N_269,N_229);
nor U561 (N_561,N_107,N_398);
and U562 (N_562,N_30,N_383);
or U563 (N_563,N_282,N_312);
nor U564 (N_564,N_12,N_284);
nand U565 (N_565,N_185,N_87);
or U566 (N_566,N_202,N_337);
and U567 (N_567,N_81,N_287);
nand U568 (N_568,N_328,N_72);
or U569 (N_569,N_446,N_465);
or U570 (N_570,N_16,N_266);
or U571 (N_571,N_158,N_451);
and U572 (N_572,N_376,N_69);
and U573 (N_573,N_181,N_357);
and U574 (N_574,N_168,N_258);
or U575 (N_575,N_278,N_221);
and U576 (N_576,N_172,N_236);
or U577 (N_577,N_247,N_10);
or U578 (N_578,N_397,N_423);
nor U579 (N_579,N_231,N_499);
nor U580 (N_580,N_208,N_339);
nand U581 (N_581,N_335,N_227);
or U582 (N_582,N_448,N_299);
nand U583 (N_583,N_161,N_365);
nor U584 (N_584,N_428,N_325);
or U585 (N_585,N_241,N_304);
nor U586 (N_586,N_207,N_362);
or U587 (N_587,N_33,N_413);
nor U588 (N_588,N_290,N_240);
and U589 (N_589,N_250,N_141);
or U590 (N_590,N_94,N_178);
and U591 (N_591,N_159,N_130);
or U592 (N_592,N_183,N_353);
nand U593 (N_593,N_102,N_379);
and U594 (N_594,N_1,N_474);
and U595 (N_595,N_149,N_184);
or U596 (N_596,N_151,N_410);
xnor U597 (N_597,N_118,N_277);
nand U598 (N_598,N_495,N_340);
or U599 (N_599,N_127,N_267);
or U600 (N_600,N_23,N_403);
and U601 (N_601,N_179,N_466);
and U602 (N_602,N_7,N_318);
and U603 (N_603,N_46,N_27);
or U604 (N_604,N_490,N_171);
nand U605 (N_605,N_25,N_21);
xor U606 (N_606,N_26,N_359);
or U607 (N_607,N_275,N_164);
nor U608 (N_608,N_93,N_440);
nor U609 (N_609,N_99,N_213);
and U610 (N_610,N_230,N_154);
or U611 (N_611,N_37,N_484);
nand U612 (N_612,N_462,N_491);
nand U613 (N_613,N_182,N_453);
and U614 (N_614,N_361,N_291);
and U615 (N_615,N_409,N_68);
nand U616 (N_616,N_323,N_334);
nor U617 (N_617,N_38,N_494);
or U618 (N_618,N_327,N_62);
nor U619 (N_619,N_404,N_177);
and U620 (N_620,N_234,N_214);
or U621 (N_621,N_407,N_420);
nand U622 (N_622,N_199,N_243);
nand U623 (N_623,N_270,N_196);
and U624 (N_624,N_389,N_64);
and U625 (N_625,N_5,N_303);
or U626 (N_626,N_224,N_369);
nor U627 (N_627,N_279,N_195);
nor U628 (N_628,N_22,N_405);
nor U629 (N_629,N_29,N_77);
or U630 (N_630,N_476,N_321);
nor U631 (N_631,N_468,N_166);
or U632 (N_632,N_48,N_219);
nand U633 (N_633,N_223,N_493);
nor U634 (N_634,N_445,N_106);
nand U635 (N_635,N_110,N_226);
or U636 (N_636,N_120,N_316);
nand U637 (N_637,N_432,N_358);
and U638 (N_638,N_496,N_373);
and U639 (N_639,N_167,N_86);
nand U640 (N_640,N_201,N_450);
and U641 (N_641,N_79,N_308);
and U642 (N_642,N_285,N_377);
nand U643 (N_643,N_482,N_9);
nand U644 (N_644,N_75,N_419);
nand U645 (N_645,N_356,N_332);
or U646 (N_646,N_438,N_53);
nor U647 (N_647,N_100,N_309);
and U648 (N_648,N_83,N_415);
or U649 (N_649,N_82,N_412);
nand U650 (N_650,N_32,N_90);
nor U651 (N_651,N_148,N_49);
or U652 (N_652,N_411,N_216);
or U653 (N_653,N_61,N_481);
and U654 (N_654,N_217,N_47);
and U655 (N_655,N_293,N_402);
nor U656 (N_656,N_265,N_105);
or U657 (N_657,N_19,N_289);
nand U658 (N_658,N_111,N_263);
or U659 (N_659,N_204,N_45);
nand U660 (N_660,N_54,N_342);
nand U661 (N_661,N_13,N_264);
and U662 (N_662,N_140,N_370);
or U663 (N_663,N_139,N_408);
or U664 (N_664,N_344,N_109);
or U665 (N_665,N_160,N_416);
and U666 (N_666,N_91,N_170);
nand U667 (N_667,N_471,N_371);
nor U668 (N_668,N_459,N_145);
and U669 (N_669,N_222,N_363);
nand U670 (N_670,N_67,N_479);
nand U671 (N_671,N_80,N_305);
and U672 (N_672,N_375,N_480);
or U673 (N_673,N_464,N_71);
nand U674 (N_674,N_147,N_57);
nand U675 (N_675,N_435,N_225);
and U676 (N_676,N_298,N_95);
and U677 (N_677,N_8,N_163);
nor U678 (N_678,N_437,N_211);
nand U679 (N_679,N_388,N_283);
or U680 (N_680,N_400,N_421);
and U681 (N_681,N_117,N_292);
nor U682 (N_682,N_249,N_78);
or U683 (N_683,N_311,N_152);
or U684 (N_684,N_255,N_256);
and U685 (N_685,N_351,N_132);
nor U686 (N_686,N_393,N_133);
and U687 (N_687,N_43,N_380);
or U688 (N_688,N_341,N_98);
nand U689 (N_689,N_281,N_271);
nand U690 (N_690,N_355,N_477);
xor U691 (N_691,N_458,N_124);
or U692 (N_692,N_165,N_478);
nand U693 (N_693,N_422,N_0);
and U694 (N_694,N_374,N_364);
xor U695 (N_695,N_242,N_317);
nand U696 (N_696,N_392,N_198);
or U697 (N_697,N_378,N_366);
and U698 (N_698,N_104,N_307);
nor U699 (N_699,N_41,N_431);
or U700 (N_700,N_162,N_206);
nand U701 (N_701,N_401,N_460);
or U702 (N_702,N_36,N_197);
or U703 (N_703,N_467,N_331);
nand U704 (N_704,N_113,N_96);
nor U705 (N_705,N_65,N_274);
nand U706 (N_706,N_301,N_390);
and U707 (N_707,N_463,N_442);
and U708 (N_708,N_252,N_144);
and U709 (N_709,N_472,N_433);
and U710 (N_710,N_212,N_187);
nand U711 (N_711,N_350,N_60);
or U712 (N_712,N_429,N_193);
and U713 (N_713,N_295,N_387);
or U714 (N_714,N_76,N_382);
or U715 (N_715,N_349,N_338);
or U716 (N_716,N_215,N_314);
nor U717 (N_717,N_439,N_441);
and U718 (N_718,N_360,N_396);
and U719 (N_719,N_156,N_310);
nand U720 (N_720,N_14,N_2);
nand U721 (N_721,N_273,N_300);
and U722 (N_722,N_452,N_417);
and U723 (N_723,N_492,N_209);
or U724 (N_724,N_333,N_367);
or U725 (N_725,N_297,N_174);
or U726 (N_726,N_128,N_191);
and U727 (N_727,N_180,N_352);
or U728 (N_728,N_238,N_485);
nand U729 (N_729,N_322,N_173);
or U730 (N_730,N_348,N_116);
nor U731 (N_731,N_406,N_319);
and U732 (N_732,N_137,N_146);
or U733 (N_733,N_424,N_313);
or U734 (N_734,N_454,N_186);
nand U735 (N_735,N_74,N_315);
and U736 (N_736,N_239,N_288);
nor U737 (N_737,N_345,N_108);
or U738 (N_738,N_210,N_103);
nand U739 (N_739,N_20,N_200);
nand U740 (N_740,N_56,N_126);
or U741 (N_741,N_101,N_436);
nand U742 (N_742,N_6,N_175);
and U743 (N_743,N_346,N_4);
and U744 (N_744,N_190,N_296);
or U745 (N_745,N_245,N_136);
nor U746 (N_746,N_320,N_153);
nor U747 (N_747,N_189,N_395);
or U748 (N_748,N_237,N_194);
or U749 (N_749,N_449,N_176);
and U750 (N_750,N_7,N_14);
or U751 (N_751,N_127,N_44);
or U752 (N_752,N_420,N_398);
nor U753 (N_753,N_63,N_453);
or U754 (N_754,N_44,N_386);
or U755 (N_755,N_225,N_463);
xor U756 (N_756,N_482,N_167);
nand U757 (N_757,N_158,N_411);
nand U758 (N_758,N_409,N_199);
nor U759 (N_759,N_84,N_308);
and U760 (N_760,N_91,N_322);
nor U761 (N_761,N_324,N_310);
and U762 (N_762,N_336,N_367);
nor U763 (N_763,N_448,N_91);
nand U764 (N_764,N_200,N_128);
nand U765 (N_765,N_476,N_299);
nor U766 (N_766,N_442,N_186);
nor U767 (N_767,N_113,N_55);
nor U768 (N_768,N_499,N_90);
nor U769 (N_769,N_460,N_490);
nand U770 (N_770,N_116,N_425);
nand U771 (N_771,N_458,N_46);
and U772 (N_772,N_356,N_413);
or U773 (N_773,N_134,N_490);
xor U774 (N_774,N_490,N_290);
nand U775 (N_775,N_230,N_491);
and U776 (N_776,N_297,N_341);
nor U777 (N_777,N_425,N_351);
or U778 (N_778,N_263,N_26);
and U779 (N_779,N_491,N_274);
and U780 (N_780,N_386,N_156);
nor U781 (N_781,N_441,N_297);
and U782 (N_782,N_272,N_141);
nor U783 (N_783,N_486,N_237);
nand U784 (N_784,N_161,N_408);
and U785 (N_785,N_195,N_9);
nor U786 (N_786,N_73,N_27);
nand U787 (N_787,N_105,N_260);
nand U788 (N_788,N_9,N_208);
nand U789 (N_789,N_300,N_158);
and U790 (N_790,N_314,N_69);
and U791 (N_791,N_197,N_462);
nand U792 (N_792,N_258,N_443);
and U793 (N_793,N_244,N_92);
nand U794 (N_794,N_303,N_217);
nand U795 (N_795,N_67,N_307);
or U796 (N_796,N_340,N_12);
and U797 (N_797,N_449,N_127);
and U798 (N_798,N_143,N_446);
and U799 (N_799,N_308,N_337);
or U800 (N_800,N_119,N_30);
or U801 (N_801,N_326,N_343);
nand U802 (N_802,N_162,N_325);
nor U803 (N_803,N_5,N_120);
and U804 (N_804,N_15,N_479);
or U805 (N_805,N_188,N_456);
nand U806 (N_806,N_374,N_35);
nor U807 (N_807,N_433,N_393);
nor U808 (N_808,N_428,N_239);
nor U809 (N_809,N_71,N_34);
and U810 (N_810,N_68,N_297);
nand U811 (N_811,N_180,N_196);
nor U812 (N_812,N_316,N_242);
nand U813 (N_813,N_364,N_209);
or U814 (N_814,N_488,N_495);
nand U815 (N_815,N_466,N_420);
and U816 (N_816,N_199,N_263);
and U817 (N_817,N_295,N_454);
nor U818 (N_818,N_426,N_370);
nor U819 (N_819,N_122,N_457);
nor U820 (N_820,N_318,N_341);
or U821 (N_821,N_462,N_256);
nor U822 (N_822,N_410,N_486);
or U823 (N_823,N_367,N_188);
xor U824 (N_824,N_423,N_281);
or U825 (N_825,N_390,N_308);
nor U826 (N_826,N_160,N_384);
nor U827 (N_827,N_430,N_285);
and U828 (N_828,N_448,N_328);
or U829 (N_829,N_436,N_377);
and U830 (N_830,N_120,N_105);
nor U831 (N_831,N_412,N_90);
or U832 (N_832,N_107,N_322);
nand U833 (N_833,N_88,N_12);
nor U834 (N_834,N_246,N_349);
nand U835 (N_835,N_22,N_6);
nor U836 (N_836,N_377,N_243);
or U837 (N_837,N_306,N_202);
or U838 (N_838,N_376,N_470);
nand U839 (N_839,N_460,N_66);
or U840 (N_840,N_134,N_473);
and U841 (N_841,N_449,N_235);
nand U842 (N_842,N_364,N_269);
or U843 (N_843,N_2,N_15);
nand U844 (N_844,N_233,N_427);
and U845 (N_845,N_336,N_334);
and U846 (N_846,N_74,N_263);
nand U847 (N_847,N_125,N_412);
nor U848 (N_848,N_306,N_73);
and U849 (N_849,N_237,N_376);
or U850 (N_850,N_461,N_156);
or U851 (N_851,N_230,N_256);
and U852 (N_852,N_380,N_187);
and U853 (N_853,N_317,N_211);
and U854 (N_854,N_125,N_279);
and U855 (N_855,N_238,N_455);
nor U856 (N_856,N_482,N_493);
nand U857 (N_857,N_372,N_252);
or U858 (N_858,N_410,N_430);
or U859 (N_859,N_236,N_200);
and U860 (N_860,N_184,N_343);
or U861 (N_861,N_61,N_306);
and U862 (N_862,N_166,N_285);
nand U863 (N_863,N_323,N_6);
or U864 (N_864,N_186,N_68);
nor U865 (N_865,N_46,N_119);
nor U866 (N_866,N_10,N_197);
or U867 (N_867,N_280,N_135);
nand U868 (N_868,N_418,N_164);
and U869 (N_869,N_398,N_177);
nor U870 (N_870,N_498,N_450);
nand U871 (N_871,N_465,N_80);
nor U872 (N_872,N_3,N_374);
and U873 (N_873,N_429,N_89);
or U874 (N_874,N_137,N_451);
nor U875 (N_875,N_337,N_310);
xnor U876 (N_876,N_295,N_400);
nand U877 (N_877,N_104,N_487);
or U878 (N_878,N_301,N_251);
nor U879 (N_879,N_402,N_141);
nor U880 (N_880,N_484,N_303);
or U881 (N_881,N_132,N_361);
nor U882 (N_882,N_353,N_9);
nand U883 (N_883,N_124,N_321);
nand U884 (N_884,N_358,N_291);
or U885 (N_885,N_142,N_211);
nand U886 (N_886,N_334,N_180);
or U887 (N_887,N_273,N_166);
nand U888 (N_888,N_362,N_321);
nand U889 (N_889,N_161,N_123);
and U890 (N_890,N_412,N_6);
nand U891 (N_891,N_200,N_136);
and U892 (N_892,N_164,N_313);
or U893 (N_893,N_472,N_113);
nand U894 (N_894,N_310,N_163);
and U895 (N_895,N_197,N_449);
nor U896 (N_896,N_108,N_386);
and U897 (N_897,N_137,N_328);
nor U898 (N_898,N_95,N_178);
nor U899 (N_899,N_287,N_53);
and U900 (N_900,N_25,N_155);
or U901 (N_901,N_495,N_402);
nand U902 (N_902,N_367,N_171);
nand U903 (N_903,N_215,N_26);
nand U904 (N_904,N_292,N_411);
and U905 (N_905,N_106,N_360);
and U906 (N_906,N_281,N_41);
or U907 (N_907,N_404,N_156);
or U908 (N_908,N_2,N_111);
or U909 (N_909,N_81,N_345);
nand U910 (N_910,N_250,N_460);
nor U911 (N_911,N_14,N_311);
nor U912 (N_912,N_498,N_476);
and U913 (N_913,N_50,N_433);
nor U914 (N_914,N_342,N_17);
nor U915 (N_915,N_379,N_253);
or U916 (N_916,N_100,N_60);
or U917 (N_917,N_254,N_150);
or U918 (N_918,N_33,N_24);
or U919 (N_919,N_166,N_496);
and U920 (N_920,N_400,N_381);
and U921 (N_921,N_177,N_203);
and U922 (N_922,N_283,N_474);
or U923 (N_923,N_303,N_190);
nor U924 (N_924,N_366,N_440);
nor U925 (N_925,N_358,N_337);
and U926 (N_926,N_173,N_117);
and U927 (N_927,N_301,N_65);
and U928 (N_928,N_68,N_358);
nand U929 (N_929,N_405,N_91);
nand U930 (N_930,N_5,N_183);
or U931 (N_931,N_483,N_374);
or U932 (N_932,N_110,N_171);
or U933 (N_933,N_25,N_233);
and U934 (N_934,N_195,N_476);
or U935 (N_935,N_301,N_414);
nor U936 (N_936,N_183,N_110);
and U937 (N_937,N_327,N_296);
and U938 (N_938,N_125,N_107);
or U939 (N_939,N_198,N_478);
or U940 (N_940,N_433,N_342);
nor U941 (N_941,N_203,N_385);
or U942 (N_942,N_309,N_461);
nand U943 (N_943,N_185,N_122);
nor U944 (N_944,N_167,N_365);
nor U945 (N_945,N_411,N_194);
nand U946 (N_946,N_97,N_463);
nand U947 (N_947,N_159,N_442);
and U948 (N_948,N_386,N_219);
or U949 (N_949,N_245,N_213);
and U950 (N_950,N_263,N_373);
nor U951 (N_951,N_310,N_359);
nand U952 (N_952,N_287,N_406);
or U953 (N_953,N_346,N_314);
and U954 (N_954,N_48,N_317);
nand U955 (N_955,N_465,N_397);
and U956 (N_956,N_104,N_448);
nor U957 (N_957,N_113,N_215);
nor U958 (N_958,N_368,N_13);
and U959 (N_959,N_424,N_20);
and U960 (N_960,N_426,N_299);
nor U961 (N_961,N_408,N_371);
nor U962 (N_962,N_39,N_206);
and U963 (N_963,N_225,N_40);
xnor U964 (N_964,N_70,N_118);
nor U965 (N_965,N_117,N_267);
or U966 (N_966,N_469,N_64);
nor U967 (N_967,N_165,N_140);
nand U968 (N_968,N_73,N_498);
nor U969 (N_969,N_385,N_114);
nand U970 (N_970,N_9,N_426);
nand U971 (N_971,N_277,N_72);
or U972 (N_972,N_434,N_202);
nor U973 (N_973,N_269,N_412);
nand U974 (N_974,N_121,N_295);
or U975 (N_975,N_175,N_190);
and U976 (N_976,N_9,N_419);
nor U977 (N_977,N_431,N_327);
nor U978 (N_978,N_345,N_85);
or U979 (N_979,N_6,N_375);
and U980 (N_980,N_72,N_1);
or U981 (N_981,N_5,N_351);
nor U982 (N_982,N_275,N_153);
nor U983 (N_983,N_313,N_416);
nand U984 (N_984,N_489,N_52);
nand U985 (N_985,N_360,N_304);
and U986 (N_986,N_301,N_81);
nor U987 (N_987,N_275,N_324);
and U988 (N_988,N_336,N_268);
and U989 (N_989,N_223,N_310);
and U990 (N_990,N_383,N_394);
and U991 (N_991,N_348,N_411);
and U992 (N_992,N_85,N_273);
nor U993 (N_993,N_155,N_12);
nand U994 (N_994,N_202,N_169);
nand U995 (N_995,N_408,N_459);
nor U996 (N_996,N_343,N_192);
nand U997 (N_997,N_234,N_208);
nor U998 (N_998,N_264,N_242);
nor U999 (N_999,N_89,N_69);
or U1000 (N_1000,N_546,N_809);
or U1001 (N_1001,N_783,N_621);
nand U1002 (N_1002,N_562,N_933);
nor U1003 (N_1003,N_626,N_799);
and U1004 (N_1004,N_939,N_634);
nor U1005 (N_1005,N_583,N_728);
or U1006 (N_1006,N_600,N_944);
nor U1007 (N_1007,N_603,N_936);
or U1008 (N_1008,N_774,N_890);
nor U1009 (N_1009,N_773,N_700);
and U1010 (N_1010,N_641,N_779);
or U1011 (N_1011,N_972,N_662);
and U1012 (N_1012,N_781,N_555);
nor U1013 (N_1013,N_958,N_599);
nor U1014 (N_1014,N_673,N_660);
and U1015 (N_1015,N_751,N_806);
nand U1016 (N_1016,N_503,N_922);
and U1017 (N_1017,N_827,N_536);
or U1018 (N_1018,N_581,N_849);
nor U1019 (N_1019,N_607,N_888);
or U1020 (N_1020,N_743,N_544);
nor U1021 (N_1021,N_689,N_740);
or U1022 (N_1022,N_990,N_545);
nand U1023 (N_1023,N_576,N_608);
and U1024 (N_1024,N_978,N_672);
nor U1025 (N_1025,N_526,N_776);
or U1026 (N_1026,N_523,N_855);
nand U1027 (N_1027,N_763,N_943);
nand U1028 (N_1028,N_693,N_816);
nor U1029 (N_1029,N_610,N_724);
or U1030 (N_1030,N_835,N_820);
or U1031 (N_1031,N_801,N_850);
and U1032 (N_1032,N_842,N_778);
and U1033 (N_1033,N_685,N_529);
or U1034 (N_1034,N_986,N_857);
nand U1035 (N_1035,N_543,N_598);
nand U1036 (N_1036,N_878,N_627);
or U1037 (N_1037,N_807,N_572);
or U1038 (N_1038,N_905,N_996);
or U1039 (N_1039,N_814,N_566);
and U1040 (N_1040,N_557,N_507);
and U1041 (N_1041,N_591,N_830);
nand U1042 (N_1042,N_585,N_993);
or U1043 (N_1043,N_559,N_860);
or U1044 (N_1044,N_615,N_937);
nand U1045 (N_1045,N_912,N_979);
nor U1046 (N_1046,N_534,N_822);
nand U1047 (N_1047,N_935,N_702);
and U1048 (N_1048,N_969,N_914);
nand U1049 (N_1049,N_926,N_881);
nor U1050 (N_1050,N_833,N_710);
nor U1051 (N_1051,N_582,N_683);
nand U1052 (N_1052,N_678,N_725);
and U1053 (N_1053,N_812,N_847);
nor U1054 (N_1054,N_690,N_705);
nand U1055 (N_1055,N_910,N_899);
and U1056 (N_1056,N_715,N_601);
or U1057 (N_1057,N_677,N_840);
and U1058 (N_1058,N_750,N_811);
nor U1059 (N_1059,N_722,N_824);
or U1060 (N_1060,N_749,N_618);
nand U1061 (N_1061,N_929,N_671);
nand U1062 (N_1062,N_864,N_647);
and U1063 (N_1063,N_755,N_942);
nand U1064 (N_1064,N_863,N_845);
xor U1065 (N_1065,N_694,N_528);
and U1066 (N_1066,N_904,N_741);
and U1067 (N_1067,N_586,N_580);
or U1068 (N_1068,N_675,N_510);
and U1069 (N_1069,N_759,N_645);
or U1070 (N_1070,N_558,N_515);
and U1071 (N_1071,N_780,N_525);
or U1072 (N_1072,N_854,N_925);
nor U1073 (N_1073,N_800,N_643);
nor U1074 (N_1074,N_839,N_887);
or U1075 (N_1075,N_718,N_719);
and U1076 (N_1076,N_974,N_602);
or U1077 (N_1077,N_819,N_731);
nand U1078 (N_1078,N_901,N_616);
nor U1079 (N_1079,N_648,N_823);
nor U1080 (N_1080,N_657,N_596);
nand U1081 (N_1081,N_885,N_846);
and U1082 (N_1082,N_575,N_636);
and U1083 (N_1083,N_777,N_518);
or U1084 (N_1084,N_551,N_549);
and U1085 (N_1085,N_737,N_637);
nand U1086 (N_1086,N_594,N_889);
nand U1087 (N_1087,N_771,N_653);
nand U1088 (N_1088,N_547,N_961);
or U1089 (N_1089,N_921,N_676);
nor U1090 (N_1090,N_656,N_630);
or U1091 (N_1091,N_620,N_955);
nand U1092 (N_1092,N_896,N_570);
nand U1093 (N_1093,N_826,N_650);
nor U1094 (N_1094,N_909,N_871);
and U1095 (N_1095,N_589,N_982);
nor U1096 (N_1096,N_697,N_511);
and U1097 (N_1097,N_924,N_617);
xor U1098 (N_1098,N_517,N_706);
nor U1099 (N_1099,N_852,N_638);
nand U1100 (N_1100,N_767,N_561);
and U1101 (N_1101,N_838,N_527);
and U1102 (N_1102,N_554,N_952);
nor U1103 (N_1103,N_894,N_913);
or U1104 (N_1104,N_761,N_975);
nor U1105 (N_1105,N_588,N_681);
or U1106 (N_1106,N_810,N_813);
nor U1107 (N_1107,N_631,N_966);
xor U1108 (N_1108,N_992,N_560);
nor U1109 (N_1109,N_506,N_713);
or U1110 (N_1110,N_739,N_917);
nand U1111 (N_1111,N_923,N_635);
nor U1112 (N_1112,N_666,N_752);
nor U1113 (N_1113,N_692,N_654);
or U1114 (N_1114,N_760,N_758);
or U1115 (N_1115,N_964,N_687);
nand U1116 (N_1116,N_918,N_744);
or U1117 (N_1117,N_768,N_735);
or U1118 (N_1118,N_742,N_565);
nand U1119 (N_1119,N_569,N_859);
nand U1120 (N_1120,N_784,N_931);
nor U1121 (N_1121,N_886,N_508);
nand U1122 (N_1122,N_729,N_699);
or U1123 (N_1123,N_629,N_766);
nor U1124 (N_1124,N_788,N_521);
nor U1125 (N_1125,N_994,N_548);
and U1126 (N_1126,N_956,N_853);
nand U1127 (N_1127,N_947,N_708);
and U1128 (N_1128,N_876,N_514);
nor U1129 (N_1129,N_532,N_727);
nand U1130 (N_1130,N_915,N_970);
and U1131 (N_1131,N_793,N_916);
nor U1132 (N_1132,N_639,N_873);
nor U1133 (N_1133,N_501,N_519);
nand U1134 (N_1134,N_999,N_791);
nor U1135 (N_1135,N_772,N_704);
nor U1136 (N_1136,N_568,N_973);
or U1137 (N_1137,N_789,N_717);
nand U1138 (N_1138,N_804,N_856);
and U1139 (N_1139,N_950,N_959);
nand U1140 (N_1140,N_714,N_651);
nor U1141 (N_1141,N_963,N_868);
nand U1142 (N_1142,N_764,N_844);
and U1143 (N_1143,N_946,N_757);
nand U1144 (N_1144,N_571,N_703);
nor U1145 (N_1145,N_664,N_795);
and U1146 (N_1146,N_892,N_948);
nand U1147 (N_1147,N_736,N_730);
or U1148 (N_1148,N_612,N_644);
nor U1149 (N_1149,N_655,N_723);
nor U1150 (N_1150,N_590,N_738);
or U1151 (N_1151,N_579,N_954);
or U1152 (N_1152,N_686,N_765);
and U1153 (N_1153,N_614,N_991);
or U1154 (N_1154,N_898,N_756);
and U1155 (N_1155,N_882,N_578);
nand U1156 (N_1156,N_817,N_977);
or U1157 (N_1157,N_530,N_997);
nor U1158 (N_1158,N_504,N_669);
nand U1159 (N_1159,N_516,N_938);
and U1160 (N_1160,N_745,N_540);
nand U1161 (N_1161,N_609,N_836);
and U1162 (N_1162,N_834,N_787);
or U1163 (N_1163,N_802,N_965);
and U1164 (N_1164,N_611,N_790);
nor U1165 (N_1165,N_985,N_762);
nand U1166 (N_1166,N_520,N_695);
and U1167 (N_1167,N_533,N_831);
nor U1168 (N_1168,N_659,N_592);
or U1169 (N_1169,N_698,N_880);
and U1170 (N_1170,N_701,N_862);
nand U1171 (N_1171,N_837,N_919);
nor U1172 (N_1172,N_584,N_535);
or U1173 (N_1173,N_577,N_897);
or U1174 (N_1174,N_874,N_747);
nor U1175 (N_1175,N_987,N_541);
nand U1176 (N_1176,N_665,N_632);
nor U1177 (N_1177,N_908,N_945);
and U1178 (N_1178,N_828,N_858);
nor U1179 (N_1179,N_649,N_861);
or U1180 (N_1180,N_622,N_754);
nor U1181 (N_1181,N_542,N_851);
or U1182 (N_1182,N_573,N_640);
nand U1183 (N_1183,N_907,N_709);
nand U1184 (N_1184,N_803,N_825);
or U1185 (N_1185,N_512,N_593);
nand U1186 (N_1186,N_866,N_895);
nor U1187 (N_1187,N_786,N_797);
nand U1188 (N_1188,N_775,N_716);
nor U1189 (N_1189,N_867,N_556);
or U1190 (N_1190,N_732,N_684);
nor U1191 (N_1191,N_870,N_829);
or U1192 (N_1192,N_875,N_769);
nor U1193 (N_1193,N_805,N_792);
or U1194 (N_1194,N_625,N_900);
nand U1195 (N_1195,N_748,N_696);
nor U1196 (N_1196,N_940,N_976);
nand U1197 (N_1197,N_531,N_891);
nor U1198 (N_1198,N_564,N_712);
and U1199 (N_1199,N_869,N_983);
and U1200 (N_1200,N_595,N_624);
and U1201 (N_1201,N_667,N_734);
nor U1202 (N_1202,N_872,N_604);
or U1203 (N_1203,N_782,N_962);
or U1204 (N_1204,N_680,N_552);
or U1205 (N_1205,N_509,N_682);
nor U1206 (N_1206,N_934,N_658);
and U1207 (N_1207,N_688,N_587);
nand U1208 (N_1208,N_623,N_911);
nor U1209 (N_1209,N_670,N_884);
nand U1210 (N_1210,N_537,N_841);
or U1211 (N_1211,N_980,N_903);
and U1212 (N_1212,N_597,N_746);
nor U1213 (N_1213,N_633,N_522);
nor U1214 (N_1214,N_843,N_539);
or U1215 (N_1215,N_998,N_613);
and U1216 (N_1216,N_574,N_538);
or U1217 (N_1217,N_928,N_988);
xor U1218 (N_1218,N_902,N_550);
nor U1219 (N_1219,N_883,N_949);
and U1220 (N_1220,N_984,N_721);
and U1221 (N_1221,N_679,N_720);
nand U1222 (N_1222,N_848,N_989);
nor U1223 (N_1223,N_502,N_818);
nand U1224 (N_1224,N_652,N_879);
or U1225 (N_1225,N_808,N_971);
nand U1226 (N_1226,N_821,N_753);
and U1227 (N_1227,N_663,N_605);
and U1228 (N_1228,N_674,N_646);
nand U1229 (N_1229,N_960,N_995);
and U1230 (N_1230,N_661,N_513);
or U1231 (N_1231,N_941,N_505);
nand U1232 (N_1232,N_981,N_619);
nand U1233 (N_1233,N_606,N_726);
nor U1234 (N_1234,N_967,N_953);
nand U1235 (N_1235,N_500,N_930);
and U1236 (N_1236,N_567,N_932);
nor U1237 (N_1237,N_785,N_815);
or U1238 (N_1238,N_733,N_642);
or U1239 (N_1239,N_865,N_707);
and U1240 (N_1240,N_968,N_877);
and U1241 (N_1241,N_906,N_957);
nor U1242 (N_1242,N_920,N_668);
or U1243 (N_1243,N_798,N_524);
and U1244 (N_1244,N_563,N_927);
nand U1245 (N_1245,N_796,N_951);
or U1246 (N_1246,N_628,N_711);
nor U1247 (N_1247,N_553,N_691);
nor U1248 (N_1248,N_794,N_832);
nor U1249 (N_1249,N_770,N_893);
nor U1250 (N_1250,N_953,N_749);
and U1251 (N_1251,N_858,N_812);
nand U1252 (N_1252,N_902,N_779);
nor U1253 (N_1253,N_901,N_758);
nor U1254 (N_1254,N_798,N_762);
or U1255 (N_1255,N_624,N_509);
and U1256 (N_1256,N_903,N_887);
or U1257 (N_1257,N_505,N_557);
nor U1258 (N_1258,N_583,N_674);
or U1259 (N_1259,N_785,N_590);
and U1260 (N_1260,N_675,N_598);
and U1261 (N_1261,N_733,N_937);
nand U1262 (N_1262,N_994,N_657);
nor U1263 (N_1263,N_732,N_654);
nor U1264 (N_1264,N_539,N_635);
nor U1265 (N_1265,N_857,N_897);
or U1266 (N_1266,N_865,N_617);
and U1267 (N_1267,N_756,N_594);
and U1268 (N_1268,N_746,N_889);
nor U1269 (N_1269,N_714,N_791);
or U1270 (N_1270,N_813,N_781);
or U1271 (N_1271,N_608,N_561);
nand U1272 (N_1272,N_847,N_917);
or U1273 (N_1273,N_820,N_934);
or U1274 (N_1274,N_562,N_690);
and U1275 (N_1275,N_704,N_777);
or U1276 (N_1276,N_575,N_743);
and U1277 (N_1277,N_958,N_868);
or U1278 (N_1278,N_864,N_718);
nand U1279 (N_1279,N_979,N_871);
and U1280 (N_1280,N_625,N_870);
and U1281 (N_1281,N_942,N_658);
nor U1282 (N_1282,N_600,N_754);
and U1283 (N_1283,N_678,N_680);
nand U1284 (N_1284,N_735,N_653);
or U1285 (N_1285,N_909,N_724);
or U1286 (N_1286,N_810,N_633);
nor U1287 (N_1287,N_602,N_554);
nand U1288 (N_1288,N_876,N_762);
nand U1289 (N_1289,N_887,N_697);
nand U1290 (N_1290,N_505,N_520);
and U1291 (N_1291,N_956,N_677);
or U1292 (N_1292,N_907,N_647);
and U1293 (N_1293,N_616,N_775);
nand U1294 (N_1294,N_673,N_565);
nor U1295 (N_1295,N_690,N_689);
nand U1296 (N_1296,N_951,N_818);
or U1297 (N_1297,N_689,N_544);
or U1298 (N_1298,N_588,N_855);
nand U1299 (N_1299,N_832,N_562);
and U1300 (N_1300,N_747,N_642);
nor U1301 (N_1301,N_675,N_774);
nor U1302 (N_1302,N_505,N_895);
or U1303 (N_1303,N_635,N_835);
or U1304 (N_1304,N_642,N_664);
or U1305 (N_1305,N_950,N_720);
and U1306 (N_1306,N_652,N_818);
nand U1307 (N_1307,N_562,N_647);
or U1308 (N_1308,N_646,N_526);
nor U1309 (N_1309,N_951,N_711);
and U1310 (N_1310,N_518,N_661);
and U1311 (N_1311,N_576,N_992);
or U1312 (N_1312,N_552,N_981);
nand U1313 (N_1313,N_811,N_970);
or U1314 (N_1314,N_950,N_669);
or U1315 (N_1315,N_947,N_849);
nand U1316 (N_1316,N_525,N_845);
and U1317 (N_1317,N_848,N_688);
or U1318 (N_1318,N_524,N_636);
nor U1319 (N_1319,N_737,N_923);
nor U1320 (N_1320,N_637,N_556);
and U1321 (N_1321,N_970,N_738);
or U1322 (N_1322,N_850,N_929);
nor U1323 (N_1323,N_708,N_629);
or U1324 (N_1324,N_879,N_634);
or U1325 (N_1325,N_602,N_783);
and U1326 (N_1326,N_888,N_640);
or U1327 (N_1327,N_651,N_854);
or U1328 (N_1328,N_605,N_742);
or U1329 (N_1329,N_835,N_768);
nand U1330 (N_1330,N_654,N_765);
or U1331 (N_1331,N_700,N_970);
or U1332 (N_1332,N_909,N_834);
nand U1333 (N_1333,N_804,N_677);
and U1334 (N_1334,N_781,N_902);
nand U1335 (N_1335,N_824,N_742);
or U1336 (N_1336,N_536,N_841);
and U1337 (N_1337,N_510,N_638);
nand U1338 (N_1338,N_824,N_523);
and U1339 (N_1339,N_509,N_795);
nor U1340 (N_1340,N_642,N_624);
nand U1341 (N_1341,N_737,N_523);
and U1342 (N_1342,N_539,N_839);
nor U1343 (N_1343,N_918,N_966);
and U1344 (N_1344,N_952,N_660);
nand U1345 (N_1345,N_577,N_671);
or U1346 (N_1346,N_866,N_574);
or U1347 (N_1347,N_600,N_503);
or U1348 (N_1348,N_708,N_720);
nand U1349 (N_1349,N_854,N_992);
nand U1350 (N_1350,N_721,N_680);
nand U1351 (N_1351,N_857,N_583);
nor U1352 (N_1352,N_823,N_952);
nor U1353 (N_1353,N_851,N_821);
and U1354 (N_1354,N_530,N_944);
nand U1355 (N_1355,N_892,N_820);
or U1356 (N_1356,N_518,N_966);
and U1357 (N_1357,N_616,N_963);
or U1358 (N_1358,N_818,N_884);
or U1359 (N_1359,N_661,N_605);
or U1360 (N_1360,N_924,N_543);
nand U1361 (N_1361,N_839,N_983);
and U1362 (N_1362,N_838,N_725);
nand U1363 (N_1363,N_545,N_773);
or U1364 (N_1364,N_885,N_859);
nand U1365 (N_1365,N_521,N_556);
nor U1366 (N_1366,N_683,N_944);
nand U1367 (N_1367,N_610,N_995);
and U1368 (N_1368,N_698,N_957);
nor U1369 (N_1369,N_675,N_574);
and U1370 (N_1370,N_786,N_982);
and U1371 (N_1371,N_557,N_670);
nor U1372 (N_1372,N_740,N_716);
nand U1373 (N_1373,N_669,N_633);
nand U1374 (N_1374,N_757,N_625);
nand U1375 (N_1375,N_740,N_598);
and U1376 (N_1376,N_889,N_774);
or U1377 (N_1377,N_704,N_987);
and U1378 (N_1378,N_630,N_811);
nand U1379 (N_1379,N_578,N_620);
nand U1380 (N_1380,N_638,N_747);
and U1381 (N_1381,N_722,N_709);
or U1382 (N_1382,N_798,N_576);
nor U1383 (N_1383,N_997,N_550);
or U1384 (N_1384,N_901,N_965);
nor U1385 (N_1385,N_660,N_566);
nor U1386 (N_1386,N_605,N_804);
or U1387 (N_1387,N_787,N_999);
or U1388 (N_1388,N_983,N_939);
and U1389 (N_1389,N_736,N_623);
and U1390 (N_1390,N_873,N_747);
or U1391 (N_1391,N_840,N_566);
nor U1392 (N_1392,N_859,N_673);
and U1393 (N_1393,N_961,N_981);
nor U1394 (N_1394,N_836,N_963);
and U1395 (N_1395,N_705,N_809);
xor U1396 (N_1396,N_510,N_535);
nand U1397 (N_1397,N_708,N_570);
or U1398 (N_1398,N_561,N_598);
and U1399 (N_1399,N_982,N_931);
and U1400 (N_1400,N_509,N_928);
nand U1401 (N_1401,N_656,N_503);
or U1402 (N_1402,N_917,N_615);
nor U1403 (N_1403,N_662,N_850);
and U1404 (N_1404,N_624,N_827);
nor U1405 (N_1405,N_826,N_876);
nand U1406 (N_1406,N_746,N_922);
and U1407 (N_1407,N_850,N_990);
nor U1408 (N_1408,N_568,N_744);
nand U1409 (N_1409,N_551,N_627);
nor U1410 (N_1410,N_936,N_701);
nor U1411 (N_1411,N_752,N_840);
nand U1412 (N_1412,N_628,N_944);
and U1413 (N_1413,N_692,N_504);
nor U1414 (N_1414,N_987,N_904);
or U1415 (N_1415,N_940,N_796);
nand U1416 (N_1416,N_969,N_866);
and U1417 (N_1417,N_694,N_663);
and U1418 (N_1418,N_801,N_524);
xnor U1419 (N_1419,N_962,N_833);
and U1420 (N_1420,N_611,N_705);
nand U1421 (N_1421,N_713,N_876);
and U1422 (N_1422,N_691,N_509);
nand U1423 (N_1423,N_925,N_885);
nor U1424 (N_1424,N_847,N_899);
nor U1425 (N_1425,N_515,N_658);
and U1426 (N_1426,N_865,N_689);
nand U1427 (N_1427,N_548,N_692);
nand U1428 (N_1428,N_769,N_755);
and U1429 (N_1429,N_783,N_914);
nor U1430 (N_1430,N_886,N_608);
and U1431 (N_1431,N_962,N_792);
nand U1432 (N_1432,N_558,N_734);
and U1433 (N_1433,N_807,N_977);
or U1434 (N_1434,N_626,N_885);
and U1435 (N_1435,N_886,N_512);
or U1436 (N_1436,N_594,N_750);
nand U1437 (N_1437,N_975,N_956);
nand U1438 (N_1438,N_792,N_586);
and U1439 (N_1439,N_524,N_506);
or U1440 (N_1440,N_997,N_762);
and U1441 (N_1441,N_562,N_521);
nor U1442 (N_1442,N_609,N_550);
and U1443 (N_1443,N_750,N_661);
nor U1444 (N_1444,N_906,N_572);
nor U1445 (N_1445,N_541,N_666);
nand U1446 (N_1446,N_976,N_954);
and U1447 (N_1447,N_637,N_752);
xnor U1448 (N_1448,N_552,N_955);
or U1449 (N_1449,N_643,N_682);
xor U1450 (N_1450,N_874,N_808);
nor U1451 (N_1451,N_513,N_704);
nor U1452 (N_1452,N_515,N_742);
and U1453 (N_1453,N_502,N_846);
nand U1454 (N_1454,N_905,N_770);
or U1455 (N_1455,N_521,N_780);
nor U1456 (N_1456,N_678,N_596);
nor U1457 (N_1457,N_693,N_987);
nand U1458 (N_1458,N_716,N_691);
nand U1459 (N_1459,N_539,N_762);
nor U1460 (N_1460,N_664,N_763);
nor U1461 (N_1461,N_614,N_663);
or U1462 (N_1462,N_782,N_773);
or U1463 (N_1463,N_938,N_848);
and U1464 (N_1464,N_784,N_701);
nor U1465 (N_1465,N_703,N_535);
nand U1466 (N_1466,N_963,N_955);
nor U1467 (N_1467,N_647,N_539);
nand U1468 (N_1468,N_593,N_985);
nor U1469 (N_1469,N_716,N_684);
nor U1470 (N_1470,N_536,N_747);
nand U1471 (N_1471,N_898,N_768);
nor U1472 (N_1472,N_653,N_749);
nor U1473 (N_1473,N_629,N_752);
and U1474 (N_1474,N_771,N_895);
and U1475 (N_1475,N_743,N_714);
and U1476 (N_1476,N_678,N_613);
or U1477 (N_1477,N_572,N_896);
nand U1478 (N_1478,N_960,N_897);
nand U1479 (N_1479,N_503,N_540);
nand U1480 (N_1480,N_650,N_864);
nor U1481 (N_1481,N_642,N_707);
nand U1482 (N_1482,N_877,N_630);
or U1483 (N_1483,N_662,N_966);
nand U1484 (N_1484,N_801,N_967);
nand U1485 (N_1485,N_867,N_821);
nor U1486 (N_1486,N_842,N_725);
and U1487 (N_1487,N_684,N_681);
xnor U1488 (N_1488,N_639,N_969);
and U1489 (N_1489,N_738,N_873);
or U1490 (N_1490,N_970,N_645);
xor U1491 (N_1491,N_506,N_642);
and U1492 (N_1492,N_889,N_601);
or U1493 (N_1493,N_727,N_794);
or U1494 (N_1494,N_608,N_962);
and U1495 (N_1495,N_884,N_618);
nand U1496 (N_1496,N_538,N_582);
nor U1497 (N_1497,N_980,N_694);
nand U1498 (N_1498,N_879,N_711);
nand U1499 (N_1499,N_525,N_889);
or U1500 (N_1500,N_1260,N_1365);
nor U1501 (N_1501,N_1085,N_1103);
or U1502 (N_1502,N_1189,N_1113);
nor U1503 (N_1503,N_1013,N_1056);
nor U1504 (N_1504,N_1356,N_1106);
or U1505 (N_1505,N_1472,N_1035);
or U1506 (N_1506,N_1053,N_1436);
or U1507 (N_1507,N_1294,N_1007);
or U1508 (N_1508,N_1425,N_1208);
or U1509 (N_1509,N_1458,N_1327);
and U1510 (N_1510,N_1027,N_1468);
and U1511 (N_1511,N_1201,N_1074);
nor U1512 (N_1512,N_1457,N_1369);
or U1513 (N_1513,N_1123,N_1387);
xor U1514 (N_1514,N_1192,N_1343);
and U1515 (N_1515,N_1128,N_1338);
nand U1516 (N_1516,N_1159,N_1291);
nor U1517 (N_1517,N_1471,N_1401);
nand U1518 (N_1518,N_1492,N_1042);
nand U1519 (N_1519,N_1317,N_1153);
or U1520 (N_1520,N_1107,N_1301);
nand U1521 (N_1521,N_1015,N_1309);
or U1522 (N_1522,N_1494,N_1202);
or U1523 (N_1523,N_1269,N_1336);
nor U1524 (N_1524,N_1377,N_1353);
nor U1525 (N_1525,N_1210,N_1285);
and U1526 (N_1526,N_1233,N_1245);
and U1527 (N_1527,N_1080,N_1034);
nor U1528 (N_1528,N_1332,N_1177);
and U1529 (N_1529,N_1479,N_1094);
and U1530 (N_1530,N_1212,N_1299);
xor U1531 (N_1531,N_1328,N_1121);
and U1532 (N_1532,N_1137,N_1429);
or U1533 (N_1533,N_1219,N_1360);
nor U1534 (N_1534,N_1049,N_1200);
or U1535 (N_1535,N_1138,N_1489);
nor U1536 (N_1536,N_1428,N_1297);
nor U1537 (N_1537,N_1061,N_1033);
and U1538 (N_1538,N_1431,N_1258);
or U1539 (N_1539,N_1131,N_1071);
nand U1540 (N_1540,N_1247,N_1079);
nand U1541 (N_1541,N_1043,N_1300);
or U1542 (N_1542,N_1312,N_1046);
or U1543 (N_1543,N_1059,N_1213);
nor U1544 (N_1544,N_1461,N_1073);
and U1545 (N_1545,N_1054,N_1198);
nor U1546 (N_1546,N_1023,N_1354);
and U1547 (N_1547,N_1286,N_1483);
or U1548 (N_1548,N_1270,N_1237);
and U1549 (N_1549,N_1382,N_1325);
nor U1550 (N_1550,N_1149,N_1413);
nand U1551 (N_1551,N_1157,N_1333);
and U1552 (N_1552,N_1124,N_1273);
nor U1553 (N_1553,N_1306,N_1344);
nand U1554 (N_1554,N_1481,N_1216);
or U1555 (N_1555,N_1319,N_1040);
nor U1556 (N_1556,N_1064,N_1257);
or U1557 (N_1557,N_1278,N_1181);
nand U1558 (N_1558,N_1199,N_1417);
and U1559 (N_1559,N_1434,N_1018);
nand U1560 (N_1560,N_1251,N_1024);
or U1561 (N_1561,N_1029,N_1437);
or U1562 (N_1562,N_1359,N_1254);
and U1563 (N_1563,N_1133,N_1112);
and U1564 (N_1564,N_1290,N_1057);
nand U1565 (N_1565,N_1229,N_1308);
nand U1566 (N_1566,N_1125,N_1261);
or U1567 (N_1567,N_1409,N_1065);
nor U1568 (N_1568,N_1069,N_1384);
or U1569 (N_1569,N_1490,N_1135);
nand U1570 (N_1570,N_1398,N_1322);
or U1571 (N_1571,N_1324,N_1364);
or U1572 (N_1572,N_1066,N_1423);
nor U1573 (N_1573,N_1185,N_1067);
or U1574 (N_1574,N_1313,N_1187);
nand U1575 (N_1575,N_1008,N_1030);
nor U1576 (N_1576,N_1321,N_1420);
nand U1577 (N_1577,N_1090,N_1218);
nor U1578 (N_1578,N_1418,N_1389);
xor U1579 (N_1579,N_1086,N_1150);
and U1580 (N_1580,N_1476,N_1039);
and U1581 (N_1581,N_1275,N_1051);
nor U1582 (N_1582,N_1170,N_1182);
or U1583 (N_1583,N_1304,N_1174);
nor U1584 (N_1584,N_1021,N_1419);
nand U1585 (N_1585,N_1371,N_1142);
and U1586 (N_1586,N_1380,N_1316);
nor U1587 (N_1587,N_1443,N_1292);
nand U1588 (N_1588,N_1412,N_1005);
and U1589 (N_1589,N_1228,N_1088);
nor U1590 (N_1590,N_1068,N_1076);
or U1591 (N_1591,N_1406,N_1209);
nand U1592 (N_1592,N_1427,N_1438);
and U1593 (N_1593,N_1224,N_1100);
and U1594 (N_1594,N_1392,N_1196);
and U1595 (N_1595,N_1102,N_1108);
nor U1596 (N_1596,N_1173,N_1156);
or U1597 (N_1597,N_1357,N_1098);
and U1598 (N_1598,N_1204,N_1063);
nor U1599 (N_1599,N_1320,N_1478);
or U1600 (N_1600,N_1404,N_1227);
or U1601 (N_1601,N_1282,N_1176);
nand U1602 (N_1602,N_1114,N_1127);
nand U1603 (N_1603,N_1161,N_1315);
nand U1604 (N_1604,N_1014,N_1310);
nand U1605 (N_1605,N_1383,N_1424);
nor U1606 (N_1606,N_1238,N_1435);
or U1607 (N_1607,N_1195,N_1462);
and U1608 (N_1608,N_1144,N_1400);
nand U1609 (N_1609,N_1330,N_1265);
nand U1610 (N_1610,N_1442,N_1239);
and U1611 (N_1611,N_1243,N_1367);
and U1612 (N_1612,N_1298,N_1263);
nor U1613 (N_1613,N_1047,N_1256);
nand U1614 (N_1614,N_1231,N_1496);
nand U1615 (N_1615,N_1140,N_1000);
and U1616 (N_1616,N_1451,N_1129);
nor U1617 (N_1617,N_1498,N_1329);
nor U1618 (N_1618,N_1197,N_1175);
or U1619 (N_1619,N_1397,N_1370);
and U1620 (N_1620,N_1183,N_1482);
or U1621 (N_1621,N_1394,N_1101);
nor U1622 (N_1622,N_1395,N_1337);
or U1623 (N_1623,N_1352,N_1342);
and U1624 (N_1624,N_1019,N_1002);
or U1625 (N_1625,N_1050,N_1164);
nand U1626 (N_1626,N_1115,N_1266);
nor U1627 (N_1627,N_1485,N_1255);
or U1628 (N_1628,N_1154,N_1178);
nor U1629 (N_1629,N_1440,N_1407);
nor U1630 (N_1630,N_1277,N_1334);
or U1631 (N_1631,N_1248,N_1465);
nand U1632 (N_1632,N_1032,N_1441);
nor U1633 (N_1633,N_1141,N_1044);
or U1634 (N_1634,N_1403,N_1143);
nor U1635 (N_1635,N_1193,N_1293);
or U1636 (N_1636,N_1408,N_1349);
nand U1637 (N_1637,N_1318,N_1460);
nor U1638 (N_1638,N_1152,N_1084);
and U1639 (N_1639,N_1411,N_1473);
or U1640 (N_1640,N_1484,N_1346);
or U1641 (N_1641,N_1022,N_1323);
nor U1642 (N_1642,N_1001,N_1048);
nor U1643 (N_1643,N_1362,N_1004);
nor U1644 (N_1644,N_1296,N_1045);
or U1645 (N_1645,N_1072,N_1388);
nand U1646 (N_1646,N_1188,N_1259);
or U1647 (N_1647,N_1486,N_1347);
and U1648 (N_1648,N_1003,N_1410);
nor U1649 (N_1649,N_1314,N_1466);
nor U1650 (N_1650,N_1405,N_1279);
nand U1651 (N_1651,N_1374,N_1130);
or U1652 (N_1652,N_1276,N_1366);
and U1653 (N_1653,N_1038,N_1117);
nor U1654 (N_1654,N_1363,N_1160);
and U1655 (N_1655,N_1455,N_1077);
nand U1656 (N_1656,N_1151,N_1017);
and U1657 (N_1657,N_1006,N_1081);
nand U1658 (N_1658,N_1381,N_1221);
nand U1659 (N_1659,N_1469,N_1093);
nand U1660 (N_1660,N_1244,N_1268);
nor U1661 (N_1661,N_1391,N_1262);
or U1662 (N_1662,N_1223,N_1126);
or U1663 (N_1663,N_1110,N_1155);
nor U1664 (N_1664,N_1163,N_1280);
or U1665 (N_1665,N_1305,N_1236);
nor U1666 (N_1666,N_1132,N_1104);
nor U1667 (N_1667,N_1497,N_1119);
or U1668 (N_1668,N_1012,N_1378);
or U1669 (N_1669,N_1096,N_1480);
nor U1670 (N_1670,N_1288,N_1186);
or U1671 (N_1671,N_1097,N_1162);
nor U1672 (N_1672,N_1295,N_1060);
or U1673 (N_1673,N_1220,N_1134);
nor U1674 (N_1674,N_1439,N_1477);
nand U1675 (N_1675,N_1241,N_1303);
and U1676 (N_1676,N_1158,N_1105);
or U1677 (N_1677,N_1272,N_1190);
or U1678 (N_1678,N_1087,N_1331);
or U1679 (N_1679,N_1009,N_1267);
or U1680 (N_1680,N_1444,N_1373);
or U1681 (N_1681,N_1368,N_1326);
nand U1682 (N_1682,N_1116,N_1399);
and U1683 (N_1683,N_1385,N_1311);
nand U1684 (N_1684,N_1414,N_1172);
and U1685 (N_1685,N_1345,N_1355);
nand U1686 (N_1686,N_1026,N_1390);
nor U1687 (N_1687,N_1205,N_1184);
and U1688 (N_1688,N_1350,N_1083);
and U1689 (N_1689,N_1148,N_1415);
nor U1690 (N_1690,N_1307,N_1230);
nor U1691 (N_1691,N_1463,N_1171);
or U1692 (N_1692,N_1448,N_1235);
nor U1693 (N_1693,N_1136,N_1372);
nor U1694 (N_1694,N_1206,N_1491);
nand U1695 (N_1695,N_1341,N_1456);
nand U1696 (N_1696,N_1445,N_1447);
and U1697 (N_1697,N_1459,N_1283);
nor U1698 (N_1698,N_1139,N_1426);
nor U1699 (N_1699,N_1335,N_1453);
and U1700 (N_1700,N_1253,N_1393);
and U1701 (N_1701,N_1433,N_1179);
nand U1702 (N_1702,N_1488,N_1055);
nand U1703 (N_1703,N_1169,N_1089);
or U1704 (N_1704,N_1240,N_1474);
nand U1705 (N_1705,N_1207,N_1339);
nor U1706 (N_1706,N_1422,N_1016);
nand U1707 (N_1707,N_1109,N_1430);
or U1708 (N_1708,N_1493,N_1416);
nand U1709 (N_1709,N_1289,N_1249);
nand U1710 (N_1710,N_1470,N_1348);
and U1711 (N_1711,N_1250,N_1284);
nor U1712 (N_1712,N_1041,N_1287);
or U1713 (N_1713,N_1421,N_1234);
nand U1714 (N_1714,N_1075,N_1215);
nor U1715 (N_1715,N_1246,N_1099);
and U1716 (N_1716,N_1180,N_1203);
nor U1717 (N_1717,N_1111,N_1225);
nand U1718 (N_1718,N_1122,N_1010);
and U1719 (N_1719,N_1052,N_1058);
and U1720 (N_1720,N_1351,N_1467);
and U1721 (N_1721,N_1464,N_1217);
or U1722 (N_1722,N_1031,N_1036);
nor U1723 (N_1723,N_1147,N_1167);
and U1724 (N_1724,N_1226,N_1062);
or U1725 (N_1725,N_1449,N_1222);
or U1726 (N_1726,N_1037,N_1450);
and U1727 (N_1727,N_1194,N_1302);
or U1728 (N_1728,N_1120,N_1487);
or U1729 (N_1729,N_1166,N_1028);
nand U1730 (N_1730,N_1242,N_1271);
or U1731 (N_1731,N_1402,N_1446);
or U1732 (N_1732,N_1214,N_1091);
nand U1733 (N_1733,N_1252,N_1211);
nor U1734 (N_1734,N_1145,N_1452);
nor U1735 (N_1735,N_1432,N_1095);
nand U1736 (N_1736,N_1025,N_1168);
or U1737 (N_1737,N_1118,N_1232);
and U1738 (N_1738,N_1376,N_1191);
nor U1739 (N_1739,N_1375,N_1165);
or U1740 (N_1740,N_1020,N_1281);
and U1741 (N_1741,N_1379,N_1495);
nand U1742 (N_1742,N_1475,N_1082);
and U1743 (N_1743,N_1386,N_1358);
nor U1744 (N_1744,N_1274,N_1264);
and U1745 (N_1745,N_1092,N_1146);
nand U1746 (N_1746,N_1070,N_1454);
nor U1747 (N_1747,N_1396,N_1011);
and U1748 (N_1748,N_1499,N_1361);
nand U1749 (N_1749,N_1340,N_1078);
and U1750 (N_1750,N_1104,N_1338);
and U1751 (N_1751,N_1166,N_1109);
nand U1752 (N_1752,N_1185,N_1333);
nor U1753 (N_1753,N_1045,N_1499);
nand U1754 (N_1754,N_1122,N_1280);
nand U1755 (N_1755,N_1389,N_1214);
or U1756 (N_1756,N_1278,N_1393);
nand U1757 (N_1757,N_1221,N_1093);
and U1758 (N_1758,N_1403,N_1012);
and U1759 (N_1759,N_1126,N_1423);
xnor U1760 (N_1760,N_1281,N_1190);
nand U1761 (N_1761,N_1432,N_1420);
or U1762 (N_1762,N_1146,N_1197);
and U1763 (N_1763,N_1450,N_1241);
nor U1764 (N_1764,N_1465,N_1327);
nor U1765 (N_1765,N_1348,N_1456);
nand U1766 (N_1766,N_1251,N_1413);
and U1767 (N_1767,N_1459,N_1369);
nor U1768 (N_1768,N_1285,N_1378);
nor U1769 (N_1769,N_1354,N_1369);
nor U1770 (N_1770,N_1376,N_1204);
or U1771 (N_1771,N_1330,N_1397);
and U1772 (N_1772,N_1256,N_1167);
or U1773 (N_1773,N_1358,N_1122);
or U1774 (N_1774,N_1444,N_1056);
or U1775 (N_1775,N_1050,N_1221);
nor U1776 (N_1776,N_1469,N_1179);
nand U1777 (N_1777,N_1138,N_1010);
or U1778 (N_1778,N_1137,N_1446);
and U1779 (N_1779,N_1045,N_1023);
or U1780 (N_1780,N_1156,N_1224);
and U1781 (N_1781,N_1069,N_1273);
nand U1782 (N_1782,N_1143,N_1242);
nor U1783 (N_1783,N_1107,N_1313);
or U1784 (N_1784,N_1489,N_1361);
nand U1785 (N_1785,N_1007,N_1385);
or U1786 (N_1786,N_1291,N_1218);
nor U1787 (N_1787,N_1206,N_1066);
or U1788 (N_1788,N_1236,N_1113);
nor U1789 (N_1789,N_1006,N_1375);
or U1790 (N_1790,N_1152,N_1176);
and U1791 (N_1791,N_1218,N_1034);
and U1792 (N_1792,N_1230,N_1030);
or U1793 (N_1793,N_1270,N_1437);
nor U1794 (N_1794,N_1444,N_1499);
and U1795 (N_1795,N_1106,N_1432);
and U1796 (N_1796,N_1230,N_1365);
nor U1797 (N_1797,N_1439,N_1127);
and U1798 (N_1798,N_1343,N_1057);
or U1799 (N_1799,N_1212,N_1286);
xor U1800 (N_1800,N_1497,N_1111);
or U1801 (N_1801,N_1144,N_1108);
nand U1802 (N_1802,N_1231,N_1340);
nand U1803 (N_1803,N_1454,N_1256);
nor U1804 (N_1804,N_1171,N_1150);
and U1805 (N_1805,N_1264,N_1425);
xnor U1806 (N_1806,N_1152,N_1486);
or U1807 (N_1807,N_1147,N_1049);
nand U1808 (N_1808,N_1379,N_1434);
and U1809 (N_1809,N_1171,N_1348);
and U1810 (N_1810,N_1430,N_1034);
nor U1811 (N_1811,N_1473,N_1162);
or U1812 (N_1812,N_1403,N_1007);
nand U1813 (N_1813,N_1491,N_1477);
nor U1814 (N_1814,N_1078,N_1311);
or U1815 (N_1815,N_1321,N_1177);
and U1816 (N_1816,N_1093,N_1293);
nand U1817 (N_1817,N_1377,N_1173);
nor U1818 (N_1818,N_1025,N_1287);
nand U1819 (N_1819,N_1329,N_1107);
nand U1820 (N_1820,N_1068,N_1386);
nand U1821 (N_1821,N_1329,N_1473);
and U1822 (N_1822,N_1215,N_1225);
nor U1823 (N_1823,N_1298,N_1306);
or U1824 (N_1824,N_1430,N_1234);
nor U1825 (N_1825,N_1237,N_1432);
nor U1826 (N_1826,N_1190,N_1194);
and U1827 (N_1827,N_1325,N_1495);
or U1828 (N_1828,N_1412,N_1392);
or U1829 (N_1829,N_1474,N_1231);
or U1830 (N_1830,N_1298,N_1408);
or U1831 (N_1831,N_1214,N_1147);
or U1832 (N_1832,N_1223,N_1162);
nand U1833 (N_1833,N_1346,N_1331);
nor U1834 (N_1834,N_1267,N_1305);
nor U1835 (N_1835,N_1347,N_1274);
nand U1836 (N_1836,N_1084,N_1258);
nand U1837 (N_1837,N_1232,N_1270);
nand U1838 (N_1838,N_1400,N_1480);
and U1839 (N_1839,N_1160,N_1337);
or U1840 (N_1840,N_1218,N_1119);
nand U1841 (N_1841,N_1112,N_1282);
or U1842 (N_1842,N_1424,N_1394);
nand U1843 (N_1843,N_1353,N_1150);
or U1844 (N_1844,N_1099,N_1108);
and U1845 (N_1845,N_1171,N_1473);
nor U1846 (N_1846,N_1451,N_1476);
and U1847 (N_1847,N_1356,N_1187);
or U1848 (N_1848,N_1220,N_1455);
or U1849 (N_1849,N_1128,N_1214);
or U1850 (N_1850,N_1054,N_1388);
and U1851 (N_1851,N_1442,N_1052);
nand U1852 (N_1852,N_1247,N_1191);
nor U1853 (N_1853,N_1432,N_1423);
nor U1854 (N_1854,N_1304,N_1055);
nor U1855 (N_1855,N_1493,N_1204);
or U1856 (N_1856,N_1249,N_1107);
nand U1857 (N_1857,N_1473,N_1228);
nor U1858 (N_1858,N_1005,N_1313);
and U1859 (N_1859,N_1193,N_1031);
or U1860 (N_1860,N_1224,N_1112);
nand U1861 (N_1861,N_1329,N_1088);
and U1862 (N_1862,N_1409,N_1401);
and U1863 (N_1863,N_1179,N_1396);
nor U1864 (N_1864,N_1444,N_1394);
nor U1865 (N_1865,N_1345,N_1485);
nor U1866 (N_1866,N_1007,N_1010);
and U1867 (N_1867,N_1409,N_1476);
nand U1868 (N_1868,N_1334,N_1032);
nor U1869 (N_1869,N_1156,N_1201);
or U1870 (N_1870,N_1233,N_1076);
nand U1871 (N_1871,N_1414,N_1002);
nor U1872 (N_1872,N_1023,N_1461);
or U1873 (N_1873,N_1014,N_1196);
or U1874 (N_1874,N_1338,N_1018);
nand U1875 (N_1875,N_1177,N_1083);
nor U1876 (N_1876,N_1143,N_1285);
nor U1877 (N_1877,N_1457,N_1449);
or U1878 (N_1878,N_1356,N_1358);
nand U1879 (N_1879,N_1424,N_1080);
or U1880 (N_1880,N_1250,N_1366);
and U1881 (N_1881,N_1138,N_1497);
and U1882 (N_1882,N_1083,N_1169);
and U1883 (N_1883,N_1307,N_1054);
or U1884 (N_1884,N_1205,N_1230);
xor U1885 (N_1885,N_1286,N_1324);
nand U1886 (N_1886,N_1273,N_1232);
nor U1887 (N_1887,N_1363,N_1278);
nor U1888 (N_1888,N_1079,N_1127);
and U1889 (N_1889,N_1421,N_1197);
and U1890 (N_1890,N_1056,N_1482);
nor U1891 (N_1891,N_1337,N_1433);
or U1892 (N_1892,N_1342,N_1098);
or U1893 (N_1893,N_1065,N_1006);
and U1894 (N_1894,N_1409,N_1455);
nor U1895 (N_1895,N_1277,N_1433);
and U1896 (N_1896,N_1480,N_1127);
nand U1897 (N_1897,N_1476,N_1230);
nor U1898 (N_1898,N_1110,N_1437);
and U1899 (N_1899,N_1299,N_1005);
nor U1900 (N_1900,N_1424,N_1466);
and U1901 (N_1901,N_1195,N_1383);
and U1902 (N_1902,N_1456,N_1200);
and U1903 (N_1903,N_1206,N_1464);
nand U1904 (N_1904,N_1289,N_1375);
or U1905 (N_1905,N_1020,N_1337);
or U1906 (N_1906,N_1036,N_1054);
nor U1907 (N_1907,N_1440,N_1169);
nand U1908 (N_1908,N_1258,N_1142);
or U1909 (N_1909,N_1306,N_1417);
and U1910 (N_1910,N_1490,N_1049);
or U1911 (N_1911,N_1055,N_1113);
nand U1912 (N_1912,N_1215,N_1259);
nand U1913 (N_1913,N_1391,N_1154);
or U1914 (N_1914,N_1364,N_1358);
nand U1915 (N_1915,N_1071,N_1201);
nor U1916 (N_1916,N_1284,N_1269);
or U1917 (N_1917,N_1063,N_1296);
nand U1918 (N_1918,N_1375,N_1272);
nor U1919 (N_1919,N_1161,N_1085);
and U1920 (N_1920,N_1005,N_1255);
or U1921 (N_1921,N_1308,N_1277);
and U1922 (N_1922,N_1451,N_1427);
nor U1923 (N_1923,N_1001,N_1487);
nand U1924 (N_1924,N_1235,N_1143);
or U1925 (N_1925,N_1099,N_1267);
nand U1926 (N_1926,N_1275,N_1157);
or U1927 (N_1927,N_1331,N_1145);
and U1928 (N_1928,N_1361,N_1098);
nor U1929 (N_1929,N_1292,N_1352);
or U1930 (N_1930,N_1351,N_1055);
and U1931 (N_1931,N_1396,N_1431);
and U1932 (N_1932,N_1219,N_1325);
nor U1933 (N_1933,N_1429,N_1086);
nand U1934 (N_1934,N_1216,N_1381);
nand U1935 (N_1935,N_1316,N_1051);
nor U1936 (N_1936,N_1439,N_1025);
nor U1937 (N_1937,N_1433,N_1128);
nand U1938 (N_1938,N_1344,N_1249);
and U1939 (N_1939,N_1267,N_1107);
and U1940 (N_1940,N_1086,N_1080);
or U1941 (N_1941,N_1227,N_1074);
or U1942 (N_1942,N_1434,N_1403);
nand U1943 (N_1943,N_1445,N_1138);
or U1944 (N_1944,N_1058,N_1486);
nor U1945 (N_1945,N_1087,N_1382);
and U1946 (N_1946,N_1447,N_1075);
and U1947 (N_1947,N_1452,N_1177);
or U1948 (N_1948,N_1108,N_1265);
or U1949 (N_1949,N_1049,N_1499);
or U1950 (N_1950,N_1430,N_1348);
nand U1951 (N_1951,N_1478,N_1232);
nand U1952 (N_1952,N_1302,N_1344);
and U1953 (N_1953,N_1158,N_1422);
and U1954 (N_1954,N_1333,N_1142);
nand U1955 (N_1955,N_1487,N_1185);
or U1956 (N_1956,N_1424,N_1396);
and U1957 (N_1957,N_1039,N_1029);
nor U1958 (N_1958,N_1325,N_1189);
and U1959 (N_1959,N_1224,N_1409);
or U1960 (N_1960,N_1047,N_1109);
nor U1961 (N_1961,N_1243,N_1286);
nor U1962 (N_1962,N_1039,N_1362);
and U1963 (N_1963,N_1037,N_1076);
nand U1964 (N_1964,N_1248,N_1173);
and U1965 (N_1965,N_1477,N_1258);
or U1966 (N_1966,N_1018,N_1040);
nor U1967 (N_1967,N_1361,N_1268);
and U1968 (N_1968,N_1338,N_1350);
nand U1969 (N_1969,N_1101,N_1465);
and U1970 (N_1970,N_1219,N_1300);
or U1971 (N_1971,N_1460,N_1132);
nand U1972 (N_1972,N_1280,N_1080);
nor U1973 (N_1973,N_1401,N_1220);
nor U1974 (N_1974,N_1341,N_1131);
nand U1975 (N_1975,N_1160,N_1066);
and U1976 (N_1976,N_1092,N_1135);
or U1977 (N_1977,N_1070,N_1094);
or U1978 (N_1978,N_1495,N_1163);
or U1979 (N_1979,N_1196,N_1225);
nand U1980 (N_1980,N_1390,N_1432);
and U1981 (N_1981,N_1241,N_1058);
or U1982 (N_1982,N_1137,N_1322);
nand U1983 (N_1983,N_1151,N_1452);
nand U1984 (N_1984,N_1244,N_1274);
nor U1985 (N_1985,N_1439,N_1364);
nand U1986 (N_1986,N_1223,N_1446);
nand U1987 (N_1987,N_1450,N_1279);
or U1988 (N_1988,N_1237,N_1488);
and U1989 (N_1989,N_1436,N_1352);
and U1990 (N_1990,N_1317,N_1236);
nand U1991 (N_1991,N_1429,N_1129);
and U1992 (N_1992,N_1466,N_1375);
and U1993 (N_1993,N_1084,N_1206);
or U1994 (N_1994,N_1251,N_1155);
and U1995 (N_1995,N_1417,N_1193);
and U1996 (N_1996,N_1237,N_1051);
and U1997 (N_1997,N_1088,N_1105);
xor U1998 (N_1998,N_1479,N_1408);
or U1999 (N_1999,N_1208,N_1420);
nor U2000 (N_2000,N_1982,N_1536);
nor U2001 (N_2001,N_1593,N_1797);
nand U2002 (N_2002,N_1796,N_1572);
nor U2003 (N_2003,N_1923,N_1583);
or U2004 (N_2004,N_1788,N_1943);
nor U2005 (N_2005,N_1612,N_1753);
nand U2006 (N_2006,N_1508,N_1743);
nand U2007 (N_2007,N_1546,N_1748);
nand U2008 (N_2008,N_1805,N_1920);
nand U2009 (N_2009,N_1847,N_1956);
nor U2010 (N_2010,N_1700,N_1927);
nor U2011 (N_2011,N_1934,N_1987);
and U2012 (N_2012,N_1651,N_1541);
nor U2013 (N_2013,N_1750,N_1878);
nor U2014 (N_2014,N_1992,N_1922);
or U2015 (N_2015,N_1532,N_1666);
nand U2016 (N_2016,N_1941,N_1655);
nor U2017 (N_2017,N_1886,N_1814);
nor U2018 (N_2018,N_1741,N_1607);
nor U2019 (N_2019,N_1798,N_1744);
and U2020 (N_2020,N_1818,N_1887);
nand U2021 (N_2021,N_1707,N_1642);
nor U2022 (N_2022,N_1527,N_1517);
nand U2023 (N_2023,N_1864,N_1767);
and U2024 (N_2024,N_1831,N_1617);
nand U2025 (N_2025,N_1795,N_1815);
and U2026 (N_2026,N_1658,N_1894);
nor U2027 (N_2027,N_1994,N_1984);
and U2028 (N_2028,N_1860,N_1513);
or U2029 (N_2029,N_1624,N_1530);
nor U2030 (N_2030,N_1812,N_1937);
nand U2031 (N_2031,N_1609,N_1938);
or U2032 (N_2032,N_1556,N_1919);
nor U2033 (N_2033,N_1697,N_1559);
nand U2034 (N_2034,N_1791,N_1543);
and U2035 (N_2035,N_1511,N_1951);
nor U2036 (N_2036,N_1710,N_1518);
or U2037 (N_2037,N_1787,N_1856);
nor U2038 (N_2038,N_1535,N_1545);
nand U2039 (N_2039,N_1998,N_1826);
or U2040 (N_2040,N_1501,N_1590);
nor U2041 (N_2041,N_1909,N_1824);
nor U2042 (N_2042,N_1936,N_1874);
or U2043 (N_2043,N_1602,N_1563);
or U2044 (N_2044,N_1865,N_1704);
nor U2045 (N_2045,N_1729,N_1686);
and U2046 (N_2046,N_1715,N_1684);
nand U2047 (N_2047,N_1505,N_1652);
and U2048 (N_2048,N_1678,N_1582);
or U2049 (N_2049,N_1544,N_1538);
nand U2050 (N_2050,N_1571,N_1746);
nor U2051 (N_2051,N_1846,N_1588);
or U2052 (N_2052,N_1575,N_1840);
nor U2053 (N_2053,N_1899,N_1755);
nand U2054 (N_2054,N_1808,N_1716);
or U2055 (N_2055,N_1876,N_1675);
nor U2056 (N_2056,N_1601,N_1599);
nor U2057 (N_2057,N_1683,N_1958);
and U2058 (N_2058,N_1685,N_1734);
and U2059 (N_2059,N_1890,N_1605);
nor U2060 (N_2060,N_1653,N_1830);
nor U2061 (N_2061,N_1529,N_1875);
nand U2062 (N_2062,N_1703,N_1918);
nand U2063 (N_2063,N_1695,N_1983);
nand U2064 (N_2064,N_1908,N_1644);
and U2065 (N_2065,N_1634,N_1576);
nor U2066 (N_2066,N_1964,N_1783);
nor U2067 (N_2067,N_1557,N_1680);
or U2068 (N_2068,N_1627,N_1589);
nor U2069 (N_2069,N_1573,N_1774);
and U2070 (N_2070,N_1647,N_1967);
nor U2071 (N_2071,N_1763,N_1821);
and U2072 (N_2072,N_1665,N_1639);
or U2073 (N_2073,N_1694,N_1502);
nor U2074 (N_2074,N_1737,N_1844);
or U2075 (N_2075,N_1528,N_1542);
or U2076 (N_2076,N_1731,N_1600);
or U2077 (N_2077,N_1777,N_1578);
and U2078 (N_2078,N_1819,N_1963);
or U2079 (N_2079,N_1570,N_1754);
nand U2080 (N_2080,N_1646,N_1628);
nor U2081 (N_2081,N_1620,N_1533);
nand U2082 (N_2082,N_1705,N_1884);
nor U2083 (N_2083,N_1671,N_1640);
or U2084 (N_2084,N_1900,N_1776);
and U2085 (N_2085,N_1650,N_1952);
and U2086 (N_2086,N_1991,N_1960);
and U2087 (N_2087,N_1801,N_1898);
nor U2088 (N_2088,N_1903,N_1577);
or U2089 (N_2089,N_1662,N_1661);
and U2090 (N_2090,N_1664,N_1891);
nor U2091 (N_2091,N_1723,N_1841);
nor U2092 (N_2092,N_1912,N_1515);
or U2093 (N_2093,N_1867,N_1550);
nand U2094 (N_2094,N_1727,N_1708);
or U2095 (N_2095,N_1955,N_1972);
or U2096 (N_2096,N_1591,N_1781);
xnor U2097 (N_2097,N_1828,N_1855);
or U2098 (N_2098,N_1782,N_1521);
nor U2099 (N_2099,N_1913,N_1523);
nand U2100 (N_2100,N_1946,N_1596);
nor U2101 (N_2101,N_1758,N_1825);
nor U2102 (N_2102,N_1733,N_1553);
or U2103 (N_2103,N_1977,N_1558);
nor U2104 (N_2104,N_1702,N_1713);
and U2105 (N_2105,N_1656,N_1822);
nor U2106 (N_2106,N_1659,N_1986);
nand U2107 (N_2107,N_1615,N_1608);
or U2108 (N_2108,N_1773,N_1693);
or U2109 (N_2109,N_1587,N_1872);
or U2110 (N_2110,N_1692,N_1929);
nand U2111 (N_2111,N_1962,N_1942);
xor U2112 (N_2112,N_1803,N_1981);
nand U2113 (N_2113,N_1949,N_1778);
nor U2114 (N_2114,N_1670,N_1806);
nand U2115 (N_2115,N_1724,N_1506);
or U2116 (N_2116,N_1722,N_1740);
or U2117 (N_2117,N_1838,N_1611);
and U2118 (N_2118,N_1732,N_1924);
nand U2119 (N_2119,N_1735,N_1745);
nor U2120 (N_2120,N_1807,N_1549);
or U2121 (N_2121,N_1638,N_1794);
or U2122 (N_2122,N_1931,N_1999);
nor U2123 (N_2123,N_1657,N_1579);
nand U2124 (N_2124,N_1779,N_1842);
and U2125 (N_2125,N_1669,N_1520);
nand U2126 (N_2126,N_1565,N_1809);
nand U2127 (N_2127,N_1827,N_1507);
and U2128 (N_2128,N_1691,N_1759);
nand U2129 (N_2129,N_1816,N_1622);
xor U2130 (N_2130,N_1548,N_1769);
and U2131 (N_2131,N_1712,N_1820);
nand U2132 (N_2132,N_1701,N_1663);
and U2133 (N_2133,N_1586,N_1711);
nor U2134 (N_2134,N_1562,N_1770);
or U2135 (N_2135,N_1630,N_1995);
nand U2136 (N_2136,N_1925,N_1973);
or U2137 (N_2137,N_1969,N_1836);
nand U2138 (N_2138,N_1585,N_1668);
or U2139 (N_2139,N_1673,N_1961);
or U2140 (N_2140,N_1682,N_1681);
and U2141 (N_2141,N_1905,N_1706);
nor U2142 (N_2142,N_1907,N_1861);
or U2143 (N_2143,N_1996,N_1643);
nand U2144 (N_2144,N_1858,N_1921);
nor U2145 (N_2145,N_1804,N_1896);
or U2146 (N_2146,N_1930,N_1749);
or U2147 (N_2147,N_1785,N_1928);
nor U2148 (N_2148,N_1954,N_1997);
nor U2149 (N_2149,N_1736,N_1793);
and U2150 (N_2150,N_1747,N_1944);
and U2151 (N_2151,N_1574,N_1833);
nand U2152 (N_2152,N_1834,N_1879);
nor U2153 (N_2153,N_1676,N_1854);
nand U2154 (N_2154,N_1771,N_1689);
nor U2155 (N_2155,N_1939,N_1568);
nand U2156 (N_2156,N_1619,N_1914);
nor U2157 (N_2157,N_1623,N_1539);
or U2158 (N_2158,N_1714,N_1728);
nor U2159 (N_2159,N_1592,N_1832);
or U2160 (N_2160,N_1613,N_1618);
and U2161 (N_2161,N_1677,N_1885);
and U2162 (N_2162,N_1957,N_1911);
nor U2163 (N_2163,N_1567,N_1947);
and U2164 (N_2164,N_1873,N_1667);
nand U2165 (N_2165,N_1742,N_1762);
and U2166 (N_2166,N_1823,N_1810);
or U2167 (N_2167,N_1635,N_1525);
and U2168 (N_2168,N_1857,N_1660);
nand U2169 (N_2169,N_1688,N_1881);
or U2170 (N_2170,N_1835,N_1730);
or U2171 (N_2171,N_1519,N_1869);
and U2172 (N_2172,N_1757,N_1817);
nor U2173 (N_2173,N_1970,N_1636);
or U2174 (N_2174,N_1641,N_1843);
nor U2175 (N_2175,N_1926,N_1719);
nand U2176 (N_2176,N_1901,N_1561);
or U2177 (N_2177,N_1540,N_1959);
nor U2178 (N_2178,N_1780,N_1564);
nor U2179 (N_2179,N_1978,N_1764);
nand U2180 (N_2180,N_1902,N_1990);
nand U2181 (N_2181,N_1569,N_1792);
or U2182 (N_2182,N_1616,N_1852);
nor U2183 (N_2183,N_1985,N_1551);
or U2184 (N_2184,N_1626,N_1880);
xnor U2185 (N_2185,N_1811,N_1637);
nand U2186 (N_2186,N_1980,N_1772);
nor U2187 (N_2187,N_1950,N_1649);
and U2188 (N_2188,N_1756,N_1603);
nor U2189 (N_2189,N_1718,N_1790);
nand U2190 (N_2190,N_1839,N_1789);
nor U2191 (N_2191,N_1514,N_1738);
nor U2192 (N_2192,N_1850,N_1849);
nand U2193 (N_2193,N_1631,N_1503);
nand U2194 (N_2194,N_1581,N_1584);
nand U2195 (N_2195,N_1910,N_1813);
or U2196 (N_2196,N_1889,N_1537);
and U2197 (N_2197,N_1524,N_1645);
nor U2198 (N_2198,N_1974,N_1766);
or U2199 (N_2199,N_1915,N_1786);
nand U2200 (N_2200,N_1953,N_1979);
nand U2201 (N_2201,N_1799,N_1721);
nand U2202 (N_2202,N_1554,N_1621);
nand U2203 (N_2203,N_1988,N_1765);
nand U2204 (N_2204,N_1866,N_1845);
nor U2205 (N_2205,N_1877,N_1848);
nand U2206 (N_2206,N_1522,N_1580);
xor U2207 (N_2207,N_1547,N_1851);
nor U2208 (N_2208,N_1853,N_1516);
or U2209 (N_2209,N_1897,N_1968);
and U2210 (N_2210,N_1690,N_1504);
nor U2211 (N_2211,N_1966,N_1906);
and U2212 (N_2212,N_1512,N_1595);
and U2213 (N_2213,N_1500,N_1837);
nand U2214 (N_2214,N_1892,N_1975);
nor U2215 (N_2215,N_1751,N_1760);
nor U2216 (N_2216,N_1610,N_1625);
nor U2217 (N_2217,N_1594,N_1859);
nor U2218 (N_2218,N_1679,N_1868);
and U2219 (N_2219,N_1560,N_1863);
or U2220 (N_2220,N_1717,N_1829);
or U2221 (N_2221,N_1629,N_1552);
and U2222 (N_2222,N_1883,N_1768);
nand U2223 (N_2223,N_1932,N_1725);
nand U2224 (N_2224,N_1761,N_1566);
xnor U2225 (N_2225,N_1989,N_1555);
and U2226 (N_2226,N_1531,N_1687);
and U2227 (N_2227,N_1784,N_1933);
nand U2228 (N_2228,N_1862,N_1775);
nor U2229 (N_2229,N_1709,N_1882);
and U2230 (N_2230,N_1752,N_1965);
and U2231 (N_2231,N_1526,N_1917);
or U2232 (N_2232,N_1976,N_1945);
and U2233 (N_2233,N_1698,N_1935);
or U2234 (N_2234,N_1606,N_1654);
and U2235 (N_2235,N_1510,N_1800);
nor U2236 (N_2236,N_1509,N_1895);
nand U2237 (N_2237,N_1871,N_1614);
or U2238 (N_2238,N_1699,N_1604);
nand U2239 (N_2239,N_1739,N_1696);
nor U2240 (N_2240,N_1916,N_1971);
nor U2241 (N_2241,N_1598,N_1726);
or U2242 (N_2242,N_1904,N_1893);
nand U2243 (N_2243,N_1993,N_1633);
nor U2244 (N_2244,N_1632,N_1888);
and U2245 (N_2245,N_1802,N_1534);
and U2246 (N_2246,N_1597,N_1870);
or U2247 (N_2247,N_1672,N_1720);
or U2248 (N_2248,N_1940,N_1948);
nor U2249 (N_2249,N_1648,N_1674);
nand U2250 (N_2250,N_1990,N_1849);
nor U2251 (N_2251,N_1730,N_1568);
nand U2252 (N_2252,N_1857,N_1887);
or U2253 (N_2253,N_1568,N_1748);
and U2254 (N_2254,N_1640,N_1589);
or U2255 (N_2255,N_1709,N_1921);
and U2256 (N_2256,N_1597,N_1517);
or U2257 (N_2257,N_1972,N_1652);
or U2258 (N_2258,N_1927,N_1755);
and U2259 (N_2259,N_1705,N_1765);
nand U2260 (N_2260,N_1964,N_1919);
and U2261 (N_2261,N_1766,N_1938);
or U2262 (N_2262,N_1660,N_1828);
nand U2263 (N_2263,N_1590,N_1672);
and U2264 (N_2264,N_1728,N_1550);
nand U2265 (N_2265,N_1729,N_1603);
xor U2266 (N_2266,N_1726,N_1959);
nand U2267 (N_2267,N_1742,N_1859);
nand U2268 (N_2268,N_1764,N_1807);
nor U2269 (N_2269,N_1833,N_1890);
or U2270 (N_2270,N_1684,N_1716);
nand U2271 (N_2271,N_1749,N_1710);
or U2272 (N_2272,N_1629,N_1541);
nor U2273 (N_2273,N_1845,N_1607);
and U2274 (N_2274,N_1872,N_1920);
nor U2275 (N_2275,N_1818,N_1546);
nor U2276 (N_2276,N_1923,N_1764);
nand U2277 (N_2277,N_1882,N_1861);
or U2278 (N_2278,N_1773,N_1904);
nand U2279 (N_2279,N_1975,N_1567);
nor U2280 (N_2280,N_1723,N_1519);
nand U2281 (N_2281,N_1845,N_1934);
nand U2282 (N_2282,N_1797,N_1544);
nor U2283 (N_2283,N_1578,N_1928);
nand U2284 (N_2284,N_1989,N_1774);
and U2285 (N_2285,N_1658,N_1907);
nand U2286 (N_2286,N_1766,N_1794);
and U2287 (N_2287,N_1889,N_1682);
nand U2288 (N_2288,N_1822,N_1602);
and U2289 (N_2289,N_1793,N_1859);
or U2290 (N_2290,N_1642,N_1645);
nor U2291 (N_2291,N_1963,N_1573);
nor U2292 (N_2292,N_1898,N_1790);
and U2293 (N_2293,N_1931,N_1864);
and U2294 (N_2294,N_1894,N_1597);
or U2295 (N_2295,N_1990,N_1723);
or U2296 (N_2296,N_1588,N_1866);
and U2297 (N_2297,N_1557,N_1634);
nor U2298 (N_2298,N_1971,N_1951);
or U2299 (N_2299,N_1532,N_1938);
and U2300 (N_2300,N_1786,N_1957);
or U2301 (N_2301,N_1659,N_1672);
nor U2302 (N_2302,N_1927,N_1825);
or U2303 (N_2303,N_1843,N_1542);
nor U2304 (N_2304,N_1927,N_1661);
and U2305 (N_2305,N_1662,N_1834);
nor U2306 (N_2306,N_1895,N_1964);
nor U2307 (N_2307,N_1784,N_1725);
nand U2308 (N_2308,N_1818,N_1698);
nor U2309 (N_2309,N_1840,N_1943);
nor U2310 (N_2310,N_1870,N_1684);
and U2311 (N_2311,N_1673,N_1960);
and U2312 (N_2312,N_1865,N_1777);
nand U2313 (N_2313,N_1792,N_1750);
xnor U2314 (N_2314,N_1973,N_1590);
and U2315 (N_2315,N_1895,N_1976);
nor U2316 (N_2316,N_1847,N_1548);
or U2317 (N_2317,N_1865,N_1939);
and U2318 (N_2318,N_1767,N_1902);
and U2319 (N_2319,N_1609,N_1913);
nor U2320 (N_2320,N_1587,N_1607);
or U2321 (N_2321,N_1894,N_1933);
nand U2322 (N_2322,N_1613,N_1786);
or U2323 (N_2323,N_1689,N_1824);
nor U2324 (N_2324,N_1869,N_1690);
nand U2325 (N_2325,N_1807,N_1737);
or U2326 (N_2326,N_1887,N_1968);
or U2327 (N_2327,N_1726,N_1929);
nand U2328 (N_2328,N_1892,N_1857);
and U2329 (N_2329,N_1535,N_1767);
nand U2330 (N_2330,N_1888,N_1977);
nand U2331 (N_2331,N_1518,N_1513);
or U2332 (N_2332,N_1777,N_1535);
or U2333 (N_2333,N_1694,N_1974);
nor U2334 (N_2334,N_1548,N_1900);
xnor U2335 (N_2335,N_1732,N_1887);
and U2336 (N_2336,N_1757,N_1530);
nand U2337 (N_2337,N_1604,N_1989);
or U2338 (N_2338,N_1858,N_1935);
nor U2339 (N_2339,N_1846,N_1516);
or U2340 (N_2340,N_1651,N_1857);
and U2341 (N_2341,N_1737,N_1892);
nor U2342 (N_2342,N_1695,N_1674);
nand U2343 (N_2343,N_1565,N_1518);
nand U2344 (N_2344,N_1882,N_1860);
or U2345 (N_2345,N_1830,N_1618);
or U2346 (N_2346,N_1659,N_1596);
nor U2347 (N_2347,N_1786,N_1505);
nor U2348 (N_2348,N_1548,N_1746);
nor U2349 (N_2349,N_1913,N_1720);
nor U2350 (N_2350,N_1909,N_1765);
nor U2351 (N_2351,N_1909,N_1859);
or U2352 (N_2352,N_1599,N_1507);
and U2353 (N_2353,N_1798,N_1945);
nor U2354 (N_2354,N_1632,N_1679);
nor U2355 (N_2355,N_1876,N_1823);
or U2356 (N_2356,N_1904,N_1831);
or U2357 (N_2357,N_1523,N_1729);
and U2358 (N_2358,N_1928,N_1613);
or U2359 (N_2359,N_1858,N_1925);
or U2360 (N_2360,N_1525,N_1831);
nand U2361 (N_2361,N_1806,N_1799);
and U2362 (N_2362,N_1794,N_1597);
nand U2363 (N_2363,N_1629,N_1971);
and U2364 (N_2364,N_1517,N_1931);
nor U2365 (N_2365,N_1826,N_1976);
and U2366 (N_2366,N_1636,N_1674);
xor U2367 (N_2367,N_1516,N_1675);
or U2368 (N_2368,N_1884,N_1887);
nand U2369 (N_2369,N_1614,N_1876);
or U2370 (N_2370,N_1770,N_1984);
and U2371 (N_2371,N_1949,N_1951);
and U2372 (N_2372,N_1964,N_1524);
or U2373 (N_2373,N_1636,N_1884);
nand U2374 (N_2374,N_1571,N_1774);
or U2375 (N_2375,N_1649,N_1825);
and U2376 (N_2376,N_1746,N_1852);
nor U2377 (N_2377,N_1957,N_1913);
nor U2378 (N_2378,N_1888,N_1604);
nand U2379 (N_2379,N_1811,N_1858);
nor U2380 (N_2380,N_1634,N_1647);
nor U2381 (N_2381,N_1859,N_1740);
nor U2382 (N_2382,N_1842,N_1593);
and U2383 (N_2383,N_1629,N_1661);
nand U2384 (N_2384,N_1655,N_1532);
nor U2385 (N_2385,N_1889,N_1749);
nand U2386 (N_2386,N_1626,N_1988);
or U2387 (N_2387,N_1807,N_1543);
nor U2388 (N_2388,N_1781,N_1933);
nand U2389 (N_2389,N_1982,N_1712);
nand U2390 (N_2390,N_1971,N_1559);
or U2391 (N_2391,N_1773,N_1915);
xor U2392 (N_2392,N_1529,N_1532);
nand U2393 (N_2393,N_1633,N_1991);
nor U2394 (N_2394,N_1815,N_1787);
and U2395 (N_2395,N_1900,N_1540);
or U2396 (N_2396,N_1641,N_1967);
nor U2397 (N_2397,N_1593,N_1952);
or U2398 (N_2398,N_1862,N_1507);
nand U2399 (N_2399,N_1618,N_1648);
or U2400 (N_2400,N_1529,N_1843);
nand U2401 (N_2401,N_1690,N_1668);
nand U2402 (N_2402,N_1603,N_1718);
nand U2403 (N_2403,N_1704,N_1923);
and U2404 (N_2404,N_1662,N_1554);
nor U2405 (N_2405,N_1999,N_1681);
nand U2406 (N_2406,N_1718,N_1687);
or U2407 (N_2407,N_1842,N_1913);
nor U2408 (N_2408,N_1949,N_1899);
or U2409 (N_2409,N_1888,N_1836);
nand U2410 (N_2410,N_1873,N_1724);
and U2411 (N_2411,N_1606,N_1710);
and U2412 (N_2412,N_1538,N_1624);
nor U2413 (N_2413,N_1910,N_1799);
nand U2414 (N_2414,N_1575,N_1959);
nand U2415 (N_2415,N_1949,N_1890);
nor U2416 (N_2416,N_1808,N_1683);
or U2417 (N_2417,N_1615,N_1585);
nand U2418 (N_2418,N_1725,N_1944);
nor U2419 (N_2419,N_1903,N_1875);
nor U2420 (N_2420,N_1604,N_1988);
nand U2421 (N_2421,N_1891,N_1756);
and U2422 (N_2422,N_1782,N_1945);
nor U2423 (N_2423,N_1924,N_1544);
nor U2424 (N_2424,N_1553,N_1628);
and U2425 (N_2425,N_1904,N_1709);
and U2426 (N_2426,N_1639,N_1886);
nor U2427 (N_2427,N_1753,N_1912);
nor U2428 (N_2428,N_1845,N_1995);
or U2429 (N_2429,N_1762,N_1703);
or U2430 (N_2430,N_1640,N_1520);
and U2431 (N_2431,N_1816,N_1641);
or U2432 (N_2432,N_1957,N_1549);
nor U2433 (N_2433,N_1907,N_1836);
and U2434 (N_2434,N_1526,N_1817);
and U2435 (N_2435,N_1726,N_1544);
or U2436 (N_2436,N_1909,N_1686);
and U2437 (N_2437,N_1514,N_1650);
nor U2438 (N_2438,N_1808,N_1883);
nand U2439 (N_2439,N_1947,N_1539);
nand U2440 (N_2440,N_1789,N_1801);
and U2441 (N_2441,N_1847,N_1671);
or U2442 (N_2442,N_1816,N_1531);
or U2443 (N_2443,N_1882,N_1713);
nor U2444 (N_2444,N_1944,N_1539);
nor U2445 (N_2445,N_1919,N_1511);
nand U2446 (N_2446,N_1985,N_1885);
nor U2447 (N_2447,N_1834,N_1734);
or U2448 (N_2448,N_1536,N_1715);
nor U2449 (N_2449,N_1554,N_1793);
and U2450 (N_2450,N_1566,N_1622);
or U2451 (N_2451,N_1851,N_1717);
nor U2452 (N_2452,N_1550,N_1760);
or U2453 (N_2453,N_1721,N_1718);
nand U2454 (N_2454,N_1919,N_1853);
or U2455 (N_2455,N_1990,N_1888);
and U2456 (N_2456,N_1914,N_1675);
or U2457 (N_2457,N_1841,N_1993);
or U2458 (N_2458,N_1806,N_1887);
nand U2459 (N_2459,N_1936,N_1527);
and U2460 (N_2460,N_1793,N_1540);
or U2461 (N_2461,N_1513,N_1585);
nor U2462 (N_2462,N_1804,N_1901);
nor U2463 (N_2463,N_1514,N_1896);
and U2464 (N_2464,N_1854,N_1782);
and U2465 (N_2465,N_1528,N_1717);
nand U2466 (N_2466,N_1582,N_1989);
and U2467 (N_2467,N_1595,N_1583);
nor U2468 (N_2468,N_1749,N_1607);
nand U2469 (N_2469,N_1974,N_1553);
nor U2470 (N_2470,N_1824,N_1899);
and U2471 (N_2471,N_1669,N_1701);
nor U2472 (N_2472,N_1858,N_1698);
and U2473 (N_2473,N_1625,N_1983);
nor U2474 (N_2474,N_1653,N_1587);
and U2475 (N_2475,N_1928,N_1914);
and U2476 (N_2476,N_1581,N_1563);
or U2477 (N_2477,N_1866,N_1873);
nor U2478 (N_2478,N_1676,N_1611);
or U2479 (N_2479,N_1955,N_1869);
nor U2480 (N_2480,N_1980,N_1655);
or U2481 (N_2481,N_1611,N_1553);
and U2482 (N_2482,N_1810,N_1758);
and U2483 (N_2483,N_1702,N_1889);
nand U2484 (N_2484,N_1643,N_1964);
nand U2485 (N_2485,N_1973,N_1645);
or U2486 (N_2486,N_1527,N_1982);
or U2487 (N_2487,N_1776,N_1763);
nor U2488 (N_2488,N_1810,N_1814);
and U2489 (N_2489,N_1957,N_1556);
or U2490 (N_2490,N_1558,N_1898);
nand U2491 (N_2491,N_1503,N_1882);
nor U2492 (N_2492,N_1618,N_1660);
xnor U2493 (N_2493,N_1660,N_1649);
nand U2494 (N_2494,N_1900,N_1918);
nand U2495 (N_2495,N_1862,N_1593);
nand U2496 (N_2496,N_1535,N_1970);
nand U2497 (N_2497,N_1783,N_1738);
nor U2498 (N_2498,N_1677,N_1689);
nand U2499 (N_2499,N_1887,N_1705);
xor U2500 (N_2500,N_2307,N_2087);
nand U2501 (N_2501,N_2104,N_2358);
nand U2502 (N_2502,N_2482,N_2077);
or U2503 (N_2503,N_2026,N_2428);
or U2504 (N_2504,N_2303,N_2300);
nand U2505 (N_2505,N_2062,N_2332);
or U2506 (N_2506,N_2465,N_2091);
or U2507 (N_2507,N_2041,N_2403);
nor U2508 (N_2508,N_2444,N_2141);
nand U2509 (N_2509,N_2000,N_2159);
and U2510 (N_2510,N_2448,N_2455);
nor U2511 (N_2511,N_2085,N_2341);
and U2512 (N_2512,N_2096,N_2458);
or U2513 (N_2513,N_2052,N_2027);
or U2514 (N_2514,N_2023,N_2427);
nor U2515 (N_2515,N_2165,N_2312);
nand U2516 (N_2516,N_2117,N_2076);
and U2517 (N_2517,N_2202,N_2366);
nand U2518 (N_2518,N_2390,N_2126);
nor U2519 (N_2519,N_2469,N_2481);
nand U2520 (N_2520,N_2274,N_2393);
or U2521 (N_2521,N_2318,N_2177);
or U2522 (N_2522,N_2146,N_2464);
or U2523 (N_2523,N_2389,N_2051);
nor U2524 (N_2524,N_2351,N_2305);
nand U2525 (N_2525,N_2098,N_2473);
and U2526 (N_2526,N_2012,N_2203);
and U2527 (N_2527,N_2240,N_2361);
or U2528 (N_2528,N_2429,N_2399);
or U2529 (N_2529,N_2217,N_2125);
and U2530 (N_2530,N_2179,N_2226);
xor U2531 (N_2531,N_2038,N_2004);
nand U2532 (N_2532,N_2426,N_2392);
nor U2533 (N_2533,N_2143,N_2235);
or U2534 (N_2534,N_2486,N_2129);
nor U2535 (N_2535,N_2266,N_2135);
or U2536 (N_2536,N_2057,N_2059);
nand U2537 (N_2537,N_2467,N_2344);
or U2538 (N_2538,N_2421,N_2063);
nand U2539 (N_2539,N_2224,N_2210);
or U2540 (N_2540,N_2437,N_2433);
nor U2541 (N_2541,N_2296,N_2102);
or U2542 (N_2542,N_2391,N_2045);
or U2543 (N_2543,N_2471,N_2174);
nand U2544 (N_2544,N_2151,N_2325);
nand U2545 (N_2545,N_2178,N_2418);
nor U2546 (N_2546,N_2396,N_2374);
or U2547 (N_2547,N_2160,N_2335);
nor U2548 (N_2548,N_2204,N_2384);
or U2549 (N_2549,N_2233,N_2331);
or U2550 (N_2550,N_2001,N_2346);
and U2551 (N_2551,N_2333,N_2212);
nor U2552 (N_2552,N_2130,N_2200);
and U2553 (N_2553,N_2169,N_2337);
nor U2554 (N_2554,N_2031,N_2083);
or U2555 (N_2555,N_2173,N_2144);
nor U2556 (N_2556,N_2449,N_2121);
and U2557 (N_2557,N_2123,N_2435);
and U2558 (N_2558,N_2443,N_2081);
nand U2559 (N_2559,N_2316,N_2199);
and U2560 (N_2560,N_2171,N_2220);
and U2561 (N_2561,N_2338,N_2231);
nor U2562 (N_2562,N_2339,N_2239);
or U2563 (N_2563,N_2357,N_2035);
and U2564 (N_2564,N_2013,N_2478);
nor U2565 (N_2565,N_2017,N_2301);
or U2566 (N_2566,N_2291,N_2075);
nand U2567 (N_2567,N_2089,N_2243);
nand U2568 (N_2568,N_2065,N_2475);
or U2569 (N_2569,N_2401,N_2133);
nand U2570 (N_2570,N_2379,N_2491);
nand U2571 (N_2571,N_2015,N_2069);
nor U2572 (N_2572,N_2356,N_2070);
nand U2573 (N_2573,N_2304,N_2453);
and U2574 (N_2574,N_2198,N_2343);
and U2575 (N_2575,N_2167,N_2056);
nand U2576 (N_2576,N_2417,N_2058);
nor U2577 (N_2577,N_2140,N_2191);
nand U2578 (N_2578,N_2474,N_2242);
nand U2579 (N_2579,N_2286,N_2328);
nand U2580 (N_2580,N_2007,N_2170);
nor U2581 (N_2581,N_2209,N_2279);
nand U2582 (N_2582,N_2251,N_2322);
nor U2583 (N_2583,N_2280,N_2313);
or U2584 (N_2584,N_2219,N_2410);
and U2585 (N_2585,N_2487,N_2252);
or U2586 (N_2586,N_2223,N_2005);
nor U2587 (N_2587,N_2131,N_2354);
nand U2588 (N_2588,N_2376,N_2009);
nor U2589 (N_2589,N_2176,N_2244);
and U2590 (N_2590,N_2257,N_2263);
nor U2591 (N_2591,N_2368,N_2398);
and U2592 (N_2592,N_2363,N_2054);
nor U2593 (N_2593,N_2461,N_2442);
or U2594 (N_2594,N_2480,N_2111);
nor U2595 (N_2595,N_2053,N_2228);
and U2596 (N_2596,N_2422,N_2414);
nand U2597 (N_2597,N_2477,N_2195);
or U2598 (N_2598,N_2405,N_2237);
nand U2599 (N_2599,N_2044,N_2373);
nor U2600 (N_2600,N_2447,N_2364);
or U2601 (N_2601,N_2306,N_2310);
nand U2602 (N_2602,N_2492,N_2214);
nor U2603 (N_2603,N_2119,N_2241);
or U2604 (N_2604,N_2105,N_2382);
nand U2605 (N_2605,N_2095,N_2362);
nor U2606 (N_2606,N_2489,N_2483);
or U2607 (N_2607,N_2342,N_2425);
nand U2608 (N_2608,N_2295,N_2147);
nand U2609 (N_2609,N_2084,N_2072);
nor U2610 (N_2610,N_2194,N_2192);
and U2611 (N_2611,N_2439,N_2079);
nor U2612 (N_2612,N_2297,N_2229);
and U2613 (N_2613,N_2024,N_2032);
nand U2614 (N_2614,N_2276,N_2459);
or U2615 (N_2615,N_2375,N_2320);
and U2616 (N_2616,N_2254,N_2016);
nand U2617 (N_2617,N_2055,N_2432);
xnor U2618 (N_2618,N_2456,N_2334);
nand U2619 (N_2619,N_2352,N_2190);
and U2620 (N_2620,N_2142,N_2247);
or U2621 (N_2621,N_2350,N_2201);
or U2622 (N_2622,N_2232,N_2476);
nand U2623 (N_2623,N_2269,N_2025);
nand U2624 (N_2624,N_2353,N_2164);
nand U2625 (N_2625,N_2182,N_2050);
and U2626 (N_2626,N_2408,N_2074);
nor U2627 (N_2627,N_2323,N_2029);
nand U2628 (N_2628,N_2175,N_2434);
nor U2629 (N_2629,N_2014,N_2088);
and U2630 (N_2630,N_2037,N_2314);
and U2631 (N_2631,N_2446,N_2246);
or U2632 (N_2632,N_2383,N_2161);
nand U2633 (N_2633,N_2168,N_2463);
or U2634 (N_2634,N_2153,N_2139);
and U2635 (N_2635,N_2213,N_2118);
nand U2636 (N_2636,N_2138,N_2260);
nor U2637 (N_2637,N_2419,N_2107);
nor U2638 (N_2638,N_2060,N_2033);
nor U2639 (N_2639,N_2340,N_2120);
and U2640 (N_2640,N_2407,N_2452);
nand U2641 (N_2641,N_2078,N_2454);
or U2642 (N_2642,N_2093,N_2385);
nand U2643 (N_2643,N_2386,N_2462);
nand U2644 (N_2644,N_2329,N_2330);
or U2645 (N_2645,N_2071,N_2430);
and U2646 (N_2646,N_2411,N_2345);
or U2647 (N_2647,N_2367,N_2282);
nor U2648 (N_2648,N_2122,N_2420);
nor U2649 (N_2649,N_2472,N_2494);
or U2650 (N_2650,N_2365,N_2048);
and U2651 (N_2651,N_2281,N_2196);
nor U2652 (N_2652,N_2094,N_2441);
nor U2653 (N_2653,N_2221,N_2166);
or U2654 (N_2654,N_2402,N_2010);
nand U2655 (N_2655,N_2436,N_2388);
nor U2656 (N_2656,N_2324,N_2137);
nor U2657 (N_2657,N_2236,N_2019);
nand U2658 (N_2658,N_2103,N_2003);
or U2659 (N_2659,N_2268,N_2127);
nand U2660 (N_2660,N_2272,N_2479);
or U2661 (N_2661,N_2068,N_2275);
nor U2662 (N_2662,N_2150,N_2114);
nor U2663 (N_2663,N_2283,N_2315);
and U2664 (N_2664,N_2238,N_2308);
and U2665 (N_2665,N_2440,N_2381);
nor U2666 (N_2666,N_2355,N_2451);
and U2667 (N_2667,N_2468,N_2180);
and U2668 (N_2668,N_2490,N_2277);
or U2669 (N_2669,N_2466,N_2293);
or U2670 (N_2670,N_2008,N_2415);
and U2671 (N_2671,N_2326,N_2205);
nor U2672 (N_2672,N_2061,N_2273);
or U2673 (N_2673,N_2485,N_2043);
and U2674 (N_2674,N_2409,N_2234);
nand U2675 (N_2675,N_2284,N_2359);
nand U2676 (N_2676,N_2360,N_2267);
and U2677 (N_2677,N_2047,N_2499);
and U2678 (N_2678,N_2309,N_2327);
and U2679 (N_2679,N_2185,N_2377);
or U2680 (N_2680,N_2259,N_2207);
or U2681 (N_2681,N_2319,N_2248);
and U2682 (N_2682,N_2034,N_2186);
xnor U2683 (N_2683,N_2271,N_2066);
and U2684 (N_2684,N_2086,N_2249);
xnor U2685 (N_2685,N_2290,N_2183);
or U2686 (N_2686,N_2299,N_2090);
or U2687 (N_2687,N_2262,N_2394);
nand U2688 (N_2688,N_2181,N_2371);
nor U2689 (N_2689,N_2387,N_2395);
and U2690 (N_2690,N_2039,N_2256);
nor U2691 (N_2691,N_2128,N_2423);
or U2692 (N_2692,N_2450,N_2124);
or U2693 (N_2693,N_2497,N_2348);
or U2694 (N_2694,N_2498,N_2424);
nand U2695 (N_2695,N_2049,N_2187);
nand U2696 (N_2696,N_2416,N_2216);
nor U2697 (N_2697,N_2347,N_2011);
or U2698 (N_2698,N_2294,N_2099);
or U2699 (N_2699,N_2154,N_2002);
nor U2700 (N_2700,N_2265,N_2149);
and U2701 (N_2701,N_2136,N_2496);
nand U2702 (N_2702,N_2080,N_2292);
or U2703 (N_2703,N_2067,N_2397);
nor U2704 (N_2704,N_2042,N_2188);
or U2705 (N_2705,N_2378,N_2431);
or U2706 (N_2706,N_2155,N_2132);
or U2707 (N_2707,N_2287,N_2109);
nor U2708 (N_2708,N_2278,N_2206);
and U2709 (N_2709,N_2211,N_2158);
nand U2710 (N_2710,N_2101,N_2064);
and U2711 (N_2711,N_2172,N_2152);
or U2712 (N_2712,N_2311,N_2116);
or U2713 (N_2713,N_2112,N_2488);
nor U2714 (N_2714,N_2189,N_2400);
nand U2715 (N_2715,N_2412,N_2245);
or U2716 (N_2716,N_2222,N_2258);
or U2717 (N_2717,N_2100,N_2145);
or U2718 (N_2718,N_2227,N_2162);
or U2719 (N_2719,N_2022,N_2030);
nand U2720 (N_2720,N_2380,N_2270);
and U2721 (N_2721,N_2208,N_2108);
nor U2722 (N_2722,N_2288,N_2113);
and U2723 (N_2723,N_2264,N_2021);
nand U2724 (N_2724,N_2372,N_2006);
nand U2725 (N_2725,N_2253,N_2134);
and U2726 (N_2726,N_2404,N_2302);
nor U2727 (N_2727,N_2321,N_2193);
and U2728 (N_2728,N_2336,N_2406);
or U2729 (N_2729,N_2218,N_2495);
or U2730 (N_2730,N_2230,N_2097);
or U2731 (N_2731,N_2285,N_2349);
nand U2732 (N_2732,N_2215,N_2225);
or U2733 (N_2733,N_2110,N_2493);
and U2734 (N_2734,N_2298,N_2250);
nor U2735 (N_2735,N_2460,N_2184);
nand U2736 (N_2736,N_2369,N_2317);
nand U2737 (N_2737,N_2157,N_2040);
or U2738 (N_2738,N_2457,N_2020);
nor U2739 (N_2739,N_2470,N_2438);
nor U2740 (N_2740,N_2445,N_2092);
nand U2741 (N_2741,N_2261,N_2255);
nor U2742 (N_2742,N_2036,N_2073);
and U2743 (N_2743,N_2018,N_2028);
or U2744 (N_2744,N_2156,N_2106);
or U2745 (N_2745,N_2413,N_2289);
nand U2746 (N_2746,N_2197,N_2370);
nand U2747 (N_2747,N_2082,N_2163);
and U2748 (N_2748,N_2148,N_2046);
nor U2749 (N_2749,N_2484,N_2115);
and U2750 (N_2750,N_2387,N_2299);
nand U2751 (N_2751,N_2091,N_2118);
and U2752 (N_2752,N_2464,N_2031);
nor U2753 (N_2753,N_2245,N_2140);
and U2754 (N_2754,N_2400,N_2204);
nor U2755 (N_2755,N_2434,N_2437);
nand U2756 (N_2756,N_2069,N_2386);
and U2757 (N_2757,N_2126,N_2389);
nand U2758 (N_2758,N_2414,N_2474);
nor U2759 (N_2759,N_2233,N_2323);
nor U2760 (N_2760,N_2247,N_2079);
nand U2761 (N_2761,N_2277,N_2295);
nor U2762 (N_2762,N_2366,N_2133);
nor U2763 (N_2763,N_2288,N_2286);
or U2764 (N_2764,N_2286,N_2040);
or U2765 (N_2765,N_2103,N_2356);
nand U2766 (N_2766,N_2050,N_2434);
nand U2767 (N_2767,N_2390,N_2414);
nand U2768 (N_2768,N_2113,N_2152);
or U2769 (N_2769,N_2088,N_2324);
nor U2770 (N_2770,N_2040,N_2433);
and U2771 (N_2771,N_2299,N_2452);
and U2772 (N_2772,N_2224,N_2229);
nor U2773 (N_2773,N_2405,N_2114);
and U2774 (N_2774,N_2367,N_2011);
nand U2775 (N_2775,N_2340,N_2205);
or U2776 (N_2776,N_2256,N_2276);
and U2777 (N_2777,N_2196,N_2399);
and U2778 (N_2778,N_2185,N_2219);
and U2779 (N_2779,N_2114,N_2093);
nor U2780 (N_2780,N_2189,N_2204);
and U2781 (N_2781,N_2020,N_2270);
or U2782 (N_2782,N_2193,N_2096);
or U2783 (N_2783,N_2114,N_2141);
and U2784 (N_2784,N_2173,N_2068);
nor U2785 (N_2785,N_2208,N_2409);
nand U2786 (N_2786,N_2255,N_2300);
nand U2787 (N_2787,N_2023,N_2441);
and U2788 (N_2788,N_2054,N_2090);
or U2789 (N_2789,N_2403,N_2133);
nor U2790 (N_2790,N_2341,N_2417);
nor U2791 (N_2791,N_2121,N_2288);
or U2792 (N_2792,N_2415,N_2472);
nand U2793 (N_2793,N_2093,N_2030);
nand U2794 (N_2794,N_2028,N_2460);
or U2795 (N_2795,N_2350,N_2295);
or U2796 (N_2796,N_2118,N_2161);
and U2797 (N_2797,N_2162,N_2353);
or U2798 (N_2798,N_2116,N_2191);
and U2799 (N_2799,N_2242,N_2327);
nor U2800 (N_2800,N_2211,N_2180);
nand U2801 (N_2801,N_2080,N_2015);
and U2802 (N_2802,N_2402,N_2416);
nand U2803 (N_2803,N_2025,N_2222);
and U2804 (N_2804,N_2067,N_2068);
nand U2805 (N_2805,N_2296,N_2433);
or U2806 (N_2806,N_2436,N_2047);
nand U2807 (N_2807,N_2292,N_2191);
nand U2808 (N_2808,N_2480,N_2254);
nand U2809 (N_2809,N_2181,N_2441);
nand U2810 (N_2810,N_2319,N_2096);
and U2811 (N_2811,N_2149,N_2419);
and U2812 (N_2812,N_2019,N_2387);
nand U2813 (N_2813,N_2303,N_2221);
and U2814 (N_2814,N_2295,N_2488);
nand U2815 (N_2815,N_2364,N_2474);
nand U2816 (N_2816,N_2038,N_2378);
and U2817 (N_2817,N_2194,N_2472);
nor U2818 (N_2818,N_2294,N_2205);
nand U2819 (N_2819,N_2246,N_2036);
or U2820 (N_2820,N_2025,N_2015);
nor U2821 (N_2821,N_2248,N_2484);
and U2822 (N_2822,N_2219,N_2045);
and U2823 (N_2823,N_2391,N_2100);
nor U2824 (N_2824,N_2252,N_2138);
and U2825 (N_2825,N_2029,N_2257);
nand U2826 (N_2826,N_2232,N_2432);
nand U2827 (N_2827,N_2265,N_2317);
nor U2828 (N_2828,N_2176,N_2317);
or U2829 (N_2829,N_2120,N_2044);
nor U2830 (N_2830,N_2246,N_2354);
nand U2831 (N_2831,N_2062,N_2074);
and U2832 (N_2832,N_2242,N_2118);
and U2833 (N_2833,N_2359,N_2087);
nand U2834 (N_2834,N_2025,N_2045);
or U2835 (N_2835,N_2255,N_2100);
or U2836 (N_2836,N_2445,N_2447);
and U2837 (N_2837,N_2032,N_2490);
and U2838 (N_2838,N_2483,N_2111);
and U2839 (N_2839,N_2253,N_2039);
and U2840 (N_2840,N_2105,N_2044);
or U2841 (N_2841,N_2427,N_2220);
nor U2842 (N_2842,N_2373,N_2145);
nor U2843 (N_2843,N_2396,N_2465);
and U2844 (N_2844,N_2246,N_2039);
and U2845 (N_2845,N_2472,N_2449);
and U2846 (N_2846,N_2008,N_2165);
nor U2847 (N_2847,N_2200,N_2024);
nor U2848 (N_2848,N_2441,N_2438);
or U2849 (N_2849,N_2449,N_2447);
or U2850 (N_2850,N_2050,N_2260);
nor U2851 (N_2851,N_2239,N_2313);
or U2852 (N_2852,N_2087,N_2295);
nand U2853 (N_2853,N_2450,N_2484);
or U2854 (N_2854,N_2023,N_2087);
nand U2855 (N_2855,N_2204,N_2331);
nand U2856 (N_2856,N_2347,N_2396);
or U2857 (N_2857,N_2086,N_2380);
nor U2858 (N_2858,N_2364,N_2438);
or U2859 (N_2859,N_2433,N_2453);
nand U2860 (N_2860,N_2261,N_2351);
or U2861 (N_2861,N_2013,N_2367);
nor U2862 (N_2862,N_2247,N_2407);
nand U2863 (N_2863,N_2284,N_2140);
nand U2864 (N_2864,N_2422,N_2248);
nor U2865 (N_2865,N_2468,N_2021);
and U2866 (N_2866,N_2308,N_2164);
or U2867 (N_2867,N_2106,N_2354);
xnor U2868 (N_2868,N_2488,N_2003);
nand U2869 (N_2869,N_2121,N_2181);
nor U2870 (N_2870,N_2290,N_2240);
or U2871 (N_2871,N_2092,N_2325);
and U2872 (N_2872,N_2258,N_2074);
nand U2873 (N_2873,N_2363,N_2193);
nand U2874 (N_2874,N_2006,N_2134);
and U2875 (N_2875,N_2355,N_2461);
or U2876 (N_2876,N_2217,N_2211);
nand U2877 (N_2877,N_2283,N_2013);
or U2878 (N_2878,N_2241,N_2235);
and U2879 (N_2879,N_2406,N_2131);
or U2880 (N_2880,N_2314,N_2102);
and U2881 (N_2881,N_2485,N_2103);
and U2882 (N_2882,N_2005,N_2092);
and U2883 (N_2883,N_2385,N_2469);
and U2884 (N_2884,N_2318,N_2202);
nor U2885 (N_2885,N_2345,N_2118);
nand U2886 (N_2886,N_2475,N_2161);
nand U2887 (N_2887,N_2256,N_2483);
and U2888 (N_2888,N_2270,N_2179);
nor U2889 (N_2889,N_2322,N_2332);
or U2890 (N_2890,N_2241,N_2337);
and U2891 (N_2891,N_2290,N_2133);
and U2892 (N_2892,N_2156,N_2439);
or U2893 (N_2893,N_2394,N_2362);
nand U2894 (N_2894,N_2125,N_2341);
nor U2895 (N_2895,N_2235,N_2021);
nand U2896 (N_2896,N_2481,N_2186);
nand U2897 (N_2897,N_2006,N_2271);
nor U2898 (N_2898,N_2281,N_2105);
and U2899 (N_2899,N_2437,N_2290);
and U2900 (N_2900,N_2270,N_2379);
nor U2901 (N_2901,N_2345,N_2020);
or U2902 (N_2902,N_2197,N_2064);
nand U2903 (N_2903,N_2139,N_2454);
or U2904 (N_2904,N_2257,N_2402);
nand U2905 (N_2905,N_2267,N_2498);
or U2906 (N_2906,N_2050,N_2151);
or U2907 (N_2907,N_2482,N_2333);
and U2908 (N_2908,N_2140,N_2221);
or U2909 (N_2909,N_2006,N_2013);
nor U2910 (N_2910,N_2406,N_2308);
or U2911 (N_2911,N_2249,N_2454);
or U2912 (N_2912,N_2107,N_2171);
or U2913 (N_2913,N_2311,N_2332);
and U2914 (N_2914,N_2349,N_2025);
and U2915 (N_2915,N_2176,N_2036);
nand U2916 (N_2916,N_2423,N_2094);
nor U2917 (N_2917,N_2298,N_2071);
or U2918 (N_2918,N_2042,N_2268);
and U2919 (N_2919,N_2058,N_2046);
nand U2920 (N_2920,N_2235,N_2266);
nand U2921 (N_2921,N_2388,N_2044);
nor U2922 (N_2922,N_2441,N_2293);
nor U2923 (N_2923,N_2422,N_2498);
nor U2924 (N_2924,N_2334,N_2344);
nor U2925 (N_2925,N_2477,N_2094);
or U2926 (N_2926,N_2213,N_2388);
or U2927 (N_2927,N_2037,N_2270);
and U2928 (N_2928,N_2291,N_2413);
nand U2929 (N_2929,N_2190,N_2144);
nand U2930 (N_2930,N_2344,N_2333);
nor U2931 (N_2931,N_2341,N_2040);
or U2932 (N_2932,N_2001,N_2273);
and U2933 (N_2933,N_2486,N_2137);
and U2934 (N_2934,N_2457,N_2461);
and U2935 (N_2935,N_2378,N_2469);
or U2936 (N_2936,N_2282,N_2278);
nand U2937 (N_2937,N_2256,N_2326);
or U2938 (N_2938,N_2392,N_2019);
or U2939 (N_2939,N_2284,N_2223);
or U2940 (N_2940,N_2306,N_2313);
nor U2941 (N_2941,N_2224,N_2296);
or U2942 (N_2942,N_2405,N_2215);
or U2943 (N_2943,N_2081,N_2260);
nor U2944 (N_2944,N_2257,N_2119);
and U2945 (N_2945,N_2076,N_2380);
nand U2946 (N_2946,N_2363,N_2293);
or U2947 (N_2947,N_2020,N_2423);
nor U2948 (N_2948,N_2257,N_2294);
and U2949 (N_2949,N_2171,N_2104);
nor U2950 (N_2950,N_2128,N_2207);
nor U2951 (N_2951,N_2169,N_2188);
nand U2952 (N_2952,N_2237,N_2189);
nand U2953 (N_2953,N_2314,N_2271);
and U2954 (N_2954,N_2226,N_2370);
nand U2955 (N_2955,N_2143,N_2418);
nor U2956 (N_2956,N_2010,N_2467);
or U2957 (N_2957,N_2248,N_2136);
or U2958 (N_2958,N_2252,N_2384);
or U2959 (N_2959,N_2217,N_2261);
xnor U2960 (N_2960,N_2023,N_2089);
nor U2961 (N_2961,N_2187,N_2169);
or U2962 (N_2962,N_2299,N_2354);
nand U2963 (N_2963,N_2455,N_2226);
or U2964 (N_2964,N_2088,N_2414);
and U2965 (N_2965,N_2444,N_2176);
and U2966 (N_2966,N_2421,N_2353);
nor U2967 (N_2967,N_2006,N_2022);
and U2968 (N_2968,N_2043,N_2468);
or U2969 (N_2969,N_2020,N_2247);
nand U2970 (N_2970,N_2420,N_2170);
or U2971 (N_2971,N_2201,N_2152);
nor U2972 (N_2972,N_2494,N_2213);
nor U2973 (N_2973,N_2258,N_2221);
nor U2974 (N_2974,N_2177,N_2358);
nand U2975 (N_2975,N_2364,N_2414);
and U2976 (N_2976,N_2237,N_2059);
nor U2977 (N_2977,N_2443,N_2157);
or U2978 (N_2978,N_2281,N_2494);
and U2979 (N_2979,N_2158,N_2180);
nand U2980 (N_2980,N_2372,N_2021);
nand U2981 (N_2981,N_2273,N_2106);
and U2982 (N_2982,N_2458,N_2477);
nor U2983 (N_2983,N_2249,N_2316);
nand U2984 (N_2984,N_2133,N_2470);
or U2985 (N_2985,N_2356,N_2280);
and U2986 (N_2986,N_2015,N_2256);
and U2987 (N_2987,N_2372,N_2183);
nand U2988 (N_2988,N_2443,N_2323);
nand U2989 (N_2989,N_2484,N_2295);
and U2990 (N_2990,N_2147,N_2106);
or U2991 (N_2991,N_2005,N_2093);
and U2992 (N_2992,N_2129,N_2485);
nor U2993 (N_2993,N_2112,N_2009);
or U2994 (N_2994,N_2341,N_2187);
nand U2995 (N_2995,N_2295,N_2127);
and U2996 (N_2996,N_2243,N_2233);
and U2997 (N_2997,N_2329,N_2246);
nor U2998 (N_2998,N_2476,N_2373);
and U2999 (N_2999,N_2379,N_2448);
nand U3000 (N_3000,N_2924,N_2729);
and U3001 (N_3001,N_2708,N_2769);
or U3002 (N_3002,N_2737,N_2801);
or U3003 (N_3003,N_2880,N_2674);
nand U3004 (N_3004,N_2915,N_2698);
nor U3005 (N_3005,N_2551,N_2962);
nand U3006 (N_3006,N_2723,N_2839);
and U3007 (N_3007,N_2894,N_2787);
and U3008 (N_3008,N_2572,N_2517);
nand U3009 (N_3009,N_2697,N_2992);
and U3010 (N_3010,N_2568,N_2726);
or U3011 (N_3011,N_2789,N_2592);
nand U3012 (N_3012,N_2805,N_2690);
nand U3013 (N_3013,N_2803,N_2521);
and U3014 (N_3014,N_2820,N_2945);
or U3015 (N_3015,N_2860,N_2902);
and U3016 (N_3016,N_2524,N_2815);
and U3017 (N_3017,N_2806,N_2986);
nor U3018 (N_3018,N_2600,N_2631);
and U3019 (N_3019,N_2622,N_2968);
nor U3020 (N_3020,N_2955,N_2620);
and U3021 (N_3021,N_2910,N_2540);
and U3022 (N_3022,N_2556,N_2740);
or U3023 (N_3023,N_2797,N_2535);
nand U3024 (N_3024,N_2874,N_2851);
or U3025 (N_3025,N_2500,N_2656);
xor U3026 (N_3026,N_2676,N_2758);
or U3027 (N_3027,N_2724,N_2651);
or U3028 (N_3028,N_2950,N_2525);
nor U3029 (N_3029,N_2505,N_2713);
and U3030 (N_3030,N_2691,N_2987);
or U3031 (N_3031,N_2781,N_2725);
or U3032 (N_3032,N_2734,N_2732);
and U3033 (N_3033,N_2934,N_2972);
nor U3034 (N_3034,N_2714,N_2558);
nor U3035 (N_3035,N_2601,N_2570);
nand U3036 (N_3036,N_2662,N_2991);
or U3037 (N_3037,N_2897,N_2811);
and U3038 (N_3038,N_2545,N_2763);
or U3039 (N_3039,N_2750,N_2864);
or U3040 (N_3040,N_2931,N_2967);
nor U3041 (N_3041,N_2964,N_2618);
nor U3042 (N_3042,N_2649,N_2786);
nand U3043 (N_3043,N_2606,N_2575);
nor U3044 (N_3044,N_2745,N_2650);
nor U3045 (N_3045,N_2644,N_2501);
nor U3046 (N_3046,N_2544,N_2585);
and U3047 (N_3047,N_2779,N_2988);
or U3048 (N_3048,N_2655,N_2928);
nand U3049 (N_3049,N_2668,N_2783);
or U3050 (N_3050,N_2835,N_2621);
nand U3051 (N_3051,N_2752,N_2716);
or U3052 (N_3052,N_2818,N_2913);
and U3053 (N_3053,N_2749,N_2583);
xor U3054 (N_3054,N_2859,N_2961);
or U3055 (N_3055,N_2626,N_2793);
and U3056 (N_3056,N_2678,N_2946);
nand U3057 (N_3057,N_2536,N_2529);
nand U3058 (N_3058,N_2994,N_2833);
and U3059 (N_3059,N_2664,N_2576);
and U3060 (N_3060,N_2559,N_2883);
nor U3061 (N_3061,N_2704,N_2981);
xor U3062 (N_3062,N_2679,N_2997);
nand U3063 (N_3063,N_2784,N_2754);
and U3064 (N_3064,N_2603,N_2628);
nand U3065 (N_3065,N_2958,N_2960);
nor U3066 (N_3066,N_2523,N_2617);
nand U3067 (N_3067,N_2586,N_2751);
nor U3068 (N_3068,N_2873,N_2895);
or U3069 (N_3069,N_2788,N_2755);
or U3070 (N_3070,N_2893,N_2736);
nor U3071 (N_3071,N_2947,N_2506);
and U3072 (N_3072,N_2966,N_2847);
and U3073 (N_3073,N_2798,N_2627);
nor U3074 (N_3074,N_2700,N_2927);
and U3075 (N_3075,N_2705,N_2827);
and U3076 (N_3076,N_2855,N_2911);
nand U3077 (N_3077,N_2999,N_2772);
and U3078 (N_3078,N_2765,N_2875);
and U3079 (N_3079,N_2825,N_2598);
and U3080 (N_3080,N_2808,N_2625);
and U3081 (N_3081,N_2905,N_2699);
nor U3082 (N_3082,N_2954,N_2744);
and U3083 (N_3083,N_2730,N_2645);
nor U3084 (N_3084,N_2854,N_2637);
or U3085 (N_3085,N_2858,N_2840);
nor U3086 (N_3086,N_2522,N_2553);
nand U3087 (N_3087,N_2990,N_2863);
or U3088 (N_3088,N_2661,N_2872);
nor U3089 (N_3089,N_2720,N_2503);
and U3090 (N_3090,N_2560,N_2879);
nor U3091 (N_3091,N_2760,N_2973);
and U3092 (N_3092,N_2543,N_2660);
and U3093 (N_3093,N_2565,N_2748);
and U3094 (N_3094,N_2799,N_2842);
nand U3095 (N_3095,N_2670,N_2581);
nor U3096 (N_3096,N_2534,N_2647);
nand U3097 (N_3097,N_2681,N_2687);
or U3098 (N_3098,N_2876,N_2666);
nor U3099 (N_3099,N_2942,N_2605);
nand U3100 (N_3100,N_2963,N_2831);
or U3101 (N_3101,N_2747,N_2926);
nand U3102 (N_3102,N_2539,N_2707);
and U3103 (N_3103,N_2982,N_2878);
or U3104 (N_3104,N_2739,N_2579);
nand U3105 (N_3105,N_2975,N_2933);
nor U3106 (N_3106,N_2980,N_2508);
nand U3107 (N_3107,N_2513,N_2908);
and U3108 (N_3108,N_2684,N_2995);
and U3109 (N_3109,N_2685,N_2871);
and U3110 (N_3110,N_2604,N_2590);
or U3111 (N_3111,N_2692,N_2596);
nor U3112 (N_3112,N_2642,N_2611);
and U3113 (N_3113,N_2721,N_2770);
and U3114 (N_3114,N_2941,N_2771);
nor U3115 (N_3115,N_2594,N_2951);
and U3116 (N_3116,N_2515,N_2904);
or U3117 (N_3117,N_2673,N_2514);
or U3118 (N_3118,N_2923,N_2722);
nor U3119 (N_3119,N_2663,N_2957);
nor U3120 (N_3120,N_2766,N_2867);
nor U3121 (N_3121,N_2925,N_2970);
nand U3122 (N_3122,N_2658,N_2978);
and U3123 (N_3123,N_2710,N_2887);
nor U3124 (N_3124,N_2917,N_2607);
or U3125 (N_3125,N_2683,N_2671);
and U3126 (N_3126,N_2949,N_2809);
and U3127 (N_3127,N_2711,N_2746);
or U3128 (N_3128,N_2757,N_2727);
nor U3129 (N_3129,N_2891,N_2566);
nand U3130 (N_3130,N_2812,N_2659);
nand U3131 (N_3131,N_2677,N_2984);
nor U3132 (N_3132,N_2906,N_2996);
nor U3133 (N_3133,N_2791,N_2584);
nor U3134 (N_3134,N_2702,N_2518);
or U3135 (N_3135,N_2686,N_2939);
xor U3136 (N_3136,N_2511,N_2824);
or U3137 (N_3137,N_2653,N_2969);
nand U3138 (N_3138,N_2567,N_2731);
nand U3139 (N_3139,N_2918,N_2853);
and U3140 (N_3140,N_2639,N_2856);
nand U3141 (N_3141,N_2993,N_2728);
or U3142 (N_3142,N_2537,N_2785);
nand U3143 (N_3143,N_2899,N_2976);
nand U3144 (N_3144,N_2709,N_2953);
nor U3145 (N_3145,N_2516,N_2948);
and U3146 (N_3146,N_2688,N_2602);
or U3147 (N_3147,N_2549,N_2810);
nor U3148 (N_3148,N_2903,N_2936);
or U3149 (N_3149,N_2777,N_2841);
and U3150 (N_3150,N_2869,N_2696);
nor U3151 (N_3151,N_2695,N_2578);
nor U3152 (N_3152,N_2944,N_2538);
nor U3153 (N_3153,N_2717,N_2907);
nand U3154 (N_3154,N_2764,N_2838);
nand U3155 (N_3155,N_2563,N_2795);
and U3156 (N_3156,N_2591,N_2921);
and U3157 (N_3157,N_2527,N_2595);
or U3158 (N_3158,N_2571,N_2857);
and U3159 (N_3159,N_2884,N_2901);
or U3160 (N_3160,N_2821,N_2519);
nand U3161 (N_3161,N_2848,N_2735);
nand U3162 (N_3162,N_2935,N_2562);
and U3163 (N_3163,N_2929,N_2998);
or U3164 (N_3164,N_2641,N_2564);
nor U3165 (N_3165,N_2956,N_2629);
xnor U3166 (N_3166,N_2657,N_2862);
nand U3167 (N_3167,N_2983,N_2733);
or U3168 (N_3168,N_2773,N_2530);
and U3169 (N_3169,N_2794,N_2623);
nor U3170 (N_3170,N_2588,N_2701);
and U3171 (N_3171,N_2640,N_2667);
and U3172 (N_3172,N_2715,N_2632);
nand U3173 (N_3173,N_2974,N_2509);
or U3174 (N_3174,N_2582,N_2814);
and U3175 (N_3175,N_2836,N_2756);
xor U3176 (N_3176,N_2738,N_2865);
and U3177 (N_3177,N_2587,N_2609);
nand U3178 (N_3178,N_2580,N_2889);
nor U3179 (N_3179,N_2742,N_2775);
nor U3180 (N_3180,N_2557,N_2554);
nor U3181 (N_3181,N_2672,N_2866);
or U3182 (N_3182,N_2550,N_2790);
or U3183 (N_3183,N_2753,N_2828);
nor U3184 (N_3184,N_2616,N_2861);
nand U3185 (N_3185,N_2914,N_2635);
nand U3186 (N_3186,N_2547,N_2512);
or U3187 (N_3187,N_2977,N_2719);
and U3188 (N_3188,N_2768,N_2816);
or U3189 (N_3189,N_2776,N_2577);
nor U3190 (N_3190,N_2900,N_2613);
nor U3191 (N_3191,N_2593,N_2533);
nand U3192 (N_3192,N_2743,N_2979);
nand U3193 (N_3193,N_2761,N_2877);
xnor U3194 (N_3194,N_2654,N_2922);
nor U3195 (N_3195,N_2898,N_2952);
nand U3196 (N_3196,N_2780,N_2909);
and U3197 (N_3197,N_2561,N_2624);
or U3198 (N_3198,N_2881,N_2919);
nand U3199 (N_3199,N_2638,N_2886);
or U3200 (N_3200,N_2502,N_2845);
nor U3201 (N_3201,N_2843,N_2504);
and U3202 (N_3202,N_2712,N_2870);
nor U3203 (N_3203,N_2665,N_2823);
or U3204 (N_3204,N_2937,N_2574);
or U3205 (N_3205,N_2703,N_2829);
nand U3206 (N_3206,N_2548,N_2694);
and U3207 (N_3207,N_2526,N_2852);
and U3208 (N_3208,N_2615,N_2693);
and U3209 (N_3209,N_2985,N_2646);
nor U3210 (N_3210,N_2938,N_2682);
nor U3211 (N_3211,N_2774,N_2612);
and U3212 (N_3212,N_2882,N_2965);
and U3213 (N_3213,N_2597,N_2680);
nor U3214 (N_3214,N_2930,N_2531);
nand U3215 (N_3215,N_2648,N_2546);
nand U3216 (N_3216,N_2767,N_2802);
or U3217 (N_3217,N_2888,N_2837);
nor U3218 (N_3218,N_2762,N_2804);
and U3219 (N_3219,N_2826,N_2971);
nand U3220 (N_3220,N_2573,N_2589);
or U3221 (N_3221,N_2541,N_2614);
nand U3222 (N_3222,N_2916,N_2555);
and U3223 (N_3223,N_2849,N_2959);
nand U3224 (N_3224,N_2759,N_2675);
or U3225 (N_3225,N_2920,N_2800);
and U3226 (N_3226,N_2796,N_2636);
xnor U3227 (N_3227,N_2542,N_2507);
and U3228 (N_3228,N_2510,N_2630);
nand U3229 (N_3229,N_2830,N_2643);
and U3230 (N_3230,N_2599,N_2520);
or U3231 (N_3231,N_2634,N_2817);
and U3232 (N_3232,N_2610,N_2741);
nor U3233 (N_3233,N_2669,N_2569);
nor U3234 (N_3234,N_2890,N_2652);
nor U3235 (N_3235,N_2850,N_2807);
nor U3236 (N_3236,N_2782,N_2689);
and U3237 (N_3237,N_2885,N_2868);
and U3238 (N_3238,N_2813,N_2778);
or U3239 (N_3239,N_2940,N_2932);
and U3240 (N_3240,N_2718,N_2943);
nand U3241 (N_3241,N_2706,N_2844);
nand U3242 (N_3242,N_2608,N_2633);
nor U3243 (N_3243,N_2846,N_2896);
or U3244 (N_3244,N_2892,N_2912);
and U3245 (N_3245,N_2532,N_2552);
nor U3246 (N_3246,N_2528,N_2819);
or U3247 (N_3247,N_2832,N_2834);
and U3248 (N_3248,N_2619,N_2989);
nand U3249 (N_3249,N_2822,N_2792);
nand U3250 (N_3250,N_2588,N_2813);
and U3251 (N_3251,N_2685,N_2667);
or U3252 (N_3252,N_2572,N_2680);
xnor U3253 (N_3253,N_2865,N_2774);
and U3254 (N_3254,N_2852,N_2982);
and U3255 (N_3255,N_2925,N_2553);
nand U3256 (N_3256,N_2963,N_2763);
nor U3257 (N_3257,N_2650,N_2779);
or U3258 (N_3258,N_2627,N_2991);
and U3259 (N_3259,N_2756,N_2986);
or U3260 (N_3260,N_2641,N_2760);
and U3261 (N_3261,N_2738,N_2513);
or U3262 (N_3262,N_2724,N_2840);
or U3263 (N_3263,N_2640,N_2853);
and U3264 (N_3264,N_2964,N_2797);
or U3265 (N_3265,N_2702,N_2937);
nor U3266 (N_3266,N_2776,N_2909);
and U3267 (N_3267,N_2687,N_2607);
nand U3268 (N_3268,N_2931,N_2650);
nand U3269 (N_3269,N_2526,N_2789);
xnor U3270 (N_3270,N_2590,N_2545);
nor U3271 (N_3271,N_2957,N_2772);
nor U3272 (N_3272,N_2538,N_2664);
or U3273 (N_3273,N_2905,N_2969);
or U3274 (N_3274,N_2516,N_2534);
nor U3275 (N_3275,N_2958,N_2554);
or U3276 (N_3276,N_2678,N_2556);
nand U3277 (N_3277,N_2823,N_2971);
nand U3278 (N_3278,N_2555,N_2500);
and U3279 (N_3279,N_2917,N_2628);
nand U3280 (N_3280,N_2541,N_2770);
or U3281 (N_3281,N_2721,N_2830);
nand U3282 (N_3282,N_2637,N_2893);
or U3283 (N_3283,N_2510,N_2651);
nand U3284 (N_3284,N_2788,N_2590);
and U3285 (N_3285,N_2871,N_2617);
nor U3286 (N_3286,N_2635,N_2897);
nand U3287 (N_3287,N_2908,N_2894);
nor U3288 (N_3288,N_2698,N_2893);
or U3289 (N_3289,N_2709,N_2594);
or U3290 (N_3290,N_2832,N_2974);
or U3291 (N_3291,N_2590,N_2829);
or U3292 (N_3292,N_2781,N_2506);
and U3293 (N_3293,N_2714,N_2664);
nor U3294 (N_3294,N_2811,N_2992);
or U3295 (N_3295,N_2729,N_2807);
nand U3296 (N_3296,N_2525,N_2632);
nand U3297 (N_3297,N_2513,N_2805);
or U3298 (N_3298,N_2707,N_2814);
nand U3299 (N_3299,N_2834,N_2983);
nand U3300 (N_3300,N_2923,N_2863);
and U3301 (N_3301,N_2960,N_2616);
or U3302 (N_3302,N_2886,N_2840);
and U3303 (N_3303,N_2515,N_2585);
nand U3304 (N_3304,N_2667,N_2613);
and U3305 (N_3305,N_2947,N_2581);
or U3306 (N_3306,N_2928,N_2607);
nor U3307 (N_3307,N_2543,N_2504);
and U3308 (N_3308,N_2774,N_2644);
or U3309 (N_3309,N_2782,N_2947);
or U3310 (N_3310,N_2605,N_2723);
or U3311 (N_3311,N_2541,N_2795);
nor U3312 (N_3312,N_2932,N_2747);
and U3313 (N_3313,N_2575,N_2807);
nor U3314 (N_3314,N_2603,N_2818);
nor U3315 (N_3315,N_2579,N_2970);
or U3316 (N_3316,N_2727,N_2574);
and U3317 (N_3317,N_2558,N_2790);
or U3318 (N_3318,N_2676,N_2612);
and U3319 (N_3319,N_2521,N_2879);
nand U3320 (N_3320,N_2987,N_2943);
or U3321 (N_3321,N_2825,N_2921);
or U3322 (N_3322,N_2520,N_2644);
nand U3323 (N_3323,N_2932,N_2979);
and U3324 (N_3324,N_2864,N_2743);
nor U3325 (N_3325,N_2697,N_2727);
nand U3326 (N_3326,N_2869,N_2546);
nand U3327 (N_3327,N_2814,N_2763);
and U3328 (N_3328,N_2896,N_2832);
nand U3329 (N_3329,N_2891,N_2542);
or U3330 (N_3330,N_2548,N_2649);
and U3331 (N_3331,N_2733,N_2671);
and U3332 (N_3332,N_2639,N_2588);
nand U3333 (N_3333,N_2603,N_2544);
and U3334 (N_3334,N_2778,N_2823);
and U3335 (N_3335,N_2802,N_2587);
and U3336 (N_3336,N_2782,N_2778);
nor U3337 (N_3337,N_2616,N_2988);
or U3338 (N_3338,N_2716,N_2877);
and U3339 (N_3339,N_2966,N_2953);
nand U3340 (N_3340,N_2870,N_2865);
nor U3341 (N_3341,N_2632,N_2722);
nor U3342 (N_3342,N_2517,N_2504);
nor U3343 (N_3343,N_2829,N_2927);
nor U3344 (N_3344,N_2888,N_2605);
and U3345 (N_3345,N_2921,N_2698);
and U3346 (N_3346,N_2550,N_2585);
and U3347 (N_3347,N_2568,N_2920);
nand U3348 (N_3348,N_2910,N_2922);
nor U3349 (N_3349,N_2753,N_2638);
and U3350 (N_3350,N_2568,N_2660);
and U3351 (N_3351,N_2524,N_2538);
and U3352 (N_3352,N_2881,N_2521);
nor U3353 (N_3353,N_2935,N_2805);
or U3354 (N_3354,N_2679,N_2673);
or U3355 (N_3355,N_2899,N_2642);
or U3356 (N_3356,N_2586,N_2923);
xnor U3357 (N_3357,N_2944,N_2812);
or U3358 (N_3358,N_2882,N_2527);
nor U3359 (N_3359,N_2552,N_2956);
nand U3360 (N_3360,N_2503,N_2827);
or U3361 (N_3361,N_2695,N_2869);
or U3362 (N_3362,N_2822,N_2767);
or U3363 (N_3363,N_2750,N_2836);
or U3364 (N_3364,N_2700,N_2975);
nand U3365 (N_3365,N_2753,N_2676);
nand U3366 (N_3366,N_2725,N_2968);
or U3367 (N_3367,N_2521,N_2874);
nor U3368 (N_3368,N_2685,N_2779);
or U3369 (N_3369,N_2886,N_2712);
nand U3370 (N_3370,N_2658,N_2708);
or U3371 (N_3371,N_2643,N_2828);
nand U3372 (N_3372,N_2594,N_2563);
nand U3373 (N_3373,N_2832,N_2610);
nor U3374 (N_3374,N_2569,N_2738);
or U3375 (N_3375,N_2927,N_2761);
or U3376 (N_3376,N_2774,N_2740);
nor U3377 (N_3377,N_2759,N_2690);
and U3378 (N_3378,N_2838,N_2863);
nand U3379 (N_3379,N_2750,N_2642);
or U3380 (N_3380,N_2706,N_2803);
nor U3381 (N_3381,N_2895,N_2820);
or U3382 (N_3382,N_2763,N_2830);
or U3383 (N_3383,N_2600,N_2970);
nor U3384 (N_3384,N_2674,N_2814);
or U3385 (N_3385,N_2963,N_2617);
and U3386 (N_3386,N_2507,N_2674);
or U3387 (N_3387,N_2524,N_2766);
nor U3388 (N_3388,N_2572,N_2643);
nor U3389 (N_3389,N_2888,N_2627);
nor U3390 (N_3390,N_2991,N_2591);
nand U3391 (N_3391,N_2784,N_2648);
nor U3392 (N_3392,N_2588,N_2865);
or U3393 (N_3393,N_2526,N_2864);
or U3394 (N_3394,N_2734,N_2720);
or U3395 (N_3395,N_2728,N_2925);
or U3396 (N_3396,N_2657,N_2787);
and U3397 (N_3397,N_2548,N_2782);
or U3398 (N_3398,N_2838,N_2840);
and U3399 (N_3399,N_2877,N_2712);
and U3400 (N_3400,N_2929,N_2561);
nor U3401 (N_3401,N_2610,N_2856);
nand U3402 (N_3402,N_2709,N_2990);
and U3403 (N_3403,N_2815,N_2520);
and U3404 (N_3404,N_2982,N_2962);
nor U3405 (N_3405,N_2585,N_2716);
and U3406 (N_3406,N_2923,N_2682);
xnor U3407 (N_3407,N_2948,N_2627);
or U3408 (N_3408,N_2743,N_2564);
or U3409 (N_3409,N_2806,N_2631);
or U3410 (N_3410,N_2889,N_2656);
nand U3411 (N_3411,N_2545,N_2694);
and U3412 (N_3412,N_2778,N_2990);
nand U3413 (N_3413,N_2924,N_2750);
or U3414 (N_3414,N_2737,N_2806);
nor U3415 (N_3415,N_2916,N_2599);
or U3416 (N_3416,N_2825,N_2696);
nand U3417 (N_3417,N_2639,N_2875);
or U3418 (N_3418,N_2530,N_2630);
nor U3419 (N_3419,N_2729,N_2599);
nand U3420 (N_3420,N_2681,N_2831);
and U3421 (N_3421,N_2510,N_2615);
nand U3422 (N_3422,N_2877,N_2789);
nand U3423 (N_3423,N_2960,N_2961);
and U3424 (N_3424,N_2630,N_2964);
or U3425 (N_3425,N_2806,N_2725);
and U3426 (N_3426,N_2554,N_2679);
or U3427 (N_3427,N_2675,N_2778);
and U3428 (N_3428,N_2769,N_2938);
and U3429 (N_3429,N_2529,N_2947);
and U3430 (N_3430,N_2510,N_2501);
nor U3431 (N_3431,N_2586,N_2939);
and U3432 (N_3432,N_2907,N_2752);
nor U3433 (N_3433,N_2846,N_2832);
and U3434 (N_3434,N_2513,N_2509);
and U3435 (N_3435,N_2745,N_2790);
and U3436 (N_3436,N_2836,N_2563);
nand U3437 (N_3437,N_2585,N_2553);
and U3438 (N_3438,N_2649,N_2537);
and U3439 (N_3439,N_2861,N_2978);
nand U3440 (N_3440,N_2845,N_2670);
nor U3441 (N_3441,N_2972,N_2601);
xor U3442 (N_3442,N_2616,N_2644);
nor U3443 (N_3443,N_2646,N_2879);
nand U3444 (N_3444,N_2792,N_2924);
nor U3445 (N_3445,N_2954,N_2521);
nand U3446 (N_3446,N_2811,N_2659);
and U3447 (N_3447,N_2788,N_2525);
and U3448 (N_3448,N_2588,N_2930);
or U3449 (N_3449,N_2802,N_2599);
or U3450 (N_3450,N_2655,N_2590);
and U3451 (N_3451,N_2653,N_2657);
and U3452 (N_3452,N_2771,N_2910);
nand U3453 (N_3453,N_2911,N_2830);
nor U3454 (N_3454,N_2641,N_2823);
nand U3455 (N_3455,N_2512,N_2606);
nor U3456 (N_3456,N_2653,N_2893);
and U3457 (N_3457,N_2926,N_2993);
and U3458 (N_3458,N_2618,N_2901);
or U3459 (N_3459,N_2983,N_2524);
nand U3460 (N_3460,N_2976,N_2760);
or U3461 (N_3461,N_2736,N_2885);
or U3462 (N_3462,N_2892,N_2832);
and U3463 (N_3463,N_2504,N_2856);
nor U3464 (N_3464,N_2590,N_2542);
or U3465 (N_3465,N_2612,N_2982);
nand U3466 (N_3466,N_2988,N_2619);
nand U3467 (N_3467,N_2684,N_2539);
and U3468 (N_3468,N_2956,N_2533);
nand U3469 (N_3469,N_2984,N_2758);
or U3470 (N_3470,N_2673,N_2825);
nand U3471 (N_3471,N_2795,N_2898);
or U3472 (N_3472,N_2668,N_2882);
and U3473 (N_3473,N_2545,N_2620);
or U3474 (N_3474,N_2696,N_2683);
nor U3475 (N_3475,N_2941,N_2775);
nor U3476 (N_3476,N_2791,N_2808);
and U3477 (N_3477,N_2965,N_2841);
and U3478 (N_3478,N_2796,N_2772);
nand U3479 (N_3479,N_2865,N_2859);
or U3480 (N_3480,N_2724,N_2936);
nor U3481 (N_3481,N_2583,N_2972);
nand U3482 (N_3482,N_2871,N_2825);
nor U3483 (N_3483,N_2857,N_2546);
nand U3484 (N_3484,N_2787,N_2548);
nor U3485 (N_3485,N_2652,N_2704);
or U3486 (N_3486,N_2904,N_2819);
nand U3487 (N_3487,N_2674,N_2882);
and U3488 (N_3488,N_2680,N_2776);
or U3489 (N_3489,N_2832,N_2768);
or U3490 (N_3490,N_2611,N_2667);
nor U3491 (N_3491,N_2705,N_2908);
nor U3492 (N_3492,N_2876,N_2796);
or U3493 (N_3493,N_2591,N_2694);
nor U3494 (N_3494,N_2946,N_2645);
or U3495 (N_3495,N_2500,N_2917);
and U3496 (N_3496,N_2703,N_2969);
nor U3497 (N_3497,N_2561,N_2522);
nand U3498 (N_3498,N_2621,N_2720);
nor U3499 (N_3499,N_2783,N_2743);
nor U3500 (N_3500,N_3344,N_3138);
nand U3501 (N_3501,N_3036,N_3490);
nor U3502 (N_3502,N_3150,N_3332);
or U3503 (N_3503,N_3272,N_3194);
or U3504 (N_3504,N_3425,N_3083);
nor U3505 (N_3505,N_3325,N_3446);
or U3506 (N_3506,N_3008,N_3279);
nand U3507 (N_3507,N_3242,N_3248);
and U3508 (N_3508,N_3256,N_3171);
nor U3509 (N_3509,N_3159,N_3497);
nand U3510 (N_3510,N_3243,N_3265);
nand U3511 (N_3511,N_3317,N_3469);
or U3512 (N_3512,N_3125,N_3476);
nor U3513 (N_3513,N_3183,N_3240);
nor U3514 (N_3514,N_3191,N_3127);
and U3515 (N_3515,N_3419,N_3372);
nor U3516 (N_3516,N_3311,N_3312);
or U3517 (N_3517,N_3299,N_3407);
nor U3518 (N_3518,N_3468,N_3361);
nor U3519 (N_3519,N_3451,N_3428);
nor U3520 (N_3520,N_3188,N_3134);
nand U3521 (N_3521,N_3306,N_3146);
nor U3522 (N_3522,N_3137,N_3432);
nor U3523 (N_3523,N_3197,N_3066);
or U3524 (N_3524,N_3026,N_3394);
or U3525 (N_3525,N_3389,N_3274);
and U3526 (N_3526,N_3293,N_3283);
nand U3527 (N_3527,N_3411,N_3478);
or U3528 (N_3528,N_3143,N_3094);
nand U3529 (N_3529,N_3148,N_3319);
nand U3530 (N_3530,N_3330,N_3464);
nor U3531 (N_3531,N_3353,N_3075);
nor U3532 (N_3532,N_3483,N_3459);
nor U3533 (N_3533,N_3069,N_3168);
and U3534 (N_3534,N_3474,N_3103);
or U3535 (N_3535,N_3487,N_3374);
and U3536 (N_3536,N_3169,N_3456);
or U3537 (N_3537,N_3135,N_3467);
nand U3538 (N_3538,N_3465,N_3124);
nor U3539 (N_3539,N_3193,N_3393);
nand U3540 (N_3540,N_3345,N_3382);
nand U3541 (N_3541,N_3049,N_3218);
nand U3542 (N_3542,N_3212,N_3209);
nand U3543 (N_3543,N_3104,N_3430);
nand U3544 (N_3544,N_3485,N_3099);
and U3545 (N_3545,N_3285,N_3268);
nor U3546 (N_3546,N_3482,N_3053);
or U3547 (N_3547,N_3184,N_3220);
or U3548 (N_3548,N_3106,N_3014);
and U3549 (N_3549,N_3131,N_3488);
or U3550 (N_3550,N_3203,N_3117);
nand U3551 (N_3551,N_3065,N_3216);
and U3552 (N_3552,N_3313,N_3080);
nor U3553 (N_3553,N_3068,N_3043);
nand U3554 (N_3554,N_3315,N_3034);
nand U3555 (N_3555,N_3149,N_3471);
nor U3556 (N_3556,N_3375,N_3381);
nor U3557 (N_3557,N_3360,N_3038);
and U3558 (N_3558,N_3016,N_3233);
nor U3559 (N_3559,N_3264,N_3009);
and U3560 (N_3560,N_3320,N_3273);
nand U3561 (N_3561,N_3115,N_3002);
and U3562 (N_3562,N_3439,N_3076);
or U3563 (N_3563,N_3051,N_3335);
nor U3564 (N_3564,N_3185,N_3229);
nor U3565 (N_3565,N_3438,N_3084);
xnor U3566 (N_3566,N_3262,N_3057);
and U3567 (N_3567,N_3296,N_3145);
nand U3568 (N_3568,N_3082,N_3436);
or U3569 (N_3569,N_3481,N_3398);
nand U3570 (N_3570,N_3277,N_3322);
nand U3571 (N_3571,N_3055,N_3028);
or U3572 (N_3572,N_3371,N_3224);
nand U3573 (N_3573,N_3199,N_3118);
nor U3574 (N_3574,N_3391,N_3221);
nand U3575 (N_3575,N_3070,N_3271);
or U3576 (N_3576,N_3037,N_3045);
or U3577 (N_3577,N_3263,N_3473);
nand U3578 (N_3578,N_3392,N_3006);
nand U3579 (N_3579,N_3295,N_3180);
and U3580 (N_3580,N_3205,N_3219);
and U3581 (N_3581,N_3350,N_3208);
nand U3582 (N_3582,N_3211,N_3161);
nand U3583 (N_3583,N_3206,N_3287);
and U3584 (N_3584,N_3093,N_3302);
or U3585 (N_3585,N_3309,N_3318);
and U3586 (N_3586,N_3058,N_3200);
and U3587 (N_3587,N_3047,N_3217);
nor U3588 (N_3588,N_3192,N_3388);
nor U3589 (N_3589,N_3499,N_3177);
nor U3590 (N_3590,N_3415,N_3112);
and U3591 (N_3591,N_3433,N_3190);
nand U3592 (N_3592,N_3426,N_3025);
nand U3593 (N_3593,N_3449,N_3241);
nand U3594 (N_3594,N_3284,N_3061);
or U3595 (N_3595,N_3020,N_3368);
nor U3596 (N_3596,N_3158,N_3307);
or U3597 (N_3597,N_3128,N_3052);
or U3598 (N_3598,N_3223,N_3342);
nand U3599 (N_3599,N_3098,N_3440);
and U3600 (N_3600,N_3427,N_3461);
nor U3601 (N_3601,N_3250,N_3097);
nand U3602 (N_3602,N_3162,N_3489);
nand U3603 (N_3603,N_3039,N_3314);
or U3604 (N_3604,N_3179,N_3442);
nand U3605 (N_3605,N_3261,N_3386);
or U3606 (N_3606,N_3405,N_3207);
and U3607 (N_3607,N_3286,N_3226);
nand U3608 (N_3608,N_3042,N_3109);
nor U3609 (N_3609,N_3362,N_3289);
nor U3610 (N_3610,N_3404,N_3136);
or U3611 (N_3611,N_3422,N_3252);
or U3612 (N_3612,N_3401,N_3095);
nand U3613 (N_3613,N_3383,N_3420);
nor U3614 (N_3614,N_3369,N_3346);
nand U3615 (N_3615,N_3329,N_3282);
or U3616 (N_3616,N_3114,N_3347);
nor U3617 (N_3617,N_3139,N_3054);
nand U3618 (N_3618,N_3395,N_3321);
nand U3619 (N_3619,N_3238,N_3331);
and U3620 (N_3620,N_3067,N_3154);
nor U3621 (N_3621,N_3107,N_3012);
nor U3622 (N_3622,N_3280,N_3380);
nor U3623 (N_3623,N_3364,N_3140);
nor U3624 (N_3624,N_3081,N_3078);
or U3625 (N_3625,N_3379,N_3035);
or U3626 (N_3626,N_3133,N_3244);
nor U3627 (N_3627,N_3495,N_3384);
nor U3628 (N_3628,N_3166,N_3044);
or U3629 (N_3629,N_3147,N_3406);
and U3630 (N_3630,N_3408,N_3215);
or U3631 (N_3631,N_3447,N_3387);
nor U3632 (N_3632,N_3003,N_3196);
and U3633 (N_3633,N_3048,N_3007);
nor U3634 (N_3634,N_3113,N_3351);
and U3635 (N_3635,N_3378,N_3290);
or U3636 (N_3636,N_3015,N_3399);
nor U3637 (N_3637,N_3018,N_3349);
and U3638 (N_3638,N_3023,N_3424);
nand U3639 (N_3639,N_3278,N_3258);
or U3640 (N_3640,N_3064,N_3298);
xor U3641 (N_3641,N_3452,N_3005);
nor U3642 (N_3642,N_3475,N_3021);
nand U3643 (N_3643,N_3308,N_3153);
and U3644 (N_3644,N_3327,N_3090);
nor U3645 (N_3645,N_3227,N_3412);
and U3646 (N_3646,N_3305,N_3431);
nor U3647 (N_3647,N_3477,N_3088);
nand U3648 (N_3648,N_3445,N_3291);
nor U3649 (N_3649,N_3297,N_3186);
nand U3650 (N_3650,N_3105,N_3496);
nand U3651 (N_3651,N_3484,N_3338);
or U3652 (N_3652,N_3120,N_3463);
or U3653 (N_3653,N_3435,N_3123);
nand U3654 (N_3654,N_3269,N_3072);
or U3655 (N_3655,N_3400,N_3071);
and U3656 (N_3656,N_3022,N_3249);
and U3657 (N_3657,N_3202,N_3413);
and U3658 (N_3658,N_3340,N_3236);
nor U3659 (N_3659,N_3175,N_3316);
nor U3660 (N_3660,N_3246,N_3418);
or U3661 (N_3661,N_3470,N_3460);
and U3662 (N_3662,N_3225,N_3050);
or U3663 (N_3663,N_3343,N_3390);
nor U3664 (N_3664,N_3234,N_3062);
nand U3665 (N_3665,N_3108,N_3195);
and U3666 (N_3666,N_3001,N_3472);
or U3667 (N_3667,N_3358,N_3030);
nor U3668 (N_3668,N_3228,N_3178);
and U3669 (N_3669,N_3356,N_3040);
nor U3670 (N_3670,N_3063,N_3181);
or U3671 (N_3671,N_3004,N_3486);
and U3672 (N_3672,N_3231,N_3152);
nor U3673 (N_3673,N_3414,N_3214);
or U3674 (N_3674,N_3276,N_3000);
nor U3675 (N_3675,N_3377,N_3174);
or U3676 (N_3676,N_3160,N_3126);
or U3677 (N_3677,N_3086,N_3434);
nand U3678 (N_3678,N_3167,N_3182);
and U3679 (N_3679,N_3100,N_3056);
nor U3680 (N_3680,N_3421,N_3450);
and U3681 (N_3681,N_3170,N_3257);
nor U3682 (N_3682,N_3232,N_3019);
and U3683 (N_3683,N_3294,N_3102);
or U3684 (N_3684,N_3443,N_3092);
nor U3685 (N_3685,N_3304,N_3101);
and U3686 (N_3686,N_3354,N_3365);
nand U3687 (N_3687,N_3033,N_3324);
or U3688 (N_3688,N_3198,N_3328);
or U3689 (N_3689,N_3089,N_3077);
nand U3690 (N_3690,N_3144,N_3011);
and U3691 (N_3691,N_3423,N_3457);
nand U3692 (N_3692,N_3010,N_3096);
and U3693 (N_3693,N_3213,N_3024);
and U3694 (N_3694,N_3275,N_3355);
and U3695 (N_3695,N_3060,N_3396);
or U3696 (N_3696,N_3245,N_3402);
nand U3697 (N_3697,N_3310,N_3156);
or U3698 (N_3698,N_3492,N_3448);
nand U3699 (N_3699,N_3336,N_3466);
or U3700 (N_3700,N_3403,N_3437);
and U3701 (N_3701,N_3441,N_3255);
and U3702 (N_3702,N_3352,N_3074);
and U3703 (N_3703,N_3480,N_3359);
xor U3704 (N_3704,N_3301,N_3046);
nand U3705 (N_3705,N_3130,N_3253);
or U3706 (N_3706,N_3363,N_3032);
nor U3707 (N_3707,N_3455,N_3087);
or U3708 (N_3708,N_3303,N_3453);
nand U3709 (N_3709,N_3172,N_3073);
or U3710 (N_3710,N_3348,N_3266);
or U3711 (N_3711,N_3454,N_3337);
nor U3712 (N_3712,N_3129,N_3479);
or U3713 (N_3713,N_3201,N_3339);
and U3714 (N_3714,N_3417,N_3121);
and U3715 (N_3715,N_3189,N_3416);
nor U3716 (N_3716,N_3119,N_3041);
nor U3717 (N_3717,N_3373,N_3357);
nand U3718 (N_3718,N_3267,N_3259);
nand U3719 (N_3719,N_3237,N_3409);
or U3720 (N_3720,N_3288,N_3085);
nand U3721 (N_3721,N_3163,N_3292);
and U3722 (N_3722,N_3164,N_3397);
or U3723 (N_3723,N_3027,N_3444);
and U3724 (N_3724,N_3251,N_3157);
nand U3725 (N_3725,N_3173,N_3410);
nand U3726 (N_3726,N_3341,N_3165);
nor U3727 (N_3727,N_3222,N_3491);
nand U3728 (N_3728,N_3210,N_3376);
nand U3729 (N_3729,N_3187,N_3132);
or U3730 (N_3730,N_3151,N_3270);
or U3731 (N_3731,N_3498,N_3116);
nor U3732 (N_3732,N_3204,N_3385);
nor U3733 (N_3733,N_3281,N_3323);
nor U3734 (N_3734,N_3111,N_3493);
and U3735 (N_3735,N_3031,N_3059);
and U3736 (N_3736,N_3013,N_3029);
nor U3737 (N_3737,N_3334,N_3458);
or U3738 (N_3738,N_3091,N_3370);
nor U3739 (N_3739,N_3110,N_3017);
xnor U3740 (N_3740,N_3235,N_3247);
and U3741 (N_3741,N_3254,N_3462);
nor U3742 (N_3742,N_3429,N_3141);
and U3743 (N_3743,N_3079,N_3230);
or U3744 (N_3744,N_3366,N_3142);
or U3745 (N_3745,N_3176,N_3333);
nor U3746 (N_3746,N_3155,N_3239);
nand U3747 (N_3747,N_3326,N_3367);
nand U3748 (N_3748,N_3494,N_3260);
nor U3749 (N_3749,N_3300,N_3122);
or U3750 (N_3750,N_3341,N_3220);
or U3751 (N_3751,N_3495,N_3338);
nand U3752 (N_3752,N_3045,N_3119);
or U3753 (N_3753,N_3220,N_3180);
nand U3754 (N_3754,N_3213,N_3365);
xnor U3755 (N_3755,N_3103,N_3269);
and U3756 (N_3756,N_3045,N_3279);
nand U3757 (N_3757,N_3270,N_3191);
xnor U3758 (N_3758,N_3490,N_3126);
nor U3759 (N_3759,N_3039,N_3499);
and U3760 (N_3760,N_3184,N_3167);
nor U3761 (N_3761,N_3058,N_3285);
or U3762 (N_3762,N_3168,N_3469);
nand U3763 (N_3763,N_3390,N_3170);
nor U3764 (N_3764,N_3463,N_3382);
nor U3765 (N_3765,N_3219,N_3156);
or U3766 (N_3766,N_3146,N_3326);
nor U3767 (N_3767,N_3172,N_3134);
or U3768 (N_3768,N_3062,N_3075);
nor U3769 (N_3769,N_3409,N_3351);
nand U3770 (N_3770,N_3333,N_3008);
or U3771 (N_3771,N_3433,N_3323);
and U3772 (N_3772,N_3036,N_3462);
and U3773 (N_3773,N_3196,N_3218);
or U3774 (N_3774,N_3342,N_3188);
and U3775 (N_3775,N_3051,N_3345);
or U3776 (N_3776,N_3291,N_3185);
nand U3777 (N_3777,N_3236,N_3232);
or U3778 (N_3778,N_3455,N_3496);
or U3779 (N_3779,N_3051,N_3418);
nor U3780 (N_3780,N_3131,N_3093);
or U3781 (N_3781,N_3109,N_3223);
or U3782 (N_3782,N_3274,N_3452);
and U3783 (N_3783,N_3328,N_3443);
nor U3784 (N_3784,N_3094,N_3412);
nor U3785 (N_3785,N_3142,N_3493);
nor U3786 (N_3786,N_3027,N_3421);
and U3787 (N_3787,N_3100,N_3458);
nor U3788 (N_3788,N_3317,N_3200);
xor U3789 (N_3789,N_3111,N_3354);
nor U3790 (N_3790,N_3122,N_3282);
or U3791 (N_3791,N_3468,N_3040);
and U3792 (N_3792,N_3055,N_3006);
nor U3793 (N_3793,N_3257,N_3247);
or U3794 (N_3794,N_3022,N_3195);
and U3795 (N_3795,N_3022,N_3393);
and U3796 (N_3796,N_3356,N_3052);
nand U3797 (N_3797,N_3009,N_3085);
nor U3798 (N_3798,N_3018,N_3001);
and U3799 (N_3799,N_3185,N_3036);
nor U3800 (N_3800,N_3407,N_3184);
or U3801 (N_3801,N_3428,N_3479);
and U3802 (N_3802,N_3052,N_3049);
or U3803 (N_3803,N_3310,N_3163);
and U3804 (N_3804,N_3371,N_3255);
or U3805 (N_3805,N_3455,N_3326);
nand U3806 (N_3806,N_3147,N_3489);
and U3807 (N_3807,N_3110,N_3207);
or U3808 (N_3808,N_3326,N_3384);
and U3809 (N_3809,N_3321,N_3241);
nor U3810 (N_3810,N_3351,N_3187);
and U3811 (N_3811,N_3217,N_3042);
and U3812 (N_3812,N_3398,N_3006);
or U3813 (N_3813,N_3077,N_3383);
nand U3814 (N_3814,N_3366,N_3133);
or U3815 (N_3815,N_3310,N_3075);
nand U3816 (N_3816,N_3120,N_3070);
nand U3817 (N_3817,N_3440,N_3428);
nor U3818 (N_3818,N_3467,N_3398);
nor U3819 (N_3819,N_3047,N_3094);
or U3820 (N_3820,N_3377,N_3284);
or U3821 (N_3821,N_3451,N_3012);
or U3822 (N_3822,N_3011,N_3424);
nand U3823 (N_3823,N_3487,N_3030);
or U3824 (N_3824,N_3025,N_3463);
xnor U3825 (N_3825,N_3346,N_3288);
and U3826 (N_3826,N_3348,N_3081);
and U3827 (N_3827,N_3301,N_3031);
or U3828 (N_3828,N_3211,N_3275);
or U3829 (N_3829,N_3101,N_3295);
nor U3830 (N_3830,N_3167,N_3175);
and U3831 (N_3831,N_3397,N_3024);
nor U3832 (N_3832,N_3495,N_3006);
nand U3833 (N_3833,N_3335,N_3407);
nor U3834 (N_3834,N_3171,N_3385);
nand U3835 (N_3835,N_3401,N_3069);
or U3836 (N_3836,N_3100,N_3480);
nand U3837 (N_3837,N_3161,N_3113);
nand U3838 (N_3838,N_3433,N_3343);
and U3839 (N_3839,N_3164,N_3314);
xor U3840 (N_3840,N_3155,N_3111);
nor U3841 (N_3841,N_3400,N_3488);
nand U3842 (N_3842,N_3413,N_3201);
nor U3843 (N_3843,N_3178,N_3444);
nor U3844 (N_3844,N_3483,N_3087);
and U3845 (N_3845,N_3015,N_3369);
nand U3846 (N_3846,N_3466,N_3107);
or U3847 (N_3847,N_3385,N_3301);
and U3848 (N_3848,N_3021,N_3271);
nor U3849 (N_3849,N_3258,N_3416);
or U3850 (N_3850,N_3414,N_3459);
nand U3851 (N_3851,N_3167,N_3278);
or U3852 (N_3852,N_3032,N_3360);
nor U3853 (N_3853,N_3351,N_3362);
nand U3854 (N_3854,N_3072,N_3238);
nand U3855 (N_3855,N_3363,N_3158);
and U3856 (N_3856,N_3023,N_3479);
or U3857 (N_3857,N_3356,N_3081);
nor U3858 (N_3858,N_3433,N_3280);
nand U3859 (N_3859,N_3315,N_3105);
nor U3860 (N_3860,N_3086,N_3081);
nand U3861 (N_3861,N_3134,N_3272);
or U3862 (N_3862,N_3390,N_3038);
nor U3863 (N_3863,N_3033,N_3363);
nor U3864 (N_3864,N_3036,N_3419);
nand U3865 (N_3865,N_3384,N_3057);
nand U3866 (N_3866,N_3464,N_3128);
and U3867 (N_3867,N_3426,N_3394);
nor U3868 (N_3868,N_3425,N_3093);
nor U3869 (N_3869,N_3221,N_3159);
nor U3870 (N_3870,N_3157,N_3095);
or U3871 (N_3871,N_3370,N_3064);
or U3872 (N_3872,N_3477,N_3300);
nor U3873 (N_3873,N_3402,N_3487);
nand U3874 (N_3874,N_3496,N_3478);
nand U3875 (N_3875,N_3149,N_3068);
nand U3876 (N_3876,N_3292,N_3138);
nor U3877 (N_3877,N_3215,N_3395);
nor U3878 (N_3878,N_3044,N_3382);
or U3879 (N_3879,N_3437,N_3343);
nand U3880 (N_3880,N_3275,N_3045);
and U3881 (N_3881,N_3167,N_3127);
or U3882 (N_3882,N_3364,N_3120);
nor U3883 (N_3883,N_3041,N_3090);
and U3884 (N_3884,N_3433,N_3491);
and U3885 (N_3885,N_3055,N_3021);
nor U3886 (N_3886,N_3157,N_3225);
or U3887 (N_3887,N_3278,N_3422);
and U3888 (N_3888,N_3039,N_3458);
or U3889 (N_3889,N_3285,N_3214);
and U3890 (N_3890,N_3078,N_3392);
nor U3891 (N_3891,N_3142,N_3152);
nand U3892 (N_3892,N_3420,N_3130);
or U3893 (N_3893,N_3028,N_3301);
and U3894 (N_3894,N_3184,N_3225);
and U3895 (N_3895,N_3145,N_3108);
nand U3896 (N_3896,N_3199,N_3442);
nor U3897 (N_3897,N_3265,N_3025);
nand U3898 (N_3898,N_3174,N_3272);
and U3899 (N_3899,N_3493,N_3490);
or U3900 (N_3900,N_3122,N_3168);
nand U3901 (N_3901,N_3026,N_3180);
nor U3902 (N_3902,N_3230,N_3161);
or U3903 (N_3903,N_3012,N_3014);
and U3904 (N_3904,N_3178,N_3247);
nor U3905 (N_3905,N_3497,N_3288);
or U3906 (N_3906,N_3455,N_3107);
and U3907 (N_3907,N_3095,N_3272);
nand U3908 (N_3908,N_3281,N_3038);
or U3909 (N_3909,N_3120,N_3452);
nand U3910 (N_3910,N_3457,N_3297);
or U3911 (N_3911,N_3296,N_3393);
nand U3912 (N_3912,N_3492,N_3498);
nand U3913 (N_3913,N_3134,N_3344);
or U3914 (N_3914,N_3303,N_3224);
and U3915 (N_3915,N_3194,N_3269);
nor U3916 (N_3916,N_3237,N_3139);
nor U3917 (N_3917,N_3138,N_3301);
or U3918 (N_3918,N_3359,N_3379);
xnor U3919 (N_3919,N_3256,N_3473);
nor U3920 (N_3920,N_3144,N_3159);
and U3921 (N_3921,N_3184,N_3195);
or U3922 (N_3922,N_3095,N_3288);
nor U3923 (N_3923,N_3339,N_3005);
and U3924 (N_3924,N_3084,N_3348);
or U3925 (N_3925,N_3065,N_3017);
and U3926 (N_3926,N_3472,N_3241);
nand U3927 (N_3927,N_3305,N_3369);
nor U3928 (N_3928,N_3098,N_3498);
and U3929 (N_3929,N_3187,N_3042);
and U3930 (N_3930,N_3118,N_3070);
nand U3931 (N_3931,N_3192,N_3316);
nor U3932 (N_3932,N_3250,N_3337);
or U3933 (N_3933,N_3004,N_3419);
nand U3934 (N_3934,N_3226,N_3088);
nand U3935 (N_3935,N_3189,N_3493);
nand U3936 (N_3936,N_3202,N_3018);
nand U3937 (N_3937,N_3486,N_3140);
and U3938 (N_3938,N_3052,N_3092);
nor U3939 (N_3939,N_3488,N_3061);
and U3940 (N_3940,N_3428,N_3437);
and U3941 (N_3941,N_3422,N_3162);
and U3942 (N_3942,N_3269,N_3082);
nand U3943 (N_3943,N_3008,N_3386);
and U3944 (N_3944,N_3291,N_3097);
nor U3945 (N_3945,N_3133,N_3246);
nor U3946 (N_3946,N_3082,N_3286);
nand U3947 (N_3947,N_3164,N_3474);
nor U3948 (N_3948,N_3437,N_3398);
nand U3949 (N_3949,N_3365,N_3352);
nand U3950 (N_3950,N_3486,N_3118);
and U3951 (N_3951,N_3195,N_3491);
nor U3952 (N_3952,N_3270,N_3222);
nand U3953 (N_3953,N_3012,N_3176);
nor U3954 (N_3954,N_3031,N_3088);
nand U3955 (N_3955,N_3425,N_3073);
nor U3956 (N_3956,N_3310,N_3479);
and U3957 (N_3957,N_3190,N_3194);
or U3958 (N_3958,N_3098,N_3315);
or U3959 (N_3959,N_3415,N_3294);
nand U3960 (N_3960,N_3245,N_3263);
nor U3961 (N_3961,N_3162,N_3367);
nor U3962 (N_3962,N_3014,N_3462);
nand U3963 (N_3963,N_3091,N_3041);
or U3964 (N_3964,N_3095,N_3170);
and U3965 (N_3965,N_3151,N_3208);
and U3966 (N_3966,N_3271,N_3019);
and U3967 (N_3967,N_3347,N_3197);
nor U3968 (N_3968,N_3232,N_3421);
and U3969 (N_3969,N_3205,N_3487);
or U3970 (N_3970,N_3295,N_3323);
and U3971 (N_3971,N_3379,N_3071);
or U3972 (N_3972,N_3031,N_3303);
or U3973 (N_3973,N_3082,N_3116);
or U3974 (N_3974,N_3045,N_3033);
or U3975 (N_3975,N_3062,N_3443);
xor U3976 (N_3976,N_3400,N_3201);
nor U3977 (N_3977,N_3099,N_3276);
and U3978 (N_3978,N_3459,N_3147);
nor U3979 (N_3979,N_3347,N_3021);
nand U3980 (N_3980,N_3246,N_3319);
nand U3981 (N_3981,N_3250,N_3164);
or U3982 (N_3982,N_3476,N_3058);
nand U3983 (N_3983,N_3158,N_3152);
nor U3984 (N_3984,N_3469,N_3458);
or U3985 (N_3985,N_3212,N_3111);
nor U3986 (N_3986,N_3333,N_3489);
nand U3987 (N_3987,N_3314,N_3098);
nor U3988 (N_3988,N_3021,N_3181);
and U3989 (N_3989,N_3197,N_3482);
or U3990 (N_3990,N_3081,N_3474);
nor U3991 (N_3991,N_3406,N_3288);
nand U3992 (N_3992,N_3060,N_3052);
xnor U3993 (N_3993,N_3484,N_3021);
nand U3994 (N_3994,N_3020,N_3393);
nor U3995 (N_3995,N_3455,N_3428);
and U3996 (N_3996,N_3420,N_3038);
and U3997 (N_3997,N_3345,N_3259);
nand U3998 (N_3998,N_3130,N_3090);
or U3999 (N_3999,N_3400,N_3240);
or U4000 (N_4000,N_3625,N_3525);
or U4001 (N_4001,N_3852,N_3799);
nand U4002 (N_4002,N_3582,N_3657);
nor U4003 (N_4003,N_3667,N_3921);
and U4004 (N_4004,N_3792,N_3930);
and U4005 (N_4005,N_3958,N_3789);
nor U4006 (N_4006,N_3669,N_3650);
nand U4007 (N_4007,N_3656,N_3658);
and U4008 (N_4008,N_3516,N_3998);
nand U4009 (N_4009,N_3855,N_3816);
nor U4010 (N_4010,N_3725,N_3660);
nor U4011 (N_4011,N_3906,N_3996);
nand U4012 (N_4012,N_3726,N_3954);
or U4013 (N_4013,N_3914,N_3812);
nand U4014 (N_4014,N_3598,N_3741);
or U4015 (N_4015,N_3808,N_3763);
nand U4016 (N_4016,N_3675,N_3963);
nor U4017 (N_4017,N_3527,N_3663);
and U4018 (N_4018,N_3857,N_3835);
nor U4019 (N_4019,N_3608,N_3715);
or U4020 (N_4020,N_3719,N_3992);
or U4021 (N_4021,N_3883,N_3563);
and U4022 (N_4022,N_3622,N_3874);
and U4023 (N_4023,N_3730,N_3579);
and U4024 (N_4024,N_3837,N_3912);
nand U4025 (N_4025,N_3793,N_3779);
or U4026 (N_4026,N_3803,N_3801);
nand U4027 (N_4027,N_3530,N_3616);
nor U4028 (N_4028,N_3588,N_3538);
nor U4029 (N_4029,N_3540,N_3897);
and U4030 (N_4030,N_3873,N_3638);
nor U4031 (N_4031,N_3981,N_3795);
or U4032 (N_4032,N_3737,N_3769);
and U4033 (N_4033,N_3811,N_3752);
nor U4034 (N_4034,N_3621,N_3768);
nand U4035 (N_4035,N_3676,N_3952);
nor U4036 (N_4036,N_3984,N_3896);
or U4037 (N_4037,N_3790,N_3871);
or U4038 (N_4038,N_3580,N_3640);
or U4039 (N_4039,N_3962,N_3888);
and U4040 (N_4040,N_3577,N_3648);
or U4041 (N_4041,N_3727,N_3970);
and U4042 (N_4042,N_3926,N_3750);
and U4043 (N_4043,N_3973,N_3544);
nor U4044 (N_4044,N_3681,N_3882);
or U4045 (N_4045,N_3806,N_3701);
nand U4046 (N_4046,N_3511,N_3546);
nor U4047 (N_4047,N_3710,N_3628);
nor U4048 (N_4048,N_3674,N_3576);
or U4049 (N_4049,N_3905,N_3629);
or U4050 (N_4050,N_3922,N_3917);
and U4051 (N_4051,N_3893,N_3673);
or U4052 (N_4052,N_3787,N_3610);
nor U4053 (N_4053,N_3594,N_3519);
or U4054 (N_4054,N_3678,N_3856);
nand U4055 (N_4055,N_3680,N_3533);
xor U4056 (N_4056,N_3743,N_3881);
or U4057 (N_4057,N_3908,N_3614);
nand U4058 (N_4058,N_3895,N_3925);
or U4059 (N_4059,N_3683,N_3612);
nand U4060 (N_4060,N_3634,N_3955);
and U4061 (N_4061,N_3771,N_3500);
or U4062 (N_4062,N_3501,N_3521);
nor U4063 (N_4063,N_3542,N_3575);
and U4064 (N_4064,N_3830,N_3786);
nor U4065 (N_4065,N_3976,N_3653);
and U4066 (N_4066,N_3817,N_3757);
and U4067 (N_4067,N_3631,N_3809);
nand U4068 (N_4068,N_3858,N_3760);
nand U4069 (N_4069,N_3553,N_3759);
or U4070 (N_4070,N_3929,N_3879);
nor U4071 (N_4071,N_3828,N_3884);
and U4072 (N_4072,N_3659,N_3554);
or U4073 (N_4073,N_3532,N_3700);
nor U4074 (N_4074,N_3581,N_3965);
nand U4075 (N_4075,N_3800,N_3911);
and U4076 (N_4076,N_3783,N_3593);
or U4077 (N_4077,N_3862,N_3744);
or U4078 (N_4078,N_3950,N_3788);
and U4079 (N_4079,N_3734,N_3875);
or U4080 (N_4080,N_3927,N_3985);
or U4081 (N_4081,N_3751,N_3724);
nor U4082 (N_4082,N_3991,N_3913);
or U4083 (N_4083,N_3565,N_3635);
and U4084 (N_4084,N_3758,N_3547);
nand U4085 (N_4085,N_3578,N_3643);
nand U4086 (N_4086,N_3765,N_3735);
nor U4087 (N_4087,N_3815,N_3591);
or U4088 (N_4088,N_3827,N_3632);
and U4089 (N_4089,N_3712,N_3961);
and U4090 (N_4090,N_3977,N_3924);
or U4091 (N_4091,N_3545,N_3587);
nand U4092 (N_4092,N_3918,N_3766);
nand U4093 (N_4093,N_3867,N_3732);
or U4094 (N_4094,N_3695,N_3604);
nor U4095 (N_4095,N_3550,N_3820);
and U4096 (N_4096,N_3601,N_3909);
and U4097 (N_4097,N_3620,N_3915);
and U4098 (N_4098,N_3818,N_3748);
and U4099 (N_4099,N_3518,N_3512);
nand U4100 (N_4100,N_3851,N_3599);
nor U4101 (N_4101,N_3987,N_3903);
nand U4102 (N_4102,N_3529,N_3507);
and U4103 (N_4103,N_3870,N_3861);
and U4104 (N_4104,N_3586,N_3574);
nand U4105 (N_4105,N_3627,N_3866);
and U4106 (N_4106,N_3777,N_3746);
nand U4107 (N_4107,N_3979,N_3933);
and U4108 (N_4108,N_3753,N_3974);
or U4109 (N_4109,N_3503,N_3729);
nor U4110 (N_4110,N_3531,N_3717);
or U4111 (N_4111,N_3824,N_3686);
nor U4112 (N_4112,N_3670,N_3953);
nand U4113 (N_4113,N_3571,N_3698);
or U4114 (N_4114,N_3931,N_3592);
nor U4115 (N_4115,N_3541,N_3975);
nand U4116 (N_4116,N_3902,N_3690);
nand U4117 (N_4117,N_3842,N_3802);
nor U4118 (N_4118,N_3754,N_3775);
nand U4119 (N_4119,N_3910,N_3891);
or U4120 (N_4120,N_3543,N_3684);
and U4121 (N_4121,N_3822,N_3968);
or U4122 (N_4122,N_3997,N_3878);
and U4123 (N_4123,N_3555,N_3739);
or U4124 (N_4124,N_3668,N_3920);
nor U4125 (N_4125,N_3615,N_3697);
and U4126 (N_4126,N_3772,N_3978);
nor U4127 (N_4127,N_3810,N_3646);
nor U4128 (N_4128,N_3645,N_3923);
nor U4129 (N_4129,N_3782,N_3679);
nand U4130 (N_4130,N_3986,N_3647);
nor U4131 (N_4131,N_3693,N_3662);
nand U4132 (N_4132,N_3943,N_3642);
and U4133 (N_4133,N_3651,N_3636);
nand U4134 (N_4134,N_3644,N_3784);
nand U4135 (N_4135,N_3585,N_3524);
and U4136 (N_4136,N_3904,N_3740);
nand U4137 (N_4137,N_3665,N_3928);
nor U4138 (N_4138,N_3664,N_3705);
or U4139 (N_4139,N_3637,N_3561);
nand U4140 (N_4140,N_3708,N_3781);
and U4141 (N_4141,N_3946,N_3590);
xor U4142 (N_4142,N_3694,N_3959);
nor U4143 (N_4143,N_3713,N_3814);
or U4144 (N_4144,N_3696,N_3773);
and U4145 (N_4145,N_3932,N_3839);
or U4146 (N_4146,N_3526,N_3890);
nand U4147 (N_4147,N_3617,N_3714);
or U4148 (N_4148,N_3687,N_3595);
and U4149 (N_4149,N_3639,N_3756);
and U4150 (N_4150,N_3600,N_3860);
or U4151 (N_4151,N_3819,N_3722);
nand U4152 (N_4152,N_3868,N_3723);
nand U4153 (N_4153,N_3682,N_3876);
nand U4154 (N_4154,N_3745,N_3613);
or U4155 (N_4155,N_3846,N_3502);
nor U4156 (N_4156,N_3887,N_3838);
nand U4157 (N_4157,N_3556,N_3564);
nand U4158 (N_4158,N_3534,N_3840);
and U4159 (N_4159,N_3559,N_3728);
nor U4160 (N_4160,N_3718,N_3654);
or U4161 (N_4161,N_3972,N_3509);
nor U4162 (N_4162,N_3843,N_3514);
nand U4163 (N_4163,N_3557,N_3520);
nand U4164 (N_4164,N_3938,N_3774);
or U4165 (N_4165,N_3731,N_3517);
or U4166 (N_4166,N_3949,N_3869);
nor U4167 (N_4167,N_3707,N_3951);
and U4168 (N_4168,N_3583,N_3900);
nand U4169 (N_4169,N_3677,N_3689);
nand U4170 (N_4170,N_3510,N_3562);
nand U4171 (N_4171,N_3649,N_3971);
nand U4172 (N_4172,N_3607,N_3834);
nand U4173 (N_4173,N_3807,N_3994);
and U4174 (N_4174,N_3692,N_3605);
or U4175 (N_4175,N_3685,N_3537);
or U4176 (N_4176,N_3894,N_3841);
nor U4177 (N_4177,N_3566,N_3848);
nand U4178 (N_4178,N_3504,N_3661);
nand U4179 (N_4179,N_3880,N_3966);
nand U4180 (N_4180,N_3936,N_3813);
and U4181 (N_4181,N_3733,N_3603);
nand U4182 (N_4182,N_3956,N_3989);
and U4183 (N_4183,N_3836,N_3889);
or U4184 (N_4184,N_3863,N_3633);
or U4185 (N_4185,N_3568,N_3791);
and U4186 (N_4186,N_3849,N_3877);
nor U4187 (N_4187,N_3854,N_3611);
or U4188 (N_4188,N_3778,N_3738);
or U4189 (N_4189,N_3691,N_3899);
or U4190 (N_4190,N_3702,N_3672);
nand U4191 (N_4191,N_3589,N_3755);
nand U4192 (N_4192,N_3780,N_3942);
nand U4193 (N_4193,N_3853,N_3859);
nor U4194 (N_4194,N_3560,N_3567);
nor U4195 (N_4195,N_3847,N_3655);
nand U4196 (N_4196,N_3845,N_3606);
nor U4197 (N_4197,N_3983,N_3990);
or U4198 (N_4198,N_3671,N_3721);
and U4199 (N_4199,N_3886,N_3624);
nor U4200 (N_4200,N_3515,N_3706);
and U4201 (N_4201,N_3941,N_3916);
nand U4202 (N_4202,N_3937,N_3865);
and U4203 (N_4203,N_3767,N_3967);
or U4204 (N_4204,N_3829,N_3513);
nand U4205 (N_4205,N_3805,N_3948);
nor U4206 (N_4206,N_3939,N_3993);
and U4207 (N_4207,N_3619,N_3919);
or U4208 (N_4208,N_3761,N_3569);
xnor U4209 (N_4209,N_3558,N_3864);
or U4210 (N_4210,N_3944,N_3764);
nand U4211 (N_4211,N_3626,N_3982);
nand U4212 (N_4212,N_3762,N_3535);
and U4213 (N_4213,N_3618,N_3506);
or U4214 (N_4214,N_3666,N_3572);
or U4215 (N_4215,N_3570,N_3548);
nand U4216 (N_4216,N_3945,N_3742);
and U4217 (N_4217,N_3823,N_3536);
nor U4218 (N_4218,N_3749,N_3797);
and U4219 (N_4219,N_3602,N_3850);
nor U4220 (N_4220,N_3747,N_3892);
and U4221 (N_4221,N_3609,N_3940);
or U4222 (N_4222,N_3833,N_3551);
nor U4223 (N_4223,N_3798,N_3804);
or U4224 (N_4224,N_3999,N_3736);
nor U4225 (N_4225,N_3539,N_3832);
nor U4226 (N_4226,N_3831,N_3885);
nor U4227 (N_4227,N_3709,N_3980);
and U4228 (N_4228,N_3825,N_3549);
or U4229 (N_4229,N_3794,N_3522);
or U4230 (N_4230,N_3703,N_3796);
nor U4231 (N_4231,N_3597,N_3960);
or U4232 (N_4232,N_3995,N_3641);
or U4233 (N_4233,N_3770,N_3630);
nor U4234 (N_4234,N_3704,N_3573);
nand U4235 (N_4235,N_3969,N_3523);
and U4236 (N_4236,N_3776,N_3821);
and U4237 (N_4237,N_3584,N_3711);
nor U4238 (N_4238,N_3699,N_3907);
nand U4239 (N_4239,N_3935,N_3957);
nand U4240 (N_4240,N_3898,N_3947);
and U4241 (N_4241,N_3964,N_3552);
nor U4242 (N_4242,N_3785,N_3901);
nor U4243 (N_4243,N_3505,N_3934);
xnor U4244 (N_4244,N_3988,N_3528);
nand U4245 (N_4245,N_3720,N_3508);
nor U4246 (N_4246,N_3623,N_3826);
or U4247 (N_4247,N_3872,N_3716);
or U4248 (N_4248,N_3596,N_3652);
nand U4249 (N_4249,N_3688,N_3844);
nor U4250 (N_4250,N_3743,N_3792);
nor U4251 (N_4251,N_3781,N_3879);
nand U4252 (N_4252,N_3925,N_3642);
nand U4253 (N_4253,N_3899,N_3618);
nand U4254 (N_4254,N_3620,N_3817);
and U4255 (N_4255,N_3769,N_3511);
nand U4256 (N_4256,N_3988,N_3710);
and U4257 (N_4257,N_3946,N_3633);
and U4258 (N_4258,N_3762,N_3998);
nor U4259 (N_4259,N_3559,N_3814);
nor U4260 (N_4260,N_3506,N_3875);
nand U4261 (N_4261,N_3851,N_3585);
nand U4262 (N_4262,N_3936,N_3772);
and U4263 (N_4263,N_3940,N_3980);
or U4264 (N_4264,N_3826,N_3941);
nand U4265 (N_4265,N_3907,N_3858);
and U4266 (N_4266,N_3790,N_3646);
or U4267 (N_4267,N_3940,N_3752);
or U4268 (N_4268,N_3984,N_3822);
nor U4269 (N_4269,N_3896,N_3878);
or U4270 (N_4270,N_3656,N_3827);
nor U4271 (N_4271,N_3946,N_3517);
and U4272 (N_4272,N_3732,N_3724);
or U4273 (N_4273,N_3661,N_3769);
or U4274 (N_4274,N_3872,N_3552);
and U4275 (N_4275,N_3558,N_3721);
nand U4276 (N_4276,N_3964,N_3690);
nor U4277 (N_4277,N_3997,N_3934);
nand U4278 (N_4278,N_3824,N_3628);
nor U4279 (N_4279,N_3811,N_3520);
nand U4280 (N_4280,N_3683,N_3555);
or U4281 (N_4281,N_3628,N_3579);
and U4282 (N_4282,N_3647,N_3626);
or U4283 (N_4283,N_3774,N_3805);
nand U4284 (N_4284,N_3941,N_3800);
and U4285 (N_4285,N_3761,N_3977);
nand U4286 (N_4286,N_3663,N_3547);
nor U4287 (N_4287,N_3895,N_3813);
nand U4288 (N_4288,N_3801,N_3815);
nor U4289 (N_4289,N_3591,N_3698);
nor U4290 (N_4290,N_3550,N_3963);
or U4291 (N_4291,N_3820,N_3605);
and U4292 (N_4292,N_3538,N_3964);
nand U4293 (N_4293,N_3891,N_3831);
nand U4294 (N_4294,N_3803,N_3906);
nand U4295 (N_4295,N_3894,N_3748);
nor U4296 (N_4296,N_3580,N_3793);
or U4297 (N_4297,N_3743,N_3920);
or U4298 (N_4298,N_3606,N_3872);
and U4299 (N_4299,N_3581,N_3507);
or U4300 (N_4300,N_3811,N_3957);
nand U4301 (N_4301,N_3613,N_3712);
and U4302 (N_4302,N_3543,N_3888);
and U4303 (N_4303,N_3641,N_3756);
xnor U4304 (N_4304,N_3926,N_3766);
or U4305 (N_4305,N_3975,N_3963);
nand U4306 (N_4306,N_3636,N_3717);
nand U4307 (N_4307,N_3631,N_3869);
and U4308 (N_4308,N_3563,N_3585);
nor U4309 (N_4309,N_3981,N_3547);
nand U4310 (N_4310,N_3832,N_3573);
nor U4311 (N_4311,N_3855,N_3945);
and U4312 (N_4312,N_3543,N_3598);
nand U4313 (N_4313,N_3883,N_3579);
nand U4314 (N_4314,N_3997,N_3699);
nor U4315 (N_4315,N_3781,N_3585);
nor U4316 (N_4316,N_3871,N_3819);
nor U4317 (N_4317,N_3868,N_3580);
nor U4318 (N_4318,N_3701,N_3593);
and U4319 (N_4319,N_3727,N_3740);
and U4320 (N_4320,N_3730,N_3934);
and U4321 (N_4321,N_3630,N_3800);
nor U4322 (N_4322,N_3712,N_3889);
nor U4323 (N_4323,N_3772,N_3754);
and U4324 (N_4324,N_3795,N_3735);
or U4325 (N_4325,N_3892,N_3970);
nor U4326 (N_4326,N_3592,N_3733);
or U4327 (N_4327,N_3568,N_3682);
or U4328 (N_4328,N_3767,N_3924);
and U4329 (N_4329,N_3783,N_3866);
nor U4330 (N_4330,N_3966,N_3917);
nand U4331 (N_4331,N_3598,N_3642);
or U4332 (N_4332,N_3894,N_3542);
nand U4333 (N_4333,N_3594,N_3740);
nor U4334 (N_4334,N_3962,N_3607);
nand U4335 (N_4335,N_3705,N_3541);
nor U4336 (N_4336,N_3991,N_3855);
and U4337 (N_4337,N_3959,N_3956);
nand U4338 (N_4338,N_3589,N_3586);
nand U4339 (N_4339,N_3901,N_3701);
and U4340 (N_4340,N_3978,N_3795);
or U4341 (N_4341,N_3742,N_3672);
and U4342 (N_4342,N_3683,N_3923);
and U4343 (N_4343,N_3628,N_3885);
and U4344 (N_4344,N_3598,N_3718);
or U4345 (N_4345,N_3521,N_3835);
nor U4346 (N_4346,N_3562,N_3932);
xnor U4347 (N_4347,N_3728,N_3750);
nand U4348 (N_4348,N_3604,N_3759);
and U4349 (N_4349,N_3841,N_3829);
nor U4350 (N_4350,N_3722,N_3659);
and U4351 (N_4351,N_3590,N_3974);
and U4352 (N_4352,N_3841,N_3975);
nor U4353 (N_4353,N_3890,N_3822);
or U4354 (N_4354,N_3763,N_3604);
nand U4355 (N_4355,N_3897,N_3766);
nand U4356 (N_4356,N_3517,N_3600);
nand U4357 (N_4357,N_3625,N_3554);
nor U4358 (N_4358,N_3532,N_3768);
and U4359 (N_4359,N_3505,N_3774);
nor U4360 (N_4360,N_3968,N_3538);
nand U4361 (N_4361,N_3505,N_3784);
or U4362 (N_4362,N_3768,N_3859);
and U4363 (N_4363,N_3885,N_3608);
nand U4364 (N_4364,N_3756,N_3947);
nor U4365 (N_4365,N_3996,N_3834);
or U4366 (N_4366,N_3676,N_3959);
nand U4367 (N_4367,N_3880,N_3720);
nor U4368 (N_4368,N_3988,N_3824);
and U4369 (N_4369,N_3974,N_3777);
or U4370 (N_4370,N_3949,N_3677);
nor U4371 (N_4371,N_3928,N_3712);
nor U4372 (N_4372,N_3705,N_3977);
nand U4373 (N_4373,N_3683,N_3783);
and U4374 (N_4374,N_3850,N_3728);
nand U4375 (N_4375,N_3576,N_3556);
or U4376 (N_4376,N_3714,N_3983);
and U4377 (N_4377,N_3584,N_3818);
and U4378 (N_4378,N_3531,N_3657);
nor U4379 (N_4379,N_3992,N_3976);
nand U4380 (N_4380,N_3758,N_3618);
nand U4381 (N_4381,N_3975,N_3643);
and U4382 (N_4382,N_3711,N_3967);
and U4383 (N_4383,N_3767,N_3566);
nor U4384 (N_4384,N_3948,N_3774);
or U4385 (N_4385,N_3844,N_3883);
and U4386 (N_4386,N_3947,N_3949);
and U4387 (N_4387,N_3532,N_3545);
and U4388 (N_4388,N_3951,N_3968);
nor U4389 (N_4389,N_3576,N_3721);
nand U4390 (N_4390,N_3712,N_3971);
nor U4391 (N_4391,N_3615,N_3846);
nand U4392 (N_4392,N_3737,N_3604);
and U4393 (N_4393,N_3602,N_3575);
and U4394 (N_4394,N_3748,N_3965);
or U4395 (N_4395,N_3797,N_3664);
nor U4396 (N_4396,N_3646,N_3569);
or U4397 (N_4397,N_3566,N_3753);
nor U4398 (N_4398,N_3854,N_3631);
or U4399 (N_4399,N_3823,N_3623);
nand U4400 (N_4400,N_3959,N_3750);
nor U4401 (N_4401,N_3757,N_3834);
and U4402 (N_4402,N_3590,N_3994);
or U4403 (N_4403,N_3811,N_3529);
nor U4404 (N_4404,N_3653,N_3983);
or U4405 (N_4405,N_3523,N_3617);
and U4406 (N_4406,N_3579,N_3564);
nor U4407 (N_4407,N_3701,N_3638);
nor U4408 (N_4408,N_3680,N_3632);
or U4409 (N_4409,N_3589,N_3672);
and U4410 (N_4410,N_3667,N_3568);
nor U4411 (N_4411,N_3723,N_3889);
and U4412 (N_4412,N_3908,N_3881);
or U4413 (N_4413,N_3589,N_3668);
or U4414 (N_4414,N_3839,N_3525);
or U4415 (N_4415,N_3843,N_3870);
and U4416 (N_4416,N_3662,N_3963);
nand U4417 (N_4417,N_3771,N_3720);
and U4418 (N_4418,N_3879,N_3540);
nand U4419 (N_4419,N_3649,N_3770);
nor U4420 (N_4420,N_3993,N_3567);
and U4421 (N_4421,N_3958,N_3704);
or U4422 (N_4422,N_3805,N_3926);
nand U4423 (N_4423,N_3667,N_3516);
nor U4424 (N_4424,N_3646,N_3627);
and U4425 (N_4425,N_3650,N_3842);
nor U4426 (N_4426,N_3907,N_3695);
nor U4427 (N_4427,N_3896,N_3686);
and U4428 (N_4428,N_3820,N_3997);
nand U4429 (N_4429,N_3713,N_3627);
and U4430 (N_4430,N_3813,N_3984);
nand U4431 (N_4431,N_3768,N_3729);
nor U4432 (N_4432,N_3826,N_3688);
or U4433 (N_4433,N_3928,N_3882);
or U4434 (N_4434,N_3959,N_3945);
or U4435 (N_4435,N_3782,N_3621);
nor U4436 (N_4436,N_3503,N_3849);
or U4437 (N_4437,N_3643,N_3823);
xor U4438 (N_4438,N_3778,N_3877);
or U4439 (N_4439,N_3555,N_3924);
xnor U4440 (N_4440,N_3938,N_3545);
or U4441 (N_4441,N_3616,N_3611);
nor U4442 (N_4442,N_3758,N_3970);
nand U4443 (N_4443,N_3866,N_3760);
nor U4444 (N_4444,N_3868,N_3841);
or U4445 (N_4445,N_3802,N_3724);
nor U4446 (N_4446,N_3729,N_3650);
or U4447 (N_4447,N_3627,N_3601);
or U4448 (N_4448,N_3749,N_3980);
nand U4449 (N_4449,N_3718,N_3710);
and U4450 (N_4450,N_3530,N_3758);
nand U4451 (N_4451,N_3544,N_3618);
or U4452 (N_4452,N_3663,N_3725);
nand U4453 (N_4453,N_3606,N_3822);
and U4454 (N_4454,N_3735,N_3971);
or U4455 (N_4455,N_3552,N_3999);
or U4456 (N_4456,N_3983,N_3552);
or U4457 (N_4457,N_3948,N_3866);
nand U4458 (N_4458,N_3822,N_3745);
nand U4459 (N_4459,N_3565,N_3563);
nor U4460 (N_4460,N_3911,N_3977);
nor U4461 (N_4461,N_3652,N_3900);
nor U4462 (N_4462,N_3684,N_3621);
or U4463 (N_4463,N_3535,N_3551);
and U4464 (N_4464,N_3862,N_3564);
and U4465 (N_4465,N_3953,N_3698);
nor U4466 (N_4466,N_3803,N_3634);
nor U4467 (N_4467,N_3952,N_3845);
or U4468 (N_4468,N_3711,N_3664);
and U4469 (N_4469,N_3860,N_3832);
nor U4470 (N_4470,N_3892,N_3602);
or U4471 (N_4471,N_3511,N_3763);
and U4472 (N_4472,N_3641,N_3884);
or U4473 (N_4473,N_3926,N_3618);
nor U4474 (N_4474,N_3844,N_3840);
nor U4475 (N_4475,N_3878,N_3593);
and U4476 (N_4476,N_3555,N_3857);
nand U4477 (N_4477,N_3598,N_3775);
nor U4478 (N_4478,N_3977,N_3848);
nor U4479 (N_4479,N_3730,N_3912);
nand U4480 (N_4480,N_3732,N_3636);
nor U4481 (N_4481,N_3842,N_3512);
or U4482 (N_4482,N_3550,N_3715);
nor U4483 (N_4483,N_3709,N_3650);
nor U4484 (N_4484,N_3853,N_3731);
nor U4485 (N_4485,N_3609,N_3725);
nor U4486 (N_4486,N_3863,N_3605);
and U4487 (N_4487,N_3579,N_3724);
nor U4488 (N_4488,N_3994,N_3537);
and U4489 (N_4489,N_3887,N_3811);
and U4490 (N_4490,N_3550,N_3676);
nand U4491 (N_4491,N_3792,N_3851);
or U4492 (N_4492,N_3965,N_3616);
or U4493 (N_4493,N_3858,N_3533);
and U4494 (N_4494,N_3864,N_3595);
or U4495 (N_4495,N_3500,N_3854);
or U4496 (N_4496,N_3786,N_3982);
and U4497 (N_4497,N_3997,N_3779);
nand U4498 (N_4498,N_3617,N_3688);
nor U4499 (N_4499,N_3608,N_3726);
nand U4500 (N_4500,N_4447,N_4276);
nand U4501 (N_4501,N_4389,N_4403);
and U4502 (N_4502,N_4405,N_4420);
and U4503 (N_4503,N_4018,N_4382);
nor U4504 (N_4504,N_4413,N_4477);
nor U4505 (N_4505,N_4460,N_4252);
nor U4506 (N_4506,N_4054,N_4033);
or U4507 (N_4507,N_4498,N_4467);
nor U4508 (N_4508,N_4422,N_4220);
nor U4509 (N_4509,N_4107,N_4112);
nor U4510 (N_4510,N_4415,N_4156);
nor U4511 (N_4511,N_4343,N_4216);
nor U4512 (N_4512,N_4211,N_4019);
and U4513 (N_4513,N_4327,N_4177);
nor U4514 (N_4514,N_4393,N_4412);
and U4515 (N_4515,N_4298,N_4170);
or U4516 (N_4516,N_4072,N_4396);
and U4517 (N_4517,N_4093,N_4416);
and U4518 (N_4518,N_4102,N_4448);
and U4519 (N_4519,N_4402,N_4058);
or U4520 (N_4520,N_4340,N_4305);
nand U4521 (N_4521,N_4330,N_4478);
or U4522 (N_4522,N_4009,N_4414);
nor U4523 (N_4523,N_4001,N_4022);
nand U4524 (N_4524,N_4334,N_4206);
and U4525 (N_4525,N_4221,N_4345);
nand U4526 (N_4526,N_4237,N_4451);
nor U4527 (N_4527,N_4264,N_4331);
nand U4528 (N_4528,N_4494,N_4065);
and U4529 (N_4529,N_4388,N_4099);
nor U4530 (N_4530,N_4372,N_4197);
or U4531 (N_4531,N_4461,N_4231);
nand U4532 (N_4532,N_4247,N_4286);
and U4533 (N_4533,N_4463,N_4351);
and U4534 (N_4534,N_4239,N_4232);
and U4535 (N_4535,N_4418,N_4049);
and U4536 (N_4536,N_4084,N_4188);
nand U4537 (N_4537,N_4470,N_4333);
and U4538 (N_4538,N_4227,N_4344);
or U4539 (N_4539,N_4245,N_4150);
nor U4540 (N_4540,N_4229,N_4496);
nand U4541 (N_4541,N_4200,N_4238);
and U4542 (N_4542,N_4214,N_4152);
or U4543 (N_4543,N_4209,N_4132);
nor U4544 (N_4544,N_4302,N_4282);
nor U4545 (N_4545,N_4445,N_4429);
nor U4546 (N_4546,N_4374,N_4387);
nor U4547 (N_4547,N_4122,N_4202);
nor U4548 (N_4548,N_4439,N_4274);
nor U4549 (N_4549,N_4249,N_4381);
or U4550 (N_4550,N_4299,N_4228);
nor U4551 (N_4551,N_4427,N_4432);
and U4552 (N_4552,N_4390,N_4142);
nor U4553 (N_4553,N_4131,N_4240);
nor U4554 (N_4554,N_4160,N_4130);
nor U4555 (N_4555,N_4198,N_4043);
or U4556 (N_4556,N_4178,N_4215);
nand U4557 (N_4557,N_4315,N_4189);
and U4558 (N_4558,N_4459,N_4092);
or U4559 (N_4559,N_4377,N_4317);
nor U4560 (N_4560,N_4184,N_4320);
and U4561 (N_4561,N_4332,N_4140);
nor U4562 (N_4562,N_4135,N_4373);
and U4563 (N_4563,N_4086,N_4095);
nor U4564 (N_4564,N_4337,N_4110);
and U4565 (N_4565,N_4485,N_4079);
nor U4566 (N_4566,N_4431,N_4201);
nand U4567 (N_4567,N_4030,N_4452);
nor U4568 (N_4568,N_4159,N_4441);
and U4569 (N_4569,N_4032,N_4279);
and U4570 (N_4570,N_4260,N_4265);
nor U4571 (N_4571,N_4123,N_4325);
and U4572 (N_4572,N_4224,N_4078);
or U4573 (N_4573,N_4134,N_4357);
nor U4574 (N_4574,N_4275,N_4400);
and U4575 (N_4575,N_4410,N_4350);
or U4576 (N_4576,N_4409,N_4246);
and U4577 (N_4577,N_4495,N_4385);
and U4578 (N_4578,N_4208,N_4081);
nand U4579 (N_4579,N_4063,N_4103);
nor U4580 (N_4580,N_4386,N_4182);
nor U4581 (N_4581,N_4354,N_4052);
or U4582 (N_4582,N_4367,N_4436);
or U4583 (N_4583,N_4404,N_4048);
and U4584 (N_4584,N_4143,N_4196);
and U4585 (N_4585,N_4244,N_4491);
or U4586 (N_4586,N_4348,N_4213);
nor U4587 (N_4587,N_4497,N_4391);
nor U4588 (N_4588,N_4195,N_4281);
and U4589 (N_4589,N_4271,N_4465);
and U4590 (N_4590,N_4269,N_4154);
xor U4591 (N_4591,N_4472,N_4044);
or U4592 (N_4592,N_4185,N_4424);
nand U4593 (N_4593,N_4219,N_4453);
nand U4594 (N_4594,N_4181,N_4155);
nor U4595 (N_4595,N_4292,N_4067);
and U4596 (N_4596,N_4443,N_4187);
nor U4597 (N_4597,N_4157,N_4426);
nor U4598 (N_4598,N_4430,N_4456);
nor U4599 (N_4599,N_4336,N_4499);
nor U4600 (N_4600,N_4450,N_4289);
or U4601 (N_4601,N_4230,N_4248);
or U4602 (N_4602,N_4487,N_4251);
and U4603 (N_4603,N_4133,N_4011);
or U4604 (N_4604,N_4149,N_4002);
or U4605 (N_4605,N_4366,N_4446);
nand U4606 (N_4606,N_4303,N_4021);
nand U4607 (N_4607,N_4218,N_4338);
and U4608 (N_4608,N_4435,N_4293);
nand U4609 (N_4609,N_4318,N_4167);
or U4610 (N_4610,N_4068,N_4458);
and U4611 (N_4611,N_4359,N_4094);
or U4612 (N_4612,N_4129,N_4027);
and U4613 (N_4613,N_4361,N_4190);
and U4614 (N_4614,N_4145,N_4000);
and U4615 (N_4615,N_4347,N_4454);
or U4616 (N_4616,N_4124,N_4346);
nand U4617 (N_4617,N_4241,N_4136);
nor U4618 (N_4618,N_4304,N_4098);
or U4619 (N_4619,N_4395,N_4356);
nand U4620 (N_4620,N_4194,N_4013);
nor U4621 (N_4621,N_4100,N_4180);
or U4622 (N_4622,N_4073,N_4006);
nand U4623 (N_4623,N_4055,N_4113);
and U4624 (N_4624,N_4365,N_4308);
nand U4625 (N_4625,N_4166,N_4226);
nor U4626 (N_4626,N_4313,N_4116);
nor U4627 (N_4627,N_4045,N_4083);
nand U4628 (N_4628,N_4088,N_4258);
nand U4629 (N_4629,N_4360,N_4162);
and U4630 (N_4630,N_4267,N_4480);
or U4631 (N_4631,N_4053,N_4203);
nor U4632 (N_4632,N_4060,N_4146);
and U4633 (N_4633,N_4121,N_4471);
or U4634 (N_4634,N_4421,N_4070);
nor U4635 (N_4635,N_4321,N_4464);
xnor U4636 (N_4636,N_4301,N_4437);
nor U4637 (N_4637,N_4310,N_4438);
nand U4638 (N_4638,N_4036,N_4031);
nor U4639 (N_4639,N_4272,N_4242);
nand U4640 (N_4640,N_4175,N_4392);
and U4641 (N_4641,N_4419,N_4141);
nand U4642 (N_4642,N_4212,N_4261);
and U4643 (N_4643,N_4139,N_4085);
nand U4644 (N_4644,N_4375,N_4349);
and U4645 (N_4645,N_4207,N_4316);
nor U4646 (N_4646,N_4089,N_4407);
or U4647 (N_4647,N_4080,N_4401);
or U4648 (N_4648,N_4128,N_4397);
nor U4649 (N_4649,N_4306,N_4341);
or U4650 (N_4650,N_4398,N_4379);
or U4651 (N_4651,N_4075,N_4172);
nand U4652 (N_4652,N_4294,N_4481);
or U4653 (N_4653,N_4369,N_4488);
nor U4654 (N_4654,N_4164,N_4257);
and U4655 (N_4655,N_4314,N_4061);
or U4656 (N_4656,N_4339,N_4004);
and U4657 (N_4657,N_4364,N_4066);
or U4658 (N_4658,N_4024,N_4176);
or U4659 (N_4659,N_4466,N_4284);
or U4660 (N_4660,N_4417,N_4479);
nor U4661 (N_4661,N_4342,N_4114);
nor U4662 (N_4662,N_4263,N_4290);
and U4663 (N_4663,N_4270,N_4191);
nor U4664 (N_4664,N_4322,N_4041);
xor U4665 (N_4665,N_4256,N_4371);
nor U4666 (N_4666,N_4362,N_4255);
nand U4667 (N_4667,N_4266,N_4101);
nor U4668 (N_4668,N_4283,N_4040);
or U4669 (N_4669,N_4090,N_4125);
and U4670 (N_4670,N_4076,N_4029);
and U4671 (N_4671,N_4425,N_4363);
and U4672 (N_4672,N_4056,N_4291);
nand U4673 (N_4673,N_4352,N_4236);
nor U4674 (N_4674,N_4297,N_4253);
and U4675 (N_4675,N_4038,N_4168);
or U4676 (N_4676,N_4111,N_4384);
or U4677 (N_4677,N_4468,N_4312);
or U4678 (N_4678,N_4469,N_4235);
or U4679 (N_4679,N_4370,N_4307);
nand U4680 (N_4680,N_4026,N_4484);
nor U4681 (N_4681,N_4428,N_4059);
or U4682 (N_4682,N_4074,N_4077);
nor U4683 (N_4683,N_4097,N_4151);
and U4684 (N_4684,N_4119,N_4295);
or U4685 (N_4685,N_4287,N_4173);
or U4686 (N_4686,N_4057,N_4309);
nand U4687 (N_4687,N_4117,N_4285);
and U4688 (N_4688,N_4126,N_4222);
nor U4689 (N_4689,N_4380,N_4474);
or U4690 (N_4690,N_4046,N_4008);
nor U4691 (N_4691,N_4169,N_4268);
nand U4692 (N_4692,N_4383,N_4475);
nor U4693 (N_4693,N_4183,N_4254);
and U4694 (N_4694,N_4288,N_4137);
and U4695 (N_4695,N_4378,N_4223);
nand U4696 (N_4696,N_4017,N_4091);
nor U4697 (N_4697,N_4442,N_4096);
and U4698 (N_4698,N_4012,N_4358);
nand U4699 (N_4699,N_4034,N_4042);
or U4700 (N_4700,N_4234,N_4051);
nand U4701 (N_4701,N_4047,N_4277);
nand U4702 (N_4702,N_4433,N_4071);
or U4703 (N_4703,N_4069,N_4174);
and U4704 (N_4704,N_4028,N_4311);
nand U4705 (N_4705,N_4104,N_4296);
or U4706 (N_4706,N_4186,N_4411);
nor U4707 (N_4707,N_4399,N_4225);
and U4708 (N_4708,N_4492,N_4493);
nand U4709 (N_4709,N_4050,N_4462);
nand U4710 (N_4710,N_4449,N_4138);
nor U4711 (N_4711,N_4106,N_4319);
and U4712 (N_4712,N_4483,N_4025);
nand U4713 (N_4713,N_4158,N_4233);
nand U4714 (N_4714,N_4250,N_4179);
nand U4715 (N_4715,N_4192,N_4408);
or U4716 (N_4716,N_4273,N_4204);
xor U4717 (N_4717,N_4376,N_4476);
or U4718 (N_4718,N_4353,N_4118);
nor U4719 (N_4719,N_4171,N_4105);
or U4720 (N_4720,N_4163,N_4482);
or U4721 (N_4721,N_4335,N_4064);
or U4722 (N_4722,N_4015,N_4217);
or U4723 (N_4723,N_4161,N_4486);
or U4724 (N_4724,N_4280,N_4210);
nand U4725 (N_4725,N_4037,N_4020);
and U4726 (N_4726,N_4005,N_4328);
and U4727 (N_4727,N_4148,N_4259);
nand U4728 (N_4728,N_4323,N_4473);
nand U4729 (N_4729,N_4368,N_4423);
nand U4730 (N_4730,N_4014,N_4355);
nor U4731 (N_4731,N_4457,N_4440);
nor U4732 (N_4732,N_4205,N_4300);
and U4733 (N_4733,N_4165,N_4035);
nand U4734 (N_4734,N_4434,N_4023);
nand U4735 (N_4735,N_4262,N_4490);
nor U4736 (N_4736,N_4153,N_4144);
nor U4737 (N_4737,N_4147,N_4329);
nor U4738 (N_4738,N_4087,N_4108);
nand U4739 (N_4739,N_4444,N_4016);
and U4740 (N_4740,N_4193,N_4489);
nand U4741 (N_4741,N_4115,N_4082);
nor U4742 (N_4742,N_4278,N_4127);
and U4743 (N_4743,N_4062,N_4010);
and U4744 (N_4744,N_4199,N_4109);
and U4745 (N_4745,N_4120,N_4394);
or U4746 (N_4746,N_4455,N_4039);
nor U4747 (N_4747,N_4406,N_4007);
and U4748 (N_4748,N_4326,N_4243);
and U4749 (N_4749,N_4324,N_4003);
or U4750 (N_4750,N_4499,N_4357);
nand U4751 (N_4751,N_4340,N_4417);
nand U4752 (N_4752,N_4496,N_4441);
nor U4753 (N_4753,N_4054,N_4347);
and U4754 (N_4754,N_4144,N_4398);
or U4755 (N_4755,N_4104,N_4185);
or U4756 (N_4756,N_4223,N_4270);
nor U4757 (N_4757,N_4088,N_4315);
or U4758 (N_4758,N_4207,N_4027);
or U4759 (N_4759,N_4287,N_4451);
or U4760 (N_4760,N_4174,N_4186);
nor U4761 (N_4761,N_4264,N_4407);
nand U4762 (N_4762,N_4067,N_4398);
nor U4763 (N_4763,N_4134,N_4069);
nor U4764 (N_4764,N_4202,N_4070);
nor U4765 (N_4765,N_4079,N_4119);
nor U4766 (N_4766,N_4181,N_4113);
nand U4767 (N_4767,N_4468,N_4059);
and U4768 (N_4768,N_4202,N_4493);
nand U4769 (N_4769,N_4331,N_4008);
nand U4770 (N_4770,N_4385,N_4445);
or U4771 (N_4771,N_4146,N_4248);
and U4772 (N_4772,N_4436,N_4389);
nor U4773 (N_4773,N_4442,N_4309);
nand U4774 (N_4774,N_4337,N_4038);
nor U4775 (N_4775,N_4063,N_4171);
nor U4776 (N_4776,N_4094,N_4430);
nor U4777 (N_4777,N_4387,N_4368);
or U4778 (N_4778,N_4046,N_4288);
nand U4779 (N_4779,N_4144,N_4427);
and U4780 (N_4780,N_4207,N_4338);
or U4781 (N_4781,N_4112,N_4467);
or U4782 (N_4782,N_4227,N_4244);
nor U4783 (N_4783,N_4241,N_4009);
nand U4784 (N_4784,N_4456,N_4141);
and U4785 (N_4785,N_4071,N_4257);
or U4786 (N_4786,N_4353,N_4281);
or U4787 (N_4787,N_4004,N_4103);
nor U4788 (N_4788,N_4168,N_4266);
or U4789 (N_4789,N_4005,N_4255);
and U4790 (N_4790,N_4411,N_4213);
and U4791 (N_4791,N_4029,N_4430);
nor U4792 (N_4792,N_4186,N_4441);
and U4793 (N_4793,N_4134,N_4203);
nand U4794 (N_4794,N_4102,N_4437);
or U4795 (N_4795,N_4361,N_4135);
or U4796 (N_4796,N_4302,N_4176);
nand U4797 (N_4797,N_4420,N_4318);
or U4798 (N_4798,N_4400,N_4051);
or U4799 (N_4799,N_4234,N_4293);
nand U4800 (N_4800,N_4219,N_4177);
nor U4801 (N_4801,N_4124,N_4178);
nor U4802 (N_4802,N_4086,N_4201);
or U4803 (N_4803,N_4115,N_4434);
and U4804 (N_4804,N_4350,N_4430);
nor U4805 (N_4805,N_4477,N_4255);
nand U4806 (N_4806,N_4496,N_4458);
and U4807 (N_4807,N_4425,N_4495);
and U4808 (N_4808,N_4129,N_4457);
or U4809 (N_4809,N_4463,N_4017);
and U4810 (N_4810,N_4277,N_4329);
nor U4811 (N_4811,N_4436,N_4365);
and U4812 (N_4812,N_4275,N_4130);
nand U4813 (N_4813,N_4474,N_4332);
and U4814 (N_4814,N_4304,N_4143);
nor U4815 (N_4815,N_4069,N_4484);
or U4816 (N_4816,N_4099,N_4162);
or U4817 (N_4817,N_4141,N_4165);
or U4818 (N_4818,N_4471,N_4384);
or U4819 (N_4819,N_4364,N_4033);
or U4820 (N_4820,N_4258,N_4202);
or U4821 (N_4821,N_4446,N_4483);
nand U4822 (N_4822,N_4228,N_4284);
or U4823 (N_4823,N_4051,N_4114);
and U4824 (N_4824,N_4392,N_4303);
nand U4825 (N_4825,N_4080,N_4290);
nand U4826 (N_4826,N_4357,N_4045);
or U4827 (N_4827,N_4429,N_4255);
or U4828 (N_4828,N_4476,N_4177);
and U4829 (N_4829,N_4385,N_4031);
or U4830 (N_4830,N_4358,N_4173);
or U4831 (N_4831,N_4138,N_4426);
nor U4832 (N_4832,N_4078,N_4441);
and U4833 (N_4833,N_4138,N_4146);
or U4834 (N_4834,N_4175,N_4115);
or U4835 (N_4835,N_4154,N_4303);
nand U4836 (N_4836,N_4399,N_4230);
nor U4837 (N_4837,N_4465,N_4330);
nor U4838 (N_4838,N_4171,N_4053);
and U4839 (N_4839,N_4347,N_4235);
nand U4840 (N_4840,N_4202,N_4246);
nand U4841 (N_4841,N_4222,N_4394);
nor U4842 (N_4842,N_4171,N_4277);
and U4843 (N_4843,N_4485,N_4002);
nand U4844 (N_4844,N_4240,N_4408);
or U4845 (N_4845,N_4489,N_4134);
or U4846 (N_4846,N_4188,N_4447);
nand U4847 (N_4847,N_4087,N_4370);
nor U4848 (N_4848,N_4277,N_4377);
and U4849 (N_4849,N_4499,N_4485);
nand U4850 (N_4850,N_4475,N_4293);
or U4851 (N_4851,N_4488,N_4272);
or U4852 (N_4852,N_4180,N_4434);
and U4853 (N_4853,N_4051,N_4205);
nor U4854 (N_4854,N_4269,N_4320);
or U4855 (N_4855,N_4326,N_4338);
nor U4856 (N_4856,N_4427,N_4480);
or U4857 (N_4857,N_4448,N_4277);
nand U4858 (N_4858,N_4356,N_4393);
nor U4859 (N_4859,N_4220,N_4425);
and U4860 (N_4860,N_4138,N_4395);
nand U4861 (N_4861,N_4161,N_4330);
nor U4862 (N_4862,N_4325,N_4099);
nor U4863 (N_4863,N_4387,N_4472);
or U4864 (N_4864,N_4250,N_4293);
and U4865 (N_4865,N_4022,N_4053);
or U4866 (N_4866,N_4127,N_4170);
nand U4867 (N_4867,N_4328,N_4204);
and U4868 (N_4868,N_4466,N_4010);
xnor U4869 (N_4869,N_4426,N_4482);
or U4870 (N_4870,N_4358,N_4061);
or U4871 (N_4871,N_4241,N_4401);
or U4872 (N_4872,N_4390,N_4092);
nand U4873 (N_4873,N_4463,N_4010);
nand U4874 (N_4874,N_4401,N_4368);
nor U4875 (N_4875,N_4116,N_4484);
nand U4876 (N_4876,N_4319,N_4003);
nor U4877 (N_4877,N_4353,N_4005);
and U4878 (N_4878,N_4066,N_4455);
nand U4879 (N_4879,N_4355,N_4317);
or U4880 (N_4880,N_4218,N_4286);
nand U4881 (N_4881,N_4189,N_4423);
nor U4882 (N_4882,N_4073,N_4165);
nand U4883 (N_4883,N_4477,N_4074);
nor U4884 (N_4884,N_4453,N_4183);
nand U4885 (N_4885,N_4071,N_4251);
or U4886 (N_4886,N_4000,N_4337);
nor U4887 (N_4887,N_4407,N_4224);
and U4888 (N_4888,N_4230,N_4396);
or U4889 (N_4889,N_4484,N_4001);
or U4890 (N_4890,N_4348,N_4053);
nor U4891 (N_4891,N_4339,N_4356);
or U4892 (N_4892,N_4432,N_4484);
or U4893 (N_4893,N_4008,N_4393);
and U4894 (N_4894,N_4090,N_4453);
or U4895 (N_4895,N_4023,N_4246);
nand U4896 (N_4896,N_4434,N_4138);
nor U4897 (N_4897,N_4350,N_4101);
or U4898 (N_4898,N_4047,N_4371);
and U4899 (N_4899,N_4381,N_4029);
nand U4900 (N_4900,N_4307,N_4282);
nor U4901 (N_4901,N_4126,N_4476);
nand U4902 (N_4902,N_4450,N_4416);
or U4903 (N_4903,N_4013,N_4379);
or U4904 (N_4904,N_4122,N_4325);
nor U4905 (N_4905,N_4193,N_4045);
or U4906 (N_4906,N_4477,N_4494);
nand U4907 (N_4907,N_4465,N_4193);
nor U4908 (N_4908,N_4303,N_4205);
nand U4909 (N_4909,N_4244,N_4230);
and U4910 (N_4910,N_4044,N_4474);
or U4911 (N_4911,N_4058,N_4288);
and U4912 (N_4912,N_4305,N_4370);
nand U4913 (N_4913,N_4062,N_4019);
and U4914 (N_4914,N_4398,N_4019);
and U4915 (N_4915,N_4391,N_4407);
nand U4916 (N_4916,N_4065,N_4397);
or U4917 (N_4917,N_4356,N_4338);
or U4918 (N_4918,N_4384,N_4072);
or U4919 (N_4919,N_4073,N_4023);
nand U4920 (N_4920,N_4481,N_4022);
nor U4921 (N_4921,N_4377,N_4222);
nand U4922 (N_4922,N_4182,N_4053);
nor U4923 (N_4923,N_4413,N_4083);
nor U4924 (N_4924,N_4284,N_4150);
nor U4925 (N_4925,N_4356,N_4337);
or U4926 (N_4926,N_4161,N_4496);
nand U4927 (N_4927,N_4003,N_4126);
nand U4928 (N_4928,N_4183,N_4141);
or U4929 (N_4929,N_4401,N_4099);
and U4930 (N_4930,N_4424,N_4499);
or U4931 (N_4931,N_4092,N_4332);
and U4932 (N_4932,N_4339,N_4293);
and U4933 (N_4933,N_4057,N_4442);
or U4934 (N_4934,N_4271,N_4475);
nor U4935 (N_4935,N_4338,N_4209);
xnor U4936 (N_4936,N_4195,N_4352);
or U4937 (N_4937,N_4112,N_4038);
nand U4938 (N_4938,N_4437,N_4406);
nand U4939 (N_4939,N_4139,N_4044);
or U4940 (N_4940,N_4177,N_4435);
or U4941 (N_4941,N_4366,N_4099);
nand U4942 (N_4942,N_4243,N_4310);
nand U4943 (N_4943,N_4114,N_4183);
or U4944 (N_4944,N_4027,N_4148);
and U4945 (N_4945,N_4382,N_4227);
nand U4946 (N_4946,N_4477,N_4312);
and U4947 (N_4947,N_4345,N_4157);
and U4948 (N_4948,N_4377,N_4243);
and U4949 (N_4949,N_4010,N_4025);
or U4950 (N_4950,N_4361,N_4081);
nor U4951 (N_4951,N_4239,N_4166);
nand U4952 (N_4952,N_4044,N_4079);
and U4953 (N_4953,N_4291,N_4025);
nand U4954 (N_4954,N_4273,N_4296);
or U4955 (N_4955,N_4436,N_4017);
nand U4956 (N_4956,N_4402,N_4241);
and U4957 (N_4957,N_4468,N_4200);
nor U4958 (N_4958,N_4088,N_4432);
or U4959 (N_4959,N_4368,N_4080);
or U4960 (N_4960,N_4118,N_4101);
or U4961 (N_4961,N_4317,N_4479);
nand U4962 (N_4962,N_4374,N_4273);
and U4963 (N_4963,N_4351,N_4257);
and U4964 (N_4964,N_4445,N_4173);
nor U4965 (N_4965,N_4414,N_4116);
and U4966 (N_4966,N_4302,N_4349);
nand U4967 (N_4967,N_4380,N_4243);
nor U4968 (N_4968,N_4309,N_4091);
or U4969 (N_4969,N_4420,N_4158);
or U4970 (N_4970,N_4370,N_4166);
nor U4971 (N_4971,N_4058,N_4112);
or U4972 (N_4972,N_4151,N_4353);
nand U4973 (N_4973,N_4491,N_4242);
and U4974 (N_4974,N_4380,N_4245);
xor U4975 (N_4975,N_4489,N_4430);
nor U4976 (N_4976,N_4007,N_4329);
nand U4977 (N_4977,N_4244,N_4138);
nor U4978 (N_4978,N_4450,N_4268);
and U4979 (N_4979,N_4421,N_4407);
and U4980 (N_4980,N_4254,N_4000);
or U4981 (N_4981,N_4392,N_4193);
nor U4982 (N_4982,N_4140,N_4153);
and U4983 (N_4983,N_4071,N_4156);
xor U4984 (N_4984,N_4335,N_4134);
or U4985 (N_4985,N_4002,N_4198);
nor U4986 (N_4986,N_4319,N_4007);
nor U4987 (N_4987,N_4124,N_4257);
nor U4988 (N_4988,N_4229,N_4271);
and U4989 (N_4989,N_4452,N_4148);
nor U4990 (N_4990,N_4294,N_4067);
or U4991 (N_4991,N_4295,N_4184);
or U4992 (N_4992,N_4149,N_4069);
nand U4993 (N_4993,N_4477,N_4270);
nand U4994 (N_4994,N_4127,N_4216);
nor U4995 (N_4995,N_4290,N_4076);
or U4996 (N_4996,N_4318,N_4230);
nor U4997 (N_4997,N_4120,N_4260);
and U4998 (N_4998,N_4146,N_4351);
nor U4999 (N_4999,N_4247,N_4142);
nand UO_0 (O_0,N_4758,N_4775);
or UO_1 (O_1,N_4957,N_4589);
or UO_2 (O_2,N_4614,N_4608);
and UO_3 (O_3,N_4568,N_4726);
and UO_4 (O_4,N_4922,N_4962);
and UO_5 (O_5,N_4664,N_4871);
nor UO_6 (O_6,N_4631,N_4791);
and UO_7 (O_7,N_4733,N_4847);
and UO_8 (O_8,N_4833,N_4683);
nand UO_9 (O_9,N_4878,N_4852);
and UO_10 (O_10,N_4604,N_4518);
nor UO_11 (O_11,N_4893,N_4676);
nand UO_12 (O_12,N_4930,N_4636);
nand UO_13 (O_13,N_4709,N_4692);
nor UO_14 (O_14,N_4932,N_4701);
or UO_15 (O_15,N_4956,N_4517);
nand UO_16 (O_16,N_4832,N_4924);
nor UO_17 (O_17,N_4675,N_4590);
or UO_18 (O_18,N_4891,N_4712);
or UO_19 (O_19,N_4974,N_4600);
nor UO_20 (O_20,N_4646,N_4633);
or UO_21 (O_21,N_4575,N_4637);
or UO_22 (O_22,N_4684,N_4897);
nor UO_23 (O_23,N_4621,N_4576);
nand UO_24 (O_24,N_4917,N_4711);
and UO_25 (O_25,N_4630,N_4725);
and UO_26 (O_26,N_4612,N_4772);
and UO_27 (O_27,N_4764,N_4741);
and UO_28 (O_28,N_4818,N_4784);
nand UO_29 (O_29,N_4815,N_4506);
and UO_30 (O_30,N_4642,N_4699);
and UO_31 (O_31,N_4953,N_4541);
xnor UO_32 (O_32,N_4990,N_4863);
or UO_33 (O_33,N_4842,N_4682);
and UO_34 (O_34,N_4916,N_4877);
and UO_35 (O_35,N_4592,N_4926);
nor UO_36 (O_36,N_4804,N_4703);
nand UO_37 (O_37,N_4963,N_4942);
and UO_38 (O_38,N_4727,N_4899);
nand UO_39 (O_39,N_4948,N_4523);
nand UO_40 (O_40,N_4807,N_4543);
or UO_41 (O_41,N_4659,N_4826);
or UO_42 (O_42,N_4892,N_4918);
nand UO_43 (O_43,N_4846,N_4509);
or UO_44 (O_44,N_4937,N_4736);
nand UO_45 (O_45,N_4879,N_4801);
or UO_46 (O_46,N_4943,N_4858);
or UO_47 (O_47,N_4613,N_4786);
and UO_48 (O_48,N_4882,N_4945);
nand UO_49 (O_49,N_4581,N_4966);
nand UO_50 (O_50,N_4588,N_4776);
or UO_51 (O_51,N_4869,N_4849);
nor UO_52 (O_52,N_4503,N_4629);
nor UO_53 (O_53,N_4920,N_4783);
and UO_54 (O_54,N_4622,N_4765);
nor UO_55 (O_55,N_4895,N_4610);
nand UO_56 (O_56,N_4658,N_4552);
and UO_57 (O_57,N_4743,N_4762);
or UO_58 (O_58,N_4752,N_4912);
or UO_59 (O_59,N_4502,N_4605);
or UO_60 (O_60,N_4619,N_4571);
and UO_61 (O_61,N_4710,N_4505);
or UO_62 (O_62,N_4848,N_4521);
or UO_63 (O_63,N_4933,N_4719);
nor UO_64 (O_64,N_4947,N_4623);
and UO_65 (O_65,N_4949,N_4841);
nand UO_66 (O_66,N_4714,N_4691);
and UO_67 (O_67,N_4678,N_4745);
and UO_68 (O_68,N_4594,N_4889);
or UO_69 (O_69,N_4564,N_4782);
or UO_70 (O_70,N_4720,N_4977);
nand UO_71 (O_71,N_4830,N_4793);
or UO_72 (O_72,N_4821,N_4811);
and UO_73 (O_73,N_4563,N_4779);
nor UO_74 (O_74,N_4655,N_4910);
nor UO_75 (O_75,N_4855,N_4615);
nor UO_76 (O_76,N_4991,N_4611);
xnor UO_77 (O_77,N_4542,N_4734);
nand UO_78 (O_78,N_4931,N_4839);
nor UO_79 (O_79,N_4723,N_4970);
nor UO_80 (O_80,N_4810,N_4875);
or UO_81 (O_81,N_4582,N_4585);
nor UO_82 (O_82,N_4984,N_4843);
nand UO_83 (O_83,N_4569,N_4750);
nor UO_84 (O_84,N_4609,N_4511);
nand UO_85 (O_85,N_4532,N_4562);
and UO_86 (O_86,N_4934,N_4737);
or UO_87 (O_87,N_4925,N_4755);
or UO_88 (O_88,N_4827,N_4886);
or UO_89 (O_89,N_4713,N_4697);
nor UO_90 (O_90,N_4995,N_4809);
and UO_91 (O_91,N_4574,N_4763);
and UO_92 (O_92,N_4620,N_4975);
nor UO_93 (O_93,N_4547,N_4767);
and UO_94 (O_94,N_4994,N_4759);
nor UO_95 (O_95,N_4520,N_4513);
or UO_96 (O_96,N_4923,N_4700);
nor UO_97 (O_97,N_4584,N_4829);
or UO_98 (O_98,N_4580,N_4989);
nor UO_99 (O_99,N_4950,N_4958);
or UO_100 (O_100,N_4721,N_4982);
nand UO_101 (O_101,N_4778,N_4706);
xor UO_102 (O_102,N_4607,N_4535);
nand UO_103 (O_103,N_4573,N_4677);
and UO_104 (O_104,N_4732,N_4694);
and UO_105 (O_105,N_4602,N_4824);
nor UO_106 (O_106,N_4883,N_4644);
nor UO_107 (O_107,N_4972,N_4819);
nor UO_108 (O_108,N_4896,N_4785);
nand UO_109 (O_109,N_4729,N_4979);
nor UO_110 (O_110,N_4999,N_4674);
or UO_111 (O_111,N_4617,N_4561);
nand UO_112 (O_112,N_4835,N_4595);
or UO_113 (O_113,N_4696,N_4993);
nand UO_114 (O_114,N_4632,N_4992);
and UO_115 (O_115,N_4671,N_4907);
and UO_116 (O_116,N_4728,N_4567);
and UO_117 (O_117,N_4967,N_4649);
nand UO_118 (O_118,N_4501,N_4794);
or UO_119 (O_119,N_4867,N_4688);
or UO_120 (O_120,N_4770,N_4544);
nand UO_121 (O_121,N_4546,N_4690);
nand UO_122 (O_122,N_4519,N_4971);
nand UO_123 (O_123,N_4853,N_4527);
and UO_124 (O_124,N_4928,N_4689);
nor UO_125 (O_125,N_4670,N_4667);
and UO_126 (O_126,N_4890,N_4618);
nor UO_127 (O_127,N_4760,N_4707);
nand UO_128 (O_128,N_4634,N_4591);
and UO_129 (O_129,N_4586,N_4840);
and UO_130 (O_130,N_4822,N_4996);
nor UO_131 (O_131,N_4978,N_4868);
nand UO_132 (O_132,N_4781,N_4663);
nor UO_133 (O_133,N_4774,N_4800);
nand UO_134 (O_134,N_4651,N_4808);
nor UO_135 (O_135,N_4685,N_4795);
xor UO_136 (O_136,N_4654,N_4645);
or UO_137 (O_137,N_4647,N_4856);
and UO_138 (O_138,N_4681,N_4859);
nor UO_139 (O_139,N_4968,N_4944);
nand UO_140 (O_140,N_4998,N_4964);
or UO_141 (O_141,N_4599,N_4587);
nand UO_142 (O_142,N_4872,N_4554);
and UO_143 (O_143,N_4813,N_4919);
or UO_144 (O_144,N_4805,N_4799);
nand UO_145 (O_145,N_4559,N_4731);
and UO_146 (O_146,N_4935,N_4792);
and UO_147 (O_147,N_4884,N_4742);
and UO_148 (O_148,N_4533,N_4909);
nor UO_149 (O_149,N_4788,N_4988);
or UO_150 (O_150,N_4865,N_4744);
and UO_151 (O_151,N_4524,N_4549);
nor UO_152 (O_152,N_4722,N_4525);
or UO_153 (O_153,N_4625,N_4851);
and UO_154 (O_154,N_4951,N_4536);
nand UO_155 (O_155,N_4624,N_4616);
and UO_156 (O_156,N_4716,N_4735);
or UO_157 (O_157,N_4705,N_4961);
or UO_158 (O_158,N_4556,N_4898);
nand UO_159 (O_159,N_4954,N_4665);
nand UO_160 (O_160,N_4927,N_4940);
and UO_161 (O_161,N_4880,N_4768);
and UO_162 (O_162,N_4717,N_4673);
xnor UO_163 (O_163,N_4531,N_4550);
and UO_164 (O_164,N_4548,N_4553);
nor UO_165 (O_165,N_4740,N_4515);
nor UO_166 (O_166,N_4572,N_4746);
nand UO_167 (O_167,N_4672,N_4959);
nand UO_168 (O_168,N_4828,N_4825);
or UO_169 (O_169,N_4946,N_4797);
or UO_170 (O_170,N_4981,N_4844);
or UO_171 (O_171,N_4769,N_4601);
nand UO_172 (O_172,N_4680,N_4638);
and UO_173 (O_173,N_4530,N_4551);
and UO_174 (O_174,N_4904,N_4598);
and UO_175 (O_175,N_4606,N_4874);
nand UO_176 (O_176,N_4695,N_4570);
nor UO_177 (O_177,N_4628,N_4860);
nor UO_178 (O_178,N_4929,N_4789);
nor UO_179 (O_179,N_4915,N_4780);
and UO_180 (O_180,N_4900,N_4526);
and UO_181 (O_181,N_4724,N_4597);
nor UO_182 (O_182,N_4749,N_4715);
and UO_183 (O_183,N_4508,N_4540);
nor UO_184 (O_184,N_4718,N_4593);
or UO_185 (O_185,N_4558,N_4565);
and UO_186 (O_186,N_4790,N_4529);
nand UO_187 (O_187,N_4911,N_4662);
nor UO_188 (O_188,N_4965,N_4698);
and UO_189 (O_189,N_4987,N_4823);
nor UO_190 (O_190,N_4850,N_4578);
nand UO_191 (O_191,N_4534,N_4861);
and UO_192 (O_192,N_4973,N_4639);
and UO_193 (O_193,N_4881,N_4908);
nor UO_194 (O_194,N_4902,N_4803);
nor UO_195 (O_195,N_4938,N_4960);
nand UO_196 (O_196,N_4652,N_4997);
or UO_197 (O_197,N_4748,N_4538);
nor UO_198 (O_198,N_4596,N_4901);
and UO_199 (O_199,N_4816,N_4812);
or UO_200 (O_200,N_4560,N_4862);
and UO_201 (O_201,N_4686,N_4983);
or UO_202 (O_202,N_4834,N_4514);
and UO_203 (O_203,N_4522,N_4566);
nand UO_204 (O_204,N_4857,N_4820);
nor UO_205 (O_205,N_4873,N_4814);
or UO_206 (O_206,N_4603,N_4738);
and UO_207 (O_207,N_4888,N_4753);
nor UO_208 (O_208,N_4507,N_4666);
nor UO_209 (O_209,N_4693,N_4854);
or UO_210 (O_210,N_4802,N_4583);
or UO_211 (O_211,N_4756,N_4657);
or UO_212 (O_212,N_4838,N_4739);
nor UO_213 (O_213,N_4866,N_4730);
and UO_214 (O_214,N_4504,N_4656);
nor UO_215 (O_215,N_4969,N_4687);
and UO_216 (O_216,N_4955,N_4557);
nand UO_217 (O_217,N_4641,N_4773);
or UO_218 (O_218,N_4577,N_4914);
nor UO_219 (O_219,N_4512,N_4650);
nand UO_220 (O_220,N_4761,N_4661);
or UO_221 (O_221,N_4806,N_4668);
or UO_222 (O_222,N_4985,N_4905);
nor UO_223 (O_223,N_4941,N_4913);
nor UO_224 (O_224,N_4980,N_4704);
nor UO_225 (O_225,N_4648,N_4796);
and UO_226 (O_226,N_4708,N_4747);
nand UO_227 (O_227,N_4643,N_4653);
and UO_228 (O_228,N_4555,N_4751);
or UO_229 (O_229,N_4921,N_4635);
and UO_230 (O_230,N_4660,N_4798);
and UO_231 (O_231,N_4836,N_4887);
or UO_232 (O_232,N_4702,N_4876);
nand UO_233 (O_233,N_4864,N_4885);
nand UO_234 (O_234,N_4952,N_4754);
and UO_235 (O_235,N_4787,N_4837);
and UO_236 (O_236,N_4936,N_4626);
and UO_237 (O_237,N_4777,N_4757);
and UO_238 (O_238,N_4528,N_4545);
nand UO_239 (O_239,N_4817,N_4831);
and UO_240 (O_240,N_4640,N_4679);
and UO_241 (O_241,N_4669,N_4500);
nand UO_242 (O_242,N_4906,N_4510);
nand UO_243 (O_243,N_4579,N_4845);
or UO_244 (O_244,N_4539,N_4766);
and UO_245 (O_245,N_4976,N_4986);
and UO_246 (O_246,N_4903,N_4537);
nor UO_247 (O_247,N_4870,N_4771);
or UO_248 (O_248,N_4939,N_4894);
nor UO_249 (O_249,N_4627,N_4516);
nand UO_250 (O_250,N_4988,N_4926);
nand UO_251 (O_251,N_4698,N_4973);
nor UO_252 (O_252,N_4997,N_4728);
and UO_253 (O_253,N_4740,N_4654);
nor UO_254 (O_254,N_4938,N_4889);
nor UO_255 (O_255,N_4653,N_4829);
or UO_256 (O_256,N_4684,N_4889);
and UO_257 (O_257,N_4711,N_4595);
and UO_258 (O_258,N_4544,N_4615);
nand UO_259 (O_259,N_4600,N_4821);
and UO_260 (O_260,N_4690,N_4683);
and UO_261 (O_261,N_4994,N_4855);
nand UO_262 (O_262,N_4858,N_4807);
xor UO_263 (O_263,N_4946,N_4890);
nor UO_264 (O_264,N_4717,N_4898);
nor UO_265 (O_265,N_4600,N_4760);
nand UO_266 (O_266,N_4627,N_4595);
and UO_267 (O_267,N_4956,N_4604);
or UO_268 (O_268,N_4810,N_4757);
or UO_269 (O_269,N_4903,N_4646);
nor UO_270 (O_270,N_4691,N_4787);
nor UO_271 (O_271,N_4807,N_4540);
and UO_272 (O_272,N_4993,N_4641);
and UO_273 (O_273,N_4841,N_4765);
or UO_274 (O_274,N_4695,N_4937);
and UO_275 (O_275,N_4828,N_4685);
nand UO_276 (O_276,N_4987,N_4641);
nand UO_277 (O_277,N_4526,N_4596);
nand UO_278 (O_278,N_4604,N_4905);
or UO_279 (O_279,N_4681,N_4843);
nand UO_280 (O_280,N_4894,N_4681);
or UO_281 (O_281,N_4698,N_4744);
or UO_282 (O_282,N_4708,N_4523);
nor UO_283 (O_283,N_4866,N_4916);
or UO_284 (O_284,N_4518,N_4540);
or UO_285 (O_285,N_4759,N_4675);
nor UO_286 (O_286,N_4554,N_4911);
or UO_287 (O_287,N_4578,N_4910);
nor UO_288 (O_288,N_4962,N_4864);
or UO_289 (O_289,N_4593,N_4972);
or UO_290 (O_290,N_4638,N_4751);
nand UO_291 (O_291,N_4683,N_4737);
or UO_292 (O_292,N_4911,N_4634);
nor UO_293 (O_293,N_4697,N_4958);
and UO_294 (O_294,N_4810,N_4600);
or UO_295 (O_295,N_4716,N_4912);
nand UO_296 (O_296,N_4707,N_4527);
nand UO_297 (O_297,N_4801,N_4828);
and UO_298 (O_298,N_4550,N_4794);
or UO_299 (O_299,N_4872,N_4580);
or UO_300 (O_300,N_4636,N_4745);
nor UO_301 (O_301,N_4708,N_4587);
nor UO_302 (O_302,N_4987,N_4707);
or UO_303 (O_303,N_4910,N_4904);
or UO_304 (O_304,N_4604,N_4503);
and UO_305 (O_305,N_4530,N_4620);
and UO_306 (O_306,N_4608,N_4825);
nor UO_307 (O_307,N_4829,N_4924);
or UO_308 (O_308,N_4925,N_4895);
and UO_309 (O_309,N_4870,N_4605);
nand UO_310 (O_310,N_4963,N_4820);
nand UO_311 (O_311,N_4796,N_4587);
or UO_312 (O_312,N_4793,N_4621);
or UO_313 (O_313,N_4732,N_4756);
nor UO_314 (O_314,N_4514,N_4939);
nand UO_315 (O_315,N_4838,N_4512);
and UO_316 (O_316,N_4919,N_4615);
nor UO_317 (O_317,N_4981,N_4851);
or UO_318 (O_318,N_4694,N_4654);
or UO_319 (O_319,N_4953,N_4632);
or UO_320 (O_320,N_4845,N_4659);
nand UO_321 (O_321,N_4859,N_4961);
nor UO_322 (O_322,N_4575,N_4926);
or UO_323 (O_323,N_4706,N_4886);
and UO_324 (O_324,N_4811,N_4503);
or UO_325 (O_325,N_4528,N_4741);
nor UO_326 (O_326,N_4538,N_4801);
or UO_327 (O_327,N_4841,N_4897);
or UO_328 (O_328,N_4605,N_4597);
or UO_329 (O_329,N_4561,N_4835);
nor UO_330 (O_330,N_4977,N_4708);
or UO_331 (O_331,N_4732,N_4959);
or UO_332 (O_332,N_4632,N_4857);
and UO_333 (O_333,N_4644,N_4768);
nor UO_334 (O_334,N_4771,N_4837);
nand UO_335 (O_335,N_4720,N_4995);
nor UO_336 (O_336,N_4636,N_4801);
and UO_337 (O_337,N_4879,N_4845);
and UO_338 (O_338,N_4845,N_4785);
and UO_339 (O_339,N_4829,N_4686);
nor UO_340 (O_340,N_4883,N_4571);
and UO_341 (O_341,N_4599,N_4831);
or UO_342 (O_342,N_4851,N_4783);
or UO_343 (O_343,N_4871,N_4941);
nor UO_344 (O_344,N_4917,N_4834);
or UO_345 (O_345,N_4624,N_4963);
or UO_346 (O_346,N_4842,N_4658);
and UO_347 (O_347,N_4549,N_4722);
nor UO_348 (O_348,N_4796,N_4631);
nand UO_349 (O_349,N_4549,N_4991);
nor UO_350 (O_350,N_4731,N_4860);
nor UO_351 (O_351,N_4908,N_4663);
nand UO_352 (O_352,N_4612,N_4633);
and UO_353 (O_353,N_4849,N_4889);
and UO_354 (O_354,N_4952,N_4672);
nand UO_355 (O_355,N_4676,N_4826);
nor UO_356 (O_356,N_4798,N_4871);
nand UO_357 (O_357,N_4597,N_4643);
nand UO_358 (O_358,N_4520,N_4510);
nand UO_359 (O_359,N_4563,N_4785);
and UO_360 (O_360,N_4756,N_4700);
nor UO_361 (O_361,N_4728,N_4935);
and UO_362 (O_362,N_4927,N_4787);
nor UO_363 (O_363,N_4810,N_4573);
or UO_364 (O_364,N_4697,N_4720);
nand UO_365 (O_365,N_4743,N_4866);
nand UO_366 (O_366,N_4759,N_4579);
or UO_367 (O_367,N_4915,N_4818);
or UO_368 (O_368,N_4609,N_4580);
nor UO_369 (O_369,N_4780,N_4937);
nor UO_370 (O_370,N_4786,N_4647);
nand UO_371 (O_371,N_4786,N_4558);
xor UO_372 (O_372,N_4633,N_4562);
and UO_373 (O_373,N_4726,N_4880);
nand UO_374 (O_374,N_4991,N_4536);
and UO_375 (O_375,N_4862,N_4882);
nor UO_376 (O_376,N_4529,N_4910);
nor UO_377 (O_377,N_4685,N_4990);
nand UO_378 (O_378,N_4527,N_4812);
and UO_379 (O_379,N_4714,N_4620);
or UO_380 (O_380,N_4742,N_4619);
or UO_381 (O_381,N_4893,N_4652);
or UO_382 (O_382,N_4527,N_4802);
nand UO_383 (O_383,N_4686,N_4680);
nor UO_384 (O_384,N_4834,N_4692);
nor UO_385 (O_385,N_4846,N_4969);
or UO_386 (O_386,N_4580,N_4765);
nand UO_387 (O_387,N_4886,N_4686);
and UO_388 (O_388,N_4678,N_4840);
and UO_389 (O_389,N_4794,N_4739);
nand UO_390 (O_390,N_4651,N_4938);
and UO_391 (O_391,N_4871,N_4953);
nand UO_392 (O_392,N_4516,N_4643);
nand UO_393 (O_393,N_4668,N_4872);
or UO_394 (O_394,N_4796,N_4857);
or UO_395 (O_395,N_4921,N_4920);
xnor UO_396 (O_396,N_4672,N_4868);
nor UO_397 (O_397,N_4524,N_4669);
xor UO_398 (O_398,N_4608,N_4828);
nor UO_399 (O_399,N_4799,N_4858);
nand UO_400 (O_400,N_4929,N_4716);
and UO_401 (O_401,N_4919,N_4890);
and UO_402 (O_402,N_4803,N_4506);
or UO_403 (O_403,N_4702,N_4766);
nor UO_404 (O_404,N_4800,N_4784);
nor UO_405 (O_405,N_4796,N_4839);
nor UO_406 (O_406,N_4709,N_4779);
nand UO_407 (O_407,N_4588,N_4882);
or UO_408 (O_408,N_4598,N_4591);
or UO_409 (O_409,N_4918,N_4543);
and UO_410 (O_410,N_4914,N_4837);
nor UO_411 (O_411,N_4988,N_4846);
or UO_412 (O_412,N_4563,N_4736);
nand UO_413 (O_413,N_4663,N_4605);
nand UO_414 (O_414,N_4841,N_4598);
xor UO_415 (O_415,N_4930,N_4656);
nor UO_416 (O_416,N_4615,N_4508);
and UO_417 (O_417,N_4525,N_4779);
nor UO_418 (O_418,N_4990,N_4744);
or UO_419 (O_419,N_4802,N_4741);
and UO_420 (O_420,N_4684,N_4765);
and UO_421 (O_421,N_4529,N_4501);
and UO_422 (O_422,N_4772,N_4608);
nand UO_423 (O_423,N_4611,N_4824);
and UO_424 (O_424,N_4779,N_4708);
or UO_425 (O_425,N_4741,N_4567);
or UO_426 (O_426,N_4719,N_4679);
and UO_427 (O_427,N_4686,N_4959);
and UO_428 (O_428,N_4710,N_4646);
nand UO_429 (O_429,N_4756,N_4508);
or UO_430 (O_430,N_4894,N_4600);
and UO_431 (O_431,N_4788,N_4941);
nand UO_432 (O_432,N_4636,N_4915);
and UO_433 (O_433,N_4559,N_4947);
or UO_434 (O_434,N_4804,N_4706);
nand UO_435 (O_435,N_4787,N_4676);
nand UO_436 (O_436,N_4927,N_4993);
or UO_437 (O_437,N_4785,N_4739);
or UO_438 (O_438,N_4657,N_4622);
nand UO_439 (O_439,N_4731,N_4510);
and UO_440 (O_440,N_4789,N_4676);
or UO_441 (O_441,N_4957,N_4826);
and UO_442 (O_442,N_4746,N_4713);
nand UO_443 (O_443,N_4549,N_4810);
xor UO_444 (O_444,N_4843,N_4551);
and UO_445 (O_445,N_4975,N_4783);
nor UO_446 (O_446,N_4596,N_4585);
or UO_447 (O_447,N_4813,N_4518);
and UO_448 (O_448,N_4607,N_4889);
or UO_449 (O_449,N_4879,N_4728);
nor UO_450 (O_450,N_4618,N_4846);
nand UO_451 (O_451,N_4925,N_4913);
xor UO_452 (O_452,N_4539,N_4815);
nor UO_453 (O_453,N_4825,N_4650);
and UO_454 (O_454,N_4701,N_4559);
nand UO_455 (O_455,N_4581,N_4533);
or UO_456 (O_456,N_4764,N_4605);
or UO_457 (O_457,N_4602,N_4621);
or UO_458 (O_458,N_4816,N_4653);
nor UO_459 (O_459,N_4626,N_4550);
and UO_460 (O_460,N_4768,N_4885);
and UO_461 (O_461,N_4980,N_4601);
and UO_462 (O_462,N_4760,N_4765);
nand UO_463 (O_463,N_4966,N_4904);
and UO_464 (O_464,N_4830,N_4930);
or UO_465 (O_465,N_4946,N_4748);
nor UO_466 (O_466,N_4825,N_4973);
or UO_467 (O_467,N_4648,N_4512);
and UO_468 (O_468,N_4807,N_4873);
nor UO_469 (O_469,N_4808,N_4954);
nor UO_470 (O_470,N_4782,N_4736);
or UO_471 (O_471,N_4990,N_4575);
or UO_472 (O_472,N_4680,N_4747);
and UO_473 (O_473,N_4994,N_4996);
nor UO_474 (O_474,N_4571,N_4961);
and UO_475 (O_475,N_4839,N_4756);
nor UO_476 (O_476,N_4647,N_4730);
nor UO_477 (O_477,N_4981,N_4801);
or UO_478 (O_478,N_4520,N_4688);
and UO_479 (O_479,N_4925,N_4964);
or UO_480 (O_480,N_4965,N_4685);
or UO_481 (O_481,N_4766,N_4528);
and UO_482 (O_482,N_4842,N_4832);
nor UO_483 (O_483,N_4501,N_4911);
nand UO_484 (O_484,N_4501,N_4759);
nand UO_485 (O_485,N_4565,N_4909);
or UO_486 (O_486,N_4546,N_4556);
or UO_487 (O_487,N_4638,N_4587);
nand UO_488 (O_488,N_4588,N_4539);
nand UO_489 (O_489,N_4922,N_4739);
and UO_490 (O_490,N_4881,N_4582);
nor UO_491 (O_491,N_4581,N_4810);
nand UO_492 (O_492,N_4775,N_4807);
or UO_493 (O_493,N_4877,N_4989);
or UO_494 (O_494,N_4945,N_4781);
nand UO_495 (O_495,N_4945,N_4584);
and UO_496 (O_496,N_4942,N_4924);
and UO_497 (O_497,N_4786,N_4664);
or UO_498 (O_498,N_4962,N_4941);
nand UO_499 (O_499,N_4627,N_4809);
nor UO_500 (O_500,N_4790,N_4598);
nor UO_501 (O_501,N_4564,N_4681);
nand UO_502 (O_502,N_4985,N_4558);
nor UO_503 (O_503,N_4844,N_4597);
and UO_504 (O_504,N_4550,N_4763);
and UO_505 (O_505,N_4780,N_4614);
or UO_506 (O_506,N_4577,N_4849);
nor UO_507 (O_507,N_4701,N_4876);
or UO_508 (O_508,N_4647,N_4741);
or UO_509 (O_509,N_4559,N_4885);
and UO_510 (O_510,N_4683,N_4579);
or UO_511 (O_511,N_4943,N_4882);
or UO_512 (O_512,N_4714,N_4663);
or UO_513 (O_513,N_4788,N_4607);
or UO_514 (O_514,N_4800,N_4791);
nor UO_515 (O_515,N_4989,N_4503);
and UO_516 (O_516,N_4864,N_4944);
and UO_517 (O_517,N_4735,N_4702);
or UO_518 (O_518,N_4980,N_4940);
and UO_519 (O_519,N_4667,N_4730);
nand UO_520 (O_520,N_4681,N_4546);
and UO_521 (O_521,N_4869,N_4880);
or UO_522 (O_522,N_4937,N_4587);
or UO_523 (O_523,N_4915,N_4813);
nor UO_524 (O_524,N_4573,N_4642);
and UO_525 (O_525,N_4814,N_4582);
nor UO_526 (O_526,N_4819,N_4722);
and UO_527 (O_527,N_4524,N_4818);
nand UO_528 (O_528,N_4541,N_4753);
or UO_529 (O_529,N_4900,N_4788);
and UO_530 (O_530,N_4835,N_4768);
or UO_531 (O_531,N_4998,N_4911);
or UO_532 (O_532,N_4753,N_4611);
nand UO_533 (O_533,N_4717,N_4986);
nand UO_534 (O_534,N_4868,N_4603);
or UO_535 (O_535,N_4655,N_4783);
and UO_536 (O_536,N_4517,N_4653);
nor UO_537 (O_537,N_4727,N_4900);
nand UO_538 (O_538,N_4552,N_4547);
nor UO_539 (O_539,N_4702,N_4906);
and UO_540 (O_540,N_4944,N_4946);
and UO_541 (O_541,N_4944,N_4994);
and UO_542 (O_542,N_4903,N_4971);
and UO_543 (O_543,N_4741,N_4525);
nand UO_544 (O_544,N_4520,N_4807);
nand UO_545 (O_545,N_4598,N_4619);
or UO_546 (O_546,N_4745,N_4808);
nand UO_547 (O_547,N_4827,N_4615);
or UO_548 (O_548,N_4659,N_4829);
and UO_549 (O_549,N_4746,N_4966);
and UO_550 (O_550,N_4731,N_4880);
nand UO_551 (O_551,N_4898,N_4950);
and UO_552 (O_552,N_4787,N_4553);
or UO_553 (O_553,N_4649,N_4858);
nand UO_554 (O_554,N_4988,N_4796);
nand UO_555 (O_555,N_4766,N_4656);
nand UO_556 (O_556,N_4902,N_4598);
nand UO_557 (O_557,N_4967,N_4972);
nand UO_558 (O_558,N_4996,N_4719);
or UO_559 (O_559,N_4516,N_4991);
nor UO_560 (O_560,N_4694,N_4995);
nor UO_561 (O_561,N_4746,N_4820);
or UO_562 (O_562,N_4533,N_4704);
or UO_563 (O_563,N_4637,N_4570);
or UO_564 (O_564,N_4637,N_4980);
nor UO_565 (O_565,N_4703,N_4743);
or UO_566 (O_566,N_4640,N_4746);
nor UO_567 (O_567,N_4588,N_4647);
or UO_568 (O_568,N_4836,N_4924);
or UO_569 (O_569,N_4772,N_4963);
nor UO_570 (O_570,N_4927,N_4629);
and UO_571 (O_571,N_4693,N_4731);
nand UO_572 (O_572,N_4710,N_4838);
and UO_573 (O_573,N_4674,N_4502);
xor UO_574 (O_574,N_4582,N_4891);
or UO_575 (O_575,N_4551,N_4677);
or UO_576 (O_576,N_4635,N_4848);
nand UO_577 (O_577,N_4833,N_4936);
or UO_578 (O_578,N_4954,N_4983);
and UO_579 (O_579,N_4968,N_4871);
and UO_580 (O_580,N_4976,N_4624);
nor UO_581 (O_581,N_4874,N_4615);
or UO_582 (O_582,N_4660,N_4572);
or UO_583 (O_583,N_4511,N_4846);
and UO_584 (O_584,N_4773,N_4531);
nand UO_585 (O_585,N_4955,N_4576);
nor UO_586 (O_586,N_4826,N_4836);
nand UO_587 (O_587,N_4776,N_4909);
nor UO_588 (O_588,N_4586,N_4639);
or UO_589 (O_589,N_4842,N_4867);
or UO_590 (O_590,N_4696,N_4880);
nor UO_591 (O_591,N_4912,N_4684);
nand UO_592 (O_592,N_4928,N_4936);
nor UO_593 (O_593,N_4935,N_4921);
or UO_594 (O_594,N_4731,N_4610);
nand UO_595 (O_595,N_4716,N_4944);
or UO_596 (O_596,N_4786,N_4936);
or UO_597 (O_597,N_4605,N_4692);
and UO_598 (O_598,N_4625,N_4534);
or UO_599 (O_599,N_4586,N_4978);
nand UO_600 (O_600,N_4583,N_4646);
nor UO_601 (O_601,N_4505,N_4789);
nand UO_602 (O_602,N_4999,N_4509);
and UO_603 (O_603,N_4965,N_4565);
or UO_604 (O_604,N_4984,N_4570);
nor UO_605 (O_605,N_4735,N_4936);
nand UO_606 (O_606,N_4881,N_4853);
nor UO_607 (O_607,N_4712,N_4874);
and UO_608 (O_608,N_4984,N_4715);
nor UO_609 (O_609,N_4614,N_4635);
nand UO_610 (O_610,N_4588,N_4517);
or UO_611 (O_611,N_4733,N_4589);
or UO_612 (O_612,N_4648,N_4556);
nand UO_613 (O_613,N_4877,N_4869);
nand UO_614 (O_614,N_4663,N_4589);
and UO_615 (O_615,N_4695,N_4913);
nand UO_616 (O_616,N_4689,N_4797);
xnor UO_617 (O_617,N_4767,N_4623);
and UO_618 (O_618,N_4751,N_4643);
nand UO_619 (O_619,N_4899,N_4974);
nor UO_620 (O_620,N_4805,N_4901);
and UO_621 (O_621,N_4779,N_4906);
or UO_622 (O_622,N_4982,N_4514);
and UO_623 (O_623,N_4657,N_4524);
and UO_624 (O_624,N_4616,N_4695);
and UO_625 (O_625,N_4700,N_4759);
nor UO_626 (O_626,N_4556,N_4863);
nor UO_627 (O_627,N_4934,N_4989);
or UO_628 (O_628,N_4655,N_4826);
and UO_629 (O_629,N_4997,N_4604);
nand UO_630 (O_630,N_4890,N_4637);
nand UO_631 (O_631,N_4697,N_4756);
nand UO_632 (O_632,N_4988,N_4559);
nor UO_633 (O_633,N_4612,N_4939);
nor UO_634 (O_634,N_4663,N_4961);
and UO_635 (O_635,N_4840,N_4519);
xor UO_636 (O_636,N_4939,N_4975);
nor UO_637 (O_637,N_4825,N_4679);
and UO_638 (O_638,N_4935,N_4780);
nand UO_639 (O_639,N_4820,N_4797);
nor UO_640 (O_640,N_4609,N_4577);
nor UO_641 (O_641,N_4805,N_4975);
and UO_642 (O_642,N_4877,N_4711);
nand UO_643 (O_643,N_4746,N_4885);
nor UO_644 (O_644,N_4806,N_4938);
nor UO_645 (O_645,N_4986,N_4752);
nor UO_646 (O_646,N_4747,N_4868);
or UO_647 (O_647,N_4980,N_4795);
nand UO_648 (O_648,N_4974,N_4681);
or UO_649 (O_649,N_4515,N_4621);
and UO_650 (O_650,N_4667,N_4543);
and UO_651 (O_651,N_4973,N_4779);
or UO_652 (O_652,N_4854,N_4862);
nand UO_653 (O_653,N_4586,N_4656);
and UO_654 (O_654,N_4765,N_4766);
or UO_655 (O_655,N_4842,N_4763);
nand UO_656 (O_656,N_4616,N_4666);
nand UO_657 (O_657,N_4681,N_4517);
nand UO_658 (O_658,N_4905,N_4867);
nor UO_659 (O_659,N_4667,N_4958);
nor UO_660 (O_660,N_4813,N_4651);
or UO_661 (O_661,N_4751,N_4639);
nand UO_662 (O_662,N_4714,N_4677);
or UO_663 (O_663,N_4802,N_4564);
nor UO_664 (O_664,N_4835,N_4765);
and UO_665 (O_665,N_4680,N_4961);
nor UO_666 (O_666,N_4688,N_4709);
xor UO_667 (O_667,N_4847,N_4854);
nor UO_668 (O_668,N_4633,N_4863);
nand UO_669 (O_669,N_4621,N_4859);
or UO_670 (O_670,N_4702,N_4858);
and UO_671 (O_671,N_4786,N_4988);
and UO_672 (O_672,N_4684,N_4995);
and UO_673 (O_673,N_4670,N_4599);
nand UO_674 (O_674,N_4752,N_4697);
or UO_675 (O_675,N_4828,N_4964);
nand UO_676 (O_676,N_4811,N_4603);
nor UO_677 (O_677,N_4667,N_4868);
or UO_678 (O_678,N_4566,N_4821);
or UO_679 (O_679,N_4576,N_4900);
or UO_680 (O_680,N_4877,N_4746);
and UO_681 (O_681,N_4946,N_4651);
nand UO_682 (O_682,N_4511,N_4861);
and UO_683 (O_683,N_4696,N_4910);
nor UO_684 (O_684,N_4985,N_4766);
and UO_685 (O_685,N_4939,N_4794);
and UO_686 (O_686,N_4698,N_4651);
nand UO_687 (O_687,N_4867,N_4793);
and UO_688 (O_688,N_4865,N_4604);
or UO_689 (O_689,N_4683,N_4717);
or UO_690 (O_690,N_4711,N_4882);
nor UO_691 (O_691,N_4962,N_4942);
nor UO_692 (O_692,N_4940,N_4965);
nand UO_693 (O_693,N_4900,N_4684);
and UO_694 (O_694,N_4580,N_4583);
and UO_695 (O_695,N_4573,N_4862);
nor UO_696 (O_696,N_4505,N_4788);
nor UO_697 (O_697,N_4514,N_4656);
or UO_698 (O_698,N_4600,N_4970);
and UO_699 (O_699,N_4814,N_4935);
nand UO_700 (O_700,N_4724,N_4951);
or UO_701 (O_701,N_4777,N_4743);
nand UO_702 (O_702,N_4567,N_4866);
and UO_703 (O_703,N_4678,N_4650);
and UO_704 (O_704,N_4535,N_4649);
xor UO_705 (O_705,N_4748,N_4627);
nor UO_706 (O_706,N_4867,N_4808);
nor UO_707 (O_707,N_4655,N_4597);
nand UO_708 (O_708,N_4772,N_4878);
or UO_709 (O_709,N_4935,N_4630);
or UO_710 (O_710,N_4513,N_4887);
nor UO_711 (O_711,N_4584,N_4515);
or UO_712 (O_712,N_4918,N_4504);
nor UO_713 (O_713,N_4557,N_4969);
and UO_714 (O_714,N_4938,N_4644);
nor UO_715 (O_715,N_4540,N_4546);
or UO_716 (O_716,N_4779,N_4857);
nand UO_717 (O_717,N_4545,N_4770);
nor UO_718 (O_718,N_4644,N_4842);
and UO_719 (O_719,N_4523,N_4681);
nand UO_720 (O_720,N_4970,N_4989);
or UO_721 (O_721,N_4671,N_4735);
and UO_722 (O_722,N_4925,N_4631);
nand UO_723 (O_723,N_4787,N_4590);
or UO_724 (O_724,N_4919,N_4852);
or UO_725 (O_725,N_4870,N_4542);
nor UO_726 (O_726,N_4544,N_4753);
and UO_727 (O_727,N_4565,N_4722);
nand UO_728 (O_728,N_4970,N_4878);
or UO_729 (O_729,N_4811,N_4756);
nand UO_730 (O_730,N_4776,N_4978);
nand UO_731 (O_731,N_4991,N_4551);
nor UO_732 (O_732,N_4809,N_4983);
nand UO_733 (O_733,N_4723,N_4762);
nand UO_734 (O_734,N_4781,N_4615);
or UO_735 (O_735,N_4764,N_4580);
and UO_736 (O_736,N_4863,N_4962);
nor UO_737 (O_737,N_4940,N_4500);
and UO_738 (O_738,N_4782,N_4630);
nor UO_739 (O_739,N_4967,N_4887);
nand UO_740 (O_740,N_4704,N_4702);
nor UO_741 (O_741,N_4720,N_4695);
nor UO_742 (O_742,N_4564,N_4604);
nor UO_743 (O_743,N_4801,N_4582);
nor UO_744 (O_744,N_4636,N_4847);
nand UO_745 (O_745,N_4560,N_4509);
nand UO_746 (O_746,N_4948,N_4854);
and UO_747 (O_747,N_4923,N_4821);
or UO_748 (O_748,N_4927,N_4809);
nand UO_749 (O_749,N_4945,N_4709);
or UO_750 (O_750,N_4587,N_4802);
or UO_751 (O_751,N_4805,N_4881);
nor UO_752 (O_752,N_4585,N_4654);
or UO_753 (O_753,N_4835,N_4776);
nand UO_754 (O_754,N_4971,N_4578);
or UO_755 (O_755,N_4905,N_4941);
and UO_756 (O_756,N_4757,N_4766);
or UO_757 (O_757,N_4920,N_4817);
nand UO_758 (O_758,N_4702,N_4728);
or UO_759 (O_759,N_4761,N_4838);
or UO_760 (O_760,N_4572,N_4522);
nor UO_761 (O_761,N_4838,N_4665);
and UO_762 (O_762,N_4792,N_4960);
and UO_763 (O_763,N_4994,N_4893);
and UO_764 (O_764,N_4681,N_4696);
and UO_765 (O_765,N_4637,N_4722);
nor UO_766 (O_766,N_4600,N_4941);
and UO_767 (O_767,N_4588,N_4723);
or UO_768 (O_768,N_4659,N_4661);
nor UO_769 (O_769,N_4824,N_4811);
and UO_770 (O_770,N_4718,N_4771);
or UO_771 (O_771,N_4522,N_4603);
and UO_772 (O_772,N_4888,N_4561);
nor UO_773 (O_773,N_4721,N_4726);
and UO_774 (O_774,N_4982,N_4642);
nand UO_775 (O_775,N_4861,N_4959);
nand UO_776 (O_776,N_4984,N_4983);
nand UO_777 (O_777,N_4816,N_4668);
nand UO_778 (O_778,N_4937,N_4863);
and UO_779 (O_779,N_4956,N_4865);
or UO_780 (O_780,N_4822,N_4542);
and UO_781 (O_781,N_4594,N_4879);
nor UO_782 (O_782,N_4588,N_4888);
nand UO_783 (O_783,N_4998,N_4694);
or UO_784 (O_784,N_4953,N_4754);
and UO_785 (O_785,N_4834,N_4847);
or UO_786 (O_786,N_4526,N_4763);
nor UO_787 (O_787,N_4597,N_4520);
nand UO_788 (O_788,N_4737,N_4619);
and UO_789 (O_789,N_4890,N_4959);
nand UO_790 (O_790,N_4617,N_4618);
and UO_791 (O_791,N_4586,N_4664);
and UO_792 (O_792,N_4510,N_4934);
or UO_793 (O_793,N_4929,N_4670);
or UO_794 (O_794,N_4907,N_4529);
nor UO_795 (O_795,N_4539,N_4616);
nand UO_796 (O_796,N_4792,N_4519);
nand UO_797 (O_797,N_4642,N_4788);
nand UO_798 (O_798,N_4696,N_4983);
or UO_799 (O_799,N_4865,N_4829);
nand UO_800 (O_800,N_4970,N_4962);
nand UO_801 (O_801,N_4713,N_4525);
or UO_802 (O_802,N_4687,N_4844);
or UO_803 (O_803,N_4901,N_4796);
and UO_804 (O_804,N_4924,N_4650);
or UO_805 (O_805,N_4815,N_4627);
nand UO_806 (O_806,N_4717,N_4663);
nor UO_807 (O_807,N_4531,N_4508);
nor UO_808 (O_808,N_4744,N_4734);
nor UO_809 (O_809,N_4966,N_4910);
and UO_810 (O_810,N_4531,N_4837);
and UO_811 (O_811,N_4974,N_4740);
nand UO_812 (O_812,N_4504,N_4601);
nand UO_813 (O_813,N_4956,N_4750);
nand UO_814 (O_814,N_4826,N_4812);
or UO_815 (O_815,N_4970,N_4900);
nand UO_816 (O_816,N_4861,N_4705);
or UO_817 (O_817,N_4584,N_4915);
nor UO_818 (O_818,N_4732,N_4866);
nand UO_819 (O_819,N_4959,N_4733);
and UO_820 (O_820,N_4888,N_4690);
and UO_821 (O_821,N_4725,N_4552);
or UO_822 (O_822,N_4718,N_4595);
nand UO_823 (O_823,N_4878,N_4877);
nor UO_824 (O_824,N_4864,N_4582);
and UO_825 (O_825,N_4631,N_4732);
and UO_826 (O_826,N_4811,N_4514);
nand UO_827 (O_827,N_4852,N_4504);
and UO_828 (O_828,N_4841,N_4880);
and UO_829 (O_829,N_4824,N_4507);
or UO_830 (O_830,N_4787,N_4816);
nor UO_831 (O_831,N_4528,N_4589);
nand UO_832 (O_832,N_4974,N_4852);
or UO_833 (O_833,N_4729,N_4969);
or UO_834 (O_834,N_4922,N_4653);
or UO_835 (O_835,N_4850,N_4550);
or UO_836 (O_836,N_4988,N_4569);
nor UO_837 (O_837,N_4881,N_4766);
nor UO_838 (O_838,N_4804,N_4554);
nor UO_839 (O_839,N_4831,N_4807);
nand UO_840 (O_840,N_4677,N_4762);
nor UO_841 (O_841,N_4625,N_4732);
or UO_842 (O_842,N_4692,N_4565);
nand UO_843 (O_843,N_4684,N_4845);
and UO_844 (O_844,N_4762,N_4505);
nand UO_845 (O_845,N_4876,N_4508);
nand UO_846 (O_846,N_4980,N_4682);
nand UO_847 (O_847,N_4550,N_4644);
nand UO_848 (O_848,N_4854,N_4821);
or UO_849 (O_849,N_4985,N_4612);
and UO_850 (O_850,N_4607,N_4696);
nand UO_851 (O_851,N_4537,N_4643);
nor UO_852 (O_852,N_4920,N_4561);
nand UO_853 (O_853,N_4661,N_4684);
and UO_854 (O_854,N_4795,N_4786);
nand UO_855 (O_855,N_4945,N_4568);
and UO_856 (O_856,N_4554,N_4617);
nand UO_857 (O_857,N_4916,N_4890);
and UO_858 (O_858,N_4764,N_4515);
nand UO_859 (O_859,N_4812,N_4967);
or UO_860 (O_860,N_4774,N_4854);
and UO_861 (O_861,N_4847,N_4590);
nor UO_862 (O_862,N_4526,N_4793);
and UO_863 (O_863,N_4710,N_4782);
or UO_864 (O_864,N_4612,N_4868);
nor UO_865 (O_865,N_4551,N_4849);
or UO_866 (O_866,N_4539,N_4917);
and UO_867 (O_867,N_4762,N_4767);
nor UO_868 (O_868,N_4649,N_4841);
or UO_869 (O_869,N_4751,N_4631);
nand UO_870 (O_870,N_4832,N_4534);
nor UO_871 (O_871,N_4736,N_4743);
or UO_872 (O_872,N_4500,N_4550);
or UO_873 (O_873,N_4864,N_4834);
nor UO_874 (O_874,N_4939,N_4936);
and UO_875 (O_875,N_4923,N_4708);
and UO_876 (O_876,N_4883,N_4874);
nor UO_877 (O_877,N_4856,N_4609);
xnor UO_878 (O_878,N_4883,N_4619);
nand UO_879 (O_879,N_4501,N_4787);
and UO_880 (O_880,N_4597,N_4522);
and UO_881 (O_881,N_4922,N_4841);
or UO_882 (O_882,N_4820,N_4736);
and UO_883 (O_883,N_4671,N_4703);
nor UO_884 (O_884,N_4539,N_4636);
or UO_885 (O_885,N_4516,N_4538);
nor UO_886 (O_886,N_4782,N_4759);
and UO_887 (O_887,N_4626,N_4877);
and UO_888 (O_888,N_4790,N_4766);
and UO_889 (O_889,N_4765,N_4647);
nor UO_890 (O_890,N_4540,N_4654);
and UO_891 (O_891,N_4842,N_4792);
nand UO_892 (O_892,N_4526,N_4770);
and UO_893 (O_893,N_4817,N_4744);
or UO_894 (O_894,N_4989,N_4530);
and UO_895 (O_895,N_4906,N_4936);
or UO_896 (O_896,N_4969,N_4676);
nand UO_897 (O_897,N_4522,N_4977);
nor UO_898 (O_898,N_4645,N_4734);
and UO_899 (O_899,N_4802,N_4961);
nor UO_900 (O_900,N_4797,N_4727);
xnor UO_901 (O_901,N_4971,N_4692);
nand UO_902 (O_902,N_4925,N_4588);
nand UO_903 (O_903,N_4722,N_4644);
nor UO_904 (O_904,N_4787,N_4594);
nand UO_905 (O_905,N_4855,N_4529);
or UO_906 (O_906,N_4936,N_4868);
nor UO_907 (O_907,N_4924,N_4790);
xnor UO_908 (O_908,N_4562,N_4655);
and UO_909 (O_909,N_4959,N_4653);
nor UO_910 (O_910,N_4909,N_4852);
or UO_911 (O_911,N_4920,N_4991);
nor UO_912 (O_912,N_4645,N_4615);
or UO_913 (O_913,N_4571,N_4676);
and UO_914 (O_914,N_4671,N_4973);
nand UO_915 (O_915,N_4888,N_4768);
and UO_916 (O_916,N_4735,N_4959);
nor UO_917 (O_917,N_4718,N_4645);
and UO_918 (O_918,N_4519,N_4712);
nand UO_919 (O_919,N_4608,N_4896);
xnor UO_920 (O_920,N_4536,N_4725);
or UO_921 (O_921,N_4771,N_4833);
and UO_922 (O_922,N_4815,N_4575);
nor UO_923 (O_923,N_4832,N_4565);
nand UO_924 (O_924,N_4698,N_4778);
nand UO_925 (O_925,N_4870,N_4515);
nand UO_926 (O_926,N_4921,N_4622);
nand UO_927 (O_927,N_4977,N_4975);
nand UO_928 (O_928,N_4733,N_4740);
or UO_929 (O_929,N_4813,N_4743);
nand UO_930 (O_930,N_4845,N_4761);
and UO_931 (O_931,N_4956,N_4856);
nand UO_932 (O_932,N_4974,N_4971);
or UO_933 (O_933,N_4808,N_4674);
or UO_934 (O_934,N_4575,N_4690);
nor UO_935 (O_935,N_4969,N_4931);
or UO_936 (O_936,N_4941,N_4890);
nor UO_937 (O_937,N_4679,N_4771);
and UO_938 (O_938,N_4936,N_4863);
nor UO_939 (O_939,N_4927,N_4714);
nand UO_940 (O_940,N_4694,N_4706);
nand UO_941 (O_941,N_4585,N_4527);
nor UO_942 (O_942,N_4578,N_4968);
and UO_943 (O_943,N_4944,N_4511);
nor UO_944 (O_944,N_4957,N_4696);
nand UO_945 (O_945,N_4640,N_4813);
and UO_946 (O_946,N_4720,N_4809);
nand UO_947 (O_947,N_4614,N_4731);
or UO_948 (O_948,N_4687,N_4799);
or UO_949 (O_949,N_4600,N_4785);
or UO_950 (O_950,N_4727,N_4774);
and UO_951 (O_951,N_4526,N_4881);
and UO_952 (O_952,N_4565,N_4712);
nor UO_953 (O_953,N_4674,N_4584);
or UO_954 (O_954,N_4837,N_4565);
nor UO_955 (O_955,N_4662,N_4687);
nand UO_956 (O_956,N_4758,N_4742);
and UO_957 (O_957,N_4736,N_4512);
nor UO_958 (O_958,N_4604,N_4509);
nand UO_959 (O_959,N_4562,N_4589);
nand UO_960 (O_960,N_4527,N_4811);
and UO_961 (O_961,N_4667,N_4942);
nand UO_962 (O_962,N_4541,N_4929);
or UO_963 (O_963,N_4856,N_4553);
or UO_964 (O_964,N_4952,N_4562);
nand UO_965 (O_965,N_4900,N_4858);
nor UO_966 (O_966,N_4704,N_4811);
nor UO_967 (O_967,N_4702,N_4695);
nand UO_968 (O_968,N_4528,N_4852);
nor UO_969 (O_969,N_4651,N_4677);
and UO_970 (O_970,N_4633,N_4597);
nor UO_971 (O_971,N_4596,N_4532);
nand UO_972 (O_972,N_4823,N_4527);
nand UO_973 (O_973,N_4742,N_4536);
or UO_974 (O_974,N_4688,N_4667);
and UO_975 (O_975,N_4629,N_4571);
and UO_976 (O_976,N_4649,N_4612);
and UO_977 (O_977,N_4971,N_4651);
and UO_978 (O_978,N_4781,N_4584);
and UO_979 (O_979,N_4661,N_4502);
nand UO_980 (O_980,N_4976,N_4532);
nor UO_981 (O_981,N_4718,N_4612);
nand UO_982 (O_982,N_4758,N_4824);
or UO_983 (O_983,N_4759,N_4586);
or UO_984 (O_984,N_4575,N_4560);
and UO_985 (O_985,N_4847,N_4805);
or UO_986 (O_986,N_4974,N_4696);
and UO_987 (O_987,N_4958,N_4776);
xnor UO_988 (O_988,N_4903,N_4580);
or UO_989 (O_989,N_4917,N_4993);
or UO_990 (O_990,N_4718,N_4755);
nand UO_991 (O_991,N_4889,N_4531);
nand UO_992 (O_992,N_4590,N_4923);
or UO_993 (O_993,N_4866,N_4582);
or UO_994 (O_994,N_4951,N_4757);
nor UO_995 (O_995,N_4675,N_4917);
and UO_996 (O_996,N_4626,N_4583);
nor UO_997 (O_997,N_4749,N_4826);
nor UO_998 (O_998,N_4947,N_4996);
or UO_999 (O_999,N_4835,N_4677);
endmodule