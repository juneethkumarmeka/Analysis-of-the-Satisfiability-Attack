module basic_3000_30000_3500_6_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
or U0 (N_0,In_1599,In_1916);
and U1 (N_1,In_2248,In_2343);
and U2 (N_2,In_411,In_1273);
or U3 (N_3,In_138,In_2521);
or U4 (N_4,In_239,In_2527);
nor U5 (N_5,In_45,In_2977);
nand U6 (N_6,In_2894,In_297);
xnor U7 (N_7,In_280,In_2062);
xnor U8 (N_8,In_2313,In_525);
nor U9 (N_9,In_2374,In_776);
nand U10 (N_10,In_2936,In_2346);
nand U11 (N_11,In_1959,In_449);
nand U12 (N_12,In_1182,In_207);
or U13 (N_13,In_1770,In_1398);
and U14 (N_14,In_891,In_1722);
xnor U15 (N_15,In_1243,In_1339);
and U16 (N_16,In_2864,In_2339);
nor U17 (N_17,In_290,In_2606);
nand U18 (N_18,In_2580,In_2481);
or U19 (N_19,In_2508,In_2239);
nand U20 (N_20,In_2445,In_2371);
nor U21 (N_21,In_491,In_711);
xnor U22 (N_22,In_2180,In_1016);
xnor U23 (N_23,In_1871,In_1221);
or U24 (N_24,In_378,In_661);
xnor U25 (N_25,In_2219,In_873);
nand U26 (N_26,In_1125,In_1235);
and U27 (N_27,In_695,In_1776);
nand U28 (N_28,In_2889,In_708);
or U29 (N_29,In_2207,In_622);
nand U30 (N_30,In_309,In_2137);
xnor U31 (N_31,In_619,In_1593);
nor U32 (N_32,In_1969,In_1992);
nor U33 (N_33,In_1910,In_2928);
xor U34 (N_34,In_166,In_398);
xnor U35 (N_35,In_2019,In_146);
and U36 (N_36,In_2910,In_2881);
or U37 (N_37,In_706,In_1848);
nor U38 (N_38,In_2483,In_83);
xor U39 (N_39,In_2042,In_1373);
nor U40 (N_40,In_1574,In_18);
and U41 (N_41,In_1086,In_1798);
nor U42 (N_42,In_1359,In_629);
and U43 (N_43,In_1923,In_1260);
and U44 (N_44,In_2751,In_782);
nor U45 (N_45,In_731,In_2170);
and U46 (N_46,In_811,In_752);
or U47 (N_47,In_2273,In_896);
xor U48 (N_48,In_2309,In_2503);
xor U49 (N_49,In_1150,In_2571);
and U50 (N_50,In_2615,In_1464);
nand U51 (N_51,In_2533,In_726);
nor U52 (N_52,In_2830,In_1090);
nand U53 (N_53,In_721,In_520);
nor U54 (N_54,In_2079,In_1606);
nand U55 (N_55,In_2603,In_203);
and U56 (N_56,In_1432,In_1516);
nand U57 (N_57,In_2496,In_1311);
nand U58 (N_58,In_2024,In_2083);
xnor U59 (N_59,In_121,In_723);
or U60 (N_60,In_2636,In_990);
xnor U61 (N_61,In_2842,In_808);
or U62 (N_62,In_155,In_1799);
or U63 (N_63,In_1056,In_1408);
nand U64 (N_64,In_2278,In_534);
nor U65 (N_65,In_668,In_2152);
nor U66 (N_66,In_202,In_1246);
nand U67 (N_67,In_28,In_74);
or U68 (N_68,In_1982,In_2310);
nor U69 (N_69,In_2944,In_2619);
or U70 (N_70,In_1586,In_1867);
nand U71 (N_71,In_2526,In_2617);
nor U72 (N_72,In_2341,In_2210);
xnor U73 (N_73,In_2632,In_1477);
nand U74 (N_74,In_246,In_565);
xnor U75 (N_75,In_2724,In_92);
nor U76 (N_76,In_1466,In_2302);
nand U77 (N_77,In_2112,In_2148);
and U78 (N_78,In_856,In_1092);
and U79 (N_79,In_876,In_601);
and U80 (N_80,In_2575,In_529);
xor U81 (N_81,In_2652,In_2014);
nor U82 (N_82,In_1116,In_2599);
xnor U83 (N_83,In_446,In_2721);
or U84 (N_84,In_278,In_184);
nand U85 (N_85,In_1225,In_122);
xnor U86 (N_86,In_263,In_1181);
or U87 (N_87,In_585,In_507);
xor U88 (N_88,In_2190,In_871);
nor U89 (N_89,In_1568,In_1201);
nand U90 (N_90,In_2337,In_807);
or U91 (N_91,In_1136,In_2450);
or U92 (N_92,In_1925,In_1860);
or U93 (N_93,In_1366,In_1229);
xnor U94 (N_94,In_167,In_2933);
nand U95 (N_95,In_1226,In_1482);
nor U96 (N_96,In_2736,In_927);
nor U97 (N_97,In_2931,In_786);
nor U98 (N_98,In_2589,In_2530);
nand U99 (N_99,In_1692,In_583);
or U100 (N_100,In_1943,In_595);
xor U101 (N_101,In_998,In_991);
or U102 (N_102,In_2631,In_2319);
nor U103 (N_103,In_432,In_527);
nand U104 (N_104,In_1906,In_1140);
nand U105 (N_105,In_2638,In_127);
xnor U106 (N_106,In_922,In_2776);
nor U107 (N_107,In_2887,In_563);
or U108 (N_108,In_2913,In_2717);
nor U109 (N_109,In_921,In_759);
or U110 (N_110,In_1750,In_2912);
and U111 (N_111,In_821,In_34);
xor U112 (N_112,In_2710,In_826);
xor U113 (N_113,In_1384,In_337);
xnor U114 (N_114,In_400,In_86);
nor U115 (N_115,In_2793,In_402);
and U116 (N_116,In_2449,In_1983);
xnor U117 (N_117,In_232,In_911);
or U118 (N_118,In_1171,In_21);
and U119 (N_119,In_1039,In_1812);
nand U120 (N_120,In_1105,In_2369);
and U121 (N_121,In_1347,In_2516);
nor U122 (N_122,In_1761,In_89);
nand U123 (N_123,In_2839,In_634);
and U124 (N_124,In_1961,In_567);
nand U125 (N_125,In_704,In_2965);
nand U126 (N_126,In_2420,In_2844);
nand U127 (N_127,In_100,In_1123);
and U128 (N_128,In_2,In_1443);
nand U129 (N_129,In_2582,In_2858);
xor U130 (N_130,In_2338,In_2493);
xnor U131 (N_131,In_114,In_195);
or U132 (N_132,In_1401,In_987);
or U133 (N_133,In_700,In_1682);
or U134 (N_134,In_2678,In_1122);
and U135 (N_135,In_956,In_1470);
or U136 (N_136,In_2029,In_1504);
nand U137 (N_137,In_2943,In_2556);
or U138 (N_138,In_1106,In_173);
and U139 (N_139,In_653,In_1327);
nor U140 (N_140,In_522,In_1188);
or U141 (N_141,In_2537,In_854);
and U142 (N_142,In_1804,In_2046);
xor U143 (N_143,In_256,In_2895);
or U144 (N_144,In_762,In_1989);
nand U145 (N_145,In_1239,In_1209);
or U146 (N_146,In_1250,In_132);
nor U147 (N_147,In_974,In_1538);
and U148 (N_148,In_2404,In_2939);
xnor U149 (N_149,In_61,In_2584);
nand U150 (N_150,In_1291,In_1011);
and U151 (N_151,In_137,In_37);
and U152 (N_152,In_1435,In_1540);
xor U153 (N_153,In_988,In_1004);
nor U154 (N_154,In_681,In_1107);
nor U155 (N_155,In_57,In_233);
or U156 (N_156,In_1375,In_1055);
or U157 (N_157,In_2090,In_660);
or U158 (N_158,In_620,In_347);
nand U159 (N_159,In_321,In_758);
and U160 (N_160,In_2455,In_2116);
nand U161 (N_161,In_2504,In_1367);
xnor U162 (N_162,In_192,In_2353);
nor U163 (N_163,In_809,In_2825);
xor U164 (N_164,In_2954,In_2154);
and U165 (N_165,In_1245,In_1721);
xnor U166 (N_166,In_1936,In_2593);
xnor U167 (N_167,In_2354,In_2654);
nand U168 (N_168,In_1218,In_2360);
nand U169 (N_169,In_790,In_2967);
and U170 (N_170,In_1614,In_5);
or U171 (N_171,In_2311,In_396);
nor U172 (N_172,In_1553,In_1180);
nor U173 (N_173,In_1383,In_2588);
or U174 (N_174,In_677,In_669);
nor U175 (N_175,In_2370,In_140);
nor U176 (N_176,In_1284,In_2733);
xnor U177 (N_177,In_2701,In_1497);
xor U178 (N_178,In_2921,In_1610);
xor U179 (N_179,In_1442,In_313);
or U180 (N_180,In_2861,In_2113);
nand U181 (N_181,In_2394,In_2845);
nand U182 (N_182,In_943,In_1619);
nor U183 (N_183,In_1753,In_171);
nand U184 (N_184,In_1364,In_2008);
or U185 (N_185,In_1036,In_32);
nor U186 (N_186,In_73,In_2513);
and U187 (N_187,In_898,In_447);
or U188 (N_188,In_46,In_191);
or U189 (N_189,In_628,In_365);
nand U190 (N_190,In_2315,In_403);
xor U191 (N_191,In_2390,In_1085);
and U192 (N_192,In_2590,In_657);
and U193 (N_193,In_2380,In_1490);
or U194 (N_194,In_993,In_1113);
xnor U195 (N_195,In_1319,In_1869);
xnor U196 (N_196,In_264,In_1095);
nand U197 (N_197,In_142,In_81);
xor U198 (N_198,In_2422,In_2809);
nand U199 (N_199,In_2897,In_36);
and U200 (N_200,In_1025,In_1353);
nor U201 (N_201,In_333,In_1087);
or U202 (N_202,In_472,In_2114);
nand U203 (N_203,In_2262,In_2209);
or U204 (N_204,In_1154,In_1533);
nor U205 (N_205,In_717,In_923);
nand U206 (N_206,In_1542,In_2110);
and U207 (N_207,In_970,In_2836);
and U208 (N_208,In_160,In_1028);
nor U209 (N_209,In_2468,In_368);
or U210 (N_210,In_2224,In_1711);
or U211 (N_211,In_967,In_2872);
xor U212 (N_212,In_957,In_474);
and U213 (N_213,In_1815,In_1927);
and U214 (N_214,In_2768,In_1792);
or U215 (N_215,In_503,In_53);
xor U216 (N_216,In_1189,In_2096);
nor U217 (N_217,In_2147,In_1978);
or U218 (N_218,In_2092,In_463);
and U219 (N_219,In_1050,In_1407);
and U220 (N_220,In_461,In_914);
xor U221 (N_221,In_2232,In_2168);
or U222 (N_222,In_1308,In_437);
nor U223 (N_223,In_2362,In_785);
and U224 (N_224,In_2326,In_64);
or U225 (N_225,In_1585,In_748);
nor U226 (N_226,In_2203,In_1826);
and U227 (N_227,In_516,In_1990);
and U228 (N_228,In_917,In_43);
or U229 (N_229,In_644,In_2192);
nor U230 (N_230,In_1083,In_1313);
and U231 (N_231,In_1270,In_1119);
xor U232 (N_232,In_2783,In_436);
nand U233 (N_233,In_1695,In_2901);
and U234 (N_234,In_554,In_1447);
xnor U235 (N_235,In_1419,In_243);
nand U236 (N_236,In_2206,In_1523);
xnor U237 (N_237,In_1775,In_765);
and U238 (N_238,In_219,In_1905);
or U239 (N_239,In_82,In_1617);
xnor U240 (N_240,In_2755,In_404);
and U241 (N_241,In_615,In_1758);
and U242 (N_242,In_1893,In_2572);
and U243 (N_243,In_1467,In_2267);
nor U244 (N_244,In_234,In_1487);
or U245 (N_245,In_2882,In_2052);
nor U246 (N_246,In_1336,In_1642);
and U247 (N_247,In_409,In_63);
nor U248 (N_248,In_1751,In_2543);
nand U249 (N_249,In_1683,In_2650);
xnor U250 (N_250,In_2061,In_2828);
and U251 (N_251,In_2460,In_274);
or U252 (N_252,In_1078,In_287);
nor U253 (N_253,In_687,In_2562);
nor U254 (N_254,In_31,In_1790);
or U255 (N_255,In_1465,In_1247);
nor U256 (N_256,In_2726,In_1794);
nand U257 (N_257,In_2271,In_1350);
nor U258 (N_258,In_330,In_2517);
or U259 (N_259,In_354,In_2667);
and U260 (N_260,In_1064,In_2005);
nand U261 (N_261,In_1628,In_2987);
xnor U262 (N_262,In_2474,In_1281);
nand U263 (N_263,In_1499,In_2205);
nand U264 (N_264,In_1963,In_1391);
nor U265 (N_265,In_1076,In_1395);
and U266 (N_266,In_569,In_1788);
or U267 (N_267,In_2485,In_1126);
and U268 (N_268,In_952,In_302);
nor U269 (N_269,In_1530,In_1445);
nor U270 (N_270,In_939,In_1605);
xor U271 (N_271,In_1479,In_1814);
xnor U272 (N_272,In_452,In_1981);
or U273 (N_273,In_2002,In_2523);
nor U274 (N_274,In_519,In_1904);
nor U275 (N_275,In_1012,In_2237);
nor U276 (N_276,In_778,In_2034);
nor U277 (N_277,In_592,In_582);
or U278 (N_278,In_584,In_1550);
and U279 (N_279,In_1747,In_1658);
or U280 (N_280,In_2214,In_2163);
xnor U281 (N_281,In_564,In_837);
and U282 (N_282,In_2738,In_707);
or U283 (N_283,In_2675,In_2452);
xor U284 (N_284,In_1731,In_1743);
and U285 (N_285,In_855,In_815);
xnor U286 (N_286,In_236,In_2056);
or U287 (N_287,In_1474,In_1724);
xor U288 (N_288,In_2094,In_1066);
nor U289 (N_289,In_479,In_1647);
nor U290 (N_290,In_817,In_1496);
nand U291 (N_291,In_295,In_2121);
nor U292 (N_292,In_2119,In_2561);
or U293 (N_293,In_2478,In_1152);
and U294 (N_294,In_2410,In_2771);
and U295 (N_295,In_1559,In_947);
xnor U296 (N_296,In_13,In_1198);
and U297 (N_297,In_2544,In_1741);
and U298 (N_298,In_1088,In_1436);
nor U299 (N_299,In_252,In_2820);
nor U300 (N_300,In_1144,In_2869);
or U301 (N_301,In_2659,In_2684);
nor U302 (N_302,In_1096,In_2649);
xor U303 (N_303,In_2447,In_33);
xnor U304 (N_304,In_869,In_300);
or U305 (N_305,In_2787,In_2679);
nor U306 (N_306,In_2653,In_1355);
and U307 (N_307,In_2323,In_1851);
nor U308 (N_308,In_1760,In_1234);
nand U309 (N_309,In_2538,In_2792);
or U310 (N_310,In_1406,In_2066);
and U311 (N_311,In_1785,In_574);
xnor U312 (N_312,In_75,In_2801);
xor U313 (N_313,In_265,In_2242);
nor U314 (N_314,In_2077,In_469);
nor U315 (N_315,In_1034,In_1681);
nand U316 (N_316,In_2378,In_307);
nor U317 (N_317,In_1303,In_2389);
and U318 (N_318,In_2236,In_2922);
xor U319 (N_319,In_1600,In_2790);
nand U320 (N_320,In_1132,In_531);
nand U321 (N_321,In_69,In_1323);
nand U322 (N_322,In_1582,In_2158);
xor U323 (N_323,In_909,In_2618);
nand U324 (N_324,In_1791,In_1588);
and U325 (N_325,In_2534,In_277);
and U326 (N_326,In_2693,In_812);
nor U327 (N_327,In_1097,In_2648);
and U328 (N_328,In_850,In_715);
and U329 (N_329,In_843,In_655);
nand U330 (N_330,In_1876,In_1891);
and U331 (N_331,In_496,In_2856);
and U332 (N_332,In_2322,In_1254);
or U333 (N_333,In_2275,In_1153);
nor U334 (N_334,In_2995,In_612);
xnor U335 (N_335,In_665,In_2863);
xor U336 (N_336,In_1163,In_2963);
and U337 (N_337,In_2662,In_1224);
nand U338 (N_338,In_1244,In_1404);
and U339 (N_339,In_296,In_1889);
nand U340 (N_340,In_2962,In_959);
nand U341 (N_341,In_1018,In_8);
nand U342 (N_342,In_2386,In_2274);
or U343 (N_343,In_2761,In_2494);
nand U344 (N_344,In_2500,In_2231);
or U345 (N_345,In_1808,In_360);
or U346 (N_346,In_2246,In_366);
and U347 (N_347,In_861,In_2876);
xnor U348 (N_348,In_1584,In_1591);
and U349 (N_349,In_1301,In_187);
and U350 (N_350,In_1040,In_1746);
nand U351 (N_351,In_1771,In_1257);
nor U352 (N_352,In_1232,In_1074);
nand U353 (N_353,In_1882,In_1809);
and U354 (N_354,In_2814,In_2959);
xnor U355 (N_355,In_678,In_1067);
nand U356 (N_356,In_2958,In_656);
and U357 (N_357,In_2752,In_1202);
nand U358 (N_358,In_1237,In_2321);
or U359 (N_359,In_1360,In_2082);
nor U360 (N_360,In_1314,In_2229);
nor U361 (N_361,In_2896,In_1897);
xnor U362 (N_362,In_903,In_124);
or U363 (N_363,In_1424,In_2695);
and U364 (N_364,In_495,In_2153);
nor U365 (N_365,In_419,In_504);
and U366 (N_366,In_2280,In_2331);
nand U367 (N_367,In_180,In_996);
nor U368 (N_368,In_1026,In_2253);
nand U369 (N_369,In_702,In_710);
nand U370 (N_370,In_487,In_1716);
nand U371 (N_371,In_1767,In_376);
or U372 (N_372,In_1537,In_1267);
nor U373 (N_373,In_129,In_1165);
or U374 (N_374,In_251,In_2157);
nor U375 (N_375,In_884,In_1615);
nand U376 (N_376,In_1577,In_2690);
and U377 (N_377,In_11,In_1370);
xnor U378 (N_378,In_1227,In_1986);
nand U379 (N_379,In_2296,In_1494);
nor U380 (N_380,In_498,In_1797);
nor U381 (N_381,In_865,In_2087);
nor U382 (N_382,In_1875,In_235);
nand U383 (N_383,In_2412,In_2796);
or U384 (N_384,In_1844,In_2874);
and U385 (N_385,In_99,In_2377);
and U386 (N_386,In_1846,In_2134);
or U387 (N_387,In_538,In_1866);
and U388 (N_388,In_214,In_2030);
and U389 (N_389,In_627,In_1390);
xnor U390 (N_390,In_1520,In_596);
or U391 (N_391,In_730,In_2713);
xor U392 (N_392,In_1361,In_2330);
nand U393 (N_393,In_1696,In_946);
and U394 (N_394,In_468,In_980);
nand U395 (N_395,In_237,In_2495);
and U396 (N_396,In_2405,In_1139);
nand U397 (N_397,In_1509,In_1024);
or U398 (N_398,In_2816,In_1156);
and U399 (N_399,In_2290,In_1623);
or U400 (N_400,In_899,In_2195);
or U401 (N_401,In_2697,In_2078);
and U402 (N_402,In_2411,In_458);
nand U403 (N_403,In_919,In_1485);
nor U404 (N_404,In_2084,In_1877);
nand U405 (N_405,In_1344,In_2502);
nor U406 (N_406,In_1999,In_908);
nand U407 (N_407,In_1885,In_2564);
xor U408 (N_408,In_728,In_285);
and U409 (N_409,In_2031,In_1899);
xnor U410 (N_410,In_2204,In_772);
nor U411 (N_411,In_1669,In_1702);
or U412 (N_412,In_887,In_2824);
and U413 (N_413,In_1149,In_2367);
or U414 (N_414,In_1703,In_1019);
nand U415 (N_415,In_2877,In_1580);
nand U416 (N_416,In_2388,In_1883);
xnor U417 (N_417,In_2391,In_868);
nand U418 (N_418,In_148,In_2202);
xnor U419 (N_419,In_892,In_2235);
xnor U420 (N_420,In_2781,In_2908);
nand U421 (N_421,In_465,In_391);
or U422 (N_422,In_176,In_679);
or U423 (N_423,In_2786,In_2174);
or U424 (N_424,In_2304,In_481);
nand U425 (N_425,In_1133,In_1423);
nand U426 (N_426,In_1694,In_2287);
nand U427 (N_427,In_1318,In_1014);
or U428 (N_428,In_1127,In_1416);
xnor U429 (N_429,In_126,In_1864);
nor U430 (N_430,In_1394,In_98);
or U431 (N_431,In_2320,In_96);
and U432 (N_432,In_261,In_1870);
nor U433 (N_433,In_1945,In_2003);
nand U434 (N_434,In_1858,In_2924);
or U435 (N_435,In_2001,In_2769);
or U436 (N_436,In_1507,In_1102);
and U437 (N_437,In_1583,In_1001);
nand U438 (N_438,In_1862,In_2990);
xor U439 (N_439,In_1389,In_802);
nand U440 (N_440,In_2841,In_2010);
nand U441 (N_441,In_2971,In_272);
and U442 (N_442,In_1434,In_51);
nor U443 (N_443,In_1680,In_65);
nand U444 (N_444,In_548,In_2283);
xnor U445 (N_445,In_2373,In_2050);
and U446 (N_446,In_188,In_1697);
or U447 (N_447,In_374,In_696);
and U448 (N_448,In_2616,In_1446);
or U449 (N_449,In_2555,In_1486);
and U450 (N_450,In_1251,In_795);
nand U451 (N_451,In_1134,In_2870);
or U452 (N_452,In_2150,In_1317);
or U453 (N_453,In_2779,In_1888);
xnor U454 (N_454,In_1324,In_838);
nand U455 (N_455,In_116,In_2162);
xnor U456 (N_456,In_1501,In_2501);
or U457 (N_457,In_1290,In_269);
nand U458 (N_458,In_1099,In_2818);
or U459 (N_459,In_1415,In_417);
nor U460 (N_460,In_1543,In_1985);
xor U461 (N_461,In_2645,In_606);
and U462 (N_462,In_2625,In_1958);
nor U463 (N_463,In_2691,In_1607);
xor U464 (N_464,In_1142,In_544);
xnor U465 (N_465,In_552,In_494);
and U466 (N_466,In_150,In_2144);
xnor U467 (N_467,In_2727,In_2525);
nor U468 (N_468,In_1135,In_1977);
and U469 (N_469,In_992,In_1670);
xor U470 (N_470,In_633,In_1100);
nand U471 (N_471,In_528,In_359);
xnor U472 (N_472,In_853,In_1739);
nand U473 (N_473,In_1939,In_1839);
or U474 (N_474,In_1428,In_1661);
and U475 (N_475,In_2393,In_2670);
and U476 (N_476,In_331,In_2417);
and U477 (N_477,In_1204,In_979);
nand U478 (N_478,In_2851,In_663);
and U479 (N_479,In_1294,In_355);
xor U480 (N_480,In_1027,In_2984);
xor U481 (N_481,In_931,In_2609);
and U482 (N_482,In_725,In_2141);
xnor U483 (N_483,In_1633,In_720);
nand U484 (N_484,In_2621,In_1675);
nand U485 (N_485,In_2750,In_1060);
xnor U486 (N_486,In_2138,In_2514);
xor U487 (N_487,In_416,In_1385);
or U488 (N_488,In_2051,In_1962);
xnor U489 (N_489,In_639,In_562);
xnor U490 (N_490,In_1616,In_152);
nor U491 (N_491,In_754,In_949);
and U492 (N_492,In_2179,In_571);
or U493 (N_493,In_2762,In_2126);
and U494 (N_494,In_1575,In_2635);
nand U495 (N_495,In_59,In_2146);
nor U496 (N_496,In_111,In_2708);
or U497 (N_497,In_2866,In_267);
and U498 (N_498,In_2676,In_835);
nor U499 (N_499,In_2840,In_1960);
nand U500 (N_500,In_1176,In_1320);
nor U501 (N_501,In_1732,In_1413);
xnor U502 (N_502,In_1873,In_1934);
and U503 (N_503,In_206,In_125);
nor U504 (N_504,In_165,In_2254);
and U505 (N_505,In_2499,In_672);
nor U506 (N_506,In_2227,In_1382);
nand U507 (N_507,In_2382,In_497);
nand U508 (N_508,In_7,In_1264);
nor U509 (N_509,In_766,In_1441);
and U510 (N_510,In_2914,In_764);
and U511 (N_511,In_460,In_1315);
or U512 (N_512,In_926,In_1884);
nor U513 (N_513,In_2479,In_16);
nand U514 (N_514,In_324,In_1548);
or U515 (N_515,In_2935,In_936);
nor U516 (N_516,In_222,In_618);
and U517 (N_517,In_1995,In_2586);
and U518 (N_518,In_154,In_2040);
nor U519 (N_519,In_2630,In_556);
nand U520 (N_520,In_1946,In_2357);
nand U521 (N_521,In_2048,In_2757);
and U522 (N_522,In_370,In_769);
nor U523 (N_523,In_561,In_1343);
and U524 (N_524,In_1725,In_70);
or U525 (N_525,In_942,In_609);
xnor U526 (N_526,In_392,In_1214);
nand U527 (N_527,In_1693,In_1994);
nor U528 (N_528,In_2563,In_1525);
nand U529 (N_529,In_1535,In_201);
nand U530 (N_530,In_1508,In_1919);
or U531 (N_531,In_553,In_1175);
xor U532 (N_532,In_2366,In_872);
xor U533 (N_533,In_836,In_1918);
and U534 (N_534,In_1953,In_1531);
and U535 (N_535,In_760,In_1381);
or U536 (N_536,In_1340,In_2039);
and U537 (N_537,In_2355,In_2469);
nand U538 (N_538,In_938,In_262);
xnor U539 (N_539,In_2688,In_2794);
xor U540 (N_540,In_2156,In_576);
and U541 (N_541,In_866,In_1268);
xnor U542 (N_542,In_2604,In_781);
nor U543 (N_543,In_117,In_10);
or U544 (N_544,In_1720,In_480);
nand U545 (N_545,In_2729,In_2865);
and U546 (N_546,In_2301,In_2443);
and U547 (N_547,In_231,In_1827);
nor U548 (N_548,In_2559,In_2926);
nor U549 (N_549,In_12,In_1093);
nand U550 (N_550,In_2597,In_1996);
nand U551 (N_551,In_2699,In_2554);
or U552 (N_552,In_1565,In_877);
nor U553 (N_553,In_1021,In_509);
and U554 (N_554,In_602,In_230);
nor U555 (N_555,In_312,In_25);
and U556 (N_556,In_1957,In_204);
nand U557 (N_557,In_2238,In_2911);
xnor U558 (N_558,In_1756,In_1688);
nor U559 (N_559,In_2013,In_2132);
xor U560 (N_560,In_2893,In_2748);
or U561 (N_561,In_2651,In_743);
nand U562 (N_562,In_2385,In_1653);
or U563 (N_563,In_2379,In_1003);
and U564 (N_564,In_1700,In_2437);
nor U565 (N_565,In_739,In_722);
nand U566 (N_566,In_250,In_2819);
or U567 (N_567,In_798,In_1045);
xnor U568 (N_568,In_273,In_1755);
nor U569 (N_569,In_2387,In_2557);
nand U570 (N_570,In_2550,In_325);
and U571 (N_571,In_1667,In_1828);
or U572 (N_572,In_1304,In_1793);
and U573 (N_573,In_2425,In_1759);
nand U574 (N_574,In_2120,In_2067);
xor U575 (N_575,In_645,In_894);
and U576 (N_576,In_2661,In_2643);
and U577 (N_577,In_275,In_2929);
nand U578 (N_578,In_2608,In_2532);
or U579 (N_579,In_1451,In_1834);
and U580 (N_580,In_603,In_1422);
and U581 (N_581,In_104,In_2065);
or U582 (N_582,In_1172,In_1645);
or U583 (N_583,In_431,In_1708);
and U584 (N_584,In_249,In_1956);
nand U585 (N_585,In_2069,In_2529);
and U586 (N_586,In_97,In_1626);
nand U587 (N_587,In_344,In_2406);
nand U588 (N_588,In_2359,In_2703);
nor U589 (N_589,In_2598,In_475);
nor U590 (N_590,In_149,In_558);
and U591 (N_591,In_1991,In_549);
nand U592 (N_592,In_1768,In_161);
nand U593 (N_593,In_1920,In_1166);
nand U594 (N_594,In_1569,In_110);
xor U595 (N_595,In_1861,In_2435);
xnor U596 (N_596,In_55,In_2988);
or U597 (N_597,In_1552,In_2160);
nand U598 (N_598,In_1216,In_2791);
and U599 (N_599,In_343,In_1555);
or U600 (N_600,In_2829,In_2536);
or U601 (N_601,In_1298,In_2183);
xor U602 (N_602,In_1627,In_845);
xor U603 (N_603,In_112,In_1345);
nand U604 (N_604,In_2444,In_2720);
nand U605 (N_605,In_1460,In_406);
xnor U606 (N_606,In_2115,In_2403);
and U607 (N_607,In_761,In_1162);
and U608 (N_608,In_1789,In_1458);
xnor U609 (N_609,In_2906,In_2172);
nand U610 (N_610,In_2418,In_2245);
and U611 (N_611,In_1964,In_473);
nor U612 (N_612,In_2139,In_2266);
nor U613 (N_613,In_2308,In_1062);
nor U614 (N_614,In_316,In_1500);
and U615 (N_615,In_1601,In_2103);
nand U616 (N_616,In_2541,In_2683);
nand U617 (N_617,In_2934,In_648);
or U618 (N_618,In_1194,In_2097);
or U619 (N_619,In_2655,In_1089);
nand U620 (N_620,In_2579,In_692);
nand U621 (N_621,In_388,In_2358);
xnor U622 (N_622,In_857,In_797);
nand U623 (N_623,In_1400,In_2602);
nand U624 (N_624,In_485,In_2558);
xnor U625 (N_625,In_317,In_433);
nand U626 (N_626,In_2409,In_2080);
and U627 (N_627,In_2324,In_1276);
xor U628 (N_628,In_2285,In_244);
nand U629 (N_629,In_1046,In_744);
or U630 (N_630,In_1310,In_1112);
nand U631 (N_631,In_1249,In_1399);
xnor U632 (N_632,In_1333,In_1222);
or U633 (N_633,In_734,In_573);
nor U634 (N_634,In_2712,In_2233);
or U635 (N_635,In_1714,In_1677);
nor U636 (N_636,In_1488,In_2250);
and U637 (N_637,In_1757,In_268);
and U638 (N_638,In_66,In_1942);
or U639 (N_639,In_2221,In_2857);
or U640 (N_640,In_2247,In_120);
or U641 (N_641,In_2798,In_2970);
nor U642 (N_642,In_1838,In_105);
xnor U643 (N_643,In_1857,In_1439);
nand U644 (N_644,In_2596,In_1726);
or U645 (N_645,In_248,In_209);
and U646 (N_646,In_1080,In_2705);
or U647 (N_647,In_513,In_2286);
and U648 (N_648,In_1796,In_842);
nand U649 (N_649,In_614,In_178);
nand U650 (N_650,In_1197,In_2361);
or U651 (N_651,In_2088,In_2299);
nand U652 (N_652,In_2879,In_91);
or U653 (N_653,In_1332,In_2476);
nand U654 (N_654,In_2813,In_830);
and U655 (N_655,In_779,In_670);
nand U656 (N_656,In_2480,In_1629);
nor U657 (N_657,In_134,In_1513);
and U658 (N_658,In_183,In_2709);
xnor U659 (N_659,In_591,In_2612);
xnor U660 (N_660,In_733,In_2277);
nand U661 (N_661,In_2151,In_2577);
and U662 (N_662,In_80,In_386);
xnor U663 (N_663,In_960,In_340);
xnor U664 (N_664,In_2327,In_883);
nor U665 (N_665,In_1881,In_1845);
xnor U666 (N_666,In_1710,In_2458);
xnor U667 (N_667,In_1968,In_162);
and U668 (N_668,In_1745,In_1524);
and U669 (N_669,In_1541,In_2737);
or U670 (N_670,In_2540,In_1115);
xor U671 (N_671,In_2256,In_1729);
xor U672 (N_672,In_693,In_740);
nand U673 (N_673,In_1967,In_2430);
nand U674 (N_674,In_2484,In_518);
nand U675 (N_675,In_1979,In_2594);
nand U676 (N_676,In_1192,In_735);
and U677 (N_677,In_1309,In_2773);
or U678 (N_678,In_1635,In_1648);
or U679 (N_679,In_1573,In_2522);
nor U680 (N_680,In_1567,In_1498);
nor U681 (N_681,In_2332,In_1058);
nand U682 (N_682,In_2788,In_578);
or U683 (N_683,In_756,In_751);
or U684 (N_684,In_26,In_954);
nand U685 (N_685,In_2487,In_2059);
nand U686 (N_686,In_2100,In_2834);
nand U687 (N_687,In_823,In_1557);
nand U688 (N_688,In_557,In_2016);
nor U689 (N_689,In_658,In_1749);
and U690 (N_690,In_1128,In_2749);
or U691 (N_691,In_1772,In_1671);
nand U692 (N_692,In_2740,In_441);
or U693 (N_693,In_2228,In_1589);
and U694 (N_694,In_2306,In_916);
or U695 (N_695,In_342,In_2334);
or U696 (N_696,In_2352,In_2823);
or U697 (N_697,In_2251,In_560);
nor U698 (N_698,In_1053,In_824);
and U699 (N_699,In_2764,In_84);
and U700 (N_700,In_2218,In_2778);
nor U701 (N_701,In_910,In_1483);
xor U702 (N_702,In_1242,In_1505);
xnor U703 (N_703,In_1829,In_1598);
xor U704 (N_704,In_2983,In_1944);
nand U705 (N_705,In_2244,In_1807);
nand U706 (N_706,In_1378,In_958);
xor U707 (N_707,In_526,In_1933);
nor U708 (N_708,In_1832,In_1576);
xnor U709 (N_709,In_816,In_2459);
xor U710 (N_710,In_2664,In_2868);
nand U711 (N_711,In_454,In_421);
nor U712 (N_712,In_210,In_1976);
xor U713 (N_713,In_819,In_286);
and U714 (N_714,In_508,In_2804);
nor U715 (N_715,In_445,In_1639);
xnor U716 (N_716,In_1689,In_2142);
nor U717 (N_717,In_420,In_789);
nor U718 (N_718,In_1377,In_2222);
or U719 (N_719,In_2509,In_2401);
or U720 (N_720,In_488,In_1230);
or U721 (N_721,In_2551,In_1010);
xnor U722 (N_722,In_1859,In_322);
nand U723 (N_723,In_1468,In_1148);
nand U724 (N_724,In_999,In_820);
xnor U725 (N_725,In_1032,In_462);
nand U726 (N_726,In_1715,In_353);
or U727 (N_727,In_1351,In_212);
and U728 (N_728,In_2838,In_363);
and U729 (N_729,In_1231,In_1481);
and U730 (N_730,In_1369,In_1203);
nor U731 (N_731,In_2880,In_1184);
nor U732 (N_732,In_1358,In_1766);
and U733 (N_733,In_1285,In_2041);
xor U734 (N_734,In_2782,In_1641);
nor U735 (N_735,In_1988,In_283);
nor U736 (N_736,In_1376,In_1277);
or U737 (N_737,In_1836,In_2743);
nand U738 (N_738,In_568,In_2581);
or U739 (N_739,In_1280,In_1342);
xor U740 (N_740,In_1802,In_2178);
nor U741 (N_741,In_1388,In_2951);
or U742 (N_742,In_890,In_900);
and U743 (N_743,In_1926,In_1274);
or U744 (N_744,In_642,In_972);
nand U745 (N_745,In_2169,In_1409);
nor U746 (N_746,In_2196,In_2365);
nor U747 (N_747,In_490,In_412);
nor U748 (N_748,In_2817,In_1833);
nor U749 (N_749,In_1579,In_271);
or U750 (N_750,In_429,In_484);
and U751 (N_751,In_2350,In_2682);
and U752 (N_752,In_17,In_1678);
nor U753 (N_753,In_2642,In_803);
or U754 (N_754,In_1660,In_1206);
or U755 (N_755,In_1630,In_773);
xor U756 (N_756,In_1974,In_141);
nand U757 (N_757,In_2601,In_716);
nand U758 (N_758,In_0,In_1069);
nor U759 (N_759,In_1440,In_303);
nor U760 (N_760,In_2191,In_2956);
nor U761 (N_761,In_1656,In_741);
nor U762 (N_762,In_540,In_1253);
xor U763 (N_763,In_2815,In_2364);
nand U764 (N_764,In_791,In_2012);
nand U765 (N_765,In_1262,In_1849);
nand U766 (N_766,In_1266,In_1632);
xnor U767 (N_767,In_2198,In_738);
nor U768 (N_768,In_1044,In_2047);
or U769 (N_769,In_2027,In_190);
nor U770 (N_770,In_1705,In_515);
and U771 (N_771,In_536,In_1178);
nand U772 (N_772,In_963,In_1137);
nor U773 (N_773,In_1602,In_962);
or U774 (N_774,In_889,In_652);
nand U775 (N_775,In_380,In_750);
or U776 (N_776,In_2085,In_2512);
xor U777 (N_777,In_937,In_2732);
nor U778 (N_778,In_1564,In_1613);
nand U779 (N_779,In_1779,In_694);
and U780 (N_780,In_1890,In_2314);
and U781 (N_781,In_2753,In_2680);
xnor U782 (N_782,In_1427,In_953);
nor U783 (N_783,In_989,In_2807);
xor U784 (N_784,In_2186,In_2873);
and U785 (N_785,In_281,In_1842);
and U786 (N_786,In_464,In_605);
nand U787 (N_787,In_2488,In_382);
xor U788 (N_788,In_2672,In_2383);
nor U789 (N_789,In_1907,In_1685);
xor U790 (N_790,In_1348,In_1837);
nor U791 (N_791,In_2099,In_2747);
nand U792 (N_792,In_2291,In_2466);
xor U793 (N_793,In_1379,In_2074);
nor U794 (N_794,In_1300,In_1556);
and U795 (N_795,In_1609,In_1472);
or U796 (N_796,In_47,In_1054);
and U797 (N_797,In_2920,In_961);
and U798 (N_798,In_2591,In_228);
and U799 (N_799,In_1975,In_288);
xor U800 (N_800,In_1554,In_1742);
xnor U801 (N_801,In_676,In_1071);
or U802 (N_802,In_67,In_2415);
nand U803 (N_803,In_1947,In_945);
or U804 (N_804,In_2072,In_15);
nand U805 (N_805,In_1396,In_1571);
or U806 (N_806,In_621,In_103);
and U807 (N_807,In_1822,In_2402);
or U808 (N_808,In_1286,In_1611);
and U809 (N_809,In_259,In_1068);
or U810 (N_810,In_2689,In_2980);
xnor U811 (N_811,In_2223,In_1806);
or U812 (N_812,In_2611,In_533);
nor U813 (N_813,In_2297,In_1042);
and U814 (N_814,In_186,In_387);
nand U815 (N_815,In_1111,In_2260);
or U816 (N_816,In_1063,In_1718);
nor U817 (N_817,In_2288,In_364);
or U818 (N_818,In_1410,In_718);
nand U819 (N_819,In_193,In_867);
nor U820 (N_820,In_1269,In_2964);
nand U821 (N_821,In_1801,In_848);
and U822 (N_822,In_1307,In_2091);
xor U823 (N_823,In_810,In_862);
and U824 (N_824,In_2565,In_27);
xor U825 (N_825,In_2806,In_2847);
nand U826 (N_826,In_467,In_1604);
xnor U827 (N_827,In_2089,In_703);
nor U828 (N_828,In_2548,In_1824);
or U829 (N_829,In_688,In_56);
nor U830 (N_830,In_1948,In_2723);
or U831 (N_831,In_2053,In_1108);
and U832 (N_832,In_1736,In_1949);
xnor U833 (N_833,In_2269,In_2883);
nor U834 (N_834,In_1013,In_1625);
and U835 (N_835,In_189,In_2294);
or U836 (N_836,In_2491,In_581);
nand U837 (N_837,In_1241,In_2938);
nor U838 (N_838,In_164,In_2744);
and U839 (N_839,In_2953,In_2968);
nor U840 (N_840,In_662,In_1065);
or U841 (N_841,In_2129,In_2725);
and U842 (N_842,In_1892,In_95);
nand U843 (N_843,In_2171,In_2431);
xnor U844 (N_844,In_1863,In_2335);
xor U845 (N_845,In_2193,In_2716);
xor U846 (N_846,In_289,In_58);
nand U847 (N_847,In_2105,In_2054);
nor U848 (N_848,In_1365,In_438);
and U849 (N_849,In_770,In_1570);
nand U850 (N_850,In_1506,In_913);
nor U851 (N_851,In_2685,In_2392);
nand U852 (N_852,In_2093,In_1393);
and U853 (N_853,In_2981,In_1402);
and U854 (N_854,In_2979,In_1914);
nand U855 (N_855,In_1282,In_1971);
nor U856 (N_856,In_2199,In_308);
nand U857 (N_857,In_997,In_1917);
or U858 (N_858,In_1493,In_1160);
or U859 (N_859,In_597,In_2421);
nand U860 (N_860,In_2043,In_1341);
xnor U861 (N_861,In_215,In_1674);
nand U862 (N_862,In_1698,In_2131);
or U863 (N_863,In_2634,In_113);
xnor U864 (N_864,In_439,In_2396);
nand U865 (N_865,In_71,In_2510);
xnor U866 (N_866,In_448,In_631);
xnor U867 (N_867,In_175,In_227);
or U868 (N_868,In_483,In_2426);
nor U869 (N_869,In_1299,In_1117);
nand U870 (N_870,In_1205,In_2104);
nand U871 (N_871,In_292,In_1357);
or U872 (N_872,In_2843,In_205);
nand U873 (N_873,In_860,In_2490);
nand U874 (N_874,In_143,In_1534);
xor U875 (N_875,In_2784,In_1529);
nand U876 (N_876,In_1208,In_1686);
and U877 (N_877,In_1754,In_1403);
and U878 (N_878,In_1091,In_2135);
and U879 (N_879,In_2498,In_2745);
nand U880 (N_880,In_2947,In_2994);
and U881 (N_881,In_935,In_2333);
nor U882 (N_882,In_2293,In_139);
xnor U883 (N_883,In_598,In_2860);
and U884 (N_884,In_2376,In_115);
nand U885 (N_885,In_2441,In_2646);
or U886 (N_886,In_1334,In_1618);
or U887 (N_887,In_551,In_128);
and U888 (N_888,In_20,In_1296);
xor U889 (N_889,In_727,In_1170);
xor U890 (N_890,In_2208,In_1433);
xnor U891 (N_891,In_145,In_2414);
xnor U892 (N_892,In_179,In_2668);
xor U893 (N_893,In_94,In_586);
nor U894 (N_894,In_1387,In_1521);
nand U895 (N_895,In_1819,In_1000);
nor U896 (N_896,In_1157,In_632);
or U897 (N_897,In_1817,In_2992);
or U898 (N_898,In_971,In_1937);
and U899 (N_899,In_2640,In_2681);
nor U900 (N_900,In_238,In_1047);
and U901 (N_901,In_2176,In_79);
or U902 (N_902,In_489,In_2182);
nand U903 (N_903,In_1595,In_1510);
or U904 (N_904,In_2687,In_185);
or U905 (N_905,In_1006,In_2408);
and U906 (N_906,In_182,In_550);
nand U907 (N_907,In_1164,In_1551);
and U908 (N_908,In_1781,In_351);
or U909 (N_909,In_2917,In_2159);
nand U910 (N_910,In_1430,In_2777);
xnor U911 (N_911,In_2647,In_478);
nor U912 (N_912,In_2128,In_68);
and U913 (N_913,In_2106,In_284);
nand U914 (N_914,In_984,In_1278);
and U915 (N_915,In_2434,In_2626);
or U916 (N_916,In_2340,In_1349);
and U917 (N_917,In_2432,In_1874);
and U918 (N_918,In_471,In_401);
nand U919 (N_919,In_572,In_24);
nor U920 (N_920,In_968,In_1728);
nand U921 (N_921,In_2850,In_2805);
or U922 (N_922,In_1813,In_613);
nand U923 (N_923,In_1129,In_2506);
or U924 (N_924,In_1841,In_2960);
xor U925 (N_925,In_2665,In_604);
nand U926 (N_926,In_1840,In_2095);
nor U927 (N_927,In_1356,In_2268);
and U928 (N_928,In_521,In_742);
xnor U929 (N_929,In_666,In_1764);
nand U930 (N_930,In_1079,In_2230);
and U931 (N_931,In_1608,In_1637);
nand U932 (N_932,In_2803,In_675);
xnor U933 (N_933,In_1321,In_2627);
or U934 (N_934,In_981,In_1455);
nor U935 (N_935,In_698,In_1643);
nand U936 (N_936,In_2578,In_690);
xor U937 (N_937,In_1514,In_2885);
xor U938 (N_938,In_1515,In_1372);
and U939 (N_939,In_1823,In_847);
nand U940 (N_940,In_732,In_792);
and U941 (N_941,In_2076,In_2989);
nand U942 (N_942,In_2071,In_2347);
nor U943 (N_943,In_385,In_315);
or U944 (N_944,In_394,In_426);
nand U945 (N_945,In_2140,In_1417);
xnor U946 (N_946,In_52,In_1454);
xor U947 (N_947,In_626,In_1654);
nor U948 (N_948,In_1921,In_1457);
xor U949 (N_949,In_2511,In_2660);
nor U950 (N_950,In_636,In_2925);
xor U951 (N_951,In_1143,In_1145);
and U952 (N_952,In_2696,In_2946);
and U953 (N_953,In_2165,In_2258);
or U954 (N_954,In_130,In_510);
nand U955 (N_955,In_169,In_879);
nand U956 (N_956,In_2583,In_2942);
xnor U957 (N_957,In_54,In_2282);
nor U958 (N_958,In_224,In_2166);
nor U959 (N_959,In_1646,In_413);
xnor U960 (N_960,In_48,In_2032);
or U961 (N_961,In_1212,In_1220);
nor U962 (N_962,In_2127,In_858);
xor U963 (N_963,In_477,In_1966);
xnor U964 (N_964,In_1463,In_794);
and U965 (N_965,In_832,In_442);
nor U966 (N_966,In_2700,In_1924);
and U967 (N_967,In_2867,In_1782);
xnor U968 (N_968,In_964,In_245);
nand U969 (N_969,In_2044,In_405);
nand U970 (N_970,In_2475,In_2891);
nand U971 (N_971,In_2212,In_326);
nand U972 (N_972,In_1072,In_14);
nand U973 (N_973,In_2549,In_1810);
and U974 (N_974,In_1219,In_1951);
nand U975 (N_975,In_673,In_985);
nor U976 (N_976,In_1652,In_434);
nand U977 (N_977,In_975,In_1297);
or U978 (N_978,In_1536,In_2318);
or U979 (N_979,In_2175,In_1843);
nor U980 (N_980,In_101,In_2811);
and U981 (N_981,In_123,In_647);
or U982 (N_982,In_2081,In_617);
or U983 (N_983,In_2770,In_2108);
nor U984 (N_984,In_2789,In_1519);
and U985 (N_985,In_2489,In_367);
and U986 (N_986,In_1452,In_2336);
nand U987 (N_987,In_1331,In_476);
or U988 (N_988,In_1031,In_944);
nor U989 (N_989,In_2060,In_40);
xor U990 (N_990,In_2461,In_2467);
and U991 (N_991,In_1811,In_1070);
nor U992 (N_992,In_349,In_2704);
or U993 (N_993,In_1147,In_745);
or U994 (N_994,In_878,In_3);
xnor U995 (N_995,In_2007,In_2780);
xnor U996 (N_996,In_685,In_410);
and U997 (N_997,In_1263,In_1305);
or U998 (N_998,In_1511,In_118);
xor U999 (N_999,In_2064,In_2023);
or U1000 (N_1000,In_2711,In_348);
xnor U1001 (N_1001,In_2033,In_2442);
or U1002 (N_1002,In_2058,In_177);
or U1003 (N_1003,In_2037,In_2948);
xnor U1004 (N_1004,In_1835,In_774);
nand U1005 (N_1005,In_805,In_638);
nand U1006 (N_1006,In_2957,In_924);
xor U1007 (N_1007,In_2772,In_415);
and U1008 (N_1008,In_156,In_1723);
and U1009 (N_1009,In_1193,In_2181);
nand U1010 (N_1010,In_377,In_1033);
nor U1011 (N_1011,In_1730,In_2909);
or U1012 (N_1012,In_1727,In_701);
or U1013 (N_1013,In_1737,In_85);
nor U1014 (N_1014,In_1717,In_1429);
and U1015 (N_1015,In_901,In_1248);
nand U1016 (N_1016,In_2049,In_338);
or U1017 (N_1017,In_918,In_2524);
xor U1018 (N_1018,In_1200,In_506);
nor U1019 (N_1019,In_542,In_306);
or U1020 (N_1020,In_2837,In_2316);
nor U1021 (N_1021,In_1084,In_450);
xor U1022 (N_1022,In_1325,In_2372);
and U1023 (N_1023,In_1326,In_2528);
or U1024 (N_1024,In_1597,In_1562);
nand U1025 (N_1025,In_144,In_863);
and U1026 (N_1026,In_1740,In_1005);
xor U1027 (N_1027,In_1592,In_2610);
and U1028 (N_1028,In_905,In_2464);
and U1029 (N_1029,In_2349,In_906);
and U1030 (N_1030,In_2574,In_1312);
nor U1031 (N_1031,In_1532,In_2399);
or U1032 (N_1032,In_1898,In_616);
and U1033 (N_1033,In_1185,In_1057);
nor U1034 (N_1034,In_486,In_76);
and U1035 (N_1035,In_2276,In_880);
nor U1036 (N_1036,In_714,In_1622);
nand U1037 (N_1037,In_1527,In_2473);
or U1038 (N_1038,In_216,In_305);
xnor U1039 (N_1039,In_2305,In_2328);
nand U1040 (N_1040,In_341,In_2945);
xor U1041 (N_1041,In_755,In_2384);
xor U1042 (N_1042,In_870,In_1973);
or U1043 (N_1043,In_1545,In_492);
or U1044 (N_1044,In_1453,In_2107);
xor U1045 (N_1045,In_199,In_713);
or U1046 (N_1046,In_1915,In_1061);
nand U1047 (N_1047,In_1167,In_977);
or U1048 (N_1048,In_2398,In_133);
xor U1049 (N_1049,In_912,In_2955);
or U1050 (N_1050,In_1258,In_2300);
nor U1051 (N_1051,In_514,In_2356);
nor U1052 (N_1052,In_1528,In_2542);
nor U1053 (N_1053,In_2257,In_1461);
nor U1054 (N_1054,In_1471,In_466);
or U1055 (N_1055,In_2111,In_1865);
nand U1056 (N_1056,In_804,In_1932);
nor U1057 (N_1057,In_623,In_424);
and U1058 (N_1058,In_2800,In_1679);
nand U1059 (N_1059,In_1478,In_994);
nor U1060 (N_1060,In_2694,In_470);
nand U1061 (N_1061,In_1522,In_1831);
or U1062 (N_1062,In_1110,In_806);
or U1063 (N_1063,In_1275,In_1512);
xor U1064 (N_1064,In_2765,In_1271);
or U1065 (N_1065,In_1158,In_1480);
or U1066 (N_1066,In_1922,In_1049);
xnor U1067 (N_1067,In_1328,In_294);
nand U1068 (N_1068,In_2216,In_1748);
and U1069 (N_1069,In_1386,In_2715);
or U1070 (N_1070,In_813,In_44);
nor U1071 (N_1071,In_2307,In_1561);
xnor U1072 (N_1072,In_749,In_1124);
and U1073 (N_1073,In_1421,In_334);
xor U1074 (N_1074,In_864,In_1972);
nor U1075 (N_1075,In_2133,In_775);
or U1076 (N_1076,In_2810,In_1261);
nand U1077 (N_1077,In_537,In_453);
and U1078 (N_1078,In_1687,In_2009);
xor U1079 (N_1079,In_30,In_532);
xor U1080 (N_1080,In_2639,In_1752);
nor U1081 (N_1081,In_799,In_875);
xnor U1082 (N_1082,In_87,In_2035);
and U1083 (N_1083,In_983,In_1186);
nor U1084 (N_1084,In_2492,In_930);
or U1085 (N_1085,In_1475,In_1329);
xnor U1086 (N_1086,In_2075,In_2068);
xnor U1087 (N_1087,In_697,In_976);
nand U1088 (N_1088,In_2201,In_2746);
nand U1089 (N_1089,In_2997,In_664);
xor U1090 (N_1090,In_2759,In_1712);
or U1091 (N_1091,In_1787,In_2472);
or U1092 (N_1092,In_2927,In_2486);
nor U1093 (N_1093,In_859,In_77);
and U1094 (N_1094,In_2622,In_147);
xor U1095 (N_1095,In_2904,In_255);
nor U1096 (N_1096,In_2758,In_831);
and U1097 (N_1097,In_2671,In_2036);
nor U1098 (N_1098,In_119,In_1940);
and U1099 (N_1099,In_2722,In_2101);
and U1100 (N_1100,In_2614,In_2312);
and U1101 (N_1101,In_1734,In_318);
nor U1102 (N_1102,In_291,In_1868);
nor U1103 (N_1103,In_2270,In_329);
and U1104 (N_1104,In_1075,In_611);
xor U1105 (N_1105,In_737,In_768);
and U1106 (N_1106,In_2261,In_2252);
xor U1107 (N_1107,In_168,In_2698);
nand U1108 (N_1108,In_546,In_2226);
xnor U1109 (N_1109,In_1029,In_2351);
and U1110 (N_1110,In_2620,In_2284);
and U1111 (N_1111,In_1699,In_1469);
xnor U1112 (N_1112,In_427,In_2595);
xor U1113 (N_1113,In_1103,In_1913);
nor U1114 (N_1114,In_1912,In_2272);
nor U1115 (N_1115,In_2011,In_1199);
nor U1116 (N_1116,In_969,In_846);
and U1117 (N_1117,In_2775,In_2941);
and U1118 (N_1118,In_1997,In_570);
nor U1119 (N_1119,In_1238,In_1664);
xnor U1120 (N_1120,In_226,In_2766);
or U1121 (N_1121,In_2570,In_500);
xor U1122 (N_1122,In_451,In_314);
or U1123 (N_1123,In_2918,In_276);
and U1124 (N_1124,In_2808,In_108);
nand U1125 (N_1125,In_2547,In_667);
and U1126 (N_1126,In_2289,In_814);
xnor U1127 (N_1127,In_1706,In_1596);
xnor U1128 (N_1128,In_940,In_159);
and U1129 (N_1129,In_2821,In_2149);
and U1130 (N_1130,In_2070,In_1236);
xnor U1131 (N_1131,In_2855,In_1450);
and U1132 (N_1132,In_1462,In_2025);
or U1133 (N_1133,In_1279,In_1362);
nor U1134 (N_1134,In_2890,In_643);
nor U1135 (N_1135,In_72,In_440);
and U1136 (N_1136,In_1289,In_1138);
and U1137 (N_1137,In_833,In_2637);
and U1138 (N_1138,In_1020,In_93);
nor U1139 (N_1139,In_327,In_1517);
xor U1140 (N_1140,In_151,In_102);
xor U1141 (N_1141,In_2795,In_157);
and U1142 (N_1142,In_1174,In_787);
nor U1143 (N_1143,In_38,In_1073);
nand U1144 (N_1144,In_851,In_1987);
nand U1145 (N_1145,In_1048,In_430);
nand U1146 (N_1146,In_389,In_523);
nand U1147 (N_1147,In_1847,In_1456);
and U1148 (N_1148,In_2996,In_547);
nor U1149 (N_1149,In_724,In_2045);
xor U1150 (N_1150,In_637,In_825);
and U1151 (N_1151,In_200,In_170);
nand U1152 (N_1152,In_1459,In_1094);
nor U1153 (N_1153,In_2255,In_986);
and U1154 (N_1154,In_310,In_282);
nor U1155 (N_1155,In_298,In_1762);
nor U1156 (N_1156,In_1363,In_1821);
xor U1157 (N_1157,In_2899,In_1786);
or U1158 (N_1158,In_2707,In_904);
xor U1159 (N_1159,In_1228,In_2535);
nor U1160 (N_1160,In_2125,In_459);
nor U1161 (N_1161,In_587,In_384);
nor U1162 (N_1162,In_1337,In_1256);
nand U1163 (N_1163,In_1007,In_1984);
nor U1164 (N_1164,In_1878,In_1109);
or U1165 (N_1165,In_2456,In_2098);
nand U1166 (N_1166,In_2259,In_2982);
and U1167 (N_1167,In_588,In_1820);
xnor U1168 (N_1168,In_2342,In_1518);
nand U1169 (N_1169,In_1190,In_2940);
and U1170 (N_1170,In_1930,In_630);
nand U1171 (N_1171,In_2978,In_1335);
and U1172 (N_1172,In_1673,In_1853);
xnor U1173 (N_1173,In_2986,In_828);
or U1174 (N_1174,In_1816,In_2991);
nor U1175 (N_1175,In_2702,In_651);
nor U1176 (N_1176,In_1902,In_1665);
or U1177 (N_1177,In_2143,In_2657);
xor U1178 (N_1178,In_1211,In_1887);
nand U1179 (N_1179,In_915,In_709);
or U1180 (N_1180,In_1850,In_2545);
and U1181 (N_1181,In_1392,In_2552);
or U1182 (N_1182,In_635,In_763);
nand U1183 (N_1183,In_1879,In_2731);
xnor U1184 (N_1184,In_1302,In_1818);
or U1185 (N_1185,In_2714,In_2117);
nand U1186 (N_1186,In_1830,In_646);
or U1187 (N_1187,In_2760,In_2937);
xnor U1188 (N_1188,In_23,In_2164);
or U1189 (N_1189,In_213,In_948);
nor U1190 (N_1190,In_1880,In_1965);
nor U1191 (N_1191,In_2249,In_689);
and U1192 (N_1192,In_1825,In_1030);
xor U1193 (N_1193,In_371,In_683);
nand U1194 (N_1194,In_253,In_1104);
or U1195 (N_1195,In_2756,In_41);
and U1196 (N_1196,In_2423,In_1155);
nor U1197 (N_1197,In_1954,In_2427);
and U1198 (N_1198,In_2871,In_2004);
nor U1199 (N_1199,In_1684,In_2518);
nand U1200 (N_1200,In_535,In_2919);
xnor U1201 (N_1201,In_2587,In_594);
xnor U1202 (N_1202,In_1292,In_1492);
nor U1203 (N_1203,In_1017,In_425);
nand U1204 (N_1204,In_1196,In_163);
xnor U1205 (N_1205,In_2686,In_2017);
nor U1206 (N_1206,In_1411,In_2507);
nand U1207 (N_1207,In_965,In_543);
and U1208 (N_1208,In_2767,In_874);
nand U1209 (N_1209,In_2576,In_357);
nor U1210 (N_1210,In_839,In_2972);
xnor U1211 (N_1211,In_1872,In_2719);
xnor U1212 (N_1212,In_2055,In_2187);
xnor U1213 (N_1213,In_375,In_2438);
nand U1214 (N_1214,In_2130,In_225);
xor U1215 (N_1215,In_2197,In_767);
nand U1216 (N_1216,In_2462,In_511);
nor U1217 (N_1217,In_1581,In_2213);
and U1218 (N_1218,In_2217,In_2666);
nand U1219 (N_1219,In_1002,In_886);
nand U1220 (N_1220,In_1735,In_2993);
nor U1221 (N_1221,In_624,In_1578);
or U1222 (N_1222,In_545,In_19);
nor U1223 (N_1223,In_705,In_1444);
nor U1224 (N_1224,In_1544,In_1041);
xnor U1225 (N_1225,In_397,In_1938);
and U1226 (N_1226,In_78,In_88);
nor U1227 (N_1227,In_1955,In_60);
xnor U1228 (N_1228,In_6,In_2735);
xnor U1229 (N_1229,In_2998,In_1624);
or U1230 (N_1230,In_2470,In_1489);
nor U1231 (N_1231,In_1037,In_1998);
nand U1232 (N_1232,In_1911,In_893);
xor U1233 (N_1233,In_610,In_320);
or U1234 (N_1234,In_369,In_345);
xor U1235 (N_1235,In_1503,In_1131);
or U1236 (N_1236,In_197,In_684);
or U1237 (N_1237,In_2633,In_1502);
nor U1238 (N_1238,In_541,In_955);
or U1239 (N_1239,In_852,In_699);
and U1240 (N_1240,In_2419,In_1666);
xor U1241 (N_1241,In_579,In_2742);
and U1242 (N_1242,In_2566,In_897);
nand U1243 (N_1243,In_1895,In_2827);
nor U1244 (N_1244,In_1051,In_2663);
nor U1245 (N_1245,In_1338,In_242);
nand U1246 (N_1246,In_929,In_973);
and U1247 (N_1247,In_1217,In_920);
nand U1248 (N_1248,In_319,In_650);
nand U1249 (N_1249,In_2453,In_2407);
nand U1250 (N_1250,In_158,In_2325);
nand U1251 (N_1251,In_457,In_1169);
nand U1252 (N_1252,In_2436,In_1023);
nor U1253 (N_1253,In_1213,In_2999);
nor U1254 (N_1254,In_1908,In_2950);
and U1255 (N_1255,In_1765,In_2605);
and U1256 (N_1256,In_1690,In_2220);
or U1257 (N_1257,In_1566,In_1177);
xnor U1258 (N_1258,In_2329,In_1644);
nand U1259 (N_1259,In_1896,In_2560);
or U1260 (N_1260,In_1191,In_2189);
nor U1261 (N_1261,In_1928,In_131);
or U1262 (N_1262,In_1431,In_1484);
or U1263 (N_1263,In_2613,In_966);
nand U1264 (N_1264,In_1371,In_2900);
nor U1265 (N_1265,In_566,In_2553);
nor U1266 (N_1266,In_2416,In_1649);
nand U1267 (N_1267,In_674,In_1293);
xor U1268 (N_1268,In_381,In_2826);
or U1269 (N_1269,In_2413,In_2884);
xnor U1270 (N_1270,In_2240,In_1476);
nor U1271 (N_1271,In_2063,In_1346);
xnor U1272 (N_1272,In_311,In_982);
nand U1273 (N_1273,In_1252,In_686);
and U1274 (N_1274,In_729,In_383);
and U1275 (N_1275,In_1405,In_2454);
and U1276 (N_1276,In_361,In_2497);
nand U1277 (N_1277,In_2739,In_2292);
xnor U1278 (N_1278,In_423,In_299);
and U1279 (N_1279,In_1738,In_2015);
or U1280 (N_1280,In_2585,In_800);
xor U1281 (N_1281,In_575,In_35);
nand U1282 (N_1282,In_2641,In_293);
xnor U1283 (N_1283,In_2471,In_746);
and U1284 (N_1284,In_1676,In_1035);
and U1285 (N_1285,In_1008,In_2674);
xnor U1286 (N_1286,In_2145,In_1784);
nand U1287 (N_1287,In_780,In_1288);
and U1288 (N_1288,In_1631,In_1546);
xor U1289 (N_1289,In_2859,In_1077);
nand U1290 (N_1290,In_2429,In_2973);
nor U1291 (N_1291,In_1473,In_1733);
and U1292 (N_1292,In_895,In_2184);
nand U1293 (N_1293,In_1620,In_260);
and U1294 (N_1294,In_22,In_2916);
nand U1295 (N_1295,In_827,In_1663);
and U1296 (N_1296,In_625,In_1970);
nor U1297 (N_1297,In_841,In_2658);
or U1298 (N_1298,In_2656,In_524);
nand U1299 (N_1299,In_1255,In_2600);
and U1300 (N_1300,In_1438,In_1121);
or U1301 (N_1301,In_2569,In_1587);
xnor U1302 (N_1302,In_372,In_2368);
xnor U1303 (N_1303,In_2022,In_2966);
xnor U1304 (N_1304,In_2439,In_2629);
and U1305 (N_1305,In_2448,In_2211);
nand U1306 (N_1306,In_2785,In_1854);
or U1307 (N_1307,In_2136,In_932);
xor U1308 (N_1308,In_2822,In_1368);
nand U1309 (N_1309,In_2932,In_818);
nor U1310 (N_1310,In_482,In_1322);
or U1311 (N_1311,In_240,In_1539);
nor U1312 (N_1312,In_1168,In_1374);
nor U1313 (N_1313,In_2298,In_2623);
nand U1314 (N_1314,In_2923,In_2799);
nor U1315 (N_1315,In_2974,In_1886);
xor U1316 (N_1316,In_1316,In_1272);
nor U1317 (N_1317,In_1560,In_2607);
xor U1318 (N_1318,In_1941,In_444);
nand U1319 (N_1319,In_680,In_2875);
xor U1320 (N_1320,In_2952,In_1187);
xor U1321 (N_1321,In_771,In_796);
nand U1322 (N_1322,In_1856,In_719);
or U1323 (N_1323,In_757,In_1397);
xnor U1324 (N_1324,In_335,In_2835);
or U1325 (N_1325,In_882,In_2930);
nand U1326 (N_1326,In_1993,In_1777);
nor U1327 (N_1327,In_1894,In_2832);
nand U1328 (N_1328,In_350,In_2812);
or U1329 (N_1329,In_691,In_2317);
xor U1330 (N_1330,In_2546,In_517);
xor U1331 (N_1331,In_559,In_399);
and U1332 (N_1332,In_2161,In_1);
or U1333 (N_1333,In_443,In_136);
nor U1334 (N_1334,In_1223,In_2854);
and U1335 (N_1335,In_2102,In_1852);
xor U1336 (N_1336,In_1448,In_659);
xor U1337 (N_1337,In_1780,In_247);
xor U1338 (N_1338,In_2188,In_822);
or U1339 (N_1339,In_783,In_793);
xor U1340 (N_1340,In_1855,In_2706);
and U1341 (N_1341,In_1795,In_1380);
nand U1342 (N_1342,In_2915,In_2155);
nor U1343 (N_1343,In_39,In_2976);
and U1344 (N_1344,In_301,In_2000);
xor U1345 (N_1345,In_907,In_358);
or U1346 (N_1346,In_2573,In_2677);
xor U1347 (N_1347,In_1952,In_352);
nor U1348 (N_1348,In_196,In_2961);
and U1349 (N_1349,In_2440,In_1330);
nor U1350 (N_1350,In_1259,In_1240);
and U1351 (N_1351,In_608,In_2234);
xor U1352 (N_1352,In_1634,In_2303);
xnor U1353 (N_1353,In_753,In_2200);
or U1354 (N_1354,In_1038,In_2734);
and U1355 (N_1355,In_29,In_2673);
xor U1356 (N_1356,In_2763,In_2038);
and U1357 (N_1357,In_1179,In_2395);
xor U1358 (N_1358,In_654,In_1931);
or U1359 (N_1359,In_198,In_925);
nand U1360 (N_1360,In_2243,In_1709);
and U1361 (N_1361,In_1547,In_2451);
and U1362 (N_1362,In_1022,In_1590);
and U1363 (N_1363,In_1929,In_2344);
xor U1364 (N_1364,In_339,In_2215);
nand U1365 (N_1365,In_2892,In_2669);
nand U1366 (N_1366,In_2457,In_62);
or U1367 (N_1367,In_1691,In_505);
nor U1368 (N_1368,In_1352,In_2177);
or U1369 (N_1369,In_1215,In_1449);
xnor U1370 (N_1370,In_1354,In_229);
xor U1371 (N_1371,In_834,In_1491);
nand U1372 (N_1372,In_2878,In_257);
or U1373 (N_1373,In_1783,In_1414);
nand U1374 (N_1374,In_1657,In_501);
nand U1375 (N_1375,In_2520,In_2465);
nor U1376 (N_1376,In_2477,In_4);
nand U1377 (N_1377,In_1412,In_2375);
or U1378 (N_1378,In_1425,In_1778);
nand U1379 (N_1379,In_1769,In_590);
xor U1380 (N_1380,In_2852,In_304);
xnor U1381 (N_1381,In_109,In_2888);
nor U1382 (N_1382,In_881,In_682);
and U1383 (N_1383,In_172,In_2400);
nor U1384 (N_1384,In_2644,In_1146);
and U1385 (N_1385,In_2628,In_208);
or U1386 (N_1386,In_2802,In_241);
nor U1387 (N_1387,In_2006,In_1636);
nand U1388 (N_1388,In_2515,In_1659);
nor U1389 (N_1389,In_1763,In_1612);
or U1390 (N_1390,In_2021,In_1426);
nand U1391 (N_1391,In_2057,In_1287);
nor U1392 (N_1392,In_736,In_1638);
and U1393 (N_1393,In_1306,In_1210);
nor U1394 (N_1394,In_950,In_332);
or U1395 (N_1395,In_1418,In_2167);
xor U1396 (N_1396,In_181,In_1980);
nand U1397 (N_1397,In_221,In_2568);
and U1398 (N_1398,In_885,In_2797);
and U1399 (N_1399,In_1800,In_395);
and U1400 (N_1400,In_379,In_2363);
nor U1401 (N_1401,In_1052,In_1081);
or U1402 (N_1402,In_2985,In_2263);
and U1403 (N_1403,In_362,In_2397);
and U1404 (N_1404,In_153,In_2073);
nand U1405 (N_1405,In_607,In_1773);
or U1406 (N_1406,In_2902,In_1161);
xnor U1407 (N_1407,In_373,In_1901);
xor U1408 (N_1408,In_1101,In_2519);
xor U1409 (N_1409,In_323,In_2898);
nand U1410 (N_1410,In_1672,In_599);
nor U1411 (N_1411,In_1655,In_1713);
nand U1412 (N_1412,In_577,In_902);
nand U1413 (N_1413,In_2886,In_2728);
and U1414 (N_1414,In_106,In_258);
xnor U1415 (N_1415,In_2592,In_2907);
nor U1416 (N_1416,In_2903,In_1935);
nand U1417 (N_1417,In_777,In_2774);
nand U1418 (N_1418,In_1195,In_223);
or U1419 (N_1419,In_2463,In_1549);
xnor U1420 (N_1420,In_1603,In_2124);
nand U1421 (N_1421,In_2446,In_1774);
or U1422 (N_1422,In_1701,In_712);
and U1423 (N_1423,In_1098,In_801);
nor U1424 (N_1424,In_1495,In_1903);
xor U1425 (N_1425,In_456,In_1118);
nand U1426 (N_1426,In_512,In_1265);
nor U1427 (N_1427,In_1141,In_279);
and U1428 (N_1428,In_2194,In_2265);
nor U1429 (N_1429,In_1159,In_393);
nand U1430 (N_1430,In_435,In_174);
nor U1431 (N_1431,In_928,In_135);
nand U1432 (N_1432,In_888,In_2424);
nand U1433 (N_1433,In_414,In_1662);
nor U1434 (N_1434,In_784,In_455);
xor U1435 (N_1435,In_499,In_589);
nand U1436 (N_1436,In_1114,In_2122);
and U1437 (N_1437,In_2692,In_1572);
nand U1438 (N_1438,In_2018,In_336);
or U1439 (N_1439,In_1707,In_539);
and U1440 (N_1440,In_502,In_1594);
nand U1441 (N_1441,In_1563,In_2846);
and U1442 (N_1442,In_600,In_640);
nand U1443 (N_1443,In_493,In_1437);
or U1444 (N_1444,In_1621,In_2505);
xor U1445 (N_1445,In_2624,In_788);
nor U1446 (N_1446,In_194,In_390);
and U1447 (N_1447,In_978,In_266);
and U1448 (N_1448,In_1668,In_1640);
xor U1449 (N_1449,In_50,In_2433);
nor U1450 (N_1450,In_2086,In_1526);
nor U1451 (N_1451,In_829,In_641);
nor U1452 (N_1452,In_2118,In_217);
nor U1453 (N_1453,In_1704,In_2718);
xnor U1454 (N_1454,In_1015,In_2028);
nand U1455 (N_1455,In_2567,In_2539);
xor U1456 (N_1456,In_270,In_1558);
xnor U1457 (N_1457,In_356,In_941);
nand U1458 (N_1458,In_849,In_42);
xnor U1459 (N_1459,In_1173,In_2862);
nor U1460 (N_1460,In_346,In_49);
or U1461 (N_1461,In_2020,In_1651);
and U1462 (N_1462,In_1233,In_2848);
nand U1463 (N_1463,In_1009,In_428);
nand U1464 (N_1464,In_2482,In_580);
nand U1465 (N_1465,In_2428,In_220);
nand U1466 (N_1466,In_1043,In_1744);
and U1467 (N_1467,In_1151,In_933);
xnor U1468 (N_1468,In_418,In_747);
nor U1469 (N_1469,In_2241,In_995);
and U1470 (N_1470,In_1283,In_555);
and U1471 (N_1471,In_2381,In_2949);
nand U1472 (N_1472,In_254,In_671);
or U1473 (N_1473,In_1207,In_2905);
nand U1474 (N_1474,In_328,In_2345);
and U1475 (N_1475,In_2173,In_2975);
and U1476 (N_1476,In_1082,In_1650);
nor U1477 (N_1477,In_1295,In_1420);
xnor U1478 (N_1478,In_1183,In_2185);
or U1479 (N_1479,In_2026,In_2264);
xnor U1480 (N_1480,In_2831,In_211);
xor U1481 (N_1481,In_218,In_1900);
xor U1482 (N_1482,In_1059,In_934);
nor U1483 (N_1483,In_1130,In_2123);
nand U1484 (N_1484,In_1805,In_90);
or U1485 (N_1485,In_2279,In_2833);
xor U1486 (N_1486,In_2348,In_1719);
xor U1487 (N_1487,In_2281,In_844);
nand U1488 (N_1488,In_1909,In_2969);
nor U1489 (N_1489,In_2730,In_840);
and U1490 (N_1490,In_2531,In_422);
nor U1491 (N_1491,In_9,In_1803);
and U1492 (N_1492,In_951,In_2741);
or U1493 (N_1493,In_2754,In_2295);
nor U1494 (N_1494,In_1950,In_408);
or U1495 (N_1495,In_2853,In_107);
xor U1496 (N_1496,In_2849,In_2109);
nand U1497 (N_1497,In_1120,In_593);
nor U1498 (N_1498,In_407,In_649);
nor U1499 (N_1499,In_2225,In_530);
nor U1500 (N_1500,In_933,In_2511);
xnor U1501 (N_1501,In_2836,In_2148);
nor U1502 (N_1502,In_2541,In_419);
nor U1503 (N_1503,In_564,In_188);
and U1504 (N_1504,In_1822,In_2224);
and U1505 (N_1505,In_1656,In_555);
nand U1506 (N_1506,In_158,In_938);
or U1507 (N_1507,In_442,In_2648);
and U1508 (N_1508,In_1462,In_527);
and U1509 (N_1509,In_2586,In_39);
xnor U1510 (N_1510,In_1036,In_1735);
xor U1511 (N_1511,In_1301,In_2302);
or U1512 (N_1512,In_1668,In_1430);
xnor U1513 (N_1513,In_1734,In_506);
and U1514 (N_1514,In_1499,In_2766);
and U1515 (N_1515,In_2829,In_503);
xor U1516 (N_1516,In_2868,In_1585);
xnor U1517 (N_1517,In_101,In_2422);
nor U1518 (N_1518,In_575,In_1385);
xnor U1519 (N_1519,In_1449,In_1878);
nor U1520 (N_1520,In_1017,In_2329);
nand U1521 (N_1521,In_1661,In_1459);
nand U1522 (N_1522,In_2006,In_1416);
xor U1523 (N_1523,In_2596,In_752);
xor U1524 (N_1524,In_1125,In_2836);
nand U1525 (N_1525,In_2399,In_676);
or U1526 (N_1526,In_2059,In_1593);
or U1527 (N_1527,In_2501,In_1710);
nor U1528 (N_1528,In_2241,In_2348);
xor U1529 (N_1529,In_1283,In_1892);
and U1530 (N_1530,In_2657,In_1296);
and U1531 (N_1531,In_2070,In_1168);
xor U1532 (N_1532,In_2129,In_1071);
nor U1533 (N_1533,In_1083,In_1697);
or U1534 (N_1534,In_1054,In_2250);
and U1535 (N_1535,In_2249,In_1603);
xnor U1536 (N_1536,In_494,In_2556);
and U1537 (N_1537,In_619,In_2299);
nor U1538 (N_1538,In_1647,In_2814);
nand U1539 (N_1539,In_828,In_2226);
and U1540 (N_1540,In_2728,In_1980);
nand U1541 (N_1541,In_2951,In_946);
or U1542 (N_1542,In_2541,In_835);
or U1543 (N_1543,In_2157,In_1852);
xor U1544 (N_1544,In_1943,In_2267);
and U1545 (N_1545,In_2804,In_1529);
nor U1546 (N_1546,In_1893,In_1587);
xor U1547 (N_1547,In_2314,In_2600);
xnor U1548 (N_1548,In_531,In_1579);
nor U1549 (N_1549,In_2508,In_747);
xor U1550 (N_1550,In_2421,In_1757);
and U1551 (N_1551,In_655,In_528);
nor U1552 (N_1552,In_1320,In_1659);
nand U1553 (N_1553,In_2588,In_671);
xnor U1554 (N_1554,In_1897,In_2103);
nor U1555 (N_1555,In_1575,In_452);
and U1556 (N_1556,In_308,In_1749);
and U1557 (N_1557,In_252,In_1821);
xor U1558 (N_1558,In_2032,In_1915);
nor U1559 (N_1559,In_2571,In_2784);
nand U1560 (N_1560,In_1917,In_878);
or U1561 (N_1561,In_972,In_1726);
nor U1562 (N_1562,In_1364,In_2168);
nand U1563 (N_1563,In_1723,In_243);
and U1564 (N_1564,In_2062,In_1951);
xnor U1565 (N_1565,In_2513,In_1554);
nand U1566 (N_1566,In_2056,In_795);
or U1567 (N_1567,In_2346,In_107);
nand U1568 (N_1568,In_1988,In_1172);
or U1569 (N_1569,In_1968,In_1936);
and U1570 (N_1570,In_1996,In_2189);
and U1571 (N_1571,In_2926,In_2075);
nand U1572 (N_1572,In_501,In_723);
xor U1573 (N_1573,In_509,In_2184);
or U1574 (N_1574,In_510,In_692);
xnor U1575 (N_1575,In_841,In_393);
and U1576 (N_1576,In_1298,In_1272);
nand U1577 (N_1577,In_1270,In_2181);
and U1578 (N_1578,In_2123,In_981);
nand U1579 (N_1579,In_1548,In_1819);
or U1580 (N_1580,In_1,In_1271);
nor U1581 (N_1581,In_670,In_2996);
xnor U1582 (N_1582,In_569,In_2878);
and U1583 (N_1583,In_1482,In_58);
nand U1584 (N_1584,In_894,In_271);
or U1585 (N_1585,In_1310,In_1064);
xnor U1586 (N_1586,In_2974,In_561);
nor U1587 (N_1587,In_859,In_255);
and U1588 (N_1588,In_97,In_1439);
nand U1589 (N_1589,In_779,In_290);
nand U1590 (N_1590,In_1271,In_2065);
xnor U1591 (N_1591,In_1731,In_2980);
nand U1592 (N_1592,In_2333,In_2829);
xnor U1593 (N_1593,In_2485,In_1370);
xnor U1594 (N_1594,In_500,In_2817);
and U1595 (N_1595,In_1612,In_2264);
nor U1596 (N_1596,In_2079,In_561);
nand U1597 (N_1597,In_80,In_294);
and U1598 (N_1598,In_1342,In_1990);
or U1599 (N_1599,In_2235,In_340);
or U1600 (N_1600,In_2361,In_1101);
or U1601 (N_1601,In_744,In_1075);
nand U1602 (N_1602,In_1503,In_2969);
and U1603 (N_1603,In_2294,In_2378);
nor U1604 (N_1604,In_1068,In_2374);
nor U1605 (N_1605,In_1036,In_2945);
or U1606 (N_1606,In_730,In_1059);
nand U1607 (N_1607,In_548,In_2251);
nand U1608 (N_1608,In_262,In_1085);
and U1609 (N_1609,In_2105,In_634);
xnor U1610 (N_1610,In_2990,In_498);
and U1611 (N_1611,In_762,In_2985);
and U1612 (N_1612,In_307,In_2285);
or U1613 (N_1613,In_466,In_2995);
nor U1614 (N_1614,In_2348,In_194);
xnor U1615 (N_1615,In_2132,In_1535);
nand U1616 (N_1616,In_1962,In_1989);
nand U1617 (N_1617,In_2702,In_295);
xor U1618 (N_1618,In_1126,In_2310);
nand U1619 (N_1619,In_1775,In_2299);
nor U1620 (N_1620,In_2165,In_2157);
nand U1621 (N_1621,In_828,In_304);
nor U1622 (N_1622,In_2554,In_2524);
or U1623 (N_1623,In_2926,In_2192);
nor U1624 (N_1624,In_1783,In_1947);
or U1625 (N_1625,In_1979,In_2377);
nor U1626 (N_1626,In_1532,In_1647);
nand U1627 (N_1627,In_831,In_306);
nand U1628 (N_1628,In_2109,In_2660);
and U1629 (N_1629,In_76,In_860);
or U1630 (N_1630,In_1362,In_2399);
or U1631 (N_1631,In_2879,In_1874);
nand U1632 (N_1632,In_819,In_2163);
and U1633 (N_1633,In_2290,In_2790);
or U1634 (N_1634,In_1865,In_1956);
and U1635 (N_1635,In_2153,In_2962);
nand U1636 (N_1636,In_2188,In_1156);
or U1637 (N_1637,In_165,In_1960);
nand U1638 (N_1638,In_62,In_2957);
nor U1639 (N_1639,In_1395,In_1569);
nand U1640 (N_1640,In_566,In_2250);
nand U1641 (N_1641,In_1603,In_1312);
or U1642 (N_1642,In_235,In_2733);
xor U1643 (N_1643,In_2501,In_1253);
nand U1644 (N_1644,In_1976,In_1707);
xnor U1645 (N_1645,In_1772,In_180);
or U1646 (N_1646,In_2352,In_2808);
nor U1647 (N_1647,In_2291,In_564);
and U1648 (N_1648,In_873,In_591);
and U1649 (N_1649,In_1173,In_2667);
nand U1650 (N_1650,In_2854,In_1319);
xor U1651 (N_1651,In_2834,In_1230);
or U1652 (N_1652,In_1203,In_1083);
or U1653 (N_1653,In_1540,In_2123);
nor U1654 (N_1654,In_2293,In_2323);
or U1655 (N_1655,In_2404,In_1054);
xnor U1656 (N_1656,In_1271,In_600);
nor U1657 (N_1657,In_1617,In_2405);
or U1658 (N_1658,In_798,In_340);
nand U1659 (N_1659,In_2413,In_1992);
nor U1660 (N_1660,In_1261,In_81);
or U1661 (N_1661,In_1811,In_2445);
nand U1662 (N_1662,In_2301,In_1657);
and U1663 (N_1663,In_1746,In_2989);
or U1664 (N_1664,In_2355,In_2850);
xor U1665 (N_1665,In_2990,In_803);
xnor U1666 (N_1666,In_776,In_1547);
and U1667 (N_1667,In_421,In_851);
or U1668 (N_1668,In_2479,In_915);
nand U1669 (N_1669,In_1386,In_1589);
and U1670 (N_1670,In_890,In_1006);
nor U1671 (N_1671,In_101,In_1701);
nand U1672 (N_1672,In_2683,In_911);
nand U1673 (N_1673,In_2194,In_2765);
nor U1674 (N_1674,In_2102,In_2987);
nand U1675 (N_1675,In_1598,In_1246);
or U1676 (N_1676,In_626,In_2946);
xnor U1677 (N_1677,In_959,In_641);
or U1678 (N_1678,In_2416,In_1091);
or U1679 (N_1679,In_616,In_2517);
nor U1680 (N_1680,In_2043,In_2230);
nand U1681 (N_1681,In_945,In_2611);
nand U1682 (N_1682,In_513,In_541);
or U1683 (N_1683,In_2192,In_2839);
and U1684 (N_1684,In_1785,In_781);
nor U1685 (N_1685,In_2866,In_561);
xnor U1686 (N_1686,In_679,In_61);
or U1687 (N_1687,In_1324,In_1840);
nand U1688 (N_1688,In_880,In_1808);
nor U1689 (N_1689,In_1401,In_2018);
or U1690 (N_1690,In_769,In_2139);
nor U1691 (N_1691,In_2274,In_1487);
and U1692 (N_1692,In_2684,In_2396);
xor U1693 (N_1693,In_2215,In_152);
or U1694 (N_1694,In_445,In_1712);
or U1695 (N_1695,In_1936,In_1274);
and U1696 (N_1696,In_2010,In_957);
or U1697 (N_1697,In_1892,In_2822);
or U1698 (N_1698,In_1377,In_1417);
nor U1699 (N_1699,In_751,In_1013);
xnor U1700 (N_1700,In_2692,In_2378);
nand U1701 (N_1701,In_69,In_988);
and U1702 (N_1702,In_2814,In_2543);
nand U1703 (N_1703,In_2748,In_1472);
xor U1704 (N_1704,In_1702,In_1960);
nor U1705 (N_1705,In_1877,In_1530);
nor U1706 (N_1706,In_447,In_832);
nand U1707 (N_1707,In_1924,In_335);
and U1708 (N_1708,In_2464,In_299);
and U1709 (N_1709,In_1246,In_1933);
and U1710 (N_1710,In_2456,In_1625);
or U1711 (N_1711,In_15,In_2627);
and U1712 (N_1712,In_2544,In_2093);
nor U1713 (N_1713,In_66,In_1589);
nand U1714 (N_1714,In_1837,In_215);
xnor U1715 (N_1715,In_1779,In_2849);
or U1716 (N_1716,In_1289,In_2078);
xnor U1717 (N_1717,In_2398,In_1946);
xnor U1718 (N_1718,In_655,In_1969);
or U1719 (N_1719,In_1949,In_1323);
nor U1720 (N_1720,In_1355,In_741);
xnor U1721 (N_1721,In_1854,In_2143);
nand U1722 (N_1722,In_2636,In_728);
nand U1723 (N_1723,In_2366,In_2438);
nand U1724 (N_1724,In_1001,In_1664);
nand U1725 (N_1725,In_618,In_1027);
and U1726 (N_1726,In_1605,In_1823);
nand U1727 (N_1727,In_1750,In_1688);
or U1728 (N_1728,In_2185,In_216);
or U1729 (N_1729,In_524,In_487);
or U1730 (N_1730,In_1727,In_1038);
and U1731 (N_1731,In_2537,In_2092);
xor U1732 (N_1732,In_651,In_638);
nor U1733 (N_1733,In_1862,In_2369);
nand U1734 (N_1734,In_2667,In_1252);
or U1735 (N_1735,In_1711,In_330);
nand U1736 (N_1736,In_2891,In_884);
xor U1737 (N_1737,In_773,In_555);
and U1738 (N_1738,In_1650,In_1145);
nor U1739 (N_1739,In_2973,In_554);
and U1740 (N_1740,In_1635,In_930);
nand U1741 (N_1741,In_765,In_965);
nand U1742 (N_1742,In_1812,In_2100);
xor U1743 (N_1743,In_1684,In_637);
or U1744 (N_1744,In_1910,In_2292);
xnor U1745 (N_1745,In_1919,In_1427);
and U1746 (N_1746,In_2979,In_2961);
xor U1747 (N_1747,In_2766,In_1330);
and U1748 (N_1748,In_1553,In_2532);
xor U1749 (N_1749,In_852,In_2051);
or U1750 (N_1750,In_76,In_1723);
nor U1751 (N_1751,In_933,In_2851);
nand U1752 (N_1752,In_23,In_1555);
xnor U1753 (N_1753,In_2948,In_1921);
nor U1754 (N_1754,In_2047,In_1281);
xnor U1755 (N_1755,In_1099,In_1060);
or U1756 (N_1756,In_1839,In_2678);
or U1757 (N_1757,In_2818,In_362);
nor U1758 (N_1758,In_672,In_2970);
xnor U1759 (N_1759,In_2913,In_916);
or U1760 (N_1760,In_286,In_1658);
xor U1761 (N_1761,In_2968,In_726);
nand U1762 (N_1762,In_2816,In_494);
nand U1763 (N_1763,In_1560,In_2133);
nor U1764 (N_1764,In_1493,In_1459);
nand U1765 (N_1765,In_1514,In_355);
or U1766 (N_1766,In_2087,In_162);
nor U1767 (N_1767,In_1932,In_482);
xor U1768 (N_1768,In_2943,In_936);
or U1769 (N_1769,In_206,In_216);
or U1770 (N_1770,In_1951,In_169);
and U1771 (N_1771,In_766,In_551);
and U1772 (N_1772,In_2361,In_667);
nor U1773 (N_1773,In_701,In_1279);
and U1774 (N_1774,In_2472,In_2717);
and U1775 (N_1775,In_2147,In_2030);
and U1776 (N_1776,In_1918,In_1578);
xor U1777 (N_1777,In_693,In_2454);
or U1778 (N_1778,In_1756,In_658);
and U1779 (N_1779,In_1116,In_2713);
nand U1780 (N_1780,In_1514,In_2575);
nand U1781 (N_1781,In_977,In_2928);
or U1782 (N_1782,In_1139,In_477);
and U1783 (N_1783,In_332,In_1558);
xor U1784 (N_1784,In_2016,In_2484);
xor U1785 (N_1785,In_1315,In_413);
xnor U1786 (N_1786,In_31,In_2948);
xnor U1787 (N_1787,In_743,In_2073);
nor U1788 (N_1788,In_2855,In_2959);
nand U1789 (N_1789,In_2735,In_1169);
or U1790 (N_1790,In_947,In_76);
nor U1791 (N_1791,In_2424,In_1926);
nand U1792 (N_1792,In_1512,In_2871);
or U1793 (N_1793,In_2339,In_1707);
xor U1794 (N_1794,In_288,In_2858);
xnor U1795 (N_1795,In_476,In_160);
nand U1796 (N_1796,In_556,In_1245);
xor U1797 (N_1797,In_1836,In_2771);
or U1798 (N_1798,In_2307,In_1122);
xnor U1799 (N_1799,In_243,In_184);
xor U1800 (N_1800,In_2192,In_1811);
or U1801 (N_1801,In_2420,In_1883);
nand U1802 (N_1802,In_2640,In_1776);
or U1803 (N_1803,In_152,In_1562);
or U1804 (N_1804,In_1,In_1739);
nand U1805 (N_1805,In_333,In_1272);
and U1806 (N_1806,In_520,In_2189);
or U1807 (N_1807,In_521,In_1827);
xor U1808 (N_1808,In_1414,In_2075);
or U1809 (N_1809,In_2785,In_165);
and U1810 (N_1810,In_754,In_2265);
and U1811 (N_1811,In_521,In_2965);
xnor U1812 (N_1812,In_2223,In_988);
and U1813 (N_1813,In_446,In_980);
and U1814 (N_1814,In_956,In_2510);
xnor U1815 (N_1815,In_890,In_2426);
nand U1816 (N_1816,In_1744,In_1308);
xnor U1817 (N_1817,In_145,In_1179);
nand U1818 (N_1818,In_1854,In_2506);
and U1819 (N_1819,In_2291,In_2268);
and U1820 (N_1820,In_1923,In_2866);
nor U1821 (N_1821,In_2236,In_2576);
xnor U1822 (N_1822,In_1941,In_998);
nand U1823 (N_1823,In_288,In_2588);
nor U1824 (N_1824,In_2530,In_1290);
nand U1825 (N_1825,In_965,In_1274);
and U1826 (N_1826,In_1950,In_1967);
or U1827 (N_1827,In_820,In_1990);
and U1828 (N_1828,In_203,In_1610);
xor U1829 (N_1829,In_1748,In_2871);
nand U1830 (N_1830,In_838,In_633);
and U1831 (N_1831,In_1951,In_843);
nand U1832 (N_1832,In_2213,In_2228);
nand U1833 (N_1833,In_863,In_612);
nor U1834 (N_1834,In_2733,In_429);
and U1835 (N_1835,In_1814,In_2944);
or U1836 (N_1836,In_1212,In_1658);
and U1837 (N_1837,In_1478,In_1393);
nand U1838 (N_1838,In_173,In_2344);
and U1839 (N_1839,In_316,In_151);
nand U1840 (N_1840,In_921,In_1470);
and U1841 (N_1841,In_1683,In_1831);
or U1842 (N_1842,In_213,In_1704);
nor U1843 (N_1843,In_1241,In_2713);
xnor U1844 (N_1844,In_999,In_1566);
nor U1845 (N_1845,In_135,In_1716);
nor U1846 (N_1846,In_1322,In_625);
or U1847 (N_1847,In_2700,In_1943);
nor U1848 (N_1848,In_2741,In_779);
xor U1849 (N_1849,In_2224,In_2667);
nand U1850 (N_1850,In_1719,In_391);
nor U1851 (N_1851,In_984,In_970);
and U1852 (N_1852,In_1495,In_693);
or U1853 (N_1853,In_1453,In_2473);
nor U1854 (N_1854,In_955,In_905);
or U1855 (N_1855,In_2005,In_239);
xnor U1856 (N_1856,In_331,In_2652);
or U1857 (N_1857,In_1085,In_2188);
nand U1858 (N_1858,In_2733,In_2085);
or U1859 (N_1859,In_255,In_827);
xnor U1860 (N_1860,In_1473,In_2841);
nand U1861 (N_1861,In_2450,In_470);
nand U1862 (N_1862,In_118,In_1755);
nor U1863 (N_1863,In_2238,In_1268);
and U1864 (N_1864,In_1294,In_2778);
or U1865 (N_1865,In_1524,In_2106);
and U1866 (N_1866,In_501,In_2398);
and U1867 (N_1867,In_1276,In_107);
nand U1868 (N_1868,In_2545,In_2862);
or U1869 (N_1869,In_1692,In_1567);
or U1870 (N_1870,In_1349,In_107);
nor U1871 (N_1871,In_334,In_2613);
and U1872 (N_1872,In_2314,In_1576);
or U1873 (N_1873,In_2671,In_1731);
nand U1874 (N_1874,In_137,In_976);
xnor U1875 (N_1875,In_104,In_2774);
nor U1876 (N_1876,In_758,In_2006);
xor U1877 (N_1877,In_2841,In_1574);
nor U1878 (N_1878,In_526,In_1791);
xnor U1879 (N_1879,In_192,In_358);
nor U1880 (N_1880,In_1392,In_1074);
nand U1881 (N_1881,In_2561,In_3);
and U1882 (N_1882,In_2610,In_933);
nor U1883 (N_1883,In_1728,In_1256);
and U1884 (N_1884,In_1554,In_2127);
or U1885 (N_1885,In_2482,In_2322);
nor U1886 (N_1886,In_830,In_1025);
nor U1887 (N_1887,In_2071,In_967);
and U1888 (N_1888,In_1969,In_403);
nand U1889 (N_1889,In_1473,In_2909);
xnor U1890 (N_1890,In_2123,In_123);
or U1891 (N_1891,In_2246,In_2689);
or U1892 (N_1892,In_989,In_2248);
or U1893 (N_1893,In_2873,In_1157);
or U1894 (N_1894,In_542,In_969);
xor U1895 (N_1895,In_2092,In_1216);
and U1896 (N_1896,In_1058,In_2780);
nand U1897 (N_1897,In_536,In_1692);
nand U1898 (N_1898,In_2416,In_531);
or U1899 (N_1899,In_2859,In_828);
xor U1900 (N_1900,In_1075,In_1868);
xor U1901 (N_1901,In_2300,In_1379);
nand U1902 (N_1902,In_1852,In_1048);
nand U1903 (N_1903,In_2824,In_499);
nand U1904 (N_1904,In_1255,In_1905);
xnor U1905 (N_1905,In_2483,In_1335);
nor U1906 (N_1906,In_648,In_1071);
nand U1907 (N_1907,In_938,In_2545);
or U1908 (N_1908,In_1931,In_174);
nand U1909 (N_1909,In_2323,In_2879);
xor U1910 (N_1910,In_1653,In_2921);
xnor U1911 (N_1911,In_420,In_2903);
nand U1912 (N_1912,In_367,In_2447);
xnor U1913 (N_1913,In_1771,In_1650);
nor U1914 (N_1914,In_1173,In_387);
nand U1915 (N_1915,In_2414,In_653);
nand U1916 (N_1916,In_1625,In_1559);
and U1917 (N_1917,In_746,In_2689);
nor U1918 (N_1918,In_1886,In_1785);
xor U1919 (N_1919,In_1349,In_164);
and U1920 (N_1920,In_1776,In_1533);
and U1921 (N_1921,In_1131,In_769);
or U1922 (N_1922,In_1053,In_2738);
or U1923 (N_1923,In_2767,In_2851);
nor U1924 (N_1924,In_665,In_2403);
nand U1925 (N_1925,In_794,In_2431);
nor U1926 (N_1926,In_1842,In_919);
and U1927 (N_1927,In_925,In_2496);
xnor U1928 (N_1928,In_2859,In_2678);
nand U1929 (N_1929,In_2878,In_969);
nand U1930 (N_1930,In_449,In_75);
nor U1931 (N_1931,In_2728,In_143);
and U1932 (N_1932,In_2290,In_1832);
nor U1933 (N_1933,In_575,In_383);
or U1934 (N_1934,In_2772,In_1795);
nor U1935 (N_1935,In_1832,In_1374);
nor U1936 (N_1936,In_2765,In_324);
and U1937 (N_1937,In_2043,In_1681);
or U1938 (N_1938,In_793,In_1888);
and U1939 (N_1939,In_578,In_4);
and U1940 (N_1940,In_1093,In_1672);
nand U1941 (N_1941,In_2206,In_852);
xnor U1942 (N_1942,In_1608,In_1393);
xor U1943 (N_1943,In_2124,In_403);
nor U1944 (N_1944,In_2204,In_893);
nor U1945 (N_1945,In_17,In_2748);
and U1946 (N_1946,In_2753,In_1026);
or U1947 (N_1947,In_892,In_2583);
nor U1948 (N_1948,In_1480,In_852);
and U1949 (N_1949,In_842,In_2682);
nand U1950 (N_1950,In_1939,In_966);
nand U1951 (N_1951,In_2033,In_2075);
and U1952 (N_1952,In_2024,In_2375);
or U1953 (N_1953,In_692,In_1527);
xnor U1954 (N_1954,In_854,In_1632);
nand U1955 (N_1955,In_1030,In_2936);
nand U1956 (N_1956,In_177,In_1053);
and U1957 (N_1957,In_2659,In_2997);
nand U1958 (N_1958,In_2870,In_555);
xor U1959 (N_1959,In_2641,In_513);
nand U1960 (N_1960,In_2336,In_1955);
xor U1961 (N_1961,In_641,In_595);
xor U1962 (N_1962,In_2413,In_2374);
nor U1963 (N_1963,In_2922,In_2535);
xnor U1964 (N_1964,In_1215,In_2213);
nand U1965 (N_1965,In_2609,In_2167);
and U1966 (N_1966,In_1939,In_29);
nand U1967 (N_1967,In_829,In_2754);
nor U1968 (N_1968,In_1091,In_1636);
and U1969 (N_1969,In_475,In_702);
xnor U1970 (N_1970,In_452,In_647);
xor U1971 (N_1971,In_2047,In_672);
nand U1972 (N_1972,In_1168,In_548);
and U1973 (N_1973,In_142,In_2522);
nand U1974 (N_1974,In_2073,In_2752);
nor U1975 (N_1975,In_12,In_1847);
and U1976 (N_1976,In_1995,In_138);
or U1977 (N_1977,In_2925,In_140);
and U1978 (N_1978,In_2460,In_1469);
nand U1979 (N_1979,In_7,In_1817);
nor U1980 (N_1980,In_908,In_2834);
nor U1981 (N_1981,In_1067,In_485);
nand U1982 (N_1982,In_2894,In_738);
or U1983 (N_1983,In_298,In_752);
or U1984 (N_1984,In_2773,In_2525);
nand U1985 (N_1985,In_253,In_954);
nand U1986 (N_1986,In_1936,In_80);
nor U1987 (N_1987,In_1086,In_1804);
or U1988 (N_1988,In_2525,In_665);
nor U1989 (N_1989,In_1186,In_870);
or U1990 (N_1990,In_1632,In_1609);
nor U1991 (N_1991,In_1869,In_1633);
nor U1992 (N_1992,In_888,In_2451);
nor U1993 (N_1993,In_451,In_1562);
xnor U1994 (N_1994,In_850,In_489);
nand U1995 (N_1995,In_476,In_1536);
or U1996 (N_1996,In_1784,In_2001);
nor U1997 (N_1997,In_2083,In_876);
and U1998 (N_1998,In_1525,In_2420);
and U1999 (N_1999,In_2521,In_45);
nor U2000 (N_2000,In_2885,In_2042);
and U2001 (N_2001,In_1919,In_2932);
nand U2002 (N_2002,In_1818,In_446);
xor U2003 (N_2003,In_1912,In_2815);
nand U2004 (N_2004,In_443,In_1444);
or U2005 (N_2005,In_2638,In_2171);
xnor U2006 (N_2006,In_1432,In_2788);
nor U2007 (N_2007,In_1369,In_1604);
or U2008 (N_2008,In_1986,In_654);
nand U2009 (N_2009,In_2587,In_561);
xor U2010 (N_2010,In_19,In_450);
and U2011 (N_2011,In_2820,In_2231);
xor U2012 (N_2012,In_2816,In_1573);
or U2013 (N_2013,In_837,In_1634);
nand U2014 (N_2014,In_906,In_28);
and U2015 (N_2015,In_1634,In_1477);
and U2016 (N_2016,In_227,In_2261);
or U2017 (N_2017,In_1893,In_2743);
or U2018 (N_2018,In_1514,In_980);
or U2019 (N_2019,In_2486,In_117);
nor U2020 (N_2020,In_1147,In_7);
nand U2021 (N_2021,In_1199,In_885);
xnor U2022 (N_2022,In_31,In_2914);
and U2023 (N_2023,In_2611,In_120);
nor U2024 (N_2024,In_11,In_396);
or U2025 (N_2025,In_2823,In_151);
nor U2026 (N_2026,In_1341,In_225);
or U2027 (N_2027,In_2076,In_30);
or U2028 (N_2028,In_397,In_505);
and U2029 (N_2029,In_2346,In_1917);
nor U2030 (N_2030,In_647,In_234);
or U2031 (N_2031,In_1284,In_2407);
and U2032 (N_2032,In_2572,In_1261);
xor U2033 (N_2033,In_1543,In_2250);
or U2034 (N_2034,In_1839,In_1352);
and U2035 (N_2035,In_1881,In_418);
nor U2036 (N_2036,In_1924,In_214);
xor U2037 (N_2037,In_22,In_2370);
or U2038 (N_2038,In_1244,In_194);
nor U2039 (N_2039,In_2795,In_1423);
nand U2040 (N_2040,In_2941,In_1866);
xor U2041 (N_2041,In_2857,In_308);
nand U2042 (N_2042,In_1775,In_2964);
nor U2043 (N_2043,In_1010,In_898);
and U2044 (N_2044,In_297,In_2073);
nand U2045 (N_2045,In_2821,In_395);
nand U2046 (N_2046,In_2025,In_83);
nor U2047 (N_2047,In_2519,In_149);
xor U2048 (N_2048,In_2719,In_373);
or U2049 (N_2049,In_558,In_2771);
xnor U2050 (N_2050,In_2961,In_1398);
nor U2051 (N_2051,In_1024,In_146);
xor U2052 (N_2052,In_2566,In_2066);
or U2053 (N_2053,In_2585,In_538);
nand U2054 (N_2054,In_232,In_954);
or U2055 (N_2055,In_2160,In_1951);
xor U2056 (N_2056,In_597,In_479);
and U2057 (N_2057,In_2802,In_1456);
and U2058 (N_2058,In_1177,In_1173);
and U2059 (N_2059,In_1730,In_2624);
nand U2060 (N_2060,In_2164,In_884);
nand U2061 (N_2061,In_2034,In_2511);
nor U2062 (N_2062,In_527,In_966);
or U2063 (N_2063,In_163,In_828);
nor U2064 (N_2064,In_963,In_994);
or U2065 (N_2065,In_520,In_247);
nand U2066 (N_2066,In_1271,In_869);
and U2067 (N_2067,In_2416,In_737);
xor U2068 (N_2068,In_1706,In_841);
nor U2069 (N_2069,In_1591,In_1372);
xor U2070 (N_2070,In_2984,In_1919);
and U2071 (N_2071,In_689,In_1600);
nor U2072 (N_2072,In_1311,In_715);
xor U2073 (N_2073,In_2464,In_1247);
nor U2074 (N_2074,In_2605,In_2078);
and U2075 (N_2075,In_345,In_154);
xnor U2076 (N_2076,In_1878,In_2403);
and U2077 (N_2077,In_715,In_957);
and U2078 (N_2078,In_1343,In_1563);
nor U2079 (N_2079,In_698,In_1295);
and U2080 (N_2080,In_130,In_1829);
xnor U2081 (N_2081,In_1912,In_1432);
nor U2082 (N_2082,In_124,In_2747);
xnor U2083 (N_2083,In_2648,In_2070);
or U2084 (N_2084,In_2629,In_2754);
nor U2085 (N_2085,In_2159,In_537);
nand U2086 (N_2086,In_2473,In_636);
or U2087 (N_2087,In_1982,In_428);
or U2088 (N_2088,In_1307,In_1251);
xnor U2089 (N_2089,In_2877,In_2091);
or U2090 (N_2090,In_739,In_1893);
and U2091 (N_2091,In_2873,In_1143);
and U2092 (N_2092,In_1400,In_1126);
nand U2093 (N_2093,In_2513,In_636);
nor U2094 (N_2094,In_1040,In_677);
nand U2095 (N_2095,In_1799,In_1592);
or U2096 (N_2096,In_972,In_98);
nor U2097 (N_2097,In_88,In_975);
nor U2098 (N_2098,In_2186,In_124);
nor U2099 (N_2099,In_2178,In_1833);
xor U2100 (N_2100,In_581,In_531);
and U2101 (N_2101,In_35,In_2449);
and U2102 (N_2102,In_2547,In_2630);
nand U2103 (N_2103,In_1123,In_1823);
and U2104 (N_2104,In_1415,In_908);
and U2105 (N_2105,In_2467,In_470);
or U2106 (N_2106,In_1706,In_757);
xor U2107 (N_2107,In_2676,In_252);
and U2108 (N_2108,In_2782,In_1915);
or U2109 (N_2109,In_1741,In_2572);
nor U2110 (N_2110,In_1931,In_1281);
nor U2111 (N_2111,In_907,In_2072);
nor U2112 (N_2112,In_2380,In_240);
or U2113 (N_2113,In_1596,In_771);
or U2114 (N_2114,In_2980,In_240);
and U2115 (N_2115,In_2033,In_1706);
nor U2116 (N_2116,In_53,In_1740);
xor U2117 (N_2117,In_396,In_1671);
xor U2118 (N_2118,In_2044,In_551);
xnor U2119 (N_2119,In_1867,In_67);
xnor U2120 (N_2120,In_2980,In_56);
or U2121 (N_2121,In_1116,In_2416);
nand U2122 (N_2122,In_2686,In_1610);
xor U2123 (N_2123,In_2076,In_1583);
xnor U2124 (N_2124,In_530,In_784);
and U2125 (N_2125,In_154,In_359);
xnor U2126 (N_2126,In_1326,In_2257);
xnor U2127 (N_2127,In_1778,In_570);
or U2128 (N_2128,In_502,In_239);
and U2129 (N_2129,In_88,In_2529);
nor U2130 (N_2130,In_2901,In_604);
xor U2131 (N_2131,In_740,In_999);
nand U2132 (N_2132,In_1461,In_2873);
xnor U2133 (N_2133,In_2278,In_202);
and U2134 (N_2134,In_1144,In_1683);
nor U2135 (N_2135,In_1795,In_1887);
nand U2136 (N_2136,In_69,In_2077);
or U2137 (N_2137,In_624,In_765);
xor U2138 (N_2138,In_1784,In_2322);
or U2139 (N_2139,In_298,In_2309);
or U2140 (N_2140,In_1270,In_1001);
nand U2141 (N_2141,In_2271,In_1540);
nor U2142 (N_2142,In_2752,In_2247);
nand U2143 (N_2143,In_2669,In_2955);
nor U2144 (N_2144,In_2944,In_1826);
nand U2145 (N_2145,In_1127,In_1877);
or U2146 (N_2146,In_2158,In_2271);
nor U2147 (N_2147,In_697,In_1063);
nor U2148 (N_2148,In_393,In_1915);
xor U2149 (N_2149,In_658,In_520);
or U2150 (N_2150,In_547,In_2115);
nor U2151 (N_2151,In_1649,In_1699);
xnor U2152 (N_2152,In_2361,In_2409);
or U2153 (N_2153,In_1097,In_177);
xnor U2154 (N_2154,In_337,In_379);
nor U2155 (N_2155,In_1956,In_2024);
or U2156 (N_2156,In_1956,In_2539);
nand U2157 (N_2157,In_658,In_1503);
nor U2158 (N_2158,In_515,In_2727);
xor U2159 (N_2159,In_2831,In_2850);
nand U2160 (N_2160,In_2655,In_271);
nor U2161 (N_2161,In_615,In_2809);
and U2162 (N_2162,In_2178,In_1158);
nor U2163 (N_2163,In_1615,In_1774);
nand U2164 (N_2164,In_1232,In_526);
nand U2165 (N_2165,In_1635,In_333);
nand U2166 (N_2166,In_1071,In_1522);
and U2167 (N_2167,In_1726,In_648);
nor U2168 (N_2168,In_249,In_2225);
or U2169 (N_2169,In_87,In_204);
and U2170 (N_2170,In_1656,In_2895);
and U2171 (N_2171,In_1482,In_1881);
or U2172 (N_2172,In_1347,In_1501);
xnor U2173 (N_2173,In_2706,In_818);
xor U2174 (N_2174,In_84,In_398);
and U2175 (N_2175,In_1611,In_2420);
xnor U2176 (N_2176,In_2327,In_870);
nand U2177 (N_2177,In_344,In_2360);
or U2178 (N_2178,In_2633,In_2288);
or U2179 (N_2179,In_2891,In_2005);
xor U2180 (N_2180,In_1418,In_2481);
nor U2181 (N_2181,In_1006,In_159);
nor U2182 (N_2182,In_865,In_2599);
or U2183 (N_2183,In_1104,In_268);
and U2184 (N_2184,In_36,In_1460);
or U2185 (N_2185,In_1228,In_981);
nor U2186 (N_2186,In_2121,In_795);
nand U2187 (N_2187,In_1474,In_583);
xnor U2188 (N_2188,In_2969,In_2836);
nor U2189 (N_2189,In_1783,In_1137);
xnor U2190 (N_2190,In_297,In_1360);
xor U2191 (N_2191,In_1863,In_2910);
nor U2192 (N_2192,In_464,In_1575);
nor U2193 (N_2193,In_1934,In_965);
xnor U2194 (N_2194,In_406,In_789);
xnor U2195 (N_2195,In_2026,In_1209);
nand U2196 (N_2196,In_1523,In_1066);
or U2197 (N_2197,In_1382,In_2574);
nand U2198 (N_2198,In_855,In_2735);
and U2199 (N_2199,In_1974,In_2519);
and U2200 (N_2200,In_1325,In_640);
nor U2201 (N_2201,In_224,In_67);
and U2202 (N_2202,In_132,In_865);
nor U2203 (N_2203,In_2509,In_394);
nor U2204 (N_2204,In_138,In_1439);
or U2205 (N_2205,In_2650,In_2281);
nand U2206 (N_2206,In_2065,In_2970);
or U2207 (N_2207,In_275,In_2423);
nand U2208 (N_2208,In_904,In_269);
and U2209 (N_2209,In_2526,In_2128);
xor U2210 (N_2210,In_507,In_1543);
xor U2211 (N_2211,In_1101,In_1183);
or U2212 (N_2212,In_182,In_2890);
or U2213 (N_2213,In_286,In_1488);
nand U2214 (N_2214,In_2585,In_2364);
and U2215 (N_2215,In_253,In_2890);
xnor U2216 (N_2216,In_242,In_2304);
or U2217 (N_2217,In_1132,In_568);
nand U2218 (N_2218,In_1329,In_2450);
xor U2219 (N_2219,In_1379,In_2460);
xor U2220 (N_2220,In_2155,In_944);
or U2221 (N_2221,In_516,In_2938);
or U2222 (N_2222,In_447,In_1537);
and U2223 (N_2223,In_402,In_1040);
xor U2224 (N_2224,In_298,In_1497);
xor U2225 (N_2225,In_1333,In_2246);
nand U2226 (N_2226,In_2091,In_2900);
and U2227 (N_2227,In_428,In_2521);
or U2228 (N_2228,In_787,In_496);
nand U2229 (N_2229,In_1763,In_2408);
nand U2230 (N_2230,In_1051,In_1759);
xor U2231 (N_2231,In_2285,In_169);
or U2232 (N_2232,In_1735,In_1450);
xor U2233 (N_2233,In_47,In_1028);
and U2234 (N_2234,In_353,In_155);
xor U2235 (N_2235,In_465,In_2299);
xor U2236 (N_2236,In_2266,In_795);
nand U2237 (N_2237,In_1154,In_1561);
or U2238 (N_2238,In_2601,In_1762);
nor U2239 (N_2239,In_2434,In_116);
xnor U2240 (N_2240,In_823,In_2930);
nand U2241 (N_2241,In_2055,In_476);
nor U2242 (N_2242,In_1806,In_513);
nand U2243 (N_2243,In_1713,In_2752);
nand U2244 (N_2244,In_2053,In_1608);
and U2245 (N_2245,In_2216,In_1007);
nor U2246 (N_2246,In_678,In_2055);
and U2247 (N_2247,In_1970,In_213);
nor U2248 (N_2248,In_569,In_429);
nand U2249 (N_2249,In_1001,In_742);
and U2250 (N_2250,In_545,In_865);
or U2251 (N_2251,In_2633,In_1050);
or U2252 (N_2252,In_2079,In_1492);
nand U2253 (N_2253,In_2261,In_1499);
xor U2254 (N_2254,In_1860,In_651);
or U2255 (N_2255,In_455,In_1107);
xor U2256 (N_2256,In_2461,In_2067);
nor U2257 (N_2257,In_2759,In_272);
nand U2258 (N_2258,In_2605,In_1146);
nor U2259 (N_2259,In_1485,In_270);
or U2260 (N_2260,In_1803,In_2270);
or U2261 (N_2261,In_2007,In_1273);
nand U2262 (N_2262,In_2462,In_1806);
xor U2263 (N_2263,In_1886,In_1666);
nand U2264 (N_2264,In_2315,In_1877);
or U2265 (N_2265,In_2139,In_554);
or U2266 (N_2266,In_402,In_2788);
xor U2267 (N_2267,In_409,In_2483);
nand U2268 (N_2268,In_2876,In_43);
or U2269 (N_2269,In_1906,In_500);
xor U2270 (N_2270,In_1718,In_277);
xnor U2271 (N_2271,In_1650,In_66);
xnor U2272 (N_2272,In_1395,In_2506);
or U2273 (N_2273,In_109,In_2055);
nor U2274 (N_2274,In_1032,In_792);
xnor U2275 (N_2275,In_2788,In_146);
nand U2276 (N_2276,In_2131,In_2599);
xnor U2277 (N_2277,In_649,In_902);
or U2278 (N_2278,In_791,In_54);
nor U2279 (N_2279,In_699,In_245);
and U2280 (N_2280,In_2549,In_2772);
and U2281 (N_2281,In_382,In_759);
and U2282 (N_2282,In_297,In_1206);
and U2283 (N_2283,In_2809,In_1771);
nand U2284 (N_2284,In_2152,In_892);
nor U2285 (N_2285,In_386,In_1516);
xnor U2286 (N_2286,In_1370,In_2789);
and U2287 (N_2287,In_384,In_667);
nand U2288 (N_2288,In_1453,In_1002);
xnor U2289 (N_2289,In_1482,In_1805);
xnor U2290 (N_2290,In_1866,In_76);
nor U2291 (N_2291,In_2041,In_1068);
nor U2292 (N_2292,In_710,In_2018);
or U2293 (N_2293,In_1436,In_2974);
xnor U2294 (N_2294,In_2944,In_2021);
nor U2295 (N_2295,In_2082,In_2513);
nor U2296 (N_2296,In_1367,In_756);
or U2297 (N_2297,In_1230,In_417);
nor U2298 (N_2298,In_1283,In_2744);
and U2299 (N_2299,In_1394,In_96);
nand U2300 (N_2300,In_1123,In_1234);
or U2301 (N_2301,In_481,In_716);
xnor U2302 (N_2302,In_2460,In_394);
xnor U2303 (N_2303,In_2638,In_1634);
nand U2304 (N_2304,In_2252,In_2678);
nor U2305 (N_2305,In_2208,In_2038);
xor U2306 (N_2306,In_1944,In_1972);
xor U2307 (N_2307,In_1883,In_2880);
nand U2308 (N_2308,In_1342,In_1461);
nand U2309 (N_2309,In_282,In_1854);
nand U2310 (N_2310,In_1231,In_1745);
or U2311 (N_2311,In_1313,In_2240);
or U2312 (N_2312,In_1958,In_869);
xnor U2313 (N_2313,In_301,In_1748);
xnor U2314 (N_2314,In_2332,In_27);
or U2315 (N_2315,In_2415,In_2335);
xor U2316 (N_2316,In_2318,In_2238);
nor U2317 (N_2317,In_225,In_2331);
and U2318 (N_2318,In_1602,In_855);
xor U2319 (N_2319,In_1669,In_1332);
nor U2320 (N_2320,In_1566,In_858);
and U2321 (N_2321,In_2544,In_2565);
or U2322 (N_2322,In_982,In_974);
nand U2323 (N_2323,In_2874,In_1642);
nand U2324 (N_2324,In_511,In_834);
xnor U2325 (N_2325,In_2614,In_691);
and U2326 (N_2326,In_1349,In_2531);
and U2327 (N_2327,In_906,In_1635);
xor U2328 (N_2328,In_390,In_1478);
or U2329 (N_2329,In_1212,In_525);
nand U2330 (N_2330,In_694,In_88);
and U2331 (N_2331,In_2624,In_206);
nor U2332 (N_2332,In_1316,In_1551);
or U2333 (N_2333,In_134,In_2788);
xor U2334 (N_2334,In_2243,In_377);
nand U2335 (N_2335,In_906,In_2983);
nor U2336 (N_2336,In_174,In_1431);
nand U2337 (N_2337,In_1459,In_360);
and U2338 (N_2338,In_2720,In_648);
and U2339 (N_2339,In_1474,In_351);
and U2340 (N_2340,In_2172,In_585);
nand U2341 (N_2341,In_2049,In_1437);
or U2342 (N_2342,In_2300,In_2126);
xor U2343 (N_2343,In_853,In_1675);
xnor U2344 (N_2344,In_573,In_2890);
and U2345 (N_2345,In_1139,In_287);
nor U2346 (N_2346,In_1776,In_593);
and U2347 (N_2347,In_1130,In_438);
or U2348 (N_2348,In_1146,In_111);
and U2349 (N_2349,In_600,In_723);
xor U2350 (N_2350,In_1375,In_842);
nor U2351 (N_2351,In_359,In_73);
xnor U2352 (N_2352,In_2683,In_2421);
nand U2353 (N_2353,In_2125,In_1903);
nor U2354 (N_2354,In_1151,In_2519);
nor U2355 (N_2355,In_2764,In_1756);
xor U2356 (N_2356,In_806,In_2759);
nor U2357 (N_2357,In_518,In_2538);
nand U2358 (N_2358,In_1404,In_1331);
xor U2359 (N_2359,In_1626,In_2972);
or U2360 (N_2360,In_2,In_889);
nand U2361 (N_2361,In_2595,In_431);
or U2362 (N_2362,In_2482,In_1177);
xor U2363 (N_2363,In_268,In_447);
nor U2364 (N_2364,In_1155,In_818);
xnor U2365 (N_2365,In_574,In_2937);
nand U2366 (N_2366,In_953,In_797);
nor U2367 (N_2367,In_2111,In_1720);
or U2368 (N_2368,In_1225,In_428);
nor U2369 (N_2369,In_1554,In_992);
nand U2370 (N_2370,In_1116,In_2234);
and U2371 (N_2371,In_2318,In_2741);
and U2372 (N_2372,In_2973,In_2330);
and U2373 (N_2373,In_1763,In_2848);
and U2374 (N_2374,In_2455,In_518);
xnor U2375 (N_2375,In_1819,In_2245);
and U2376 (N_2376,In_709,In_906);
nor U2377 (N_2377,In_2058,In_1972);
nor U2378 (N_2378,In_879,In_1889);
or U2379 (N_2379,In_474,In_2715);
and U2380 (N_2380,In_2334,In_1307);
and U2381 (N_2381,In_2497,In_2188);
nor U2382 (N_2382,In_1569,In_1303);
and U2383 (N_2383,In_418,In_2025);
nand U2384 (N_2384,In_2010,In_610);
nand U2385 (N_2385,In_2425,In_2642);
nor U2386 (N_2386,In_526,In_2606);
nand U2387 (N_2387,In_731,In_186);
nand U2388 (N_2388,In_1041,In_253);
nor U2389 (N_2389,In_683,In_448);
and U2390 (N_2390,In_178,In_216);
nand U2391 (N_2391,In_2700,In_488);
xor U2392 (N_2392,In_659,In_923);
nor U2393 (N_2393,In_1819,In_967);
xor U2394 (N_2394,In_2604,In_303);
or U2395 (N_2395,In_1167,In_1145);
nand U2396 (N_2396,In_1096,In_1331);
nand U2397 (N_2397,In_2820,In_1707);
nand U2398 (N_2398,In_141,In_2231);
nand U2399 (N_2399,In_2331,In_2987);
and U2400 (N_2400,In_2206,In_2872);
xnor U2401 (N_2401,In_1857,In_1869);
or U2402 (N_2402,In_2791,In_349);
xor U2403 (N_2403,In_492,In_68);
and U2404 (N_2404,In_1891,In_2683);
nand U2405 (N_2405,In_1163,In_1189);
nor U2406 (N_2406,In_1426,In_2884);
or U2407 (N_2407,In_2986,In_2658);
xnor U2408 (N_2408,In_2937,In_1886);
and U2409 (N_2409,In_183,In_343);
or U2410 (N_2410,In_24,In_982);
and U2411 (N_2411,In_944,In_1035);
xnor U2412 (N_2412,In_1743,In_65);
nor U2413 (N_2413,In_2723,In_2588);
nor U2414 (N_2414,In_581,In_1594);
xor U2415 (N_2415,In_2563,In_1677);
nor U2416 (N_2416,In_1380,In_2822);
nor U2417 (N_2417,In_1946,In_2680);
or U2418 (N_2418,In_1525,In_1657);
and U2419 (N_2419,In_68,In_2375);
xnor U2420 (N_2420,In_249,In_2092);
nand U2421 (N_2421,In_2171,In_485);
nand U2422 (N_2422,In_1027,In_2359);
nand U2423 (N_2423,In_2225,In_473);
xnor U2424 (N_2424,In_2447,In_2390);
and U2425 (N_2425,In_2267,In_2652);
nor U2426 (N_2426,In_1172,In_1292);
or U2427 (N_2427,In_2230,In_1505);
and U2428 (N_2428,In_642,In_2903);
and U2429 (N_2429,In_717,In_2604);
xnor U2430 (N_2430,In_2193,In_320);
nor U2431 (N_2431,In_2549,In_964);
nand U2432 (N_2432,In_2002,In_1991);
and U2433 (N_2433,In_2849,In_973);
nor U2434 (N_2434,In_55,In_1443);
nor U2435 (N_2435,In_188,In_2432);
and U2436 (N_2436,In_1575,In_1181);
and U2437 (N_2437,In_934,In_57);
or U2438 (N_2438,In_1662,In_957);
nand U2439 (N_2439,In_1986,In_244);
and U2440 (N_2440,In_1311,In_2478);
xor U2441 (N_2441,In_2585,In_1595);
or U2442 (N_2442,In_377,In_1382);
nand U2443 (N_2443,In_2819,In_2329);
and U2444 (N_2444,In_1828,In_1569);
nor U2445 (N_2445,In_2848,In_221);
or U2446 (N_2446,In_136,In_945);
or U2447 (N_2447,In_1116,In_372);
xnor U2448 (N_2448,In_1693,In_1162);
nor U2449 (N_2449,In_392,In_206);
and U2450 (N_2450,In_1525,In_413);
and U2451 (N_2451,In_2492,In_292);
xor U2452 (N_2452,In_2812,In_2887);
nand U2453 (N_2453,In_2873,In_1730);
nor U2454 (N_2454,In_1163,In_2358);
nor U2455 (N_2455,In_1516,In_2973);
xnor U2456 (N_2456,In_2095,In_2758);
xor U2457 (N_2457,In_2676,In_1398);
nor U2458 (N_2458,In_1320,In_822);
nor U2459 (N_2459,In_344,In_2162);
xor U2460 (N_2460,In_2222,In_2882);
nor U2461 (N_2461,In_857,In_476);
xor U2462 (N_2462,In_1748,In_2162);
nor U2463 (N_2463,In_909,In_2631);
xor U2464 (N_2464,In_2925,In_1971);
xnor U2465 (N_2465,In_2387,In_865);
or U2466 (N_2466,In_1577,In_1665);
nor U2467 (N_2467,In_1576,In_1496);
or U2468 (N_2468,In_2809,In_1253);
xnor U2469 (N_2469,In_659,In_1836);
or U2470 (N_2470,In_1639,In_1650);
or U2471 (N_2471,In_682,In_1615);
nand U2472 (N_2472,In_2824,In_1384);
and U2473 (N_2473,In_592,In_2674);
xnor U2474 (N_2474,In_1150,In_767);
xnor U2475 (N_2475,In_1374,In_2841);
and U2476 (N_2476,In_1831,In_1602);
xnor U2477 (N_2477,In_103,In_977);
or U2478 (N_2478,In_2017,In_1284);
and U2479 (N_2479,In_156,In_574);
or U2480 (N_2480,In_2448,In_1120);
or U2481 (N_2481,In_124,In_1688);
nand U2482 (N_2482,In_1638,In_2528);
nor U2483 (N_2483,In_2446,In_955);
nand U2484 (N_2484,In_2255,In_2755);
and U2485 (N_2485,In_761,In_2906);
or U2486 (N_2486,In_1919,In_2768);
nand U2487 (N_2487,In_214,In_173);
or U2488 (N_2488,In_1128,In_1596);
and U2489 (N_2489,In_354,In_2621);
xnor U2490 (N_2490,In_1125,In_1691);
nor U2491 (N_2491,In_1579,In_2902);
xor U2492 (N_2492,In_1676,In_2211);
xor U2493 (N_2493,In_223,In_2472);
nor U2494 (N_2494,In_1218,In_1773);
and U2495 (N_2495,In_239,In_2397);
or U2496 (N_2496,In_1608,In_2839);
nand U2497 (N_2497,In_1191,In_1252);
xnor U2498 (N_2498,In_991,In_664);
nor U2499 (N_2499,In_1225,In_2135);
xor U2500 (N_2500,In_1015,In_2991);
and U2501 (N_2501,In_1666,In_666);
or U2502 (N_2502,In_2239,In_452);
nand U2503 (N_2503,In_2197,In_141);
nand U2504 (N_2504,In_733,In_1969);
xnor U2505 (N_2505,In_1479,In_989);
or U2506 (N_2506,In_628,In_1404);
nor U2507 (N_2507,In_402,In_332);
nand U2508 (N_2508,In_485,In_462);
and U2509 (N_2509,In_1597,In_1908);
xor U2510 (N_2510,In_2683,In_1933);
or U2511 (N_2511,In_1720,In_2628);
or U2512 (N_2512,In_968,In_1676);
xnor U2513 (N_2513,In_744,In_1785);
xnor U2514 (N_2514,In_2355,In_1780);
and U2515 (N_2515,In_446,In_1856);
nand U2516 (N_2516,In_1112,In_941);
or U2517 (N_2517,In_737,In_1504);
and U2518 (N_2518,In_557,In_1238);
or U2519 (N_2519,In_2163,In_2437);
xor U2520 (N_2520,In_781,In_2001);
xnor U2521 (N_2521,In_1046,In_909);
nand U2522 (N_2522,In_1442,In_2475);
and U2523 (N_2523,In_2029,In_270);
nand U2524 (N_2524,In_2040,In_560);
nor U2525 (N_2525,In_721,In_2524);
and U2526 (N_2526,In_6,In_330);
xor U2527 (N_2527,In_2777,In_589);
or U2528 (N_2528,In_324,In_1685);
xnor U2529 (N_2529,In_277,In_1794);
xor U2530 (N_2530,In_1169,In_393);
and U2531 (N_2531,In_926,In_1068);
xor U2532 (N_2532,In_2700,In_2849);
xnor U2533 (N_2533,In_1351,In_1533);
xor U2534 (N_2534,In_90,In_828);
or U2535 (N_2535,In_1497,In_509);
and U2536 (N_2536,In_1446,In_1092);
and U2537 (N_2537,In_1999,In_2271);
and U2538 (N_2538,In_351,In_874);
nand U2539 (N_2539,In_717,In_2288);
or U2540 (N_2540,In_428,In_2700);
nand U2541 (N_2541,In_306,In_1641);
and U2542 (N_2542,In_1365,In_1765);
xor U2543 (N_2543,In_2422,In_372);
nor U2544 (N_2544,In_1340,In_1776);
and U2545 (N_2545,In_875,In_1484);
nor U2546 (N_2546,In_2475,In_2073);
xnor U2547 (N_2547,In_119,In_1316);
and U2548 (N_2548,In_2526,In_580);
or U2549 (N_2549,In_576,In_2888);
xnor U2550 (N_2550,In_523,In_871);
nand U2551 (N_2551,In_756,In_2565);
nand U2552 (N_2552,In_239,In_2179);
and U2553 (N_2553,In_1260,In_768);
nand U2554 (N_2554,In_1493,In_2550);
xnor U2555 (N_2555,In_441,In_2066);
nand U2556 (N_2556,In_1472,In_2341);
nand U2557 (N_2557,In_2008,In_853);
nand U2558 (N_2558,In_1498,In_2802);
nor U2559 (N_2559,In_755,In_972);
nor U2560 (N_2560,In_107,In_1972);
nand U2561 (N_2561,In_998,In_1594);
and U2562 (N_2562,In_929,In_1932);
nor U2563 (N_2563,In_2536,In_892);
nand U2564 (N_2564,In_189,In_1284);
nand U2565 (N_2565,In_1778,In_666);
and U2566 (N_2566,In_1380,In_1286);
xnor U2567 (N_2567,In_626,In_1004);
nand U2568 (N_2568,In_1889,In_1747);
xnor U2569 (N_2569,In_1095,In_853);
and U2570 (N_2570,In_141,In_1040);
nand U2571 (N_2571,In_834,In_2828);
or U2572 (N_2572,In_413,In_740);
nand U2573 (N_2573,In_811,In_2037);
nand U2574 (N_2574,In_1827,In_2450);
xor U2575 (N_2575,In_565,In_2747);
nor U2576 (N_2576,In_2981,In_2584);
nand U2577 (N_2577,In_2013,In_2008);
xor U2578 (N_2578,In_2292,In_771);
nand U2579 (N_2579,In_1861,In_405);
and U2580 (N_2580,In_2849,In_1101);
nor U2581 (N_2581,In_2526,In_457);
nand U2582 (N_2582,In_1259,In_593);
nor U2583 (N_2583,In_2325,In_1131);
xnor U2584 (N_2584,In_2330,In_1326);
or U2585 (N_2585,In_1036,In_1372);
and U2586 (N_2586,In_106,In_689);
nand U2587 (N_2587,In_2127,In_1986);
and U2588 (N_2588,In_2318,In_2598);
or U2589 (N_2589,In_2727,In_2883);
nand U2590 (N_2590,In_2742,In_1015);
xnor U2591 (N_2591,In_2500,In_1003);
nor U2592 (N_2592,In_1173,In_2440);
nor U2593 (N_2593,In_1251,In_2247);
or U2594 (N_2594,In_1755,In_2698);
nor U2595 (N_2595,In_195,In_204);
nor U2596 (N_2596,In_2814,In_453);
or U2597 (N_2597,In_674,In_2013);
xor U2598 (N_2598,In_2542,In_1908);
nand U2599 (N_2599,In_160,In_415);
and U2600 (N_2600,In_1886,In_167);
xnor U2601 (N_2601,In_2686,In_466);
nor U2602 (N_2602,In_2269,In_2248);
nor U2603 (N_2603,In_2488,In_1966);
or U2604 (N_2604,In_355,In_2792);
nand U2605 (N_2605,In_2290,In_2775);
nand U2606 (N_2606,In_471,In_2522);
xnor U2607 (N_2607,In_2024,In_173);
nor U2608 (N_2608,In_353,In_1522);
or U2609 (N_2609,In_1847,In_2595);
and U2610 (N_2610,In_167,In_1345);
nor U2611 (N_2611,In_2407,In_2460);
nor U2612 (N_2612,In_2351,In_1365);
nor U2613 (N_2613,In_1134,In_155);
xnor U2614 (N_2614,In_609,In_1596);
or U2615 (N_2615,In_1242,In_2297);
xnor U2616 (N_2616,In_921,In_2823);
nand U2617 (N_2617,In_2210,In_459);
nor U2618 (N_2618,In_2530,In_1384);
nand U2619 (N_2619,In_183,In_76);
and U2620 (N_2620,In_621,In_742);
xnor U2621 (N_2621,In_1777,In_2513);
nand U2622 (N_2622,In_2587,In_1784);
nand U2623 (N_2623,In_494,In_2871);
nand U2624 (N_2624,In_598,In_388);
xnor U2625 (N_2625,In_2554,In_1505);
and U2626 (N_2626,In_646,In_24);
nor U2627 (N_2627,In_1542,In_116);
and U2628 (N_2628,In_1580,In_1291);
and U2629 (N_2629,In_2304,In_1447);
or U2630 (N_2630,In_1794,In_472);
xor U2631 (N_2631,In_1142,In_2534);
nand U2632 (N_2632,In_1327,In_2559);
nand U2633 (N_2633,In_577,In_144);
and U2634 (N_2634,In_82,In_454);
nand U2635 (N_2635,In_1512,In_1569);
nor U2636 (N_2636,In_653,In_2681);
or U2637 (N_2637,In_651,In_2384);
and U2638 (N_2638,In_242,In_1028);
nor U2639 (N_2639,In_2750,In_2463);
or U2640 (N_2640,In_2367,In_2457);
nor U2641 (N_2641,In_242,In_219);
xnor U2642 (N_2642,In_605,In_1543);
xnor U2643 (N_2643,In_246,In_1673);
and U2644 (N_2644,In_405,In_2580);
or U2645 (N_2645,In_764,In_2700);
nor U2646 (N_2646,In_1466,In_1089);
nand U2647 (N_2647,In_1827,In_529);
or U2648 (N_2648,In_1818,In_1296);
and U2649 (N_2649,In_2872,In_2986);
xnor U2650 (N_2650,In_1976,In_154);
and U2651 (N_2651,In_2127,In_2380);
nor U2652 (N_2652,In_2623,In_524);
or U2653 (N_2653,In_2516,In_495);
nor U2654 (N_2654,In_1431,In_2720);
or U2655 (N_2655,In_1004,In_1461);
nand U2656 (N_2656,In_2508,In_354);
xor U2657 (N_2657,In_1671,In_2867);
and U2658 (N_2658,In_2235,In_1612);
nor U2659 (N_2659,In_846,In_2696);
xor U2660 (N_2660,In_2680,In_2785);
or U2661 (N_2661,In_1967,In_2263);
or U2662 (N_2662,In_1927,In_2578);
or U2663 (N_2663,In_971,In_1786);
and U2664 (N_2664,In_1471,In_2688);
nor U2665 (N_2665,In_165,In_1167);
or U2666 (N_2666,In_1662,In_2194);
xnor U2667 (N_2667,In_62,In_2387);
xor U2668 (N_2668,In_465,In_2646);
xor U2669 (N_2669,In_2262,In_552);
or U2670 (N_2670,In_988,In_904);
xnor U2671 (N_2671,In_1127,In_847);
nand U2672 (N_2672,In_1730,In_877);
nor U2673 (N_2673,In_2464,In_2627);
xnor U2674 (N_2674,In_739,In_2431);
or U2675 (N_2675,In_1155,In_715);
nor U2676 (N_2676,In_1692,In_2352);
nor U2677 (N_2677,In_1609,In_1015);
and U2678 (N_2678,In_2307,In_1161);
nor U2679 (N_2679,In_2391,In_2477);
nand U2680 (N_2680,In_1864,In_334);
or U2681 (N_2681,In_1776,In_1632);
or U2682 (N_2682,In_2373,In_2781);
nor U2683 (N_2683,In_1086,In_2597);
xor U2684 (N_2684,In_861,In_2761);
or U2685 (N_2685,In_1316,In_1716);
or U2686 (N_2686,In_942,In_2588);
nor U2687 (N_2687,In_1453,In_1975);
or U2688 (N_2688,In_1050,In_1039);
nand U2689 (N_2689,In_200,In_887);
and U2690 (N_2690,In_374,In_1299);
xnor U2691 (N_2691,In_61,In_2347);
xnor U2692 (N_2692,In_214,In_2962);
nand U2693 (N_2693,In_2010,In_1575);
and U2694 (N_2694,In_703,In_1341);
nand U2695 (N_2695,In_2374,In_2559);
and U2696 (N_2696,In_1340,In_1855);
nor U2697 (N_2697,In_1846,In_1589);
and U2698 (N_2698,In_1196,In_331);
nand U2699 (N_2699,In_1817,In_1409);
nand U2700 (N_2700,In_1698,In_1314);
xor U2701 (N_2701,In_1815,In_865);
nor U2702 (N_2702,In_988,In_2449);
and U2703 (N_2703,In_1526,In_1097);
and U2704 (N_2704,In_1597,In_656);
or U2705 (N_2705,In_237,In_8);
and U2706 (N_2706,In_448,In_2671);
or U2707 (N_2707,In_2600,In_1717);
nor U2708 (N_2708,In_261,In_1225);
nand U2709 (N_2709,In_1498,In_1649);
nand U2710 (N_2710,In_2931,In_38);
and U2711 (N_2711,In_2981,In_1884);
xor U2712 (N_2712,In_1720,In_2287);
nand U2713 (N_2713,In_645,In_574);
or U2714 (N_2714,In_2146,In_1547);
xor U2715 (N_2715,In_2278,In_1257);
or U2716 (N_2716,In_551,In_2800);
or U2717 (N_2717,In_1097,In_981);
nand U2718 (N_2718,In_2179,In_278);
and U2719 (N_2719,In_462,In_1345);
nand U2720 (N_2720,In_2324,In_1804);
and U2721 (N_2721,In_1231,In_1017);
nand U2722 (N_2722,In_2105,In_1860);
or U2723 (N_2723,In_302,In_2964);
nand U2724 (N_2724,In_1566,In_2674);
xor U2725 (N_2725,In_2319,In_1282);
nor U2726 (N_2726,In_2016,In_527);
or U2727 (N_2727,In_937,In_2938);
or U2728 (N_2728,In_1154,In_2964);
nor U2729 (N_2729,In_661,In_685);
nand U2730 (N_2730,In_2414,In_501);
nor U2731 (N_2731,In_79,In_1114);
and U2732 (N_2732,In_907,In_1321);
nand U2733 (N_2733,In_537,In_1712);
nor U2734 (N_2734,In_1030,In_812);
xor U2735 (N_2735,In_970,In_2087);
or U2736 (N_2736,In_2334,In_1993);
nor U2737 (N_2737,In_1703,In_535);
nor U2738 (N_2738,In_1191,In_2713);
and U2739 (N_2739,In_2331,In_1425);
xnor U2740 (N_2740,In_2206,In_2150);
xor U2741 (N_2741,In_1836,In_2830);
nor U2742 (N_2742,In_1522,In_2092);
nor U2743 (N_2743,In_2644,In_2280);
and U2744 (N_2744,In_515,In_1299);
nand U2745 (N_2745,In_438,In_2317);
nor U2746 (N_2746,In_2652,In_1023);
nor U2747 (N_2747,In_677,In_2276);
nand U2748 (N_2748,In_2899,In_2157);
xor U2749 (N_2749,In_2719,In_616);
or U2750 (N_2750,In_325,In_2710);
or U2751 (N_2751,In_127,In_1022);
nor U2752 (N_2752,In_2913,In_1633);
nor U2753 (N_2753,In_2246,In_2017);
nand U2754 (N_2754,In_1266,In_207);
and U2755 (N_2755,In_2257,In_2522);
nor U2756 (N_2756,In_1900,In_1710);
and U2757 (N_2757,In_102,In_839);
or U2758 (N_2758,In_1184,In_168);
and U2759 (N_2759,In_2011,In_1387);
and U2760 (N_2760,In_679,In_300);
xnor U2761 (N_2761,In_2478,In_1655);
xor U2762 (N_2762,In_145,In_703);
xor U2763 (N_2763,In_1119,In_150);
nor U2764 (N_2764,In_2271,In_1928);
nand U2765 (N_2765,In_1786,In_2139);
nand U2766 (N_2766,In_1303,In_438);
xnor U2767 (N_2767,In_1957,In_684);
and U2768 (N_2768,In_2090,In_1578);
xnor U2769 (N_2769,In_2774,In_623);
nand U2770 (N_2770,In_2703,In_2542);
nor U2771 (N_2771,In_1732,In_1164);
or U2772 (N_2772,In_1795,In_121);
xnor U2773 (N_2773,In_1986,In_1783);
or U2774 (N_2774,In_796,In_2804);
xor U2775 (N_2775,In_2616,In_2895);
nand U2776 (N_2776,In_143,In_2125);
or U2777 (N_2777,In_2367,In_38);
nand U2778 (N_2778,In_2977,In_2171);
and U2779 (N_2779,In_2505,In_2814);
or U2780 (N_2780,In_2492,In_1063);
or U2781 (N_2781,In_2356,In_2561);
xnor U2782 (N_2782,In_1895,In_2110);
xor U2783 (N_2783,In_393,In_2654);
xor U2784 (N_2784,In_1999,In_2208);
and U2785 (N_2785,In_288,In_2310);
or U2786 (N_2786,In_1677,In_78);
and U2787 (N_2787,In_2518,In_2601);
or U2788 (N_2788,In_1496,In_2826);
or U2789 (N_2789,In_1504,In_1411);
nand U2790 (N_2790,In_192,In_265);
nor U2791 (N_2791,In_2539,In_1272);
and U2792 (N_2792,In_509,In_2621);
xnor U2793 (N_2793,In_2139,In_2024);
or U2794 (N_2794,In_2479,In_121);
or U2795 (N_2795,In_1179,In_2491);
xor U2796 (N_2796,In_2108,In_1377);
xor U2797 (N_2797,In_78,In_37);
or U2798 (N_2798,In_1423,In_2031);
nor U2799 (N_2799,In_1085,In_526);
nor U2800 (N_2800,In_399,In_1387);
or U2801 (N_2801,In_2146,In_844);
and U2802 (N_2802,In_1359,In_2020);
and U2803 (N_2803,In_408,In_718);
and U2804 (N_2804,In_1625,In_2830);
nand U2805 (N_2805,In_2245,In_2156);
and U2806 (N_2806,In_2437,In_1226);
nor U2807 (N_2807,In_584,In_2874);
nor U2808 (N_2808,In_2185,In_307);
and U2809 (N_2809,In_2213,In_1158);
and U2810 (N_2810,In_1082,In_2671);
xor U2811 (N_2811,In_2667,In_732);
or U2812 (N_2812,In_2687,In_2109);
nor U2813 (N_2813,In_2518,In_1147);
xnor U2814 (N_2814,In_328,In_2999);
nor U2815 (N_2815,In_220,In_767);
xor U2816 (N_2816,In_1472,In_742);
nor U2817 (N_2817,In_1787,In_449);
xnor U2818 (N_2818,In_683,In_1995);
nor U2819 (N_2819,In_2878,In_1979);
and U2820 (N_2820,In_212,In_1010);
and U2821 (N_2821,In_169,In_632);
or U2822 (N_2822,In_2801,In_2899);
nand U2823 (N_2823,In_839,In_2362);
and U2824 (N_2824,In_1173,In_538);
nor U2825 (N_2825,In_2440,In_617);
nand U2826 (N_2826,In_2252,In_2612);
nand U2827 (N_2827,In_192,In_2611);
nor U2828 (N_2828,In_2610,In_1996);
nand U2829 (N_2829,In_1098,In_674);
or U2830 (N_2830,In_2834,In_185);
and U2831 (N_2831,In_1391,In_2356);
xnor U2832 (N_2832,In_2441,In_984);
xor U2833 (N_2833,In_2474,In_2703);
and U2834 (N_2834,In_889,In_1778);
xor U2835 (N_2835,In_270,In_1846);
nand U2836 (N_2836,In_2890,In_346);
xor U2837 (N_2837,In_2908,In_1431);
and U2838 (N_2838,In_1654,In_1033);
or U2839 (N_2839,In_430,In_1752);
nor U2840 (N_2840,In_2912,In_1768);
xnor U2841 (N_2841,In_284,In_1551);
nand U2842 (N_2842,In_1086,In_935);
or U2843 (N_2843,In_913,In_219);
nor U2844 (N_2844,In_2221,In_1124);
nand U2845 (N_2845,In_1597,In_86);
xnor U2846 (N_2846,In_664,In_1341);
and U2847 (N_2847,In_887,In_2794);
xor U2848 (N_2848,In_873,In_24);
and U2849 (N_2849,In_318,In_494);
or U2850 (N_2850,In_278,In_43);
nand U2851 (N_2851,In_2348,In_1838);
xnor U2852 (N_2852,In_2054,In_2460);
nor U2853 (N_2853,In_2117,In_2017);
nand U2854 (N_2854,In_2746,In_2005);
nor U2855 (N_2855,In_2474,In_1777);
and U2856 (N_2856,In_1281,In_1014);
or U2857 (N_2857,In_2134,In_2532);
nor U2858 (N_2858,In_1563,In_8);
or U2859 (N_2859,In_1,In_700);
or U2860 (N_2860,In_1944,In_1592);
or U2861 (N_2861,In_2376,In_2325);
nor U2862 (N_2862,In_174,In_708);
xor U2863 (N_2863,In_407,In_258);
nand U2864 (N_2864,In_1773,In_1285);
nand U2865 (N_2865,In_2941,In_2720);
xnor U2866 (N_2866,In_2326,In_970);
nand U2867 (N_2867,In_317,In_2557);
nor U2868 (N_2868,In_1719,In_1810);
nor U2869 (N_2869,In_1981,In_1097);
nor U2870 (N_2870,In_1811,In_2494);
nor U2871 (N_2871,In_2964,In_804);
and U2872 (N_2872,In_697,In_2925);
nor U2873 (N_2873,In_703,In_2329);
nand U2874 (N_2874,In_589,In_649);
or U2875 (N_2875,In_797,In_296);
nor U2876 (N_2876,In_1243,In_498);
nand U2877 (N_2877,In_1870,In_977);
or U2878 (N_2878,In_7,In_591);
or U2879 (N_2879,In_1972,In_1019);
nand U2880 (N_2880,In_1984,In_1414);
or U2881 (N_2881,In_389,In_249);
or U2882 (N_2882,In_268,In_2854);
nand U2883 (N_2883,In_464,In_523);
or U2884 (N_2884,In_2686,In_1779);
nand U2885 (N_2885,In_654,In_1078);
nand U2886 (N_2886,In_2699,In_1119);
or U2887 (N_2887,In_2890,In_1910);
xor U2888 (N_2888,In_1210,In_537);
or U2889 (N_2889,In_907,In_1997);
and U2890 (N_2890,In_1655,In_1487);
xnor U2891 (N_2891,In_2506,In_2166);
and U2892 (N_2892,In_2992,In_1810);
nand U2893 (N_2893,In_2441,In_2745);
nand U2894 (N_2894,In_292,In_2465);
and U2895 (N_2895,In_47,In_864);
or U2896 (N_2896,In_497,In_2287);
xnor U2897 (N_2897,In_1257,In_576);
nor U2898 (N_2898,In_353,In_2552);
nand U2899 (N_2899,In_2992,In_2383);
and U2900 (N_2900,In_1181,In_681);
nor U2901 (N_2901,In_2325,In_560);
nand U2902 (N_2902,In_2267,In_2797);
or U2903 (N_2903,In_2893,In_2656);
nor U2904 (N_2904,In_1404,In_2062);
nor U2905 (N_2905,In_1787,In_2544);
xnor U2906 (N_2906,In_2158,In_2179);
and U2907 (N_2907,In_1789,In_596);
nand U2908 (N_2908,In_2466,In_510);
xnor U2909 (N_2909,In_2679,In_455);
xnor U2910 (N_2910,In_1000,In_1745);
nand U2911 (N_2911,In_285,In_1549);
or U2912 (N_2912,In_5,In_912);
nand U2913 (N_2913,In_2622,In_1599);
and U2914 (N_2914,In_2216,In_1571);
and U2915 (N_2915,In_437,In_1519);
xnor U2916 (N_2916,In_1413,In_2897);
xor U2917 (N_2917,In_80,In_1912);
and U2918 (N_2918,In_448,In_1890);
nor U2919 (N_2919,In_1155,In_1104);
and U2920 (N_2920,In_2228,In_1424);
nand U2921 (N_2921,In_2533,In_63);
nor U2922 (N_2922,In_103,In_573);
and U2923 (N_2923,In_1940,In_2318);
or U2924 (N_2924,In_284,In_1606);
and U2925 (N_2925,In_366,In_230);
nand U2926 (N_2926,In_343,In_1073);
nand U2927 (N_2927,In_2278,In_625);
nand U2928 (N_2928,In_2519,In_2737);
nor U2929 (N_2929,In_251,In_2904);
and U2930 (N_2930,In_2175,In_2472);
nand U2931 (N_2931,In_1395,In_2330);
xnor U2932 (N_2932,In_782,In_1421);
or U2933 (N_2933,In_2513,In_601);
or U2934 (N_2934,In_765,In_247);
nand U2935 (N_2935,In_2288,In_2348);
or U2936 (N_2936,In_2261,In_2230);
and U2937 (N_2937,In_1294,In_2011);
or U2938 (N_2938,In_436,In_1471);
nor U2939 (N_2939,In_82,In_388);
nor U2940 (N_2940,In_1398,In_1892);
nor U2941 (N_2941,In_0,In_2776);
nor U2942 (N_2942,In_2614,In_1863);
or U2943 (N_2943,In_1577,In_159);
xnor U2944 (N_2944,In_2193,In_1171);
and U2945 (N_2945,In_2496,In_2579);
xor U2946 (N_2946,In_1983,In_426);
nor U2947 (N_2947,In_574,In_1733);
nor U2948 (N_2948,In_1487,In_2433);
and U2949 (N_2949,In_1009,In_1862);
xor U2950 (N_2950,In_2111,In_1911);
or U2951 (N_2951,In_2731,In_1590);
and U2952 (N_2952,In_1206,In_396);
nand U2953 (N_2953,In_1678,In_541);
xor U2954 (N_2954,In_108,In_1881);
xor U2955 (N_2955,In_2530,In_2123);
or U2956 (N_2956,In_1899,In_2823);
nand U2957 (N_2957,In_1196,In_883);
xor U2958 (N_2958,In_559,In_330);
xor U2959 (N_2959,In_257,In_967);
or U2960 (N_2960,In_2297,In_2031);
nor U2961 (N_2961,In_2569,In_2628);
xor U2962 (N_2962,In_606,In_2247);
xnor U2963 (N_2963,In_1948,In_2221);
or U2964 (N_2964,In_656,In_2166);
nor U2965 (N_2965,In_959,In_954);
or U2966 (N_2966,In_2763,In_507);
and U2967 (N_2967,In_1483,In_2742);
nor U2968 (N_2968,In_2795,In_16);
nand U2969 (N_2969,In_1347,In_2882);
and U2970 (N_2970,In_399,In_2473);
and U2971 (N_2971,In_1713,In_36);
or U2972 (N_2972,In_2099,In_1129);
and U2973 (N_2973,In_135,In_1491);
and U2974 (N_2974,In_1298,In_427);
xnor U2975 (N_2975,In_1386,In_651);
nand U2976 (N_2976,In_1985,In_1174);
or U2977 (N_2977,In_1264,In_345);
xnor U2978 (N_2978,In_548,In_460);
and U2979 (N_2979,In_905,In_2978);
or U2980 (N_2980,In_2777,In_919);
and U2981 (N_2981,In_2721,In_2464);
xnor U2982 (N_2982,In_1025,In_37);
xnor U2983 (N_2983,In_232,In_2700);
nand U2984 (N_2984,In_444,In_2939);
nand U2985 (N_2985,In_773,In_2634);
and U2986 (N_2986,In_1109,In_1349);
or U2987 (N_2987,In_626,In_31);
xnor U2988 (N_2988,In_1672,In_2981);
xor U2989 (N_2989,In_1011,In_1822);
and U2990 (N_2990,In_881,In_1857);
and U2991 (N_2991,In_776,In_748);
and U2992 (N_2992,In_2984,In_942);
or U2993 (N_2993,In_2637,In_2397);
nor U2994 (N_2994,In_2971,In_241);
nand U2995 (N_2995,In_261,In_1925);
and U2996 (N_2996,In_2660,In_1913);
xor U2997 (N_2997,In_65,In_447);
or U2998 (N_2998,In_1865,In_2922);
or U2999 (N_2999,In_1001,In_2074);
and U3000 (N_3000,In_1830,In_986);
xnor U3001 (N_3001,In_2807,In_1569);
nand U3002 (N_3002,In_530,In_1589);
nand U3003 (N_3003,In_91,In_436);
nor U3004 (N_3004,In_2617,In_1532);
and U3005 (N_3005,In_1895,In_2564);
or U3006 (N_3006,In_2005,In_1275);
nor U3007 (N_3007,In_1100,In_1038);
xor U3008 (N_3008,In_1075,In_801);
xnor U3009 (N_3009,In_657,In_2358);
or U3010 (N_3010,In_1311,In_1707);
xnor U3011 (N_3011,In_747,In_2517);
nand U3012 (N_3012,In_2119,In_1683);
or U3013 (N_3013,In_2228,In_2645);
nor U3014 (N_3014,In_1078,In_1373);
nor U3015 (N_3015,In_800,In_850);
or U3016 (N_3016,In_1537,In_782);
nand U3017 (N_3017,In_2007,In_875);
nor U3018 (N_3018,In_2218,In_2724);
or U3019 (N_3019,In_986,In_2151);
or U3020 (N_3020,In_2488,In_2820);
and U3021 (N_3021,In_2594,In_1114);
nor U3022 (N_3022,In_2545,In_1392);
nor U3023 (N_3023,In_217,In_2857);
or U3024 (N_3024,In_199,In_2773);
xnor U3025 (N_3025,In_550,In_1284);
nor U3026 (N_3026,In_412,In_1044);
xor U3027 (N_3027,In_50,In_2872);
nor U3028 (N_3028,In_2672,In_1529);
or U3029 (N_3029,In_1250,In_1684);
nor U3030 (N_3030,In_2075,In_2310);
and U3031 (N_3031,In_2330,In_2765);
xor U3032 (N_3032,In_1014,In_1715);
nor U3033 (N_3033,In_1008,In_1799);
or U3034 (N_3034,In_1060,In_1753);
nor U3035 (N_3035,In_1425,In_2209);
and U3036 (N_3036,In_1697,In_2977);
or U3037 (N_3037,In_2722,In_2681);
and U3038 (N_3038,In_2436,In_2440);
or U3039 (N_3039,In_1611,In_237);
xor U3040 (N_3040,In_310,In_1131);
nor U3041 (N_3041,In_1964,In_1881);
nand U3042 (N_3042,In_1028,In_1832);
xnor U3043 (N_3043,In_1874,In_2679);
nor U3044 (N_3044,In_952,In_28);
nor U3045 (N_3045,In_887,In_547);
nand U3046 (N_3046,In_2371,In_2564);
nand U3047 (N_3047,In_514,In_1104);
and U3048 (N_3048,In_1048,In_705);
nor U3049 (N_3049,In_842,In_1752);
or U3050 (N_3050,In_549,In_144);
nor U3051 (N_3051,In_2641,In_686);
or U3052 (N_3052,In_1700,In_559);
nand U3053 (N_3053,In_405,In_2507);
xor U3054 (N_3054,In_1220,In_2330);
and U3055 (N_3055,In_1500,In_952);
and U3056 (N_3056,In_297,In_2410);
xor U3057 (N_3057,In_1440,In_969);
xnor U3058 (N_3058,In_362,In_768);
xnor U3059 (N_3059,In_2071,In_982);
nor U3060 (N_3060,In_2080,In_1250);
nand U3061 (N_3061,In_358,In_1798);
or U3062 (N_3062,In_2261,In_945);
and U3063 (N_3063,In_6,In_2247);
nand U3064 (N_3064,In_23,In_1391);
nand U3065 (N_3065,In_602,In_2287);
or U3066 (N_3066,In_2076,In_2244);
or U3067 (N_3067,In_221,In_1595);
nand U3068 (N_3068,In_1503,In_2786);
xnor U3069 (N_3069,In_1359,In_477);
and U3070 (N_3070,In_122,In_1643);
nor U3071 (N_3071,In_628,In_2309);
or U3072 (N_3072,In_2966,In_1035);
or U3073 (N_3073,In_2605,In_2968);
and U3074 (N_3074,In_2829,In_1156);
nand U3075 (N_3075,In_2816,In_1911);
or U3076 (N_3076,In_1509,In_2477);
or U3077 (N_3077,In_1595,In_2524);
or U3078 (N_3078,In_1325,In_629);
nor U3079 (N_3079,In_1244,In_2636);
or U3080 (N_3080,In_1167,In_2417);
or U3081 (N_3081,In_2545,In_408);
nand U3082 (N_3082,In_1499,In_1907);
xor U3083 (N_3083,In_2991,In_2782);
xor U3084 (N_3084,In_2904,In_326);
nand U3085 (N_3085,In_1722,In_2966);
or U3086 (N_3086,In_2241,In_1199);
xnor U3087 (N_3087,In_1040,In_1951);
and U3088 (N_3088,In_1802,In_1396);
nand U3089 (N_3089,In_611,In_624);
or U3090 (N_3090,In_2805,In_2370);
nand U3091 (N_3091,In_2244,In_714);
and U3092 (N_3092,In_119,In_2043);
or U3093 (N_3093,In_391,In_1016);
and U3094 (N_3094,In_726,In_2370);
xnor U3095 (N_3095,In_2938,In_413);
and U3096 (N_3096,In_2066,In_836);
or U3097 (N_3097,In_1823,In_956);
nor U3098 (N_3098,In_2903,In_2673);
nand U3099 (N_3099,In_2108,In_2435);
nor U3100 (N_3100,In_497,In_254);
nor U3101 (N_3101,In_221,In_832);
xnor U3102 (N_3102,In_1753,In_2534);
and U3103 (N_3103,In_2412,In_2472);
or U3104 (N_3104,In_2439,In_282);
xor U3105 (N_3105,In_1395,In_1298);
nor U3106 (N_3106,In_942,In_2431);
or U3107 (N_3107,In_1990,In_301);
or U3108 (N_3108,In_2238,In_1315);
nor U3109 (N_3109,In_1725,In_1557);
nand U3110 (N_3110,In_312,In_1494);
xnor U3111 (N_3111,In_1823,In_2124);
nand U3112 (N_3112,In_1795,In_1557);
nor U3113 (N_3113,In_472,In_613);
nand U3114 (N_3114,In_1453,In_1841);
or U3115 (N_3115,In_2585,In_1123);
nand U3116 (N_3116,In_43,In_390);
and U3117 (N_3117,In_644,In_2246);
nand U3118 (N_3118,In_366,In_532);
nor U3119 (N_3119,In_460,In_528);
nand U3120 (N_3120,In_2736,In_282);
xor U3121 (N_3121,In_27,In_2142);
or U3122 (N_3122,In_1556,In_2558);
nand U3123 (N_3123,In_2566,In_2002);
xor U3124 (N_3124,In_665,In_1386);
and U3125 (N_3125,In_2952,In_1397);
nand U3126 (N_3126,In_1179,In_168);
or U3127 (N_3127,In_1260,In_1601);
nor U3128 (N_3128,In_277,In_1309);
nor U3129 (N_3129,In_1923,In_655);
xor U3130 (N_3130,In_1717,In_1803);
or U3131 (N_3131,In_1322,In_1278);
nor U3132 (N_3132,In_1778,In_2777);
and U3133 (N_3133,In_1705,In_495);
nor U3134 (N_3134,In_357,In_269);
nand U3135 (N_3135,In_2051,In_740);
xor U3136 (N_3136,In_589,In_110);
and U3137 (N_3137,In_204,In_663);
nand U3138 (N_3138,In_2236,In_2173);
nor U3139 (N_3139,In_2233,In_1313);
xnor U3140 (N_3140,In_2823,In_2522);
nor U3141 (N_3141,In_1671,In_2718);
nand U3142 (N_3142,In_829,In_2324);
or U3143 (N_3143,In_357,In_1936);
nand U3144 (N_3144,In_271,In_1089);
nand U3145 (N_3145,In_543,In_1337);
nand U3146 (N_3146,In_2322,In_932);
nand U3147 (N_3147,In_2439,In_1240);
nand U3148 (N_3148,In_1319,In_841);
and U3149 (N_3149,In_286,In_719);
and U3150 (N_3150,In_133,In_933);
and U3151 (N_3151,In_1772,In_85);
nor U3152 (N_3152,In_2857,In_2895);
nor U3153 (N_3153,In_2363,In_322);
nor U3154 (N_3154,In_1683,In_32);
xor U3155 (N_3155,In_652,In_2637);
nand U3156 (N_3156,In_2977,In_2659);
nor U3157 (N_3157,In_97,In_2706);
nor U3158 (N_3158,In_1815,In_1739);
and U3159 (N_3159,In_999,In_1014);
nor U3160 (N_3160,In_857,In_2566);
or U3161 (N_3161,In_1705,In_2745);
nor U3162 (N_3162,In_2188,In_2849);
nand U3163 (N_3163,In_2880,In_2896);
xor U3164 (N_3164,In_1994,In_1688);
nor U3165 (N_3165,In_335,In_2723);
or U3166 (N_3166,In_68,In_1954);
and U3167 (N_3167,In_371,In_2618);
xnor U3168 (N_3168,In_2321,In_1955);
or U3169 (N_3169,In_363,In_1509);
or U3170 (N_3170,In_1469,In_672);
and U3171 (N_3171,In_440,In_908);
nor U3172 (N_3172,In_2364,In_2570);
and U3173 (N_3173,In_2236,In_1583);
or U3174 (N_3174,In_1059,In_2144);
nand U3175 (N_3175,In_1882,In_2694);
or U3176 (N_3176,In_147,In_2649);
nand U3177 (N_3177,In_1322,In_639);
xor U3178 (N_3178,In_2441,In_24);
and U3179 (N_3179,In_1821,In_2436);
and U3180 (N_3180,In_325,In_927);
nor U3181 (N_3181,In_198,In_2060);
nand U3182 (N_3182,In_1672,In_2912);
nand U3183 (N_3183,In_2554,In_1127);
nor U3184 (N_3184,In_1138,In_2002);
xor U3185 (N_3185,In_42,In_1120);
and U3186 (N_3186,In_1792,In_217);
nand U3187 (N_3187,In_763,In_2414);
or U3188 (N_3188,In_2979,In_2711);
nor U3189 (N_3189,In_1682,In_2824);
nand U3190 (N_3190,In_1450,In_1417);
xnor U3191 (N_3191,In_1045,In_2903);
nor U3192 (N_3192,In_1573,In_2659);
nand U3193 (N_3193,In_1215,In_8);
nor U3194 (N_3194,In_2447,In_2741);
nand U3195 (N_3195,In_2472,In_1403);
nor U3196 (N_3196,In_2019,In_648);
and U3197 (N_3197,In_2509,In_1041);
nor U3198 (N_3198,In_1324,In_1085);
or U3199 (N_3199,In_405,In_2176);
nand U3200 (N_3200,In_880,In_1730);
nand U3201 (N_3201,In_2965,In_536);
or U3202 (N_3202,In_356,In_1726);
nor U3203 (N_3203,In_1613,In_60);
nor U3204 (N_3204,In_2096,In_1003);
nor U3205 (N_3205,In_806,In_1662);
xor U3206 (N_3206,In_489,In_2290);
nor U3207 (N_3207,In_2553,In_1424);
nand U3208 (N_3208,In_1215,In_2308);
nor U3209 (N_3209,In_158,In_505);
and U3210 (N_3210,In_1335,In_2412);
nor U3211 (N_3211,In_1877,In_2860);
nor U3212 (N_3212,In_414,In_1633);
xnor U3213 (N_3213,In_1280,In_362);
and U3214 (N_3214,In_719,In_2840);
nand U3215 (N_3215,In_2504,In_2250);
or U3216 (N_3216,In_636,In_273);
and U3217 (N_3217,In_890,In_981);
or U3218 (N_3218,In_1405,In_1088);
xor U3219 (N_3219,In_2763,In_271);
xor U3220 (N_3220,In_1362,In_2645);
xnor U3221 (N_3221,In_1994,In_3);
nand U3222 (N_3222,In_1493,In_2659);
nor U3223 (N_3223,In_2942,In_1528);
or U3224 (N_3224,In_2905,In_1560);
xor U3225 (N_3225,In_2049,In_1945);
nor U3226 (N_3226,In_788,In_1342);
and U3227 (N_3227,In_999,In_2775);
nor U3228 (N_3228,In_362,In_2616);
nor U3229 (N_3229,In_986,In_1085);
xor U3230 (N_3230,In_2539,In_2244);
xor U3231 (N_3231,In_382,In_726);
xor U3232 (N_3232,In_2145,In_2857);
and U3233 (N_3233,In_2721,In_2225);
xnor U3234 (N_3234,In_1470,In_867);
or U3235 (N_3235,In_2605,In_1026);
xnor U3236 (N_3236,In_1055,In_2279);
nand U3237 (N_3237,In_2043,In_2508);
nand U3238 (N_3238,In_1359,In_1447);
nor U3239 (N_3239,In_948,In_2607);
nor U3240 (N_3240,In_2760,In_2236);
or U3241 (N_3241,In_2262,In_362);
or U3242 (N_3242,In_556,In_1117);
nor U3243 (N_3243,In_171,In_1010);
xor U3244 (N_3244,In_1197,In_403);
and U3245 (N_3245,In_1736,In_1998);
xnor U3246 (N_3246,In_1748,In_29);
nand U3247 (N_3247,In_2809,In_2571);
xnor U3248 (N_3248,In_1220,In_1975);
xnor U3249 (N_3249,In_2999,In_267);
or U3250 (N_3250,In_236,In_339);
nand U3251 (N_3251,In_71,In_1546);
or U3252 (N_3252,In_1620,In_1095);
nor U3253 (N_3253,In_2111,In_353);
or U3254 (N_3254,In_1588,In_2745);
nand U3255 (N_3255,In_479,In_1212);
or U3256 (N_3256,In_793,In_1406);
xnor U3257 (N_3257,In_2665,In_1034);
and U3258 (N_3258,In_901,In_112);
nand U3259 (N_3259,In_241,In_2801);
nor U3260 (N_3260,In_1913,In_413);
nor U3261 (N_3261,In_965,In_833);
nand U3262 (N_3262,In_401,In_2113);
or U3263 (N_3263,In_1767,In_601);
nor U3264 (N_3264,In_2143,In_1246);
or U3265 (N_3265,In_943,In_1832);
nand U3266 (N_3266,In_1792,In_1741);
nor U3267 (N_3267,In_2288,In_746);
nor U3268 (N_3268,In_412,In_2704);
xor U3269 (N_3269,In_971,In_1231);
or U3270 (N_3270,In_2405,In_2075);
nor U3271 (N_3271,In_828,In_2363);
nand U3272 (N_3272,In_1317,In_2840);
nand U3273 (N_3273,In_2393,In_2651);
or U3274 (N_3274,In_2810,In_17);
nand U3275 (N_3275,In_542,In_189);
and U3276 (N_3276,In_1084,In_2174);
nand U3277 (N_3277,In_2903,In_1844);
and U3278 (N_3278,In_2478,In_2590);
nand U3279 (N_3279,In_1995,In_2484);
nand U3280 (N_3280,In_2241,In_2239);
xnor U3281 (N_3281,In_1482,In_134);
nand U3282 (N_3282,In_2292,In_2350);
and U3283 (N_3283,In_1773,In_1923);
and U3284 (N_3284,In_1648,In_1681);
nand U3285 (N_3285,In_2348,In_163);
or U3286 (N_3286,In_2731,In_1760);
nand U3287 (N_3287,In_907,In_2566);
nand U3288 (N_3288,In_2191,In_2045);
xor U3289 (N_3289,In_1383,In_2734);
xnor U3290 (N_3290,In_737,In_1657);
xnor U3291 (N_3291,In_1728,In_1049);
or U3292 (N_3292,In_2942,In_1752);
xor U3293 (N_3293,In_836,In_1555);
nor U3294 (N_3294,In_380,In_770);
nor U3295 (N_3295,In_2041,In_2088);
nand U3296 (N_3296,In_2793,In_2539);
or U3297 (N_3297,In_2794,In_2405);
xor U3298 (N_3298,In_2932,In_1354);
xnor U3299 (N_3299,In_1997,In_1186);
nand U3300 (N_3300,In_1315,In_186);
nand U3301 (N_3301,In_701,In_1067);
xnor U3302 (N_3302,In_2122,In_1710);
and U3303 (N_3303,In_530,In_1270);
and U3304 (N_3304,In_2634,In_2492);
xnor U3305 (N_3305,In_727,In_1778);
nor U3306 (N_3306,In_541,In_2455);
xor U3307 (N_3307,In_2790,In_392);
or U3308 (N_3308,In_2776,In_2519);
xnor U3309 (N_3309,In_102,In_2908);
nand U3310 (N_3310,In_2552,In_104);
and U3311 (N_3311,In_421,In_1284);
or U3312 (N_3312,In_1169,In_1858);
or U3313 (N_3313,In_247,In_761);
xor U3314 (N_3314,In_1450,In_1685);
and U3315 (N_3315,In_180,In_1329);
xor U3316 (N_3316,In_1043,In_57);
nand U3317 (N_3317,In_782,In_933);
nand U3318 (N_3318,In_2821,In_912);
or U3319 (N_3319,In_880,In_1755);
or U3320 (N_3320,In_191,In_2776);
nor U3321 (N_3321,In_1154,In_2551);
xor U3322 (N_3322,In_403,In_2920);
and U3323 (N_3323,In_307,In_1670);
or U3324 (N_3324,In_1534,In_958);
xor U3325 (N_3325,In_2057,In_2694);
or U3326 (N_3326,In_157,In_932);
nor U3327 (N_3327,In_2118,In_988);
nor U3328 (N_3328,In_247,In_107);
nand U3329 (N_3329,In_889,In_725);
or U3330 (N_3330,In_226,In_2399);
xor U3331 (N_3331,In_2435,In_2493);
nand U3332 (N_3332,In_1140,In_1808);
xor U3333 (N_3333,In_2318,In_600);
and U3334 (N_3334,In_2074,In_2989);
nand U3335 (N_3335,In_288,In_1939);
nor U3336 (N_3336,In_2861,In_1451);
xnor U3337 (N_3337,In_1695,In_868);
xor U3338 (N_3338,In_2102,In_1102);
and U3339 (N_3339,In_2778,In_1232);
xnor U3340 (N_3340,In_2115,In_1035);
xnor U3341 (N_3341,In_301,In_564);
nor U3342 (N_3342,In_876,In_2477);
nand U3343 (N_3343,In_2978,In_1520);
xnor U3344 (N_3344,In_2369,In_455);
and U3345 (N_3345,In_846,In_2987);
nor U3346 (N_3346,In_2721,In_2637);
and U3347 (N_3347,In_553,In_2681);
or U3348 (N_3348,In_1722,In_2681);
and U3349 (N_3349,In_31,In_1846);
xor U3350 (N_3350,In_858,In_1769);
nor U3351 (N_3351,In_2250,In_215);
nand U3352 (N_3352,In_390,In_2137);
xor U3353 (N_3353,In_2574,In_2826);
or U3354 (N_3354,In_2026,In_2622);
or U3355 (N_3355,In_829,In_2454);
and U3356 (N_3356,In_997,In_1993);
xnor U3357 (N_3357,In_2301,In_1929);
nor U3358 (N_3358,In_1698,In_2213);
or U3359 (N_3359,In_138,In_1863);
and U3360 (N_3360,In_2757,In_2268);
and U3361 (N_3361,In_1013,In_615);
or U3362 (N_3362,In_769,In_2847);
xnor U3363 (N_3363,In_526,In_552);
nor U3364 (N_3364,In_319,In_2417);
nor U3365 (N_3365,In_2684,In_282);
nor U3366 (N_3366,In_1208,In_2820);
nand U3367 (N_3367,In_2955,In_2988);
xor U3368 (N_3368,In_2891,In_135);
or U3369 (N_3369,In_384,In_1179);
nor U3370 (N_3370,In_2888,In_2373);
and U3371 (N_3371,In_2807,In_813);
or U3372 (N_3372,In_1419,In_2244);
and U3373 (N_3373,In_796,In_1935);
or U3374 (N_3374,In_46,In_1191);
nor U3375 (N_3375,In_2623,In_678);
xnor U3376 (N_3376,In_1541,In_2731);
or U3377 (N_3377,In_1594,In_1859);
and U3378 (N_3378,In_1222,In_2915);
and U3379 (N_3379,In_533,In_2945);
nand U3380 (N_3380,In_2245,In_1806);
or U3381 (N_3381,In_1460,In_1047);
xnor U3382 (N_3382,In_1910,In_321);
xor U3383 (N_3383,In_1619,In_2022);
nor U3384 (N_3384,In_2440,In_606);
or U3385 (N_3385,In_204,In_2854);
and U3386 (N_3386,In_714,In_2045);
nand U3387 (N_3387,In_2562,In_1999);
nor U3388 (N_3388,In_2554,In_1604);
xnor U3389 (N_3389,In_359,In_2298);
nand U3390 (N_3390,In_2140,In_2160);
or U3391 (N_3391,In_335,In_2873);
xnor U3392 (N_3392,In_164,In_546);
nor U3393 (N_3393,In_2082,In_1358);
and U3394 (N_3394,In_1493,In_1813);
or U3395 (N_3395,In_971,In_1096);
or U3396 (N_3396,In_635,In_1278);
nand U3397 (N_3397,In_1159,In_1540);
xnor U3398 (N_3398,In_2188,In_2129);
and U3399 (N_3399,In_2762,In_1176);
and U3400 (N_3400,In_1801,In_837);
or U3401 (N_3401,In_2850,In_2975);
xor U3402 (N_3402,In_7,In_2354);
nor U3403 (N_3403,In_873,In_1411);
nor U3404 (N_3404,In_878,In_998);
xor U3405 (N_3405,In_2772,In_540);
xnor U3406 (N_3406,In_1185,In_2538);
nand U3407 (N_3407,In_855,In_1657);
nor U3408 (N_3408,In_870,In_438);
nor U3409 (N_3409,In_2391,In_728);
nor U3410 (N_3410,In_1494,In_2771);
nand U3411 (N_3411,In_150,In_2072);
nand U3412 (N_3412,In_1544,In_2106);
nand U3413 (N_3413,In_962,In_1798);
nand U3414 (N_3414,In_2868,In_866);
nand U3415 (N_3415,In_1993,In_1504);
xor U3416 (N_3416,In_938,In_1624);
nand U3417 (N_3417,In_1460,In_2154);
nor U3418 (N_3418,In_1456,In_2008);
or U3419 (N_3419,In_333,In_200);
and U3420 (N_3420,In_1065,In_1687);
nor U3421 (N_3421,In_2298,In_1203);
nand U3422 (N_3422,In_1191,In_882);
xnor U3423 (N_3423,In_1661,In_1872);
nand U3424 (N_3424,In_2653,In_427);
xor U3425 (N_3425,In_2510,In_2218);
xor U3426 (N_3426,In_1688,In_2748);
nand U3427 (N_3427,In_736,In_831);
xnor U3428 (N_3428,In_2095,In_1426);
nor U3429 (N_3429,In_632,In_2511);
or U3430 (N_3430,In_2140,In_2114);
xnor U3431 (N_3431,In_1636,In_2116);
nand U3432 (N_3432,In_2861,In_2332);
and U3433 (N_3433,In_1506,In_2586);
and U3434 (N_3434,In_1626,In_821);
nand U3435 (N_3435,In_2667,In_984);
or U3436 (N_3436,In_679,In_2935);
and U3437 (N_3437,In_198,In_417);
nor U3438 (N_3438,In_1312,In_2291);
or U3439 (N_3439,In_1073,In_2503);
xnor U3440 (N_3440,In_2461,In_401);
and U3441 (N_3441,In_1002,In_2124);
nand U3442 (N_3442,In_906,In_2982);
nand U3443 (N_3443,In_1074,In_2880);
and U3444 (N_3444,In_280,In_2767);
and U3445 (N_3445,In_2829,In_775);
nand U3446 (N_3446,In_173,In_1658);
nor U3447 (N_3447,In_1583,In_505);
and U3448 (N_3448,In_594,In_915);
xor U3449 (N_3449,In_1108,In_677);
nand U3450 (N_3450,In_2484,In_2321);
and U3451 (N_3451,In_2011,In_2653);
nand U3452 (N_3452,In_1320,In_817);
nor U3453 (N_3453,In_357,In_2941);
and U3454 (N_3454,In_1043,In_1706);
xor U3455 (N_3455,In_2573,In_501);
or U3456 (N_3456,In_2140,In_2464);
xnor U3457 (N_3457,In_2408,In_2228);
xor U3458 (N_3458,In_481,In_887);
nor U3459 (N_3459,In_2409,In_2257);
xnor U3460 (N_3460,In_2396,In_2390);
or U3461 (N_3461,In_2180,In_358);
or U3462 (N_3462,In_1103,In_560);
xnor U3463 (N_3463,In_2910,In_1077);
nand U3464 (N_3464,In_2636,In_2480);
nand U3465 (N_3465,In_191,In_1704);
xnor U3466 (N_3466,In_2572,In_2748);
or U3467 (N_3467,In_258,In_2815);
or U3468 (N_3468,In_2589,In_1578);
xnor U3469 (N_3469,In_10,In_2197);
or U3470 (N_3470,In_754,In_1179);
and U3471 (N_3471,In_295,In_2953);
nand U3472 (N_3472,In_1462,In_2055);
or U3473 (N_3473,In_1130,In_1283);
nand U3474 (N_3474,In_2729,In_904);
nand U3475 (N_3475,In_2402,In_1477);
or U3476 (N_3476,In_1165,In_2971);
and U3477 (N_3477,In_2216,In_793);
xnor U3478 (N_3478,In_789,In_1285);
and U3479 (N_3479,In_841,In_2726);
or U3480 (N_3480,In_446,In_898);
and U3481 (N_3481,In_567,In_2102);
or U3482 (N_3482,In_876,In_2675);
nor U3483 (N_3483,In_2282,In_14);
xor U3484 (N_3484,In_2338,In_2583);
or U3485 (N_3485,In_1920,In_2178);
or U3486 (N_3486,In_490,In_692);
nand U3487 (N_3487,In_2203,In_930);
xnor U3488 (N_3488,In_616,In_828);
nand U3489 (N_3489,In_2246,In_857);
xnor U3490 (N_3490,In_992,In_2186);
and U3491 (N_3491,In_1540,In_2830);
and U3492 (N_3492,In_2760,In_2568);
nor U3493 (N_3493,In_185,In_1189);
nand U3494 (N_3494,In_728,In_2414);
xnor U3495 (N_3495,In_1424,In_2857);
xor U3496 (N_3496,In_519,In_1251);
or U3497 (N_3497,In_264,In_292);
xnor U3498 (N_3498,In_1467,In_660);
or U3499 (N_3499,In_1136,In_1521);
nand U3500 (N_3500,In_384,In_1786);
xnor U3501 (N_3501,In_1338,In_2574);
or U3502 (N_3502,In_1215,In_266);
xnor U3503 (N_3503,In_2660,In_1413);
or U3504 (N_3504,In_2138,In_411);
xor U3505 (N_3505,In_629,In_1919);
or U3506 (N_3506,In_845,In_2500);
or U3507 (N_3507,In_2464,In_30);
or U3508 (N_3508,In_2540,In_1821);
or U3509 (N_3509,In_273,In_1202);
or U3510 (N_3510,In_730,In_952);
xnor U3511 (N_3511,In_1415,In_1792);
nand U3512 (N_3512,In_1943,In_1260);
and U3513 (N_3513,In_1062,In_2767);
nor U3514 (N_3514,In_296,In_188);
nand U3515 (N_3515,In_775,In_800);
or U3516 (N_3516,In_1863,In_2437);
nand U3517 (N_3517,In_374,In_1309);
xor U3518 (N_3518,In_1700,In_1259);
nand U3519 (N_3519,In_2076,In_972);
and U3520 (N_3520,In_2789,In_2277);
xor U3521 (N_3521,In_2929,In_1955);
nand U3522 (N_3522,In_2765,In_1229);
xor U3523 (N_3523,In_1971,In_2719);
nor U3524 (N_3524,In_555,In_1056);
nor U3525 (N_3525,In_1722,In_592);
nor U3526 (N_3526,In_849,In_1871);
nand U3527 (N_3527,In_1932,In_2610);
or U3528 (N_3528,In_249,In_668);
or U3529 (N_3529,In_1503,In_444);
nor U3530 (N_3530,In_369,In_1550);
and U3531 (N_3531,In_13,In_2849);
and U3532 (N_3532,In_326,In_2886);
or U3533 (N_3533,In_284,In_1558);
and U3534 (N_3534,In_322,In_424);
nor U3535 (N_3535,In_693,In_442);
or U3536 (N_3536,In_630,In_1499);
nor U3537 (N_3537,In_1014,In_2473);
nor U3538 (N_3538,In_2920,In_2971);
and U3539 (N_3539,In_2567,In_1264);
or U3540 (N_3540,In_929,In_1582);
nor U3541 (N_3541,In_2305,In_1469);
xor U3542 (N_3542,In_2749,In_728);
nor U3543 (N_3543,In_296,In_128);
and U3544 (N_3544,In_1756,In_2187);
xnor U3545 (N_3545,In_2076,In_1145);
or U3546 (N_3546,In_2199,In_1682);
nand U3547 (N_3547,In_105,In_1641);
or U3548 (N_3548,In_1286,In_265);
or U3549 (N_3549,In_1272,In_51);
nor U3550 (N_3550,In_982,In_2935);
nand U3551 (N_3551,In_2584,In_749);
or U3552 (N_3552,In_782,In_717);
nor U3553 (N_3553,In_2761,In_2408);
xnor U3554 (N_3554,In_2717,In_532);
nand U3555 (N_3555,In_763,In_2819);
and U3556 (N_3556,In_2244,In_2980);
nor U3557 (N_3557,In_1218,In_1312);
xnor U3558 (N_3558,In_449,In_50);
or U3559 (N_3559,In_2217,In_1081);
nor U3560 (N_3560,In_2472,In_2805);
nor U3561 (N_3561,In_910,In_2575);
xor U3562 (N_3562,In_2619,In_1878);
nor U3563 (N_3563,In_1470,In_2426);
and U3564 (N_3564,In_984,In_1254);
or U3565 (N_3565,In_2888,In_2389);
xor U3566 (N_3566,In_2343,In_1066);
nor U3567 (N_3567,In_12,In_1067);
xnor U3568 (N_3568,In_1221,In_2658);
or U3569 (N_3569,In_2355,In_25);
nor U3570 (N_3570,In_508,In_1181);
and U3571 (N_3571,In_1200,In_2995);
or U3572 (N_3572,In_400,In_461);
nand U3573 (N_3573,In_2121,In_1582);
xor U3574 (N_3574,In_1840,In_2412);
nand U3575 (N_3575,In_2770,In_252);
or U3576 (N_3576,In_1515,In_535);
xor U3577 (N_3577,In_1249,In_2147);
nor U3578 (N_3578,In_282,In_2872);
nand U3579 (N_3579,In_328,In_1384);
or U3580 (N_3580,In_1204,In_1306);
nand U3581 (N_3581,In_1559,In_23);
nand U3582 (N_3582,In_73,In_2162);
nor U3583 (N_3583,In_257,In_1178);
or U3584 (N_3584,In_2876,In_1493);
or U3585 (N_3585,In_493,In_992);
nor U3586 (N_3586,In_1313,In_1348);
nand U3587 (N_3587,In_400,In_2718);
nor U3588 (N_3588,In_2675,In_1388);
nand U3589 (N_3589,In_288,In_2472);
nor U3590 (N_3590,In_1136,In_877);
nor U3591 (N_3591,In_645,In_1895);
xnor U3592 (N_3592,In_1408,In_2246);
or U3593 (N_3593,In_2612,In_1729);
xor U3594 (N_3594,In_370,In_250);
or U3595 (N_3595,In_2391,In_2454);
xnor U3596 (N_3596,In_2530,In_129);
xor U3597 (N_3597,In_1752,In_330);
nor U3598 (N_3598,In_198,In_983);
and U3599 (N_3599,In_1340,In_957);
or U3600 (N_3600,In_837,In_762);
or U3601 (N_3601,In_2112,In_1095);
nor U3602 (N_3602,In_1686,In_665);
nor U3603 (N_3603,In_707,In_749);
and U3604 (N_3604,In_698,In_2711);
nand U3605 (N_3605,In_2105,In_1352);
nand U3606 (N_3606,In_2204,In_1878);
nand U3607 (N_3607,In_1809,In_1566);
and U3608 (N_3608,In_2817,In_1778);
or U3609 (N_3609,In_1489,In_2290);
nor U3610 (N_3610,In_2469,In_2006);
or U3611 (N_3611,In_431,In_209);
and U3612 (N_3612,In_2358,In_118);
xor U3613 (N_3613,In_227,In_2953);
or U3614 (N_3614,In_1943,In_272);
or U3615 (N_3615,In_1288,In_1620);
nand U3616 (N_3616,In_2258,In_2069);
and U3617 (N_3617,In_919,In_1875);
xor U3618 (N_3618,In_2604,In_2922);
nor U3619 (N_3619,In_271,In_1427);
or U3620 (N_3620,In_68,In_1540);
nor U3621 (N_3621,In_303,In_2805);
nand U3622 (N_3622,In_2121,In_2949);
xor U3623 (N_3623,In_2402,In_2748);
nor U3624 (N_3624,In_2688,In_2340);
nand U3625 (N_3625,In_1765,In_1034);
nand U3626 (N_3626,In_2912,In_2875);
nand U3627 (N_3627,In_1760,In_462);
and U3628 (N_3628,In_2282,In_973);
nor U3629 (N_3629,In_1628,In_231);
and U3630 (N_3630,In_1285,In_192);
or U3631 (N_3631,In_1020,In_2018);
or U3632 (N_3632,In_2053,In_1949);
xor U3633 (N_3633,In_828,In_562);
xor U3634 (N_3634,In_2494,In_2459);
nand U3635 (N_3635,In_2791,In_1870);
xnor U3636 (N_3636,In_2813,In_497);
xnor U3637 (N_3637,In_2189,In_101);
nand U3638 (N_3638,In_2309,In_1532);
xnor U3639 (N_3639,In_1085,In_454);
and U3640 (N_3640,In_2756,In_629);
xor U3641 (N_3641,In_630,In_1839);
xnor U3642 (N_3642,In_304,In_2722);
nand U3643 (N_3643,In_2771,In_443);
nor U3644 (N_3644,In_2034,In_2412);
xor U3645 (N_3645,In_1819,In_1652);
and U3646 (N_3646,In_72,In_1900);
nand U3647 (N_3647,In_2369,In_984);
nor U3648 (N_3648,In_1479,In_541);
nand U3649 (N_3649,In_1719,In_219);
xnor U3650 (N_3650,In_2075,In_2650);
xor U3651 (N_3651,In_1433,In_662);
and U3652 (N_3652,In_1088,In_2660);
and U3653 (N_3653,In_1065,In_1244);
nor U3654 (N_3654,In_1982,In_2317);
and U3655 (N_3655,In_2582,In_1513);
or U3656 (N_3656,In_1864,In_2593);
or U3657 (N_3657,In_2565,In_2285);
and U3658 (N_3658,In_1792,In_57);
nand U3659 (N_3659,In_1507,In_2130);
xor U3660 (N_3660,In_1383,In_2848);
xnor U3661 (N_3661,In_1390,In_2206);
or U3662 (N_3662,In_2013,In_1284);
or U3663 (N_3663,In_2490,In_1907);
nor U3664 (N_3664,In_1388,In_2306);
nor U3665 (N_3665,In_2195,In_1253);
nand U3666 (N_3666,In_1807,In_674);
nor U3667 (N_3667,In_1652,In_851);
and U3668 (N_3668,In_2033,In_1096);
nand U3669 (N_3669,In_1609,In_2085);
or U3670 (N_3670,In_324,In_2213);
and U3671 (N_3671,In_884,In_2680);
or U3672 (N_3672,In_2220,In_720);
xnor U3673 (N_3673,In_2239,In_1111);
nor U3674 (N_3674,In_1769,In_2679);
and U3675 (N_3675,In_2490,In_420);
and U3676 (N_3676,In_2076,In_638);
nor U3677 (N_3677,In_2986,In_178);
xnor U3678 (N_3678,In_2082,In_637);
or U3679 (N_3679,In_564,In_510);
or U3680 (N_3680,In_1000,In_1633);
or U3681 (N_3681,In_277,In_1944);
nand U3682 (N_3682,In_1472,In_794);
or U3683 (N_3683,In_1795,In_1286);
nor U3684 (N_3684,In_454,In_817);
nor U3685 (N_3685,In_2663,In_145);
or U3686 (N_3686,In_1761,In_1298);
or U3687 (N_3687,In_1395,In_2675);
or U3688 (N_3688,In_2352,In_754);
nor U3689 (N_3689,In_1804,In_2232);
xnor U3690 (N_3690,In_2943,In_1786);
nand U3691 (N_3691,In_109,In_2199);
nor U3692 (N_3692,In_1831,In_297);
and U3693 (N_3693,In_18,In_921);
or U3694 (N_3694,In_2563,In_520);
and U3695 (N_3695,In_2652,In_2322);
xor U3696 (N_3696,In_2123,In_1394);
nand U3697 (N_3697,In_2967,In_2163);
xnor U3698 (N_3698,In_86,In_2461);
nand U3699 (N_3699,In_2693,In_507);
nand U3700 (N_3700,In_1642,In_461);
nor U3701 (N_3701,In_1251,In_1379);
nand U3702 (N_3702,In_375,In_1614);
nand U3703 (N_3703,In_289,In_26);
nand U3704 (N_3704,In_21,In_2607);
nand U3705 (N_3705,In_1316,In_1611);
nor U3706 (N_3706,In_2305,In_63);
or U3707 (N_3707,In_2343,In_1506);
or U3708 (N_3708,In_2302,In_2403);
or U3709 (N_3709,In_2531,In_2144);
and U3710 (N_3710,In_738,In_72);
nor U3711 (N_3711,In_784,In_1559);
and U3712 (N_3712,In_2896,In_1397);
nor U3713 (N_3713,In_2812,In_486);
nand U3714 (N_3714,In_2291,In_1685);
and U3715 (N_3715,In_1935,In_1762);
or U3716 (N_3716,In_1299,In_1767);
or U3717 (N_3717,In_2603,In_1578);
xnor U3718 (N_3718,In_75,In_1664);
nand U3719 (N_3719,In_1126,In_440);
nand U3720 (N_3720,In_1519,In_855);
nand U3721 (N_3721,In_2368,In_1238);
xor U3722 (N_3722,In_766,In_925);
and U3723 (N_3723,In_2524,In_2276);
nor U3724 (N_3724,In_1183,In_970);
xnor U3725 (N_3725,In_1169,In_2699);
or U3726 (N_3726,In_2413,In_2741);
and U3727 (N_3727,In_2482,In_1385);
xor U3728 (N_3728,In_766,In_291);
and U3729 (N_3729,In_1872,In_1835);
or U3730 (N_3730,In_2514,In_1867);
xnor U3731 (N_3731,In_2040,In_1834);
or U3732 (N_3732,In_2576,In_1842);
or U3733 (N_3733,In_2419,In_1781);
xnor U3734 (N_3734,In_477,In_245);
nor U3735 (N_3735,In_2047,In_1965);
xnor U3736 (N_3736,In_156,In_1683);
xor U3737 (N_3737,In_1355,In_2591);
and U3738 (N_3738,In_1492,In_917);
or U3739 (N_3739,In_2844,In_1607);
xor U3740 (N_3740,In_2979,In_580);
or U3741 (N_3741,In_2066,In_1683);
xnor U3742 (N_3742,In_1142,In_88);
nand U3743 (N_3743,In_482,In_1238);
and U3744 (N_3744,In_278,In_1918);
and U3745 (N_3745,In_2043,In_1186);
and U3746 (N_3746,In_1797,In_400);
and U3747 (N_3747,In_1608,In_1451);
xor U3748 (N_3748,In_1466,In_877);
and U3749 (N_3749,In_2770,In_2460);
nor U3750 (N_3750,In_1358,In_2001);
or U3751 (N_3751,In_765,In_934);
xor U3752 (N_3752,In_1094,In_2333);
nor U3753 (N_3753,In_2117,In_1498);
nor U3754 (N_3754,In_745,In_911);
nand U3755 (N_3755,In_2447,In_857);
or U3756 (N_3756,In_2530,In_1425);
and U3757 (N_3757,In_1307,In_1500);
nand U3758 (N_3758,In_2329,In_395);
nor U3759 (N_3759,In_563,In_697);
nand U3760 (N_3760,In_663,In_307);
nand U3761 (N_3761,In_2011,In_1362);
and U3762 (N_3762,In_2558,In_422);
xor U3763 (N_3763,In_2018,In_2494);
nor U3764 (N_3764,In_1792,In_1051);
xnor U3765 (N_3765,In_472,In_11);
nor U3766 (N_3766,In_2952,In_1636);
and U3767 (N_3767,In_1086,In_2385);
and U3768 (N_3768,In_1426,In_1471);
or U3769 (N_3769,In_1561,In_978);
and U3770 (N_3770,In_1711,In_710);
xnor U3771 (N_3771,In_2762,In_939);
nand U3772 (N_3772,In_2065,In_304);
nand U3773 (N_3773,In_620,In_1727);
and U3774 (N_3774,In_596,In_2756);
xor U3775 (N_3775,In_1566,In_1018);
and U3776 (N_3776,In_2582,In_2971);
or U3777 (N_3777,In_2985,In_1225);
and U3778 (N_3778,In_2946,In_2446);
nor U3779 (N_3779,In_2054,In_2923);
or U3780 (N_3780,In_1063,In_149);
xnor U3781 (N_3781,In_437,In_1889);
or U3782 (N_3782,In_2547,In_2197);
xor U3783 (N_3783,In_2321,In_425);
xnor U3784 (N_3784,In_1458,In_2224);
nand U3785 (N_3785,In_9,In_2179);
nand U3786 (N_3786,In_2495,In_352);
nor U3787 (N_3787,In_2928,In_462);
xor U3788 (N_3788,In_2061,In_930);
or U3789 (N_3789,In_618,In_1608);
xnor U3790 (N_3790,In_369,In_2524);
or U3791 (N_3791,In_1557,In_41);
nor U3792 (N_3792,In_1958,In_2483);
xnor U3793 (N_3793,In_41,In_449);
and U3794 (N_3794,In_553,In_1832);
and U3795 (N_3795,In_363,In_1102);
nand U3796 (N_3796,In_2609,In_2220);
nor U3797 (N_3797,In_187,In_431);
nand U3798 (N_3798,In_1655,In_2367);
nor U3799 (N_3799,In_565,In_1126);
nor U3800 (N_3800,In_1561,In_1510);
or U3801 (N_3801,In_1729,In_468);
and U3802 (N_3802,In_1269,In_2781);
or U3803 (N_3803,In_1106,In_1741);
nor U3804 (N_3804,In_2815,In_1721);
nand U3805 (N_3805,In_1735,In_457);
nand U3806 (N_3806,In_186,In_1601);
or U3807 (N_3807,In_2239,In_2245);
and U3808 (N_3808,In_783,In_1743);
nand U3809 (N_3809,In_1225,In_1828);
and U3810 (N_3810,In_2959,In_2345);
nor U3811 (N_3811,In_1557,In_422);
xnor U3812 (N_3812,In_1403,In_696);
or U3813 (N_3813,In_2577,In_409);
and U3814 (N_3814,In_23,In_878);
xnor U3815 (N_3815,In_2945,In_2217);
nand U3816 (N_3816,In_2925,In_1722);
nor U3817 (N_3817,In_1735,In_130);
nor U3818 (N_3818,In_2871,In_738);
and U3819 (N_3819,In_332,In_1965);
nand U3820 (N_3820,In_1429,In_2377);
and U3821 (N_3821,In_2116,In_2918);
or U3822 (N_3822,In_2429,In_2034);
nor U3823 (N_3823,In_1988,In_2686);
nand U3824 (N_3824,In_1261,In_2748);
and U3825 (N_3825,In_858,In_1971);
nor U3826 (N_3826,In_311,In_57);
or U3827 (N_3827,In_1125,In_399);
xor U3828 (N_3828,In_2400,In_87);
xor U3829 (N_3829,In_602,In_1612);
nand U3830 (N_3830,In_2886,In_585);
or U3831 (N_3831,In_1583,In_2573);
and U3832 (N_3832,In_1236,In_714);
and U3833 (N_3833,In_1550,In_1572);
xor U3834 (N_3834,In_1922,In_510);
or U3835 (N_3835,In_386,In_2792);
and U3836 (N_3836,In_1041,In_2800);
or U3837 (N_3837,In_255,In_2270);
nor U3838 (N_3838,In_2555,In_1072);
or U3839 (N_3839,In_1216,In_2300);
and U3840 (N_3840,In_1606,In_2023);
and U3841 (N_3841,In_2001,In_2230);
xnor U3842 (N_3842,In_819,In_2807);
xnor U3843 (N_3843,In_1050,In_2898);
or U3844 (N_3844,In_314,In_512);
xnor U3845 (N_3845,In_2803,In_1743);
and U3846 (N_3846,In_252,In_2426);
nand U3847 (N_3847,In_1833,In_877);
nor U3848 (N_3848,In_888,In_2611);
and U3849 (N_3849,In_579,In_319);
xor U3850 (N_3850,In_1018,In_2144);
nand U3851 (N_3851,In_351,In_1653);
xor U3852 (N_3852,In_889,In_1234);
nand U3853 (N_3853,In_1515,In_1868);
and U3854 (N_3854,In_2993,In_319);
xnor U3855 (N_3855,In_542,In_1705);
xnor U3856 (N_3856,In_1109,In_2937);
or U3857 (N_3857,In_2312,In_818);
and U3858 (N_3858,In_1026,In_2579);
or U3859 (N_3859,In_338,In_943);
xor U3860 (N_3860,In_2941,In_1014);
and U3861 (N_3861,In_2566,In_1823);
nand U3862 (N_3862,In_2854,In_1841);
xnor U3863 (N_3863,In_972,In_1784);
or U3864 (N_3864,In_1960,In_1580);
and U3865 (N_3865,In_2069,In_1387);
nand U3866 (N_3866,In_2288,In_2010);
nor U3867 (N_3867,In_1534,In_2677);
xnor U3868 (N_3868,In_611,In_2470);
xor U3869 (N_3869,In_2110,In_1250);
and U3870 (N_3870,In_2353,In_2766);
nor U3871 (N_3871,In_1205,In_2465);
or U3872 (N_3872,In_2304,In_1345);
nor U3873 (N_3873,In_1403,In_2689);
and U3874 (N_3874,In_1464,In_2731);
and U3875 (N_3875,In_633,In_1694);
xor U3876 (N_3876,In_968,In_1406);
nor U3877 (N_3877,In_1218,In_1000);
and U3878 (N_3878,In_955,In_670);
and U3879 (N_3879,In_2826,In_2910);
nor U3880 (N_3880,In_1594,In_435);
nor U3881 (N_3881,In_1079,In_2704);
and U3882 (N_3882,In_2926,In_266);
or U3883 (N_3883,In_1792,In_998);
xnor U3884 (N_3884,In_1375,In_2360);
nor U3885 (N_3885,In_1859,In_64);
xnor U3886 (N_3886,In_2184,In_2453);
nor U3887 (N_3887,In_1069,In_2133);
xor U3888 (N_3888,In_2946,In_1150);
and U3889 (N_3889,In_1782,In_2611);
xnor U3890 (N_3890,In_2497,In_2332);
or U3891 (N_3891,In_945,In_470);
and U3892 (N_3892,In_1202,In_348);
and U3893 (N_3893,In_2742,In_549);
and U3894 (N_3894,In_1920,In_1263);
or U3895 (N_3895,In_216,In_2143);
or U3896 (N_3896,In_2454,In_2002);
or U3897 (N_3897,In_25,In_1509);
or U3898 (N_3898,In_15,In_908);
or U3899 (N_3899,In_1691,In_1527);
nor U3900 (N_3900,In_2606,In_1481);
nand U3901 (N_3901,In_198,In_2119);
and U3902 (N_3902,In_2113,In_457);
nor U3903 (N_3903,In_2949,In_1455);
xor U3904 (N_3904,In_712,In_1104);
nand U3905 (N_3905,In_1454,In_1256);
and U3906 (N_3906,In_1263,In_865);
nor U3907 (N_3907,In_1781,In_1032);
xnor U3908 (N_3908,In_2413,In_2281);
nand U3909 (N_3909,In_2752,In_1008);
and U3910 (N_3910,In_1739,In_1072);
nor U3911 (N_3911,In_1737,In_41);
nor U3912 (N_3912,In_233,In_576);
xor U3913 (N_3913,In_1495,In_1759);
nand U3914 (N_3914,In_2180,In_225);
or U3915 (N_3915,In_2500,In_1040);
or U3916 (N_3916,In_548,In_977);
nor U3917 (N_3917,In_454,In_2631);
or U3918 (N_3918,In_476,In_2609);
and U3919 (N_3919,In_825,In_428);
nor U3920 (N_3920,In_2179,In_1542);
nor U3921 (N_3921,In_2815,In_2115);
or U3922 (N_3922,In_574,In_2169);
nand U3923 (N_3923,In_446,In_284);
and U3924 (N_3924,In_1936,In_435);
nand U3925 (N_3925,In_2203,In_1353);
and U3926 (N_3926,In_2198,In_2791);
and U3927 (N_3927,In_924,In_2319);
xnor U3928 (N_3928,In_2165,In_729);
and U3929 (N_3929,In_1310,In_1270);
nor U3930 (N_3930,In_1793,In_1729);
xor U3931 (N_3931,In_1447,In_2681);
nand U3932 (N_3932,In_583,In_505);
nand U3933 (N_3933,In_1493,In_1562);
xnor U3934 (N_3934,In_1726,In_1493);
nand U3935 (N_3935,In_1677,In_2617);
and U3936 (N_3936,In_2413,In_1826);
or U3937 (N_3937,In_1105,In_135);
xor U3938 (N_3938,In_572,In_884);
nor U3939 (N_3939,In_1649,In_118);
nand U3940 (N_3940,In_1080,In_2957);
nor U3941 (N_3941,In_2078,In_637);
and U3942 (N_3942,In_1598,In_1273);
xnor U3943 (N_3943,In_2809,In_2015);
nand U3944 (N_3944,In_1622,In_2317);
and U3945 (N_3945,In_2542,In_2772);
nor U3946 (N_3946,In_1263,In_2876);
and U3947 (N_3947,In_1814,In_2464);
nand U3948 (N_3948,In_2383,In_906);
and U3949 (N_3949,In_1433,In_1473);
nand U3950 (N_3950,In_1529,In_1272);
or U3951 (N_3951,In_109,In_2062);
xor U3952 (N_3952,In_2321,In_1270);
nor U3953 (N_3953,In_557,In_1013);
nand U3954 (N_3954,In_682,In_1373);
xnor U3955 (N_3955,In_1723,In_2527);
xnor U3956 (N_3956,In_2626,In_2181);
and U3957 (N_3957,In_931,In_711);
and U3958 (N_3958,In_1141,In_1965);
nand U3959 (N_3959,In_2432,In_1355);
or U3960 (N_3960,In_2571,In_962);
nor U3961 (N_3961,In_385,In_2935);
or U3962 (N_3962,In_1669,In_1987);
nand U3963 (N_3963,In_2528,In_199);
nor U3964 (N_3964,In_1002,In_1512);
nand U3965 (N_3965,In_837,In_2099);
xnor U3966 (N_3966,In_544,In_2725);
and U3967 (N_3967,In_1239,In_575);
xor U3968 (N_3968,In_1252,In_2403);
and U3969 (N_3969,In_249,In_2795);
nand U3970 (N_3970,In_2038,In_1427);
and U3971 (N_3971,In_2230,In_741);
or U3972 (N_3972,In_1876,In_764);
and U3973 (N_3973,In_1727,In_302);
or U3974 (N_3974,In_256,In_269);
or U3975 (N_3975,In_133,In_1792);
nor U3976 (N_3976,In_142,In_1987);
nor U3977 (N_3977,In_2183,In_938);
nand U3978 (N_3978,In_174,In_503);
nor U3979 (N_3979,In_2468,In_2232);
or U3980 (N_3980,In_2848,In_2234);
xnor U3981 (N_3981,In_2015,In_2164);
and U3982 (N_3982,In_126,In_1346);
xnor U3983 (N_3983,In_2675,In_1811);
or U3984 (N_3984,In_2757,In_2043);
nand U3985 (N_3985,In_2131,In_1012);
xnor U3986 (N_3986,In_1848,In_79);
and U3987 (N_3987,In_1893,In_1151);
nand U3988 (N_3988,In_1551,In_1457);
nor U3989 (N_3989,In_2971,In_1552);
or U3990 (N_3990,In_958,In_451);
and U3991 (N_3991,In_2310,In_559);
and U3992 (N_3992,In_1639,In_1688);
nor U3993 (N_3993,In_156,In_1026);
and U3994 (N_3994,In_731,In_2959);
nor U3995 (N_3995,In_745,In_2487);
nor U3996 (N_3996,In_2637,In_2287);
and U3997 (N_3997,In_947,In_1120);
nor U3998 (N_3998,In_1296,In_2090);
nand U3999 (N_3999,In_298,In_1648);
or U4000 (N_4000,In_2906,In_864);
nand U4001 (N_4001,In_774,In_1086);
nor U4002 (N_4002,In_1946,In_968);
and U4003 (N_4003,In_2828,In_122);
nand U4004 (N_4004,In_1971,In_738);
xnor U4005 (N_4005,In_2335,In_2569);
nor U4006 (N_4006,In_61,In_2781);
nor U4007 (N_4007,In_2333,In_2547);
and U4008 (N_4008,In_1427,In_2689);
nand U4009 (N_4009,In_1388,In_1490);
or U4010 (N_4010,In_2471,In_539);
xnor U4011 (N_4011,In_2406,In_2007);
xnor U4012 (N_4012,In_2150,In_756);
and U4013 (N_4013,In_2879,In_2328);
and U4014 (N_4014,In_1789,In_1669);
nor U4015 (N_4015,In_2908,In_206);
nor U4016 (N_4016,In_506,In_2713);
or U4017 (N_4017,In_768,In_1010);
or U4018 (N_4018,In_2189,In_937);
xnor U4019 (N_4019,In_323,In_254);
and U4020 (N_4020,In_2328,In_594);
xor U4021 (N_4021,In_1031,In_646);
and U4022 (N_4022,In_1364,In_2072);
nor U4023 (N_4023,In_2260,In_5);
and U4024 (N_4024,In_1054,In_1550);
or U4025 (N_4025,In_1166,In_334);
or U4026 (N_4026,In_2322,In_2261);
nand U4027 (N_4027,In_2235,In_1662);
nand U4028 (N_4028,In_373,In_1899);
nor U4029 (N_4029,In_320,In_2015);
nor U4030 (N_4030,In_1537,In_547);
nand U4031 (N_4031,In_2375,In_2121);
nor U4032 (N_4032,In_2852,In_2107);
and U4033 (N_4033,In_2324,In_1262);
nand U4034 (N_4034,In_639,In_368);
xnor U4035 (N_4035,In_403,In_1192);
nor U4036 (N_4036,In_588,In_636);
xnor U4037 (N_4037,In_1342,In_269);
or U4038 (N_4038,In_2747,In_2097);
nand U4039 (N_4039,In_29,In_1619);
or U4040 (N_4040,In_374,In_2301);
or U4041 (N_4041,In_1403,In_602);
nand U4042 (N_4042,In_1571,In_630);
nand U4043 (N_4043,In_1068,In_320);
and U4044 (N_4044,In_1126,In_2168);
xnor U4045 (N_4045,In_994,In_235);
nand U4046 (N_4046,In_1671,In_1847);
nand U4047 (N_4047,In_2349,In_454);
xor U4048 (N_4048,In_1422,In_784);
nor U4049 (N_4049,In_2554,In_1900);
or U4050 (N_4050,In_1697,In_1031);
xnor U4051 (N_4051,In_2459,In_1324);
nor U4052 (N_4052,In_221,In_1964);
nor U4053 (N_4053,In_2080,In_1697);
nand U4054 (N_4054,In_2789,In_1304);
and U4055 (N_4055,In_1086,In_920);
or U4056 (N_4056,In_795,In_2154);
and U4057 (N_4057,In_1227,In_1370);
or U4058 (N_4058,In_2440,In_1608);
nor U4059 (N_4059,In_2621,In_1945);
nor U4060 (N_4060,In_1391,In_2561);
and U4061 (N_4061,In_1203,In_1144);
nor U4062 (N_4062,In_2918,In_1811);
nor U4063 (N_4063,In_1887,In_721);
or U4064 (N_4064,In_696,In_1252);
or U4065 (N_4065,In_2277,In_2250);
nand U4066 (N_4066,In_1426,In_1878);
nand U4067 (N_4067,In_774,In_1070);
nor U4068 (N_4068,In_1650,In_885);
nand U4069 (N_4069,In_1610,In_2586);
xor U4070 (N_4070,In_2033,In_779);
xnor U4071 (N_4071,In_613,In_616);
nand U4072 (N_4072,In_1527,In_2398);
and U4073 (N_4073,In_1237,In_1426);
nor U4074 (N_4074,In_2980,In_2538);
and U4075 (N_4075,In_81,In_216);
and U4076 (N_4076,In_2452,In_2873);
nand U4077 (N_4077,In_1297,In_1040);
nand U4078 (N_4078,In_2764,In_31);
xor U4079 (N_4079,In_2571,In_2545);
and U4080 (N_4080,In_966,In_1072);
nand U4081 (N_4081,In_617,In_2445);
nor U4082 (N_4082,In_1699,In_1422);
nand U4083 (N_4083,In_2852,In_1430);
and U4084 (N_4084,In_2437,In_200);
or U4085 (N_4085,In_2205,In_77);
or U4086 (N_4086,In_929,In_84);
nand U4087 (N_4087,In_435,In_790);
xnor U4088 (N_4088,In_2885,In_2298);
nor U4089 (N_4089,In_150,In_772);
and U4090 (N_4090,In_2496,In_2982);
xnor U4091 (N_4091,In_2557,In_1013);
or U4092 (N_4092,In_1642,In_2051);
nor U4093 (N_4093,In_129,In_2156);
or U4094 (N_4094,In_1119,In_653);
or U4095 (N_4095,In_643,In_122);
xor U4096 (N_4096,In_1053,In_1373);
and U4097 (N_4097,In_2327,In_2736);
nand U4098 (N_4098,In_1094,In_2514);
and U4099 (N_4099,In_107,In_573);
or U4100 (N_4100,In_1297,In_1039);
nand U4101 (N_4101,In_2114,In_2384);
or U4102 (N_4102,In_108,In_2801);
nor U4103 (N_4103,In_2110,In_1717);
nand U4104 (N_4104,In_720,In_2633);
nand U4105 (N_4105,In_750,In_2142);
xnor U4106 (N_4106,In_1481,In_729);
nand U4107 (N_4107,In_2051,In_1188);
nand U4108 (N_4108,In_416,In_1399);
or U4109 (N_4109,In_834,In_1159);
xor U4110 (N_4110,In_2980,In_210);
or U4111 (N_4111,In_1833,In_2463);
xor U4112 (N_4112,In_11,In_1478);
xor U4113 (N_4113,In_847,In_1224);
xor U4114 (N_4114,In_820,In_1479);
xor U4115 (N_4115,In_2041,In_2927);
and U4116 (N_4116,In_453,In_2809);
and U4117 (N_4117,In_2400,In_910);
or U4118 (N_4118,In_2305,In_2843);
nand U4119 (N_4119,In_1632,In_229);
xnor U4120 (N_4120,In_1332,In_1151);
or U4121 (N_4121,In_2575,In_2890);
and U4122 (N_4122,In_1244,In_1715);
or U4123 (N_4123,In_1153,In_2462);
nand U4124 (N_4124,In_1176,In_1657);
and U4125 (N_4125,In_1797,In_2732);
nand U4126 (N_4126,In_2732,In_2761);
nand U4127 (N_4127,In_917,In_1678);
nor U4128 (N_4128,In_1677,In_1878);
nor U4129 (N_4129,In_1480,In_723);
nand U4130 (N_4130,In_2572,In_2658);
and U4131 (N_4131,In_1452,In_1802);
nor U4132 (N_4132,In_2923,In_1438);
or U4133 (N_4133,In_543,In_1398);
xnor U4134 (N_4134,In_1798,In_943);
xnor U4135 (N_4135,In_2807,In_2164);
and U4136 (N_4136,In_1409,In_2556);
or U4137 (N_4137,In_124,In_889);
or U4138 (N_4138,In_2579,In_956);
nand U4139 (N_4139,In_1082,In_1268);
nand U4140 (N_4140,In_1564,In_1790);
nor U4141 (N_4141,In_1963,In_881);
nor U4142 (N_4142,In_18,In_1908);
or U4143 (N_4143,In_2079,In_1966);
and U4144 (N_4144,In_2098,In_2185);
or U4145 (N_4145,In_2501,In_417);
nand U4146 (N_4146,In_776,In_1548);
or U4147 (N_4147,In_616,In_55);
xnor U4148 (N_4148,In_2403,In_1490);
nor U4149 (N_4149,In_427,In_2422);
or U4150 (N_4150,In_863,In_320);
nor U4151 (N_4151,In_1322,In_2352);
nand U4152 (N_4152,In_317,In_1799);
and U4153 (N_4153,In_1191,In_1485);
nor U4154 (N_4154,In_357,In_321);
or U4155 (N_4155,In_590,In_1083);
xor U4156 (N_4156,In_686,In_1824);
and U4157 (N_4157,In_1587,In_2469);
or U4158 (N_4158,In_2358,In_663);
xor U4159 (N_4159,In_660,In_2825);
nor U4160 (N_4160,In_1173,In_754);
and U4161 (N_4161,In_140,In_2641);
nor U4162 (N_4162,In_2963,In_808);
and U4163 (N_4163,In_2720,In_2838);
and U4164 (N_4164,In_1463,In_1755);
xnor U4165 (N_4165,In_2027,In_390);
xor U4166 (N_4166,In_108,In_266);
xnor U4167 (N_4167,In_1461,In_1547);
or U4168 (N_4168,In_2507,In_2053);
nor U4169 (N_4169,In_1209,In_31);
nand U4170 (N_4170,In_2657,In_1660);
nand U4171 (N_4171,In_14,In_2801);
and U4172 (N_4172,In_2401,In_181);
and U4173 (N_4173,In_213,In_2993);
and U4174 (N_4174,In_1194,In_1802);
or U4175 (N_4175,In_1855,In_2542);
nor U4176 (N_4176,In_1334,In_1035);
nand U4177 (N_4177,In_2320,In_195);
or U4178 (N_4178,In_2673,In_856);
nand U4179 (N_4179,In_985,In_1978);
nor U4180 (N_4180,In_863,In_696);
xnor U4181 (N_4181,In_2968,In_1961);
nand U4182 (N_4182,In_1071,In_59);
nand U4183 (N_4183,In_1486,In_1090);
or U4184 (N_4184,In_1939,In_754);
nand U4185 (N_4185,In_1816,In_2688);
xnor U4186 (N_4186,In_454,In_419);
nand U4187 (N_4187,In_990,In_1020);
and U4188 (N_4188,In_714,In_2518);
and U4189 (N_4189,In_599,In_279);
nand U4190 (N_4190,In_2629,In_777);
and U4191 (N_4191,In_2403,In_1242);
xor U4192 (N_4192,In_1197,In_1413);
nand U4193 (N_4193,In_1633,In_1399);
or U4194 (N_4194,In_872,In_2769);
nand U4195 (N_4195,In_2701,In_2032);
nand U4196 (N_4196,In_2087,In_1968);
or U4197 (N_4197,In_1552,In_1682);
xor U4198 (N_4198,In_1257,In_2067);
nand U4199 (N_4199,In_311,In_643);
nor U4200 (N_4200,In_1455,In_729);
or U4201 (N_4201,In_1280,In_462);
nand U4202 (N_4202,In_625,In_1810);
and U4203 (N_4203,In_792,In_2013);
nor U4204 (N_4204,In_2690,In_716);
nand U4205 (N_4205,In_491,In_2483);
and U4206 (N_4206,In_548,In_2220);
and U4207 (N_4207,In_1998,In_1333);
xnor U4208 (N_4208,In_229,In_1087);
and U4209 (N_4209,In_2886,In_1498);
nor U4210 (N_4210,In_318,In_2870);
xor U4211 (N_4211,In_894,In_2181);
or U4212 (N_4212,In_1043,In_1511);
nand U4213 (N_4213,In_892,In_1816);
or U4214 (N_4214,In_2991,In_1661);
and U4215 (N_4215,In_1063,In_336);
nor U4216 (N_4216,In_832,In_892);
xnor U4217 (N_4217,In_1726,In_1097);
nor U4218 (N_4218,In_2752,In_1572);
nor U4219 (N_4219,In_526,In_1053);
nor U4220 (N_4220,In_2160,In_1369);
and U4221 (N_4221,In_857,In_1022);
nor U4222 (N_4222,In_710,In_436);
xor U4223 (N_4223,In_1258,In_486);
nor U4224 (N_4224,In_882,In_45);
xnor U4225 (N_4225,In_780,In_2324);
nand U4226 (N_4226,In_1286,In_540);
nand U4227 (N_4227,In_1564,In_334);
xor U4228 (N_4228,In_126,In_1305);
nor U4229 (N_4229,In_1689,In_2265);
nand U4230 (N_4230,In_2383,In_2497);
nand U4231 (N_4231,In_1010,In_2479);
nor U4232 (N_4232,In_1790,In_487);
xnor U4233 (N_4233,In_2806,In_889);
and U4234 (N_4234,In_1920,In_345);
xor U4235 (N_4235,In_953,In_1280);
and U4236 (N_4236,In_1035,In_2402);
xor U4237 (N_4237,In_2682,In_188);
xnor U4238 (N_4238,In_2593,In_1485);
nand U4239 (N_4239,In_199,In_1414);
and U4240 (N_4240,In_2172,In_574);
xnor U4241 (N_4241,In_2723,In_2624);
nand U4242 (N_4242,In_871,In_1407);
xor U4243 (N_4243,In_1531,In_1752);
xnor U4244 (N_4244,In_1641,In_544);
or U4245 (N_4245,In_2407,In_1372);
nor U4246 (N_4246,In_2313,In_1314);
nand U4247 (N_4247,In_1002,In_2514);
nor U4248 (N_4248,In_397,In_2221);
nor U4249 (N_4249,In_2738,In_2937);
xor U4250 (N_4250,In_2354,In_495);
nand U4251 (N_4251,In_1614,In_2407);
nor U4252 (N_4252,In_634,In_1789);
or U4253 (N_4253,In_869,In_164);
or U4254 (N_4254,In_2362,In_1729);
and U4255 (N_4255,In_925,In_1100);
and U4256 (N_4256,In_996,In_2917);
nor U4257 (N_4257,In_1125,In_461);
xnor U4258 (N_4258,In_2457,In_2522);
and U4259 (N_4259,In_1530,In_545);
nand U4260 (N_4260,In_205,In_1094);
nor U4261 (N_4261,In_2203,In_934);
xnor U4262 (N_4262,In_2414,In_372);
nand U4263 (N_4263,In_1474,In_1350);
and U4264 (N_4264,In_1246,In_243);
and U4265 (N_4265,In_278,In_2891);
nand U4266 (N_4266,In_2493,In_1709);
and U4267 (N_4267,In_1856,In_557);
or U4268 (N_4268,In_2896,In_860);
or U4269 (N_4269,In_957,In_2583);
or U4270 (N_4270,In_2540,In_1673);
xor U4271 (N_4271,In_919,In_2427);
and U4272 (N_4272,In_1920,In_2297);
and U4273 (N_4273,In_283,In_1342);
and U4274 (N_4274,In_421,In_119);
xnor U4275 (N_4275,In_2009,In_558);
xnor U4276 (N_4276,In_1827,In_291);
nand U4277 (N_4277,In_1176,In_1397);
xor U4278 (N_4278,In_563,In_2454);
or U4279 (N_4279,In_1725,In_2540);
xor U4280 (N_4280,In_796,In_2805);
or U4281 (N_4281,In_2073,In_2612);
or U4282 (N_4282,In_2948,In_478);
or U4283 (N_4283,In_2092,In_2808);
and U4284 (N_4284,In_864,In_2943);
and U4285 (N_4285,In_2628,In_2408);
nand U4286 (N_4286,In_2492,In_2571);
or U4287 (N_4287,In_1580,In_1903);
nand U4288 (N_4288,In_1759,In_1747);
xor U4289 (N_4289,In_1607,In_2899);
nand U4290 (N_4290,In_3,In_1952);
nand U4291 (N_4291,In_456,In_2458);
xnor U4292 (N_4292,In_1997,In_1277);
xor U4293 (N_4293,In_291,In_1698);
or U4294 (N_4294,In_2353,In_580);
nor U4295 (N_4295,In_1916,In_623);
xnor U4296 (N_4296,In_829,In_606);
nand U4297 (N_4297,In_2495,In_1712);
and U4298 (N_4298,In_1190,In_1685);
nor U4299 (N_4299,In_560,In_1143);
nand U4300 (N_4300,In_285,In_26);
or U4301 (N_4301,In_529,In_2424);
and U4302 (N_4302,In_1035,In_1609);
nor U4303 (N_4303,In_1903,In_1366);
or U4304 (N_4304,In_383,In_1732);
xor U4305 (N_4305,In_567,In_729);
nand U4306 (N_4306,In_1669,In_1445);
nor U4307 (N_4307,In_2111,In_158);
or U4308 (N_4308,In_2798,In_2600);
or U4309 (N_4309,In_2767,In_1366);
and U4310 (N_4310,In_204,In_2989);
nand U4311 (N_4311,In_1432,In_2134);
nor U4312 (N_4312,In_2350,In_836);
nand U4313 (N_4313,In_1030,In_1807);
and U4314 (N_4314,In_675,In_2118);
nor U4315 (N_4315,In_2558,In_740);
xnor U4316 (N_4316,In_1045,In_1353);
nor U4317 (N_4317,In_1761,In_2666);
nor U4318 (N_4318,In_1551,In_1122);
nand U4319 (N_4319,In_1742,In_1571);
nor U4320 (N_4320,In_1299,In_1760);
nor U4321 (N_4321,In_1794,In_1877);
or U4322 (N_4322,In_2371,In_1018);
and U4323 (N_4323,In_482,In_1408);
xnor U4324 (N_4324,In_1727,In_311);
or U4325 (N_4325,In_746,In_2164);
nor U4326 (N_4326,In_11,In_1857);
xnor U4327 (N_4327,In_280,In_1256);
xor U4328 (N_4328,In_2173,In_605);
nand U4329 (N_4329,In_1028,In_1228);
nand U4330 (N_4330,In_2532,In_148);
or U4331 (N_4331,In_2808,In_1309);
nor U4332 (N_4332,In_1952,In_1060);
or U4333 (N_4333,In_2690,In_994);
nor U4334 (N_4334,In_1930,In_2672);
nand U4335 (N_4335,In_847,In_2226);
xor U4336 (N_4336,In_448,In_787);
xor U4337 (N_4337,In_450,In_2304);
xor U4338 (N_4338,In_2335,In_2305);
or U4339 (N_4339,In_1863,In_591);
and U4340 (N_4340,In_1640,In_1549);
nor U4341 (N_4341,In_1524,In_2279);
or U4342 (N_4342,In_2700,In_842);
nor U4343 (N_4343,In_297,In_2174);
xor U4344 (N_4344,In_2839,In_2028);
and U4345 (N_4345,In_2398,In_2001);
xor U4346 (N_4346,In_1769,In_966);
nand U4347 (N_4347,In_100,In_564);
xor U4348 (N_4348,In_1563,In_1819);
xnor U4349 (N_4349,In_1023,In_2769);
nand U4350 (N_4350,In_2667,In_308);
xor U4351 (N_4351,In_56,In_236);
nor U4352 (N_4352,In_1856,In_2948);
and U4353 (N_4353,In_665,In_378);
xor U4354 (N_4354,In_1737,In_58);
xor U4355 (N_4355,In_1844,In_1998);
xor U4356 (N_4356,In_1240,In_231);
or U4357 (N_4357,In_2802,In_1676);
xor U4358 (N_4358,In_2739,In_2816);
nand U4359 (N_4359,In_1216,In_2478);
nand U4360 (N_4360,In_702,In_1362);
or U4361 (N_4361,In_1586,In_2790);
and U4362 (N_4362,In_450,In_578);
or U4363 (N_4363,In_2757,In_1308);
nand U4364 (N_4364,In_1169,In_1381);
xor U4365 (N_4365,In_435,In_2607);
nand U4366 (N_4366,In_2922,In_882);
xor U4367 (N_4367,In_2174,In_2998);
nand U4368 (N_4368,In_12,In_1187);
nand U4369 (N_4369,In_1298,In_2558);
nand U4370 (N_4370,In_353,In_827);
or U4371 (N_4371,In_2873,In_238);
nor U4372 (N_4372,In_1057,In_2188);
or U4373 (N_4373,In_1644,In_1924);
xnor U4374 (N_4374,In_293,In_1521);
xnor U4375 (N_4375,In_437,In_2250);
nor U4376 (N_4376,In_1527,In_268);
and U4377 (N_4377,In_2382,In_2691);
nand U4378 (N_4378,In_176,In_2295);
or U4379 (N_4379,In_1400,In_2713);
and U4380 (N_4380,In_782,In_1583);
and U4381 (N_4381,In_1035,In_2334);
and U4382 (N_4382,In_866,In_1912);
xor U4383 (N_4383,In_2164,In_1177);
or U4384 (N_4384,In_1547,In_2996);
xor U4385 (N_4385,In_2479,In_1468);
and U4386 (N_4386,In_1152,In_401);
nor U4387 (N_4387,In_2934,In_1458);
nand U4388 (N_4388,In_164,In_1854);
xnor U4389 (N_4389,In_554,In_2251);
or U4390 (N_4390,In_1792,In_2136);
and U4391 (N_4391,In_2056,In_1870);
and U4392 (N_4392,In_1458,In_1709);
and U4393 (N_4393,In_257,In_2479);
and U4394 (N_4394,In_194,In_2583);
xnor U4395 (N_4395,In_939,In_2394);
or U4396 (N_4396,In_1529,In_1974);
xnor U4397 (N_4397,In_2265,In_2319);
nand U4398 (N_4398,In_2861,In_2540);
nand U4399 (N_4399,In_1289,In_2763);
nor U4400 (N_4400,In_1712,In_435);
or U4401 (N_4401,In_2072,In_2090);
or U4402 (N_4402,In_2839,In_2190);
and U4403 (N_4403,In_2623,In_362);
and U4404 (N_4404,In_471,In_1202);
nor U4405 (N_4405,In_2048,In_2101);
nand U4406 (N_4406,In_1570,In_955);
xnor U4407 (N_4407,In_630,In_68);
nand U4408 (N_4408,In_1177,In_144);
and U4409 (N_4409,In_2099,In_70);
or U4410 (N_4410,In_827,In_2672);
and U4411 (N_4411,In_217,In_1407);
nor U4412 (N_4412,In_2222,In_2651);
nor U4413 (N_4413,In_2898,In_2493);
or U4414 (N_4414,In_1770,In_1938);
nand U4415 (N_4415,In_1654,In_311);
xor U4416 (N_4416,In_2573,In_1451);
xnor U4417 (N_4417,In_2463,In_70);
and U4418 (N_4418,In_239,In_1075);
xnor U4419 (N_4419,In_2705,In_950);
and U4420 (N_4420,In_1492,In_2701);
nand U4421 (N_4421,In_2507,In_1315);
and U4422 (N_4422,In_599,In_658);
nor U4423 (N_4423,In_300,In_1330);
and U4424 (N_4424,In_1633,In_544);
and U4425 (N_4425,In_1035,In_891);
xnor U4426 (N_4426,In_745,In_201);
xor U4427 (N_4427,In_318,In_1750);
nand U4428 (N_4428,In_518,In_2614);
nand U4429 (N_4429,In_1534,In_611);
xor U4430 (N_4430,In_173,In_2503);
nor U4431 (N_4431,In_2491,In_1884);
xor U4432 (N_4432,In_1744,In_2590);
or U4433 (N_4433,In_2416,In_1866);
and U4434 (N_4434,In_910,In_1043);
and U4435 (N_4435,In_1177,In_2089);
nand U4436 (N_4436,In_2079,In_2601);
or U4437 (N_4437,In_2034,In_2853);
or U4438 (N_4438,In_864,In_781);
and U4439 (N_4439,In_2944,In_1120);
nand U4440 (N_4440,In_2568,In_2447);
and U4441 (N_4441,In_2377,In_1835);
nor U4442 (N_4442,In_2357,In_853);
or U4443 (N_4443,In_770,In_1399);
xnor U4444 (N_4444,In_1072,In_2549);
xor U4445 (N_4445,In_722,In_457);
nand U4446 (N_4446,In_1253,In_1236);
nand U4447 (N_4447,In_328,In_595);
and U4448 (N_4448,In_2150,In_2639);
or U4449 (N_4449,In_1478,In_147);
and U4450 (N_4450,In_118,In_2343);
or U4451 (N_4451,In_1219,In_2482);
xnor U4452 (N_4452,In_377,In_624);
nor U4453 (N_4453,In_2227,In_2739);
and U4454 (N_4454,In_483,In_1195);
xnor U4455 (N_4455,In_1328,In_155);
or U4456 (N_4456,In_61,In_1163);
or U4457 (N_4457,In_2797,In_840);
nor U4458 (N_4458,In_24,In_1465);
and U4459 (N_4459,In_499,In_1754);
and U4460 (N_4460,In_400,In_504);
nand U4461 (N_4461,In_944,In_798);
nand U4462 (N_4462,In_2800,In_1808);
nor U4463 (N_4463,In_1343,In_35);
or U4464 (N_4464,In_2702,In_888);
nor U4465 (N_4465,In_2782,In_814);
nor U4466 (N_4466,In_2281,In_874);
and U4467 (N_4467,In_2549,In_27);
or U4468 (N_4468,In_1897,In_2373);
or U4469 (N_4469,In_1709,In_1038);
and U4470 (N_4470,In_2990,In_2813);
nand U4471 (N_4471,In_391,In_2236);
nand U4472 (N_4472,In_1590,In_280);
or U4473 (N_4473,In_251,In_2728);
nor U4474 (N_4474,In_2777,In_1984);
and U4475 (N_4475,In_380,In_1201);
xor U4476 (N_4476,In_2840,In_1617);
or U4477 (N_4477,In_2544,In_1057);
nand U4478 (N_4478,In_467,In_351);
nand U4479 (N_4479,In_792,In_2156);
nor U4480 (N_4480,In_579,In_1528);
or U4481 (N_4481,In_2519,In_990);
nor U4482 (N_4482,In_1852,In_311);
nand U4483 (N_4483,In_1317,In_1788);
or U4484 (N_4484,In_121,In_1849);
or U4485 (N_4485,In_1897,In_2372);
and U4486 (N_4486,In_8,In_332);
nor U4487 (N_4487,In_2629,In_2095);
or U4488 (N_4488,In_2552,In_510);
nor U4489 (N_4489,In_406,In_857);
xnor U4490 (N_4490,In_1848,In_444);
or U4491 (N_4491,In_1979,In_20);
nand U4492 (N_4492,In_2916,In_2043);
or U4493 (N_4493,In_283,In_160);
or U4494 (N_4494,In_1377,In_1813);
nor U4495 (N_4495,In_2022,In_1797);
or U4496 (N_4496,In_581,In_1325);
and U4497 (N_4497,In_2517,In_1264);
and U4498 (N_4498,In_2601,In_2241);
nor U4499 (N_4499,In_2654,In_34);
or U4500 (N_4500,In_1579,In_703);
xnor U4501 (N_4501,In_2477,In_1856);
nand U4502 (N_4502,In_1560,In_1979);
nand U4503 (N_4503,In_529,In_511);
or U4504 (N_4504,In_1571,In_22);
or U4505 (N_4505,In_1472,In_1706);
nor U4506 (N_4506,In_1434,In_527);
nand U4507 (N_4507,In_1130,In_2486);
nor U4508 (N_4508,In_97,In_1720);
nor U4509 (N_4509,In_1354,In_2886);
nand U4510 (N_4510,In_1667,In_497);
nand U4511 (N_4511,In_2709,In_1331);
xnor U4512 (N_4512,In_133,In_11);
nor U4513 (N_4513,In_1290,In_963);
xor U4514 (N_4514,In_2547,In_2346);
xor U4515 (N_4515,In_674,In_1290);
and U4516 (N_4516,In_2945,In_872);
xor U4517 (N_4517,In_1487,In_2259);
xnor U4518 (N_4518,In_1661,In_1264);
and U4519 (N_4519,In_1169,In_2882);
nand U4520 (N_4520,In_924,In_2004);
or U4521 (N_4521,In_856,In_443);
nand U4522 (N_4522,In_2137,In_2484);
nand U4523 (N_4523,In_2632,In_666);
nor U4524 (N_4524,In_513,In_1996);
nor U4525 (N_4525,In_616,In_967);
nand U4526 (N_4526,In_2515,In_1960);
and U4527 (N_4527,In_1454,In_2359);
nand U4528 (N_4528,In_690,In_1262);
or U4529 (N_4529,In_178,In_2080);
xor U4530 (N_4530,In_1040,In_894);
nand U4531 (N_4531,In_2671,In_807);
nand U4532 (N_4532,In_741,In_1310);
nand U4533 (N_4533,In_1325,In_1976);
xnor U4534 (N_4534,In_555,In_1761);
or U4535 (N_4535,In_2792,In_947);
nor U4536 (N_4536,In_278,In_1510);
xor U4537 (N_4537,In_2390,In_544);
xor U4538 (N_4538,In_947,In_2565);
or U4539 (N_4539,In_2474,In_478);
nor U4540 (N_4540,In_960,In_1438);
xnor U4541 (N_4541,In_308,In_801);
and U4542 (N_4542,In_254,In_2441);
xnor U4543 (N_4543,In_858,In_1879);
nor U4544 (N_4544,In_181,In_935);
or U4545 (N_4545,In_575,In_1601);
and U4546 (N_4546,In_1634,In_1762);
nand U4547 (N_4547,In_2755,In_379);
and U4548 (N_4548,In_2381,In_2263);
xor U4549 (N_4549,In_2578,In_2704);
or U4550 (N_4550,In_1199,In_270);
nand U4551 (N_4551,In_1989,In_34);
nor U4552 (N_4552,In_2281,In_1860);
or U4553 (N_4553,In_647,In_416);
and U4554 (N_4554,In_430,In_512);
nor U4555 (N_4555,In_2526,In_2190);
and U4556 (N_4556,In_90,In_899);
xor U4557 (N_4557,In_711,In_849);
xnor U4558 (N_4558,In_1931,In_139);
xor U4559 (N_4559,In_2174,In_645);
nand U4560 (N_4560,In_2468,In_2163);
or U4561 (N_4561,In_2996,In_219);
or U4562 (N_4562,In_422,In_297);
nor U4563 (N_4563,In_2682,In_1349);
nor U4564 (N_4564,In_2875,In_871);
xor U4565 (N_4565,In_569,In_1995);
xnor U4566 (N_4566,In_1021,In_2744);
or U4567 (N_4567,In_379,In_1925);
or U4568 (N_4568,In_2493,In_1001);
nor U4569 (N_4569,In_1426,In_972);
xnor U4570 (N_4570,In_2605,In_2110);
nor U4571 (N_4571,In_1366,In_2570);
xnor U4572 (N_4572,In_176,In_1299);
xor U4573 (N_4573,In_2388,In_1319);
and U4574 (N_4574,In_582,In_1523);
nand U4575 (N_4575,In_2502,In_368);
nand U4576 (N_4576,In_1929,In_2800);
and U4577 (N_4577,In_1105,In_1241);
or U4578 (N_4578,In_2077,In_2220);
nor U4579 (N_4579,In_635,In_2425);
nand U4580 (N_4580,In_2145,In_1512);
xnor U4581 (N_4581,In_2175,In_2590);
and U4582 (N_4582,In_2151,In_1075);
xnor U4583 (N_4583,In_2173,In_2687);
and U4584 (N_4584,In_455,In_2578);
xnor U4585 (N_4585,In_697,In_1401);
and U4586 (N_4586,In_2927,In_2973);
nor U4587 (N_4587,In_70,In_2342);
xor U4588 (N_4588,In_254,In_2290);
and U4589 (N_4589,In_2082,In_113);
nor U4590 (N_4590,In_2700,In_839);
nor U4591 (N_4591,In_580,In_2130);
nor U4592 (N_4592,In_1511,In_1873);
nand U4593 (N_4593,In_1672,In_2639);
xnor U4594 (N_4594,In_1439,In_21);
and U4595 (N_4595,In_2488,In_1439);
nor U4596 (N_4596,In_2093,In_2420);
or U4597 (N_4597,In_513,In_1208);
and U4598 (N_4598,In_2611,In_1110);
and U4599 (N_4599,In_2585,In_2747);
nand U4600 (N_4600,In_2527,In_2830);
nor U4601 (N_4601,In_388,In_2936);
nor U4602 (N_4602,In_1820,In_2779);
and U4603 (N_4603,In_2170,In_391);
and U4604 (N_4604,In_149,In_28);
nand U4605 (N_4605,In_587,In_2473);
nand U4606 (N_4606,In_1101,In_426);
xnor U4607 (N_4607,In_2685,In_964);
nor U4608 (N_4608,In_2240,In_1061);
or U4609 (N_4609,In_2472,In_1104);
nand U4610 (N_4610,In_966,In_1812);
nand U4611 (N_4611,In_232,In_1630);
nand U4612 (N_4612,In_342,In_1820);
and U4613 (N_4613,In_2314,In_1799);
or U4614 (N_4614,In_1920,In_2708);
or U4615 (N_4615,In_2970,In_650);
nand U4616 (N_4616,In_2981,In_785);
and U4617 (N_4617,In_1005,In_2856);
and U4618 (N_4618,In_877,In_2205);
and U4619 (N_4619,In_2048,In_782);
or U4620 (N_4620,In_2310,In_418);
nand U4621 (N_4621,In_2530,In_694);
xor U4622 (N_4622,In_541,In_864);
nand U4623 (N_4623,In_768,In_1767);
or U4624 (N_4624,In_2004,In_1864);
nor U4625 (N_4625,In_1548,In_2989);
and U4626 (N_4626,In_2012,In_228);
nor U4627 (N_4627,In_2044,In_1893);
or U4628 (N_4628,In_2410,In_1281);
nand U4629 (N_4629,In_2025,In_2566);
xnor U4630 (N_4630,In_2404,In_410);
nand U4631 (N_4631,In_1854,In_2419);
and U4632 (N_4632,In_1017,In_782);
nand U4633 (N_4633,In_1325,In_292);
and U4634 (N_4634,In_997,In_2830);
nor U4635 (N_4635,In_1168,In_920);
and U4636 (N_4636,In_1406,In_822);
or U4637 (N_4637,In_1072,In_157);
nand U4638 (N_4638,In_750,In_984);
xor U4639 (N_4639,In_879,In_1355);
nand U4640 (N_4640,In_1437,In_2965);
or U4641 (N_4641,In_2861,In_1056);
nand U4642 (N_4642,In_1499,In_1094);
xnor U4643 (N_4643,In_1935,In_793);
nor U4644 (N_4644,In_1890,In_2078);
or U4645 (N_4645,In_1744,In_1703);
or U4646 (N_4646,In_1699,In_2707);
nand U4647 (N_4647,In_1070,In_1265);
nor U4648 (N_4648,In_1146,In_2063);
nand U4649 (N_4649,In_238,In_2833);
nand U4650 (N_4650,In_1656,In_1008);
nand U4651 (N_4651,In_1801,In_30);
and U4652 (N_4652,In_1236,In_1678);
nand U4653 (N_4653,In_305,In_1713);
or U4654 (N_4654,In_1591,In_623);
nor U4655 (N_4655,In_2155,In_2130);
and U4656 (N_4656,In_2467,In_970);
and U4657 (N_4657,In_2424,In_1612);
and U4658 (N_4658,In_1414,In_2678);
nor U4659 (N_4659,In_1832,In_1202);
and U4660 (N_4660,In_2130,In_2984);
xnor U4661 (N_4661,In_173,In_2600);
nand U4662 (N_4662,In_1838,In_2601);
nor U4663 (N_4663,In_2056,In_2655);
xnor U4664 (N_4664,In_1590,In_814);
xor U4665 (N_4665,In_453,In_71);
nand U4666 (N_4666,In_857,In_1677);
nor U4667 (N_4667,In_2289,In_1336);
nor U4668 (N_4668,In_1299,In_2927);
and U4669 (N_4669,In_134,In_1920);
nor U4670 (N_4670,In_777,In_1032);
and U4671 (N_4671,In_1507,In_2402);
or U4672 (N_4672,In_1136,In_436);
or U4673 (N_4673,In_819,In_781);
xnor U4674 (N_4674,In_899,In_2081);
xor U4675 (N_4675,In_2637,In_2909);
or U4676 (N_4676,In_66,In_974);
nand U4677 (N_4677,In_899,In_2841);
and U4678 (N_4678,In_674,In_1182);
or U4679 (N_4679,In_2065,In_1699);
xor U4680 (N_4680,In_1232,In_2921);
and U4681 (N_4681,In_2616,In_2642);
nor U4682 (N_4682,In_0,In_1254);
or U4683 (N_4683,In_1457,In_324);
and U4684 (N_4684,In_2231,In_2294);
or U4685 (N_4685,In_2857,In_2892);
xor U4686 (N_4686,In_60,In_708);
or U4687 (N_4687,In_2585,In_2215);
nand U4688 (N_4688,In_2939,In_2505);
and U4689 (N_4689,In_2040,In_1923);
xor U4690 (N_4690,In_601,In_205);
nand U4691 (N_4691,In_1525,In_367);
or U4692 (N_4692,In_2132,In_1366);
and U4693 (N_4693,In_2147,In_775);
nand U4694 (N_4694,In_1515,In_809);
xnor U4695 (N_4695,In_827,In_740);
or U4696 (N_4696,In_2460,In_281);
xnor U4697 (N_4697,In_1128,In_1597);
or U4698 (N_4698,In_1500,In_919);
xor U4699 (N_4699,In_1018,In_1410);
or U4700 (N_4700,In_676,In_469);
and U4701 (N_4701,In_1230,In_2579);
nand U4702 (N_4702,In_191,In_142);
nand U4703 (N_4703,In_2107,In_574);
nand U4704 (N_4704,In_2052,In_1973);
xnor U4705 (N_4705,In_2657,In_248);
and U4706 (N_4706,In_263,In_1275);
nand U4707 (N_4707,In_2250,In_1803);
nor U4708 (N_4708,In_2276,In_1792);
and U4709 (N_4709,In_867,In_2875);
xnor U4710 (N_4710,In_2824,In_2483);
nor U4711 (N_4711,In_2206,In_1072);
or U4712 (N_4712,In_2052,In_2939);
xor U4713 (N_4713,In_165,In_2174);
nor U4714 (N_4714,In_1928,In_328);
nand U4715 (N_4715,In_2936,In_1463);
xor U4716 (N_4716,In_2424,In_54);
and U4717 (N_4717,In_675,In_1902);
or U4718 (N_4718,In_1508,In_1700);
and U4719 (N_4719,In_658,In_2453);
xor U4720 (N_4720,In_196,In_600);
nor U4721 (N_4721,In_2836,In_1722);
or U4722 (N_4722,In_2192,In_1067);
or U4723 (N_4723,In_2412,In_1477);
nor U4724 (N_4724,In_282,In_2154);
nand U4725 (N_4725,In_2596,In_2400);
xor U4726 (N_4726,In_1893,In_1697);
nand U4727 (N_4727,In_2764,In_1098);
nor U4728 (N_4728,In_2998,In_2218);
nand U4729 (N_4729,In_2597,In_225);
nand U4730 (N_4730,In_1048,In_1405);
xor U4731 (N_4731,In_220,In_377);
nor U4732 (N_4732,In_2762,In_2342);
or U4733 (N_4733,In_2961,In_2806);
and U4734 (N_4734,In_2669,In_1628);
xnor U4735 (N_4735,In_1146,In_723);
or U4736 (N_4736,In_1673,In_65);
or U4737 (N_4737,In_600,In_1235);
nor U4738 (N_4738,In_2996,In_2421);
and U4739 (N_4739,In_1521,In_391);
nand U4740 (N_4740,In_1805,In_2922);
nor U4741 (N_4741,In_680,In_33);
nor U4742 (N_4742,In_1245,In_909);
xnor U4743 (N_4743,In_2900,In_1992);
nand U4744 (N_4744,In_1686,In_1786);
nor U4745 (N_4745,In_1635,In_1951);
and U4746 (N_4746,In_1419,In_229);
xor U4747 (N_4747,In_934,In_85);
nand U4748 (N_4748,In_65,In_2696);
and U4749 (N_4749,In_560,In_112);
and U4750 (N_4750,In_1009,In_889);
or U4751 (N_4751,In_850,In_1055);
nor U4752 (N_4752,In_202,In_1194);
nand U4753 (N_4753,In_2850,In_750);
nor U4754 (N_4754,In_2476,In_2960);
or U4755 (N_4755,In_2730,In_564);
xnor U4756 (N_4756,In_598,In_1598);
or U4757 (N_4757,In_2542,In_2685);
nor U4758 (N_4758,In_692,In_209);
nand U4759 (N_4759,In_1152,In_2300);
nand U4760 (N_4760,In_2123,In_0);
nor U4761 (N_4761,In_894,In_671);
or U4762 (N_4762,In_2757,In_2299);
xnor U4763 (N_4763,In_1174,In_77);
xnor U4764 (N_4764,In_1085,In_762);
or U4765 (N_4765,In_153,In_149);
nand U4766 (N_4766,In_1264,In_269);
nand U4767 (N_4767,In_918,In_379);
nand U4768 (N_4768,In_58,In_2835);
or U4769 (N_4769,In_1864,In_2575);
nor U4770 (N_4770,In_1930,In_935);
xnor U4771 (N_4771,In_1949,In_157);
or U4772 (N_4772,In_2266,In_316);
and U4773 (N_4773,In_110,In_395);
or U4774 (N_4774,In_2033,In_146);
nand U4775 (N_4775,In_2082,In_1089);
nor U4776 (N_4776,In_2262,In_897);
nand U4777 (N_4777,In_1085,In_751);
and U4778 (N_4778,In_1187,In_265);
nand U4779 (N_4779,In_1416,In_904);
nor U4780 (N_4780,In_988,In_2865);
nand U4781 (N_4781,In_2281,In_2017);
and U4782 (N_4782,In_2282,In_378);
or U4783 (N_4783,In_2678,In_93);
xnor U4784 (N_4784,In_429,In_2108);
nand U4785 (N_4785,In_1376,In_1486);
or U4786 (N_4786,In_1054,In_178);
nor U4787 (N_4787,In_2496,In_1002);
nand U4788 (N_4788,In_1753,In_1582);
nand U4789 (N_4789,In_0,In_2443);
nor U4790 (N_4790,In_981,In_2629);
or U4791 (N_4791,In_1419,In_2355);
xnor U4792 (N_4792,In_615,In_2956);
nand U4793 (N_4793,In_2902,In_1910);
nand U4794 (N_4794,In_2715,In_2705);
nand U4795 (N_4795,In_1368,In_1651);
and U4796 (N_4796,In_2376,In_2846);
xor U4797 (N_4797,In_2095,In_1363);
xnor U4798 (N_4798,In_190,In_1245);
nand U4799 (N_4799,In_426,In_2947);
nand U4800 (N_4800,In_1808,In_2414);
nor U4801 (N_4801,In_1595,In_1410);
or U4802 (N_4802,In_2078,In_1351);
and U4803 (N_4803,In_2193,In_976);
or U4804 (N_4804,In_924,In_662);
or U4805 (N_4805,In_2199,In_2625);
nand U4806 (N_4806,In_2711,In_591);
nand U4807 (N_4807,In_1946,In_777);
or U4808 (N_4808,In_1970,In_1473);
nand U4809 (N_4809,In_2246,In_2837);
or U4810 (N_4810,In_792,In_1083);
and U4811 (N_4811,In_1691,In_548);
and U4812 (N_4812,In_1940,In_1356);
or U4813 (N_4813,In_398,In_364);
nor U4814 (N_4814,In_1225,In_1745);
or U4815 (N_4815,In_1205,In_762);
nand U4816 (N_4816,In_870,In_2148);
xnor U4817 (N_4817,In_1155,In_2425);
nor U4818 (N_4818,In_2494,In_127);
xnor U4819 (N_4819,In_676,In_896);
xnor U4820 (N_4820,In_1316,In_2960);
and U4821 (N_4821,In_2861,In_879);
nand U4822 (N_4822,In_2258,In_2474);
nor U4823 (N_4823,In_809,In_1952);
or U4824 (N_4824,In_1048,In_163);
and U4825 (N_4825,In_2570,In_2909);
or U4826 (N_4826,In_2618,In_868);
nor U4827 (N_4827,In_848,In_1234);
nor U4828 (N_4828,In_576,In_466);
xor U4829 (N_4829,In_2331,In_2647);
and U4830 (N_4830,In_2631,In_838);
or U4831 (N_4831,In_724,In_2777);
nand U4832 (N_4832,In_549,In_1728);
xnor U4833 (N_4833,In_1510,In_1325);
xor U4834 (N_4834,In_1060,In_1691);
nand U4835 (N_4835,In_2243,In_1350);
xnor U4836 (N_4836,In_1358,In_1636);
or U4837 (N_4837,In_2977,In_695);
nor U4838 (N_4838,In_1389,In_2539);
nor U4839 (N_4839,In_944,In_1457);
nand U4840 (N_4840,In_581,In_2672);
xor U4841 (N_4841,In_332,In_383);
and U4842 (N_4842,In_2457,In_1508);
nand U4843 (N_4843,In_2442,In_2749);
and U4844 (N_4844,In_1979,In_419);
and U4845 (N_4845,In_2385,In_2168);
or U4846 (N_4846,In_916,In_1379);
nand U4847 (N_4847,In_2708,In_774);
and U4848 (N_4848,In_183,In_663);
nand U4849 (N_4849,In_419,In_2345);
xor U4850 (N_4850,In_1133,In_1820);
or U4851 (N_4851,In_2066,In_1996);
or U4852 (N_4852,In_578,In_2603);
or U4853 (N_4853,In_732,In_2089);
nor U4854 (N_4854,In_753,In_1847);
xnor U4855 (N_4855,In_1883,In_2060);
or U4856 (N_4856,In_1389,In_862);
nor U4857 (N_4857,In_2797,In_1895);
xnor U4858 (N_4858,In_2037,In_618);
or U4859 (N_4859,In_1795,In_799);
or U4860 (N_4860,In_1044,In_2181);
xor U4861 (N_4861,In_830,In_1893);
xor U4862 (N_4862,In_1305,In_1437);
nand U4863 (N_4863,In_2733,In_1704);
xor U4864 (N_4864,In_1042,In_2875);
xor U4865 (N_4865,In_2227,In_1271);
and U4866 (N_4866,In_262,In_2455);
and U4867 (N_4867,In_1856,In_2288);
and U4868 (N_4868,In_2660,In_1774);
or U4869 (N_4869,In_668,In_2226);
and U4870 (N_4870,In_820,In_1027);
nand U4871 (N_4871,In_2588,In_1514);
and U4872 (N_4872,In_159,In_2519);
nand U4873 (N_4873,In_2936,In_1467);
nand U4874 (N_4874,In_2114,In_1275);
or U4875 (N_4875,In_597,In_1086);
and U4876 (N_4876,In_616,In_661);
or U4877 (N_4877,In_2106,In_2999);
xnor U4878 (N_4878,In_198,In_679);
xor U4879 (N_4879,In_2015,In_863);
and U4880 (N_4880,In_1945,In_1910);
nor U4881 (N_4881,In_2514,In_378);
xnor U4882 (N_4882,In_1837,In_2770);
nor U4883 (N_4883,In_2015,In_2765);
or U4884 (N_4884,In_1853,In_2472);
nand U4885 (N_4885,In_1733,In_2041);
and U4886 (N_4886,In_2388,In_362);
or U4887 (N_4887,In_1387,In_199);
or U4888 (N_4888,In_198,In_1069);
and U4889 (N_4889,In_359,In_574);
and U4890 (N_4890,In_488,In_2591);
xor U4891 (N_4891,In_2048,In_1637);
or U4892 (N_4892,In_1631,In_540);
xnor U4893 (N_4893,In_925,In_2696);
nor U4894 (N_4894,In_1565,In_925);
nand U4895 (N_4895,In_2944,In_1070);
and U4896 (N_4896,In_2101,In_2619);
or U4897 (N_4897,In_438,In_2640);
xor U4898 (N_4898,In_897,In_2449);
nand U4899 (N_4899,In_2463,In_2078);
nor U4900 (N_4900,In_795,In_2486);
nor U4901 (N_4901,In_2100,In_1929);
and U4902 (N_4902,In_2912,In_1168);
xnor U4903 (N_4903,In_2864,In_2284);
or U4904 (N_4904,In_1838,In_2147);
and U4905 (N_4905,In_2944,In_196);
and U4906 (N_4906,In_1592,In_674);
and U4907 (N_4907,In_644,In_1207);
or U4908 (N_4908,In_1343,In_1653);
nor U4909 (N_4909,In_2324,In_2065);
or U4910 (N_4910,In_1956,In_1001);
nand U4911 (N_4911,In_1293,In_699);
nand U4912 (N_4912,In_2130,In_937);
or U4913 (N_4913,In_2476,In_2903);
nand U4914 (N_4914,In_740,In_1439);
and U4915 (N_4915,In_1034,In_1604);
nor U4916 (N_4916,In_1074,In_961);
and U4917 (N_4917,In_1076,In_2537);
or U4918 (N_4918,In_1593,In_845);
nand U4919 (N_4919,In_1563,In_862);
xnor U4920 (N_4920,In_1945,In_2544);
nand U4921 (N_4921,In_2945,In_695);
nor U4922 (N_4922,In_2810,In_2150);
nor U4923 (N_4923,In_13,In_522);
xnor U4924 (N_4924,In_1388,In_2605);
and U4925 (N_4925,In_2870,In_2553);
and U4926 (N_4926,In_309,In_2097);
xnor U4927 (N_4927,In_2429,In_2335);
nand U4928 (N_4928,In_719,In_2142);
nor U4929 (N_4929,In_479,In_1171);
and U4930 (N_4930,In_1962,In_330);
or U4931 (N_4931,In_373,In_2829);
nand U4932 (N_4932,In_199,In_2081);
or U4933 (N_4933,In_2771,In_268);
or U4934 (N_4934,In_2065,In_2597);
xnor U4935 (N_4935,In_2263,In_2610);
xor U4936 (N_4936,In_1904,In_2916);
nand U4937 (N_4937,In_794,In_2575);
or U4938 (N_4938,In_1978,In_527);
xor U4939 (N_4939,In_550,In_1963);
and U4940 (N_4940,In_1534,In_2777);
xnor U4941 (N_4941,In_1127,In_1431);
nand U4942 (N_4942,In_522,In_796);
xnor U4943 (N_4943,In_1419,In_295);
nor U4944 (N_4944,In_2569,In_1310);
xor U4945 (N_4945,In_139,In_1174);
or U4946 (N_4946,In_1532,In_1903);
and U4947 (N_4947,In_329,In_1919);
nor U4948 (N_4948,In_1587,In_2722);
nor U4949 (N_4949,In_1822,In_1513);
xnor U4950 (N_4950,In_2596,In_1411);
and U4951 (N_4951,In_2969,In_1199);
nor U4952 (N_4952,In_1643,In_1975);
nand U4953 (N_4953,In_2301,In_1427);
nand U4954 (N_4954,In_921,In_2679);
nand U4955 (N_4955,In_2779,In_73);
nand U4956 (N_4956,In_2609,In_871);
or U4957 (N_4957,In_2610,In_361);
nand U4958 (N_4958,In_82,In_2941);
and U4959 (N_4959,In_1621,In_1215);
or U4960 (N_4960,In_2742,In_1149);
and U4961 (N_4961,In_2154,In_2447);
or U4962 (N_4962,In_2471,In_779);
nand U4963 (N_4963,In_2978,In_1053);
nor U4964 (N_4964,In_1925,In_956);
and U4965 (N_4965,In_2589,In_295);
or U4966 (N_4966,In_841,In_2605);
nand U4967 (N_4967,In_2054,In_1639);
or U4968 (N_4968,In_1948,In_1239);
nand U4969 (N_4969,In_132,In_1900);
nor U4970 (N_4970,In_1455,In_32);
or U4971 (N_4971,In_1575,In_906);
nor U4972 (N_4972,In_1769,In_2625);
or U4973 (N_4973,In_2997,In_588);
and U4974 (N_4974,In_2610,In_1464);
nor U4975 (N_4975,In_187,In_1146);
xnor U4976 (N_4976,In_2194,In_725);
and U4977 (N_4977,In_2139,In_1869);
xor U4978 (N_4978,In_1759,In_2009);
nand U4979 (N_4979,In_2384,In_2645);
xnor U4980 (N_4980,In_833,In_1957);
nand U4981 (N_4981,In_812,In_632);
or U4982 (N_4982,In_1199,In_2367);
nor U4983 (N_4983,In_649,In_2424);
nor U4984 (N_4984,In_1844,In_1464);
nor U4985 (N_4985,In_2206,In_1816);
or U4986 (N_4986,In_317,In_2531);
or U4987 (N_4987,In_276,In_888);
nor U4988 (N_4988,In_2893,In_1870);
nor U4989 (N_4989,In_2420,In_39);
nand U4990 (N_4990,In_1779,In_452);
nand U4991 (N_4991,In_2003,In_2990);
xnor U4992 (N_4992,In_2911,In_2063);
or U4993 (N_4993,In_1920,In_567);
nor U4994 (N_4994,In_1856,In_1060);
and U4995 (N_4995,In_438,In_2182);
and U4996 (N_4996,In_2583,In_2340);
nand U4997 (N_4997,In_1593,In_2611);
and U4998 (N_4998,In_2957,In_350);
nor U4999 (N_4999,In_1620,In_2444);
or U5000 (N_5000,N_2600,N_298);
nand U5001 (N_5001,N_3746,N_252);
or U5002 (N_5002,N_1697,N_779);
nor U5003 (N_5003,N_1287,N_1925);
xnor U5004 (N_5004,N_4574,N_1542);
or U5005 (N_5005,N_2087,N_4415);
nor U5006 (N_5006,N_3922,N_2203);
nand U5007 (N_5007,N_3755,N_3056);
nor U5008 (N_5008,N_4303,N_1225);
nand U5009 (N_5009,N_1465,N_2903);
nor U5010 (N_5010,N_1122,N_3582);
or U5011 (N_5011,N_2367,N_344);
and U5012 (N_5012,N_1301,N_2052);
and U5013 (N_5013,N_559,N_3046);
xor U5014 (N_5014,N_1099,N_1018);
xor U5015 (N_5015,N_4254,N_2125);
xor U5016 (N_5016,N_625,N_3917);
and U5017 (N_5017,N_2807,N_2599);
nand U5018 (N_5018,N_1083,N_2827);
and U5019 (N_5019,N_3790,N_2047);
xnor U5020 (N_5020,N_3331,N_712);
and U5021 (N_5021,N_3739,N_4359);
xor U5022 (N_5022,N_4457,N_2794);
and U5023 (N_5023,N_1919,N_2665);
xor U5024 (N_5024,N_4585,N_2050);
or U5025 (N_5025,N_2431,N_4403);
or U5026 (N_5026,N_642,N_498);
nand U5027 (N_5027,N_576,N_4396);
nand U5028 (N_5028,N_304,N_973);
xnor U5029 (N_5029,N_2967,N_3016);
or U5030 (N_5030,N_2963,N_4862);
nand U5031 (N_5031,N_362,N_1050);
or U5032 (N_5032,N_1551,N_2057);
nand U5033 (N_5033,N_1887,N_1505);
xor U5034 (N_5034,N_1516,N_3152);
nand U5035 (N_5035,N_4888,N_1853);
and U5036 (N_5036,N_2316,N_2675);
nor U5037 (N_5037,N_4247,N_1237);
xnor U5038 (N_5038,N_2091,N_721);
and U5039 (N_5039,N_4795,N_3212);
and U5040 (N_5040,N_2915,N_674);
nand U5041 (N_5041,N_2005,N_4905);
nand U5042 (N_5042,N_81,N_554);
or U5043 (N_5043,N_4262,N_3261);
and U5044 (N_5044,N_600,N_832);
or U5045 (N_5045,N_4,N_862);
xor U5046 (N_5046,N_341,N_3438);
xnor U5047 (N_5047,N_3565,N_3224);
and U5048 (N_5048,N_3829,N_2575);
xnor U5049 (N_5049,N_1259,N_1860);
nand U5050 (N_5050,N_651,N_3504);
nor U5051 (N_5051,N_4335,N_2064);
xor U5052 (N_5052,N_164,N_4987);
nor U5053 (N_5053,N_3428,N_3758);
xnor U5054 (N_5054,N_1147,N_2760);
nand U5055 (N_5055,N_3168,N_3411);
or U5056 (N_5056,N_4828,N_3809);
nor U5057 (N_5057,N_3815,N_3656);
nor U5058 (N_5058,N_1052,N_3867);
and U5059 (N_5059,N_4505,N_2448);
or U5060 (N_5060,N_450,N_3921);
or U5061 (N_5061,N_3419,N_3886);
xnor U5062 (N_5062,N_1833,N_1086);
or U5063 (N_5063,N_123,N_3734);
nor U5064 (N_5064,N_620,N_3812);
xnor U5065 (N_5065,N_3130,N_242);
xnor U5066 (N_5066,N_3598,N_352);
nand U5067 (N_5067,N_162,N_301);
and U5068 (N_5068,N_283,N_2364);
nor U5069 (N_5069,N_2116,N_328);
nor U5070 (N_5070,N_4044,N_2099);
nand U5071 (N_5071,N_3410,N_438);
or U5072 (N_5072,N_1514,N_4410);
or U5073 (N_5073,N_4842,N_4550);
nor U5074 (N_5074,N_2,N_1213);
nand U5075 (N_5075,N_1377,N_2202);
nor U5076 (N_5076,N_1474,N_813);
nor U5077 (N_5077,N_4840,N_3024);
nor U5078 (N_5078,N_4789,N_3554);
xor U5079 (N_5079,N_4437,N_4409);
nor U5080 (N_5080,N_3021,N_2508);
and U5081 (N_5081,N_4259,N_3763);
and U5082 (N_5082,N_4418,N_3521);
nand U5083 (N_5083,N_4204,N_1778);
nor U5084 (N_5084,N_349,N_2013);
nor U5085 (N_5085,N_2654,N_3690);
nor U5086 (N_5086,N_756,N_1023);
or U5087 (N_5087,N_4103,N_4826);
nand U5088 (N_5088,N_1262,N_4628);
and U5089 (N_5089,N_2918,N_1317);
and U5090 (N_5090,N_1995,N_4273);
and U5091 (N_5091,N_1634,N_639);
nand U5092 (N_5092,N_1340,N_59);
xor U5093 (N_5093,N_811,N_2400);
or U5094 (N_5094,N_4343,N_4730);
xor U5095 (N_5095,N_3696,N_1970);
nor U5096 (N_5096,N_2892,N_87);
nor U5097 (N_5097,N_2060,N_4707);
xnor U5098 (N_5098,N_3463,N_1762);
or U5099 (N_5099,N_901,N_595);
or U5100 (N_5100,N_983,N_3707);
and U5101 (N_5101,N_1600,N_4600);
and U5102 (N_5102,N_4670,N_1367);
or U5103 (N_5103,N_4007,N_1884);
nand U5104 (N_5104,N_2983,N_696);
nand U5105 (N_5105,N_3190,N_4733);
nor U5106 (N_5106,N_3450,N_999);
nand U5107 (N_5107,N_68,N_4200);
or U5108 (N_5108,N_2185,N_4294);
nand U5109 (N_5109,N_2233,N_2707);
xnor U5110 (N_5110,N_4079,N_214);
or U5111 (N_5111,N_2289,N_4560);
nand U5112 (N_5112,N_4006,N_3742);
nand U5113 (N_5113,N_4025,N_4414);
nand U5114 (N_5114,N_2608,N_1700);
and U5115 (N_5115,N_556,N_4228);
and U5116 (N_5116,N_2634,N_1628);
or U5117 (N_5117,N_3091,N_4784);
or U5118 (N_5118,N_1299,N_3782);
and U5119 (N_5119,N_53,N_4356);
xor U5120 (N_5120,N_951,N_3013);
and U5121 (N_5121,N_1011,N_1730);
nand U5122 (N_5122,N_3377,N_241);
nand U5123 (N_5123,N_2257,N_2811);
xor U5124 (N_5124,N_1092,N_4990);
nor U5125 (N_5125,N_515,N_157);
nor U5126 (N_5126,N_1771,N_3749);
or U5127 (N_5127,N_3292,N_546);
or U5128 (N_5128,N_1358,N_1321);
or U5129 (N_5129,N_3641,N_1392);
xnor U5130 (N_5130,N_1246,N_4351);
and U5131 (N_5131,N_2616,N_4774);
or U5132 (N_5132,N_3165,N_3219);
nand U5133 (N_5133,N_3811,N_3381);
and U5134 (N_5134,N_1175,N_1531);
xor U5135 (N_5135,N_1777,N_3630);
or U5136 (N_5136,N_1654,N_3129);
and U5137 (N_5137,N_3394,N_4700);
xor U5138 (N_5138,N_2721,N_2861);
and U5139 (N_5139,N_4704,N_1934);
nand U5140 (N_5140,N_3706,N_264);
xnor U5141 (N_5141,N_1360,N_2279);
or U5142 (N_5142,N_4357,N_219);
nand U5143 (N_5143,N_1864,N_259);
and U5144 (N_5144,N_4684,N_329);
nand U5145 (N_5145,N_930,N_2323);
and U5146 (N_5146,N_3629,N_3184);
nor U5147 (N_5147,N_4541,N_3638);
or U5148 (N_5148,N_1624,N_711);
nand U5149 (N_5149,N_158,N_2979);
and U5150 (N_5150,N_2375,N_2399);
or U5151 (N_5151,N_1565,N_3666);
and U5152 (N_5152,N_2831,N_695);
nor U5153 (N_5153,N_1193,N_3540);
and U5154 (N_5154,N_955,N_3857);
nand U5155 (N_5155,N_413,N_824);
nor U5156 (N_5156,N_4520,N_1732);
nor U5157 (N_5157,N_3273,N_3303);
nand U5158 (N_5158,N_1064,N_3090);
and U5159 (N_5159,N_24,N_874);
xnor U5160 (N_5160,N_3290,N_3839);
nand U5161 (N_5161,N_3341,N_3532);
and U5162 (N_5162,N_1486,N_4597);
xnor U5163 (N_5163,N_2026,N_322);
xor U5164 (N_5164,N_4101,N_4782);
or U5165 (N_5165,N_2871,N_3388);
xor U5166 (N_5166,N_309,N_3076);
xor U5167 (N_5167,N_3316,N_3467);
nand U5168 (N_5168,N_927,N_466);
or U5169 (N_5169,N_2998,N_3126);
nand U5170 (N_5170,N_79,N_4720);
and U5171 (N_5171,N_452,N_4102);
and U5172 (N_5172,N_2914,N_2816);
and U5173 (N_5173,N_631,N_4408);
xor U5174 (N_5174,N_2910,N_3896);
nand U5175 (N_5175,N_1570,N_3157);
and U5176 (N_5176,N_1649,N_4321);
and U5177 (N_5177,N_3835,N_43);
nand U5178 (N_5178,N_2336,N_3110);
or U5179 (N_5179,N_1578,N_3133);
xor U5180 (N_5180,N_111,N_4794);
nor U5181 (N_5181,N_2950,N_1170);
and U5182 (N_5182,N_3553,N_3893);
and U5183 (N_5183,N_4918,N_869);
and U5184 (N_5184,N_3300,N_1047);
nand U5185 (N_5185,N_4275,N_4093);
nand U5186 (N_5186,N_240,N_3193);
nor U5187 (N_5187,N_1110,N_2614);
nor U5188 (N_5188,N_1524,N_110);
and U5189 (N_5189,N_4646,N_3862);
nand U5190 (N_5190,N_211,N_3607);
or U5191 (N_5191,N_4923,N_3201);
and U5192 (N_5192,N_2456,N_1491);
xor U5193 (N_5193,N_4516,N_3590);
xor U5194 (N_5194,N_4999,N_4014);
nand U5195 (N_5195,N_2775,N_3564);
xor U5196 (N_5196,N_655,N_4711);
nor U5197 (N_5197,N_2247,N_589);
xor U5198 (N_5198,N_98,N_1822);
and U5199 (N_5199,N_212,N_2096);
and U5200 (N_5200,N_3580,N_2529);
xnor U5201 (N_5201,N_1109,N_1717);
xor U5202 (N_5202,N_3938,N_1209);
nor U5203 (N_5203,N_582,N_2045);
nor U5204 (N_5204,N_1954,N_3485);
xnor U5205 (N_5205,N_4757,N_3055);
nand U5206 (N_5206,N_13,N_3964);
nand U5207 (N_5207,N_3744,N_3628);
or U5208 (N_5208,N_4816,N_4120);
or U5209 (N_5209,N_2261,N_4345);
or U5210 (N_5210,N_2221,N_2120);
nand U5211 (N_5211,N_2539,N_4797);
nand U5212 (N_5212,N_665,N_4777);
and U5213 (N_5213,N_688,N_4282);
nand U5214 (N_5214,N_1585,N_16);
and U5215 (N_5215,N_1966,N_1855);
xor U5216 (N_5216,N_3900,N_4595);
xor U5217 (N_5217,N_1346,N_3894);
and U5218 (N_5218,N_3956,N_3285);
nand U5219 (N_5219,N_2660,N_2768);
xnor U5220 (N_5220,N_2516,N_1810);
nand U5221 (N_5221,N_3669,N_4703);
nor U5222 (N_5222,N_2882,N_691);
or U5223 (N_5223,N_1280,N_1488);
nand U5224 (N_5224,N_2372,N_161);
xor U5225 (N_5225,N_464,N_1245);
or U5226 (N_5226,N_4189,N_2310);
xor U5227 (N_5227,N_1386,N_3724);
and U5228 (N_5228,N_1057,N_2236);
xor U5229 (N_5229,N_4499,N_2278);
and U5230 (N_5230,N_3281,N_1710);
and U5231 (N_5231,N_825,N_1535);
nand U5232 (N_5232,N_1908,N_147);
xnor U5233 (N_5233,N_3636,N_2497);
and U5234 (N_5234,N_2685,N_3716);
xnor U5235 (N_5235,N_4253,N_4504);
nand U5236 (N_5236,N_202,N_3328);
nor U5237 (N_5237,N_3041,N_1418);
nand U5238 (N_5238,N_3246,N_3537);
nor U5239 (N_5239,N_2636,N_3032);
nor U5240 (N_5240,N_2752,N_3362);
and U5241 (N_5241,N_1435,N_960);
and U5242 (N_5242,N_4592,N_1338);
or U5243 (N_5243,N_1160,N_1759);
nand U5244 (N_5244,N_1638,N_3748);
xor U5245 (N_5245,N_117,N_3351);
nor U5246 (N_5246,N_1070,N_4121);
nor U5247 (N_5247,N_2897,N_2063);
nor U5248 (N_5248,N_4953,N_1823);
xnor U5249 (N_5249,N_412,N_3353);
nor U5250 (N_5250,N_3405,N_1029);
or U5251 (N_5251,N_3586,N_2702);
xor U5252 (N_5252,N_166,N_2435);
xnor U5253 (N_5253,N_47,N_4696);
or U5254 (N_5254,N_45,N_947);
or U5255 (N_5255,N_2952,N_3712);
xor U5256 (N_5256,N_2040,N_1967);
or U5257 (N_5257,N_4822,N_1081);
nand U5258 (N_5258,N_3287,N_4274);
xnor U5259 (N_5259,N_2444,N_4448);
and U5260 (N_5260,N_2075,N_2533);
or U5261 (N_5261,N_3806,N_2422);
and U5262 (N_5262,N_4861,N_1827);
and U5263 (N_5263,N_4658,N_1623);
and U5264 (N_5264,N_424,N_4529);
xnor U5265 (N_5265,N_1519,N_1975);
or U5266 (N_5266,N_565,N_4665);
xor U5267 (N_5267,N_2281,N_1767);
or U5268 (N_5268,N_2568,N_1492);
nor U5269 (N_5269,N_3196,N_3665);
or U5270 (N_5270,N_4527,N_4683);
and U5271 (N_5271,N_3169,N_2962);
and U5272 (N_5272,N_2157,N_2274);
nand U5273 (N_5273,N_3424,N_4366);
or U5274 (N_5274,N_933,N_4232);
nor U5275 (N_5275,N_2839,N_2030);
or U5276 (N_5276,N_1063,N_4059);
nor U5277 (N_5277,N_1243,N_1330);
or U5278 (N_5278,N_577,N_1879);
and U5279 (N_5279,N_4019,N_1312);
xor U5280 (N_5280,N_2085,N_3167);
nand U5281 (N_5281,N_28,N_611);
and U5282 (N_5282,N_4399,N_988);
or U5283 (N_5283,N_4258,N_566);
nand U5284 (N_5284,N_932,N_4892);
or U5285 (N_5285,N_397,N_2392);
xnor U5286 (N_5286,N_4444,N_4779);
nor U5287 (N_5287,N_4545,N_2272);
xnor U5288 (N_5288,N_1438,N_1441);
and U5289 (N_5289,N_3144,N_2813);
or U5290 (N_5290,N_3530,N_1460);
or U5291 (N_5291,N_492,N_4713);
and U5292 (N_5292,N_4113,N_1252);
nand U5293 (N_5293,N_3510,N_2517);
nor U5294 (N_5294,N_1998,N_1690);
or U5295 (N_5295,N_431,N_2264);
xnor U5296 (N_5296,N_2408,N_463);
xor U5297 (N_5297,N_2809,N_1475);
or U5298 (N_5298,N_3158,N_4078);
xnor U5299 (N_5299,N_4706,N_2713);
xnor U5300 (N_5300,N_1283,N_2668);
or U5301 (N_5301,N_3124,N_3087);
nor U5302 (N_5302,N_3545,N_261);
nor U5303 (N_5303,N_1261,N_529);
xnor U5304 (N_5304,N_1899,N_3804);
and U5305 (N_5305,N_4949,N_539);
xor U5306 (N_5306,N_1150,N_3721);
nand U5307 (N_5307,N_1674,N_4559);
nor U5308 (N_5308,N_1646,N_2416);
nor U5309 (N_5309,N_2450,N_4947);
xnor U5310 (N_5310,N_3408,N_1381);
nand U5311 (N_5311,N_3719,N_135);
xnor U5312 (N_5312,N_2232,N_4391);
or U5313 (N_5313,N_912,N_1902);
nand U5314 (N_5314,N_3093,N_3741);
nor U5315 (N_5315,N_1764,N_2669);
xnor U5316 (N_5316,N_975,N_3766);
xnor U5317 (N_5317,N_590,N_4344);
or U5318 (N_5318,N_4490,N_3258);
nor U5319 (N_5319,N_1727,N_4593);
xor U5320 (N_5320,N_1288,N_942);
nor U5321 (N_5321,N_3198,N_680);
xnor U5322 (N_5322,N_3,N_2094);
xnor U5323 (N_5323,N_3154,N_4518);
xnor U5324 (N_5324,N_1640,N_3538);
and U5325 (N_5325,N_4970,N_734);
or U5326 (N_5326,N_150,N_2856);
nand U5327 (N_5327,N_4625,N_258);
xnor U5328 (N_5328,N_3709,N_1276);
nor U5329 (N_5329,N_2391,N_3670);
nand U5330 (N_5330,N_4034,N_3795);
nor U5331 (N_5331,N_1477,N_2119);
or U5332 (N_5332,N_2231,N_1819);
and U5333 (N_5333,N_4161,N_2701);
xor U5334 (N_5334,N_1635,N_1856);
nor U5335 (N_5335,N_101,N_2546);
or U5336 (N_5336,N_3703,N_200);
and U5337 (N_5337,N_2987,N_993);
nand U5338 (N_5338,N_1247,N_414);
and U5339 (N_5339,N_1053,N_4802);
nand U5340 (N_5340,N_808,N_44);
nor U5341 (N_5341,N_3904,N_4249);
and U5342 (N_5342,N_4526,N_3616);
xnor U5343 (N_5343,N_1561,N_1801);
xor U5344 (N_5344,N_550,N_303);
and U5345 (N_5345,N_4914,N_1873);
or U5346 (N_5346,N_83,N_1537);
xor U5347 (N_5347,N_3478,N_1625);
nand U5348 (N_5348,N_4417,N_2420);
nand U5349 (N_5349,N_3653,N_382);
nor U5350 (N_5350,N_4839,N_2465);
and U5351 (N_5351,N_953,N_3652);
nor U5352 (N_5352,N_686,N_3720);
xnor U5353 (N_5353,N_1036,N_802);
nor U5354 (N_5354,N_18,N_4089);
nor U5355 (N_5355,N_1374,N_536);
nand U5356 (N_5356,N_1756,N_745);
and U5357 (N_5357,N_1719,N_1667);
xnor U5358 (N_5358,N_3054,N_286);
or U5359 (N_5359,N_3067,N_588);
nand U5360 (N_5360,N_3883,N_1458);
or U5361 (N_5361,N_4023,N_4623);
or U5362 (N_5362,N_4199,N_1498);
nand U5363 (N_5363,N_3606,N_4884);
xnor U5364 (N_5364,N_2691,N_1007);
or U5365 (N_5365,N_3191,N_3939);
or U5366 (N_5366,N_1398,N_1355);
and U5367 (N_5367,N_4219,N_3033);
and U5368 (N_5368,N_204,N_1111);
nor U5369 (N_5369,N_1645,N_2425);
and U5370 (N_5370,N_2581,N_694);
or U5371 (N_5371,N_185,N_501);
or U5372 (N_5372,N_1353,N_1877);
and U5373 (N_5373,N_3026,N_127);
and U5374 (N_5374,N_1878,N_4786);
or U5375 (N_5375,N_2540,N_1597);
or U5376 (N_5376,N_2102,N_3363);
nor U5377 (N_5377,N_4296,N_3177);
or U5378 (N_5378,N_2787,N_2081);
xor U5379 (N_5379,N_2960,N_4459);
xnor U5380 (N_5380,N_4156,N_1790);
nand U5381 (N_5381,N_4866,N_2156);
nand U5382 (N_5382,N_4252,N_1294);
nand U5383 (N_5383,N_3955,N_1861);
nor U5384 (N_5384,N_2490,N_4570);
nor U5385 (N_5385,N_3282,N_4354);
nor U5386 (N_5386,N_4511,N_2250);
or U5387 (N_5387,N_3242,N_1348);
nand U5388 (N_5388,N_4233,N_2637);
nor U5389 (N_5389,N_3671,N_614);
and U5390 (N_5390,N_3000,N_4844);
or U5391 (N_5391,N_2349,N_959);
xnor U5392 (N_5392,N_1760,N_2718);
xor U5393 (N_5393,N_2525,N_2511);
or U5394 (N_5394,N_1071,N_4361);
nand U5395 (N_5395,N_3830,N_4744);
or U5396 (N_5396,N_2303,N_1862);
nor U5397 (N_5397,N_3047,N_2282);
xor U5398 (N_5398,N_3966,N_2379);
nor U5399 (N_5399,N_1728,N_2783);
and U5400 (N_5400,N_3983,N_377);
or U5401 (N_5401,N_752,N_4917);
nor U5402 (N_5402,N_648,N_4770);
or U5403 (N_5403,N_3311,N_3761);
nand U5404 (N_5404,N_3950,N_2321);
nand U5405 (N_5405,N_3718,N_3914);
and U5406 (N_5406,N_1757,N_3953);
xor U5407 (N_5407,N_3988,N_421);
or U5408 (N_5408,N_1114,N_4179);
nand U5409 (N_5409,N_1464,N_2758);
xnor U5410 (N_5410,N_2471,N_4146);
and U5411 (N_5411,N_4738,N_524);
and U5412 (N_5412,N_1747,N_2716);
and U5413 (N_5413,N_3488,N_3278);
and U5414 (N_5414,N_1978,N_1944);
and U5415 (N_5415,N_4198,N_2108);
nand U5416 (N_5416,N_4238,N_4154);
nand U5417 (N_5417,N_1858,N_894);
nor U5418 (N_5418,N_4435,N_2981);
nor U5419 (N_5419,N_3361,N_1372);
or U5420 (N_5420,N_4629,N_4454);
or U5421 (N_5421,N_2890,N_1324);
xnor U5422 (N_5422,N_388,N_4358);
nor U5423 (N_5423,N_1712,N_1075);
nor U5424 (N_5424,N_3289,N_1829);
or U5425 (N_5425,N_383,N_2534);
nand U5426 (N_5426,N_1562,N_1680);
nor U5427 (N_5427,N_357,N_425);
or U5428 (N_5428,N_2409,N_2936);
and U5429 (N_5429,N_2693,N_3350);
nor U5430 (N_5430,N_4185,N_271);
and U5431 (N_5431,N_2252,N_3837);
nor U5432 (N_5432,N_350,N_4763);
xnor U5433 (N_5433,N_1388,N_4279);
and U5434 (N_5434,N_4697,N_2615);
and U5435 (N_5435,N_1490,N_4988);
xnor U5436 (N_5436,N_48,N_2470);
xor U5437 (N_5437,N_3063,N_3615);
and U5438 (N_5438,N_3573,N_3708);
or U5439 (N_5439,N_1553,N_3188);
nand U5440 (N_5440,N_4220,N_2583);
xnor U5441 (N_5441,N_1511,N_3853);
or U5442 (N_5442,N_1972,N_2748);
xor U5443 (N_5443,N_1688,N_3004);
nand U5444 (N_5444,N_2510,N_941);
or U5445 (N_5445,N_21,N_4663);
nand U5446 (N_5446,N_4227,N_2891);
xnor U5447 (N_5447,N_4631,N_669);
nand U5448 (N_5448,N_664,N_2907);
nand U5449 (N_5449,N_364,N_2661);
nor U5450 (N_5450,N_4677,N_4687);
and U5451 (N_5451,N_1315,N_63);
nand U5452 (N_5452,N_2451,N_4612);
xnor U5453 (N_5453,N_472,N_4656);
and U5454 (N_5454,N_175,N_4169);
and U5455 (N_5455,N_2082,N_1940);
xor U5456 (N_5456,N_4695,N_4710);
nand U5457 (N_5457,N_906,N_1955);
nor U5458 (N_5458,N_1826,N_3107);
or U5459 (N_5459,N_861,N_3392);
nor U5460 (N_5460,N_3912,N_1274);
xnor U5461 (N_5461,N_2507,N_4648);
xnor U5462 (N_5462,N_229,N_914);
xnor U5463 (N_5463,N_2629,N_2369);
xor U5464 (N_5464,N_3946,N_544);
nand U5465 (N_5465,N_3619,N_4264);
or U5466 (N_5466,N_2595,N_4458);
or U5467 (N_5467,N_1238,N_4756);
xor U5468 (N_5468,N_621,N_3413);
nor U5469 (N_5469,N_1154,N_635);
or U5470 (N_5470,N_1200,N_867);
nand U5471 (N_5471,N_3116,N_2219);
and U5472 (N_5472,N_2841,N_629);
nor U5473 (N_5473,N_2774,N_3880);
or U5474 (N_5474,N_3396,N_3379);
nand U5475 (N_5475,N_2046,N_2577);
nor U5476 (N_5476,N_3737,N_3018);
nor U5477 (N_5477,N_108,N_2756);
and U5478 (N_5478,N_2277,N_3434);
and U5479 (N_5479,N_3860,N_902);
xnor U5480 (N_5480,N_657,N_2441);
nor U5481 (N_5481,N_1314,N_3385);
nand U5482 (N_5482,N_1334,N_1617);
xnor U5483 (N_5483,N_4465,N_3557);
xor U5484 (N_5484,N_4742,N_4024);
or U5485 (N_5485,N_4685,N_800);
nor U5486 (N_5486,N_1085,N_1987);
xnor U5487 (N_5487,N_475,N_172);
xor U5488 (N_5488,N_2896,N_2217);
nand U5489 (N_5489,N_2836,N_1736);
nand U5490 (N_5490,N_78,N_2295);
xnor U5491 (N_5491,N_1117,N_967);
xnor U5492 (N_5492,N_1959,N_786);
or U5493 (N_5493,N_4251,N_1532);
and U5494 (N_5494,N_1067,N_2260);
nor U5495 (N_5495,N_34,N_4012);
nor U5496 (N_5496,N_3484,N_3338);
and U5497 (N_5497,N_4525,N_1073);
or U5498 (N_5498,N_1179,N_4290);
or U5499 (N_5499,N_4611,N_3773);
and U5500 (N_5500,N_426,N_2246);
and U5501 (N_5501,N_765,N_1042);
xnor U5502 (N_5502,N_2909,N_4136);
xnor U5503 (N_5503,N_3643,N_2906);
and U5504 (N_5504,N_3108,N_1241);
and U5505 (N_5505,N_587,N_340);
nor U5506 (N_5506,N_4008,N_3050);
and U5507 (N_5507,N_1824,N_4446);
nand U5508 (N_5508,N_3135,N_718);
nor U5509 (N_5509,N_4421,N_3065);
nand U5510 (N_5510,N_2528,N_1630);
and U5511 (N_5511,N_4891,N_4661);
nor U5512 (N_5512,N_2114,N_1841);
or U5513 (N_5513,N_2405,N_516);
or U5514 (N_5514,N_2664,N_1707);
xnor U5515 (N_5515,N_3100,N_3585);
and U5516 (N_5516,N_46,N_3407);
nor U5517 (N_5517,N_2368,N_4659);
and U5518 (N_5518,N_2273,N_1738);
nor U5519 (N_5519,N_1663,N_3502);
xor U5520 (N_5520,N_434,N_2789);
and U5521 (N_5521,N_4666,N_3728);
and U5522 (N_5522,N_3226,N_979);
nand U5523 (N_5523,N_2308,N_2016);
nand U5524 (N_5524,N_3603,N_3997);
and U5525 (N_5525,N_113,N_4157);
nor U5526 (N_5526,N_1415,N_4618);
or U5527 (N_5527,N_1817,N_4478);
nor U5528 (N_5528,N_4747,N_1668);
and U5529 (N_5529,N_2878,N_484);
nor U5530 (N_5530,N_1120,N_4466);
nand U5531 (N_5531,N_26,N_4176);
xnor U5532 (N_5532,N_1506,N_1297);
and U5533 (N_5533,N_1788,N_1813);
nor U5534 (N_5534,N_4474,N_1407);
or U5535 (N_5535,N_3518,N_4981);
nand U5536 (N_5536,N_3094,N_3241);
and U5537 (N_5537,N_1422,N_2346);
and U5538 (N_5538,N_3057,N_3496);
or U5539 (N_5539,N_3142,N_3444);
nand U5540 (N_5540,N_1931,N_814);
nor U5541 (N_5541,N_2711,N_1669);
and U5542 (N_5542,N_1366,N_1921);
nor U5543 (N_5543,N_567,N_920);
and U5544 (N_5544,N_650,N_1142);
nand U5545 (N_5545,N_4578,N_4484);
or U5546 (N_5546,N_109,N_2875);
or U5547 (N_5547,N_427,N_3500);
and U5548 (N_5548,N_3317,N_542);
xor U5549 (N_5549,N_183,N_1195);
and U5550 (N_5550,N_2551,N_875);
nor U5551 (N_5551,N_2543,N_3805);
nor U5552 (N_5552,N_850,N_888);
nor U5553 (N_5553,N_1108,N_1761);
nor U5554 (N_5554,N_2797,N_3717);
xor U5555 (N_5555,N_4750,N_4671);
nor U5556 (N_5556,N_4371,N_2710);
and U5557 (N_5557,N_675,N_3725);
nor U5558 (N_5558,N_1410,N_792);
and U5559 (N_5559,N_2199,N_3910);
xor U5560 (N_5560,N_1322,N_659);
nand U5561 (N_5561,N_224,N_307);
and U5562 (N_5562,N_4614,N_2982);
and U5563 (N_5563,N_249,N_4235);
and U5564 (N_5564,N_3451,N_2648);
nand U5565 (N_5565,N_436,N_2220);
xnor U5566 (N_5566,N_2776,N_4376);
nor U5567 (N_5567,N_2862,N_4536);
nor U5568 (N_5568,N_2175,N_4422);
nand U5569 (N_5569,N_1780,N_1417);
or U5570 (N_5570,N_3421,N_3775);
nor U5571 (N_5571,N_4548,N_3913);
or U5572 (N_5572,N_4431,N_3730);
and U5573 (N_5573,N_159,N_2329);
nand U5574 (N_5574,N_1876,N_4186);
or U5575 (N_5575,N_457,N_3695);
or U5576 (N_5576,N_3624,N_3890);
and U5577 (N_5577,N_830,N_1402);
nor U5578 (N_5578,N_1157,N_1319);
xnor U5579 (N_5579,N_4082,N_190);
xor U5580 (N_5580,N_2653,N_3617);
xnor U5581 (N_5581,N_1503,N_302);
and U5582 (N_5582,N_772,N_514);
xor U5583 (N_5583,N_4476,N_2443);
nand U5584 (N_5584,N_2976,N_2178);
nor U5585 (N_5585,N_1981,N_4995);
nor U5586 (N_5586,N_4921,N_3263);
nor U5587 (N_5587,N_3141,N_4904);
nand U5588 (N_5588,N_1389,N_4134);
and U5589 (N_5589,N_1681,N_3465);
xor U5590 (N_5590,N_881,N_3227);
xor U5591 (N_5591,N_4002,N_2644);
and U5592 (N_5592,N_3757,N_2620);
xnor U5593 (N_5593,N_2306,N_2638);
or U5594 (N_5594,N_3260,N_1560);
or U5595 (N_5595,N_3733,N_1397);
or U5596 (N_5596,N_936,N_4834);
or U5597 (N_5597,N_160,N_176);
nor U5598 (N_5598,N_2421,N_1889);
xor U5599 (N_5599,N_2335,N_3824);
xnor U5600 (N_5600,N_4330,N_4272);
or U5601 (N_5601,N_1576,N_3254);
nor U5602 (N_5602,N_3920,N_744);
nand U5603 (N_5603,N_3214,N_1345);
xnor U5604 (N_5604,N_1748,N_981);
nand U5605 (N_5605,N_4755,N_337);
nor U5606 (N_5606,N_2782,N_2384);
and U5607 (N_5607,N_905,N_3848);
or U5608 (N_5608,N_456,N_822);
xnor U5609 (N_5609,N_3210,N_2522);
nand U5610 (N_5610,N_917,N_3314);
nor U5611 (N_5611,N_4605,N_3694);
and U5612 (N_5612,N_67,N_3503);
or U5613 (N_5613,N_289,N_876);
xor U5614 (N_5614,N_994,N_1948);
or U5615 (N_5615,N_3240,N_964);
or U5616 (N_5616,N_2006,N_9);
xor U5617 (N_5617,N_1615,N_3003);
nor U5618 (N_5618,N_1173,N_3497);
or U5619 (N_5619,N_1912,N_3614);
nor U5620 (N_5620,N_1375,N_2239);
and U5621 (N_5621,N_1504,N_3931);
xnor U5622 (N_5622,N_3280,N_1337);
nand U5623 (N_5623,N_3499,N_1468);
nor U5624 (N_5624,N_1868,N_4523);
or U5625 (N_5625,N_593,N_2412);
nor U5626 (N_5626,N_4615,N_3916);
or U5627 (N_5627,N_504,N_1033);
nand U5628 (N_5628,N_856,N_1497);
nand U5629 (N_5629,N_4063,N_4876);
and U5630 (N_5630,N_4311,N_1009);
nor U5631 (N_5631,N_701,N_3870);
and U5632 (N_5632,N_1880,N_1385);
nor U5633 (N_5633,N_230,N_2212);
nand U5634 (N_5634,N_2442,N_2194);
xnor U5635 (N_5635,N_2537,N_2518);
nand U5636 (N_5636,N_49,N_3963);
xor U5637 (N_5637,N_753,N_2673);
or U5638 (N_5638,N_3877,N_4741);
nand U5639 (N_5639,N_3967,N_2925);
or U5640 (N_5640,N_1942,N_2506);
xnor U5641 (N_5641,N_857,N_2449);
nor U5642 (N_5642,N_3323,N_4727);
xor U5643 (N_5643,N_3233,N_1229);
and U5644 (N_5644,N_4040,N_1469);
and U5645 (N_5645,N_1356,N_995);
xnor U5646 (N_5646,N_4630,N_4966);
nor U5647 (N_5647,N_3810,N_2988);
xor U5648 (N_5648,N_810,N_1545);
xor U5649 (N_5649,N_165,N_1359);
or U5650 (N_5650,N_1686,N_1515);
nor U5651 (N_5651,N_4875,N_4669);
nand U5652 (N_5652,N_509,N_2739);
xor U5653 (N_5653,N_496,N_3044);
and U5654 (N_5654,N_312,N_4401);
nor U5655 (N_5655,N_2196,N_592);
nand U5656 (N_5656,N_612,N_564);
xor U5657 (N_5657,N_277,N_978);
and U5658 (N_5658,N_4651,N_2704);
xnor U5659 (N_5659,N_798,N_460);
nand U5660 (N_5660,N_3899,N_4248);
nor U5661 (N_5661,N_459,N_2851);
xor U5662 (N_5662,N_3661,N_4698);
and U5663 (N_5663,N_666,N_4682);
xnor U5664 (N_5664,N_2937,N_3312);
nand U5665 (N_5665,N_2164,N_2330);
nor U5666 (N_5666,N_739,N_2818);
or U5667 (N_5667,N_3705,N_2848);
nand U5668 (N_5668,N_2955,N_3199);
xnor U5669 (N_5669,N_1723,N_3683);
nor U5670 (N_5670,N_4976,N_4653);
nand U5671 (N_5671,N_296,N_2424);
nor U5672 (N_5672,N_1041,N_2358);
nor U5673 (N_5673,N_3442,N_1239);
xnor U5674 (N_5674,N_3722,N_946);
and U5675 (N_5675,N_2863,N_189);
and U5676 (N_5676,N_191,N_1079);
nand U5677 (N_5677,N_4026,N_3461);
or U5678 (N_5678,N_3172,N_1189);
and U5679 (N_5679,N_4948,N_1846);
nand U5680 (N_5680,N_239,N_1898);
nor U5681 (N_5681,N_998,N_1284);
and U5682 (N_5682,N_1892,N_2975);
and U5683 (N_5683,N_4144,N_3387);
xor U5684 (N_5684,N_2961,N_4688);
xnor U5685 (N_5685,N_2751,N_1834);
nor U5686 (N_5686,N_3230,N_2759);
xor U5687 (N_5687,N_991,N_1566);
and U5688 (N_5688,N_2843,N_2345);
nand U5689 (N_5689,N_2800,N_549);
nor U5690 (N_5690,N_3994,N_4020);
or U5691 (N_5691,N_2554,N_4564);
and U5692 (N_5692,N_4353,N_637);
or U5693 (N_5693,N_2024,N_1370);
nor U5694 (N_5694,N_3527,N_885);
xnor U5695 (N_5695,N_661,N_803);
nor U5696 (N_5696,N_4568,N_134);
and U5697 (N_5697,N_3180,N_787);
or U5698 (N_5698,N_3092,N_3678);
nand U5699 (N_5699,N_2560,N_523);
xnor U5700 (N_5700,N_36,N_4289);
nor U5701 (N_5701,N_1687,N_645);
and U5702 (N_5702,N_1820,N_789);
nor U5703 (N_5703,N_1273,N_1500);
and U5704 (N_5704,N_247,N_2900);
nor U5705 (N_5705,N_4334,N_2187);
nand U5706 (N_5706,N_145,N_3513);
nand U5707 (N_5707,N_1791,N_3845);
or U5708 (N_5708,N_4563,N_2304);
nor U5709 (N_5709,N_2366,N_3928);
nand U5710 (N_5710,N_3459,N_1509);
xor U5711 (N_5711,N_154,N_3774);
nand U5712 (N_5712,N_3647,N_2163);
xor U5713 (N_5713,N_1850,N_171);
or U5714 (N_5714,N_2754,N_2908);
nand U5715 (N_5715,N_2055,N_3416);
and U5716 (N_5716,N_2285,N_94);
and U5717 (N_5717,N_4127,N_4028);
nor U5718 (N_5718,N_3367,N_740);
and U5719 (N_5719,N_1002,N_3555);
and U5720 (N_5720,N_1296,N_2567);
xnor U5721 (N_5721,N_3238,N_1089);
nand U5722 (N_5722,N_1088,N_2823);
nor U5723 (N_5723,N_2170,N_31);
and U5724 (N_5724,N_3901,N_892);
or U5725 (N_5725,N_4881,N_2487);
nor U5726 (N_5726,N_2136,N_4734);
or U5727 (N_5727,N_429,N_2240);
or U5728 (N_5728,N_780,N_461);
xnor U5729 (N_5729,N_1447,N_996);
nor U5730 (N_5730,N_1320,N_4462);
xnor U5731 (N_5731,N_3211,N_4717);
nand U5732 (N_5732,N_543,N_2307);
xnor U5733 (N_5733,N_2858,N_817);
nor U5734 (N_5734,N_3059,N_1106);
or U5735 (N_5735,N_922,N_4880);
xnor U5736 (N_5736,N_181,N_2749);
nand U5737 (N_5737,N_4168,N_652);
xor U5738 (N_5738,N_2418,N_507);
and U5739 (N_5739,N_385,N_816);
nor U5740 (N_5740,N_2184,N_3034);
nor U5741 (N_5741,N_2901,N_3014);
and U5742 (N_5742,N_1405,N_4853);
or U5743 (N_5743,N_1499,N_2724);
xor U5744 (N_5744,N_4236,N_215);
nor U5745 (N_5745,N_1413,N_131);
nor U5746 (N_5746,N_2572,N_580);
or U5747 (N_5747,N_4114,N_1161);
or U5748 (N_5748,N_2017,N_1607);
nand U5749 (N_5749,N_3574,N_144);
nor U5750 (N_5750,N_3911,N_2027);
and U5751 (N_5751,N_1199,N_4911);
nand U5752 (N_5752,N_2684,N_1648);
and U5753 (N_5753,N_761,N_141);
nand U5754 (N_5754,N_3476,N_1832);
or U5755 (N_5755,N_3173,N_3511);
or U5756 (N_5756,N_3159,N_3128);
or U5757 (N_5757,N_3864,N_4230);
and U5758 (N_5758,N_3464,N_778);
or U5759 (N_5759,N_1091,N_4626);
nand U5760 (N_5760,N_2167,N_4908);
nand U5761 (N_5761,N_3945,N_598);
or U5762 (N_5762,N_3828,N_4373);
xor U5763 (N_5763,N_882,N_923);
xnor U5764 (N_5764,N_3854,N_2779);
nand U5765 (N_5765,N_4445,N_3395);
and U5766 (N_5766,N_4314,N_3618);
nor U5767 (N_5767,N_2688,N_1804);
or U5768 (N_5768,N_2312,N_2645);
nor U5769 (N_5769,N_3267,N_4799);
and U5770 (N_5770,N_179,N_4142);
xor U5771 (N_5771,N_877,N_1512);
or U5772 (N_5772,N_1336,N_2762);
or U5773 (N_5773,N_4573,N_226);
or U5774 (N_5774,N_2945,N_4443);
nand U5775 (N_5775,N_790,N_508);
nor U5776 (N_5776,N_4318,N_2757);
xor U5777 (N_5777,N_262,N_4302);
xnor U5778 (N_5778,N_479,N_4419);
xor U5779 (N_5779,N_3972,N_2244);
nor U5780 (N_5780,N_2249,N_4620);
and U5781 (N_5781,N_2717,N_3941);
and U5782 (N_5782,N_768,N_2213);
nor U5783 (N_5783,N_2147,N_1941);
xor U5784 (N_5784,N_962,N_4216);
nand U5785 (N_5785,N_2207,N_1129);
nand U5786 (N_5786,N_4170,N_847);
nor U5787 (N_5787,N_1478,N_1439);
nor U5788 (N_5788,N_1655,N_4110);
xor U5789 (N_5789,N_1292,N_4740);
or U5790 (N_5790,N_974,N_903);
and U5791 (N_5791,N_4450,N_2073);
nand U5792 (N_5792,N_1731,N_112);
xor U5793 (N_5793,N_4363,N_4978);
xor U5794 (N_5794,N_1310,N_596);
or U5795 (N_5795,N_2715,N_2491);
or U5796 (N_5796,N_2512,N_3355);
nand U5797 (N_5797,N_3452,N_2576);
or U5798 (N_5798,N_3084,N_4393);
and U5799 (N_5799,N_186,N_820);
nor U5800 (N_5800,N_2662,N_2302);
or U5801 (N_5801,N_3365,N_3898);
xnor U5802 (N_5802,N_2803,N_4694);
and U5803 (N_5803,N_4297,N_2829);
or U5804 (N_5804,N_4480,N_2447);
or U5805 (N_5805,N_4494,N_4257);
nand U5806 (N_5806,N_4920,N_1222);
nor U5807 (N_5807,N_4108,N_519);
nand U5808 (N_5808,N_3635,N_1390);
and U5809 (N_5809,N_2270,N_1734);
and U5810 (N_5810,N_3935,N_3404);
and U5811 (N_5811,N_2564,N_2509);
nand U5812 (N_5812,N_4725,N_1613);
xor U5813 (N_5813,N_1101,N_4991);
nor U5814 (N_5814,N_3759,N_281);
or U5815 (N_5815,N_1105,N_4922);
or U5816 (N_5816,N_1963,N_2018);
xnor U5817 (N_5817,N_4832,N_4107);
nor U5818 (N_5818,N_4714,N_4223);
or U5819 (N_5819,N_2838,N_1947);
and U5820 (N_5820,N_345,N_317);
nor U5821 (N_5821,N_2611,N_3366);
and U5822 (N_5822,N_1019,N_4060);
and U5823 (N_5823,N_1165,N_129);
or U5824 (N_5824,N_3244,N_2857);
xnor U5825 (N_5825,N_699,N_1235);
and U5826 (N_5826,N_1391,N_4339);
or U5827 (N_5827,N_4737,N_783);
nor U5828 (N_5828,N_4105,N_2430);
nor U5829 (N_5829,N_1694,N_3480);
or U5830 (N_5830,N_1765,N_2709);
or U5831 (N_5831,N_2459,N_2895);
nor U5832 (N_5832,N_3391,N_2341);
and U5833 (N_5833,N_2627,N_1132);
xnor U5834 (N_5834,N_3253,N_3711);
or U5835 (N_5835,N_732,N_678);
or U5836 (N_5836,N_4122,N_2269);
nor U5837 (N_5837,N_1031,N_3610);
nor U5838 (N_5838,N_1493,N_1641);
nor U5839 (N_5839,N_3702,N_644);
nor U5840 (N_5840,N_985,N_4174);
nand U5841 (N_5841,N_2182,N_1496);
xor U5842 (N_5842,N_403,N_2842);
or U5843 (N_5843,N_4287,N_91);
nor U5844 (N_5844,N_4850,N_4601);
and U5845 (N_5845,N_1128,N_4680);
xor U5846 (N_5846,N_3505,N_1768);
xor U5847 (N_5847,N_325,N_1119);
nand U5848 (N_5848,N_2493,N_2647);
or U5849 (N_5849,N_759,N_169);
nor U5850 (N_5850,N_3787,N_93);
and U5851 (N_5851,N_2174,N_2917);
and U5852 (N_5852,N_2394,N_2297);
and U5853 (N_5853,N_4992,N_1440);
nand U5854 (N_5854,N_931,N_3551);
nor U5855 (N_5855,N_3072,N_1895);
nand U5856 (N_5856,N_2530,N_2056);
xor U5857 (N_5857,N_3023,N_1443);
nand U5858 (N_5858,N_3794,N_846);
nor U5859 (N_5859,N_2245,N_3992);
nand U5860 (N_5860,N_2997,N_3097);
xnor U5861 (N_5861,N_3878,N_2744);
xor U5862 (N_5862,N_1933,N_310);
nor U5863 (N_5863,N_323,N_819);
xnor U5864 (N_5864,N_662,N_3559);
or U5865 (N_5865,N_2965,N_738);
nor U5866 (N_5866,N_4411,N_4109);
nand U5867 (N_5867,N_2294,N_2160);
xor U5868 (N_5868,N_1080,N_4365);
xnor U5869 (N_5869,N_4551,N_3176);
nand U5870 (N_5870,N_1046,N_73);
xnor U5871 (N_5871,N_4292,N_4085);
nor U5872 (N_5872,N_1582,N_4263);
and U5873 (N_5873,N_4164,N_3036);
or U5874 (N_5874,N_4218,N_2650);
xor U5875 (N_5875,N_3822,N_3727);
xor U5876 (N_5876,N_2318,N_153);
and U5877 (N_5877,N_890,N_1543);
nor U5878 (N_5878,N_3823,N_2678);
or U5879 (N_5879,N_2681,N_4509);
and U5880 (N_5880,N_1755,N_4364);
nand U5881 (N_5881,N_2872,N_2259);
and U5882 (N_5882,N_2419,N_395);
nor U5883 (N_5883,N_3548,N_3827);
or U5884 (N_5884,N_4382,N_2031);
and U5885 (N_5885,N_1382,N_3275);
xor U5886 (N_5886,N_4196,N_1996);
nor U5887 (N_5887,N_2482,N_1722);
xnor U5888 (N_5888,N_2773,N_4394);
nand U5889 (N_5889,N_4958,N_3600);
nand U5890 (N_5890,N_2873,N_4942);
and U5891 (N_5891,N_3909,N_4097);
and U5892 (N_5892,N_3506,N_4413);
and U5893 (N_5893,N_4213,N_3881);
nand U5894 (N_5894,N_4087,N_1068);
xor U5895 (N_5895,N_1609,N_1932);
or U5896 (N_5896,N_152,N_1016);
nand U5897 (N_5897,N_3457,N_1168);
xnor U5898 (N_5898,N_2847,N_940);
xnor U5899 (N_5899,N_4472,N_3369);
nand U5900 (N_5900,N_2532,N_2352);
nand U5901 (N_5901,N_3027,N_3571);
xor U5902 (N_5902,N_1298,N_796);
and U5903 (N_5903,N_855,N_2049);
and U5904 (N_5904,N_265,N_3639);
and U5905 (N_5905,N_4293,N_4469);
nor U5906 (N_5906,N_3106,N_1171);
or U5907 (N_5907,N_2161,N_4860);
and U5908 (N_5908,N_4455,N_710);
or U5909 (N_5909,N_442,N_3146);
nor U5910 (N_5910,N_1442,N_2395);
nor U5911 (N_5911,N_1185,N_604);
nor U5912 (N_5912,N_122,N_1784);
or U5913 (N_5913,N_4129,N_1701);
nor U5914 (N_5914,N_628,N_3693);
and U5915 (N_5915,N_2989,N_705);
xor U5916 (N_5916,N_4820,N_4075);
xnor U5917 (N_5917,N_4873,N_1266);
nor U5918 (N_5918,N_997,N_1689);
nor U5919 (N_5919,N_2154,N_3460);
xnor U5920 (N_5920,N_140,N_4406);
nand U5921 (N_5921,N_4760,N_1893);
or U5922 (N_5922,N_3778,N_653);
or U5923 (N_5923,N_1204,N_3301);
xor U5924 (N_5924,N_3262,N_250);
and U5925 (N_5925,N_2667,N_2846);
xnor U5926 (N_5926,N_439,N_681);
or U5927 (N_5927,N_2879,N_1594);
or U5928 (N_5928,N_1242,N_771);
or U5929 (N_5929,N_2104,N_880);
xor U5930 (N_5930,N_2569,N_3987);
nor U5931 (N_5931,N_4647,N_2361);
nand U5932 (N_5932,N_853,N_4438);
and U5933 (N_5933,N_4115,N_2033);
or U5934 (N_5934,N_3284,N_3688);
xor U5935 (N_5935,N_1865,N_1614);
and U5936 (N_5936,N_2864,N_4402);
or U5937 (N_5937,N_2191,N_2224);
xor U5938 (N_5938,N_3685,N_4284);
or U5939 (N_5939,N_2433,N_2602);
nand U5940 (N_5940,N_3102,N_4691);
nor U5941 (N_5941,N_2649,N_597);
or U5942 (N_5942,N_2401,N_749);
or U5943 (N_5943,N_1485,N_831);
xnor U5944 (N_5944,N_1212,N_4046);
or U5945 (N_5945,N_1573,N_3197);
nor U5946 (N_5946,N_2271,N_3820);
and U5947 (N_5947,N_1622,N_1683);
nor U5948 (N_5948,N_4907,N_1177);
nor U5949 (N_5949,N_4208,N_3649);
and U5950 (N_5950,N_3482,N_4798);
or U5951 (N_5951,N_2772,N_2780);
xor U5952 (N_5952,N_1121,N_1432);
nand U5953 (N_5953,N_1773,N_1051);
nor U5954 (N_5954,N_2792,N_3789);
or U5955 (N_5955,N_1233,N_2978);
xor U5956 (N_5956,N_2039,N_1584);
or U5957 (N_5957,N_3892,N_3940);
nor U5958 (N_5958,N_1426,N_3223);
xnor U5959 (N_5959,N_10,N_4057);
or U5960 (N_5960,N_2402,N_2437);
nor U5961 (N_5961,N_3111,N_916);
and U5962 (N_5962,N_943,N_4926);
nor U5963 (N_5963,N_3577,N_971);
and U5964 (N_5964,N_1642,N_1644);
or U5965 (N_5965,N_4900,N_2299);
and U5966 (N_5966,N_42,N_1675);
nand U5967 (N_5967,N_4111,N_3597);
nor U5968 (N_5968,N_441,N_418);
nor U5969 (N_5969,N_3856,N_2298);
and U5970 (N_5970,N_180,N_90);
or U5971 (N_5971,N_4519,N_3654);
or U5972 (N_5972,N_480,N_3216);
nor U5973 (N_5973,N_294,N_1992);
nor U5974 (N_5974,N_1267,N_667);
nand U5975 (N_5975,N_2396,N_1540);
and U5976 (N_5976,N_2954,N_3121);
nand U5977 (N_5977,N_2682,N_3228);
nand U5978 (N_5978,N_2397,N_2284);
nand U5979 (N_5979,N_4539,N_3960);
and U5980 (N_5980,N_522,N_2432);
or U5981 (N_5981,N_3792,N_2188);
or U5982 (N_5982,N_4893,N_65);
or U5983 (N_5983,N_76,N_2089);
nand U5984 (N_5984,N_3676,N_206);
nor U5985 (N_5985,N_1557,N_1807);
nand U5986 (N_5986,N_2573,N_368);
or U5987 (N_5987,N_4201,N_1221);
or U5988 (N_5988,N_1281,N_1618);
or U5989 (N_5989,N_2825,N_4897);
nand U5990 (N_5990,N_3692,N_4849);
or U5991 (N_5991,N_2038,N_2698);
nand U5992 (N_5992,N_3637,N_1006);
xnor U5993 (N_5993,N_453,N_3252);
nand U5994 (N_5994,N_7,N_4855);
or U5995 (N_5995,N_3433,N_3583);
or U5996 (N_5996,N_3006,N_2686);
and U5997 (N_5997,N_2995,N_2557);
or U5998 (N_5998,N_4183,N_4400);
nor U5999 (N_5999,N_2458,N_4652);
xor U6000 (N_6000,N_2778,N_555);
nor U6001 (N_6001,N_3089,N_3780);
nor U6002 (N_6002,N_3347,N_3578);
xor U6003 (N_6003,N_2556,N_342);
nand U6004 (N_6004,N_4800,N_4368);
or U6005 (N_6005,N_297,N_1685);
xor U6006 (N_6006,N_1412,N_2025);
and U6007 (N_6007,N_4890,N_2727);
and U6008 (N_6008,N_4018,N_3704);
nand U6009 (N_6009,N_3243,N_4439);
and U6010 (N_6010,N_1751,N_256);
and U6011 (N_6011,N_305,N_2286);
nand U6012 (N_6012,N_2584,N_3436);
or U6013 (N_6013,N_2835,N_228);
or U6014 (N_6014,N_1095,N_4668);
and U6015 (N_6015,N_2000,N_2932);
nor U6016 (N_6016,N_649,N_4412);
or U6017 (N_6017,N_1226,N_2130);
or U6018 (N_6018,N_4496,N_616);
nand U6019 (N_6019,N_4180,N_4342);
nand U6020 (N_6020,N_900,N_105);
nor U6021 (N_6021,N_272,N_1344);
nand U6022 (N_6022,N_3078,N_3508);
and U6023 (N_6023,N_568,N_3028);
and U6024 (N_6024,N_2536,N_1999);
or U6025 (N_6025,N_3625,N_3813);
or U6026 (N_6026,N_2300,N_915);
nand U6027 (N_6027,N_3234,N_3677);
and U6028 (N_6028,N_3753,N_3891);
or U6029 (N_6029,N_1339,N_4946);
or U6030 (N_6030,N_1803,N_4718);
and U6031 (N_6031,N_957,N_1770);
xor U6032 (N_6032,N_2035,N_4867);
nor U6033 (N_6033,N_4543,N_2374);
and U6034 (N_6034,N_4133,N_4544);
nor U6035 (N_6035,N_707,N_1352);
nand U6036 (N_6036,N_3686,N_3118);
or U6037 (N_6037,N_3112,N_399);
xnor U6038 (N_6038,N_3349,N_1331);
nand U6039 (N_6039,N_1517,N_3104);
or U6040 (N_6040,N_483,N_4690);
nand U6041 (N_6041,N_3535,N_4848);
nor U6042 (N_6042,N_4487,N_2192);
nor U6043 (N_6043,N_3971,N_1816);
nand U6044 (N_6044,N_2406,N_4546);
xor U6045 (N_6045,N_2206,N_102);
or U6046 (N_6046,N_4767,N_2942);
and U6047 (N_6047,N_1979,N_2690);
xnor U6048 (N_6048,N_3786,N_3874);
nor U6049 (N_6049,N_1365,N_3415);
and U6050 (N_6050,N_2582,N_3271);
or U6051 (N_6051,N_3441,N_896);
nor U6052 (N_6052,N_1587,N_815);
nor U6053 (N_6053,N_4181,N_2964);
or U6054 (N_6054,N_3466,N_2538);
xnor U6055 (N_6055,N_4906,N_1102);
and U6056 (N_6056,N_4068,N_2381);
xnor U6057 (N_6057,N_538,N_3579);
and U6058 (N_6058,N_3403,N_1155);
nand U6059 (N_6059,N_4955,N_1643);
or U6060 (N_6060,N_1672,N_4610);
nand U6061 (N_6061,N_3453,N_766);
nor U6062 (N_6062,N_2359,N_4486);
nand U6063 (N_6063,N_1416,N_2805);
and U6064 (N_6064,N_2211,N_4977);
and U6065 (N_6065,N_3066,N_1141);
nand U6066 (N_6066,N_4250,N_913);
and U6067 (N_6067,N_3329,N_2747);
and U6068 (N_6068,N_633,N_868);
and U6069 (N_6069,N_918,N_1796);
xor U6070 (N_6070,N_1411,N_291);
xor U6071 (N_6071,N_1918,N_513);
xnor U6072 (N_6072,N_95,N_4736);
or U6073 (N_6073,N_69,N_3339);
or U6074 (N_6074,N_2957,N_1632);
and U6075 (N_6075,N_4788,N_1039);
xnor U6076 (N_6076,N_4776,N_3529);
nand U6077 (N_6077,N_2383,N_1393);
or U6078 (N_6078,N_3373,N_3589);
xor U6079 (N_6079,N_4212,N_3207);
and U6080 (N_6080,N_1676,N_1842);
nand U6081 (N_6081,N_3592,N_1277);
and U6082 (N_6082,N_4765,N_3754);
xor U6083 (N_6083,N_1692,N_1357);
nor U6084 (N_6084,N_4116,N_2552);
nor U6085 (N_6085,N_205,N_408);
nand U6086 (N_6086,N_3031,N_2905);
nor U6087 (N_6087,N_4607,N_1347);
nand U6088 (N_6088,N_1539,N_4432);
nor U6089 (N_6089,N_4962,N_3357);
or U6090 (N_6090,N_4094,N_4731);
nor U6091 (N_6091,N_4173,N_3113);
or U6092 (N_6092,N_4531,N_3469);
or U6093 (N_6093,N_39,N_1178);
and U6094 (N_6094,N_3443,N_2630);
xnor U6095 (N_6095,N_2112,N_1268);
xor U6096 (N_6096,N_4370,N_4596);
xor U6097 (N_6097,N_558,N_671);
nor U6098 (N_6098,N_2777,N_2028);
or U6099 (N_6099,N_2524,N_502);
nand U6100 (N_6100,N_89,N_2946);
nor U6101 (N_6101,N_3767,N_415);
nor U6102 (N_6102,N_1232,N_236);
nand U6103 (N_6103,N_511,N_3309);
nand U6104 (N_6104,N_2631,N_4925);
nand U6105 (N_6105,N_4043,N_1845);
and U6106 (N_6106,N_468,N_4267);
nor U6107 (N_6107,N_949,N_2820);
nand U6108 (N_6108,N_873,N_125);
xor U6109 (N_6109,N_1708,N_1112);
nand U6110 (N_6110,N_1203,N_4859);
xnor U6111 (N_6111,N_506,N_2548);
and U6112 (N_6112,N_601,N_2501);
nor U6113 (N_6113,N_2585,N_3248);
or U6114 (N_6114,N_4305,N_1580);
and U6115 (N_6115,N_1550,N_3332);
nor U6116 (N_6116,N_2658,N_3430);
xor U6117 (N_6117,N_2521,N_1705);
xnor U6118 (N_6118,N_2596,N_2417);
nor U6119 (N_6119,N_3483,N_883);
and U6120 (N_6120,N_2834,N_713);
or U6121 (N_6121,N_4634,N_2118);
and U6122 (N_6122,N_1660,N_1126);
nor U6123 (N_6123,N_4604,N_1911);
xor U6124 (N_6124,N_4561,N_3587);
xor U6125 (N_6125,N_3069,N_4118);
nand U6126 (N_6126,N_4870,N_4182);
xnor U6127 (N_6127,N_1169,N_1423);
nor U6128 (N_6128,N_2695,N_392);
nand U6129 (N_6129,N_4473,N_2354);
xnor U6130 (N_6130,N_2015,N_1049);
nand U6131 (N_6131,N_1134,N_736);
nand U6132 (N_6132,N_1448,N_2009);
nor U6133 (N_6133,N_2305,N_2208);
nand U6134 (N_6134,N_2483,N_1230);
and U6135 (N_6135,N_3611,N_535);
nand U6136 (N_6136,N_3030,N_1696);
nor U6137 (N_6137,N_405,N_1571);
or U6138 (N_6138,N_1037,N_518);
xnor U6139 (N_6139,N_1341,N_4440);
nand U6140 (N_6140,N_3161,N_1335);
nand U6141 (N_6141,N_3977,N_1709);
and U6142 (N_6142,N_4705,N_2183);
or U6143 (N_6143,N_1923,N_3675);
xnor U6144 (N_6144,N_520,N_899);
or U6145 (N_6145,N_4299,N_1387);
xnor U6146 (N_6146,N_2943,N_4300);
nand U6147 (N_6147,N_2598,N_318);
xnor U6148 (N_6148,N_2023,N_1702);
nand U6149 (N_6149,N_3148,N_3310);
nand U6150 (N_6150,N_4032,N_4793);
xnor U6151 (N_6151,N_3563,N_2480);
nand U6152 (N_6152,N_1882,N_3123);
and U6153 (N_6153,N_4824,N_2228);
xnor U6154 (N_6154,N_643,N_3337);
or U6155 (N_6155,N_2888,N_2755);
nand U6156 (N_6156,N_1404,N_1013);
nor U6157 (N_6157,N_232,N_4968);
or U6158 (N_6158,N_1802,N_2726);
nor U6159 (N_6159,N_2764,N_1139);
nor U6160 (N_6160,N_55,N_1008);
nand U6161 (N_6161,N_2676,N_196);
xnor U6162 (N_6162,N_703,N_1103);
and U6163 (N_6163,N_3064,N_2166);
nor U6164 (N_6164,N_2474,N_3470);
xnor U6165 (N_6165,N_130,N_1351);
and U6166 (N_6166,N_2689,N_4868);
xnor U6167 (N_6167,N_1135,N_4392);
or U6168 (N_6168,N_4338,N_4673);
or U6169 (N_6169,N_2586,N_2763);
or U6170 (N_6170,N_334,N_3035);
nor U6171 (N_6171,N_4553,N_1769);
or U6172 (N_6172,N_3844,N_4679);
xor U6173 (N_6173,N_3221,N_4986);
or U6174 (N_6174,N_2423,N_115);
nor U6175 (N_6175,N_1210,N_2410);
nand U6176 (N_6176,N_4762,N_2884);
or U6177 (N_6177,N_4586,N_2326);
and U6178 (N_6178,N_2876,N_2931);
xnor U6179 (N_6179,N_64,N_1703);
nand U6180 (N_6180,N_2376,N_2469);
or U6181 (N_6181,N_3489,N_545);
or U6182 (N_6182,N_2309,N_2229);
nand U6183 (N_6183,N_928,N_0);
nand U6184 (N_6184,N_3884,N_2770);
nand U6185 (N_6185,N_143,N_1590);
nand U6186 (N_6186,N_1704,N_2874);
nand U6187 (N_6187,N_4759,N_2993);
xnor U6188 (N_6188,N_4963,N_2290);
and U6189 (N_6189,N_4166,N_3858);
and U6190 (N_6190,N_1146,N_2795);
xor U6191 (N_6191,N_3869,N_22);
xnor U6192 (N_6192,N_3947,N_2131);
nor U6193 (N_6193,N_4827,N_330);
nor U6194 (N_6194,N_2495,N_4433);
and U6195 (N_6195,N_4031,N_2348);
nand U6196 (N_6196,N_1295,N_3875);
or U6197 (N_6197,N_3304,N_167);
nand U6198 (N_6198,N_1215,N_2659);
xor U6199 (N_6199,N_2061,N_1034);
xnor U6200 (N_6200,N_3550,N_3581);
xor U6201 (N_6201,N_3325,N_4163);
or U6202 (N_6202,N_327,N_1371);
nor U6203 (N_6203,N_4224,N_4427);
nand U6204 (N_6204,N_32,N_3492);
xnor U6205 (N_6205,N_3495,N_2387);
and U6206 (N_6206,N_1020,N_88);
xor U6207 (N_6207,N_4701,N_4477);
or U6208 (N_6208,N_579,N_4621);
and U6209 (N_6209,N_1659,N_2266);
nand U6210 (N_6210,N_3490,N_2020);
and U6211 (N_6211,N_3846,N_741);
or U6212 (N_6212,N_1082,N_3372);
nand U6213 (N_6213,N_1429,N_2652);
nand U6214 (N_6214,N_448,N_4372);
nor U6215 (N_6215,N_1436,N_4814);
nor U6216 (N_6216,N_1907,N_4771);
xor U6217 (N_6217,N_311,N_3915);
or U6218 (N_6218,N_1446,N_4090);
and U6219 (N_6219,N_4769,N_3750);
or U6220 (N_6220,N_2671,N_378);
nand U6221 (N_6221,N_4655,N_2173);
nand U6222 (N_6222,N_2218,N_422);
nor U6223 (N_6223,N_561,N_194);
nor U6224 (N_6224,N_826,N_1406);
nor U6225 (N_6225,N_4158,N_3777);
or U6226 (N_6226,N_854,N_3926);
nand U6227 (N_6227,N_446,N_2609);
xor U6228 (N_6228,N_3455,N_3796);
or U6229 (N_6229,N_1508,N_4745);
nor U6230 (N_6230,N_3051,N_4001);
xor U6231 (N_6231,N_2996,N_4577);
or U6232 (N_6232,N_3764,N_3163);
nor U6233 (N_6233,N_1848,N_4933);
xor U6234 (N_6234,N_3194,N_2750);
xor U6235 (N_6235,N_3534,N_2930);
or U6236 (N_6236,N_4719,N_4805);
and U6237 (N_6237,N_3927,N_3608);
or U6238 (N_6238,N_3114,N_4728);
xor U6239 (N_6239,N_2327,N_4320);
xnor U6240 (N_6240,N_1482,N_1836);
nor U6241 (N_6241,N_4954,N_1706);
nor U6242 (N_6242,N_656,N_245);
nor U6243 (N_6243,N_3826,N_253);
xnor U6244 (N_6244,N_581,N_267);
nor U6245 (N_6245,N_4716,N_2127);
xnor U6246 (N_6246,N_4938,N_373);
or U6247 (N_6247,N_1577,N_391);
nor U6248 (N_6248,N_4936,N_1510);
nor U6249 (N_6249,N_3544,N_3448);
nand U6250 (N_6250,N_4197,N_474);
or U6251 (N_6251,N_4993,N_3383);
nand U6252 (N_6252,N_1307,N_2806);
xor U6253 (N_6253,N_4241,N_797);
or U6254 (N_6254,N_3474,N_2254);
xnor U6255 (N_6255,N_2189,N_605);
nor U6256 (N_6256,N_3576,N_1938);
nor U6257 (N_6257,N_533,N_121);
and U6258 (N_6258,N_2137,N_3962);
and U6259 (N_6259,N_827,N_1926);
xnor U6260 (N_6260,N_2201,N_1749);
nand U6261 (N_6261,N_499,N_4743);
xnor U6262 (N_6262,N_3235,N_2951);
and U6263 (N_6263,N_871,N_3556);
nor U6264 (N_6264,N_4808,N_2844);
nor U6265 (N_6265,N_1656,N_38);
nand U6266 (N_6266,N_4269,N_2109);
or U6267 (N_6267,N_801,N_1217);
or U6268 (N_6268,N_1969,N_4205);
and U6269 (N_6269,N_4362,N_1990);
nor U6270 (N_6270,N_679,N_2855);
nand U6271 (N_6271,N_3838,N_386);
nand U6272 (N_6272,N_371,N_4817);
nor U6273 (N_6273,N_2481,N_747);
xnor U6274 (N_6274,N_3756,N_2738);
xor U6275 (N_6275,N_2563,N_4092);
xnor U6276 (N_6276,N_1004,N_3701);
xnor U6277 (N_6277,N_3368,N_4722);
and U6278 (N_6278,N_440,N_3179);
xnor U6279 (N_6279,N_1564,N_3213);
xnor U6280 (N_6280,N_708,N_2004);
or U6281 (N_6281,N_4245,N_1449);
xor U6282 (N_6282,N_1131,N_3334);
or U6283 (N_6283,N_2134,N_4050);
and U6284 (N_6284,N_2985,N_3876);
or U6285 (N_6285,N_293,N_4837);
and U6286 (N_6286,N_1502,N_4746);
and U6287 (N_6287,N_4436,N_3797);
nor U6288 (N_6288,N_1798,N_2940);
nand U6289 (N_6289,N_3924,N_3897);
nand U6290 (N_6290,N_2703,N_723);
nand U6291 (N_6291,N_1883,N_2140);
xor U6292 (N_6292,N_1333,N_1219);
nor U6293 (N_6293,N_1124,N_1462);
nor U6294 (N_6294,N_2144,N_2205);
xnor U6295 (N_6295,N_1753,N_4633);
xor U6296 (N_6296,N_1104,N_2927);
nor U6297 (N_6297,N_2991,N_838);
nor U6298 (N_6298,N_4613,N_3398);
xor U6299 (N_6299,N_3566,N_2058);
xor U6300 (N_6300,N_1530,N_722);
and U6301 (N_6301,N_3250,N_2626);
and U6302 (N_6302,N_4945,N_2617);
xor U6303 (N_6303,N_1797,N_2360);
xor U6304 (N_6304,N_3745,N_4148);
nor U6305 (N_6305,N_3048,N_2722);
nor U6306 (N_6306,N_3723,N_50);
and U6307 (N_6307,N_1285,N_3420);
nor U6308 (N_6308,N_4715,N_4112);
or U6309 (N_6309,N_4062,N_4086);
and U6310 (N_6310,N_1024,N_1032);
or U6311 (N_6311,N_132,N_4535);
and U6312 (N_6312,N_3673,N_2427);
nand U6313 (N_6313,N_3991,N_617);
and U6314 (N_6314,N_3109,N_4471);
nand U6315 (N_6315,N_2193,N_3936);
xor U6316 (N_6316,N_3370,N_2445);
xor U6317 (N_6317,N_2728,N_1935);
xnor U6318 (N_6318,N_1743,N_4562);
and U6319 (N_6319,N_1896,N_1087);
and U6320 (N_6320,N_4780,N_2472);
xnor U6321 (N_6321,N_1946,N_2622);
nand U6322 (N_6322,N_4483,N_2158);
nor U6323 (N_6323,N_3042,N_818);
and U6324 (N_6324,N_1453,N_4654);
xor U6325 (N_6325,N_4481,N_1289);
xnor U6326 (N_6326,N_3793,N_2561);
xor U6327 (N_6327,N_3800,N_4304);
or U6328 (N_6328,N_3274,N_3402);
and U6329 (N_6329,N_3321,N_4485);
or U6330 (N_6330,N_4309,N_3923);
or U6331 (N_6331,N_4463,N_834);
and U6332 (N_6332,N_4785,N_4886);
or U6333 (N_6333,N_1107,N_4841);
and U6334 (N_6334,N_4347,N_1254);
and U6335 (N_6335,N_1840,N_2815);
and U6336 (N_6336,N_2683,N_2343);
xnor U6337 (N_6337,N_3153,N_1136);
and U6338 (N_6338,N_1742,N_3814);
nor U6339 (N_6339,N_1651,N_1716);
nor U6340 (N_6340,N_754,N_346);
nor U6341 (N_6341,N_3684,N_1197);
xnor U6342 (N_6342,N_632,N_4584);
and U6343 (N_6343,N_2845,N_1616);
xnor U6344 (N_6344,N_353,N_1494);
and U6345 (N_6345,N_3020,N_1373);
and U6346 (N_6346,N_3519,N_3079);
nand U6347 (N_6347,N_2115,N_583);
xnor U6348 (N_6348,N_2970,N_1118);
xor U6349 (N_6349,N_2210,N_4796);
nor U6350 (N_6350,N_4277,N_4405);
nand U6351 (N_6351,N_1604,N_2382);
or U6352 (N_6352,N_4310,N_416);
or U6353 (N_6353,N_4831,N_4187);
nand U6354 (N_6354,N_3029,N_3333);
xor U6355 (N_6355,N_3454,N_4407);
xor U6356 (N_6356,N_4327,N_3077);
or U6357 (N_6357,N_921,N_4932);
xor U6358 (N_6358,N_1787,N_821);
xnor U6359 (N_6359,N_2014,N_4838);
xor U6360 (N_6360,N_840,N_485);
nand U6361 (N_6361,N_208,N_4619);
and U6362 (N_6362,N_682,N_4676);
nand U6363 (N_6363,N_1750,N_3412);
or U6364 (N_6364,N_2558,N_3522);
xor U6365 (N_6365,N_527,N_3239);
and U6366 (N_6366,N_4775,N_1951);
nand U6367 (N_6367,N_4131,N_2869);
nor U6368 (N_6368,N_1872,N_2850);
xnor U6369 (N_6369,N_471,N_578);
nor U6370 (N_6370,N_1775,N_2107);
or U6371 (N_6371,N_246,N_3217);
or U6372 (N_6372,N_1470,N_4151);
nand U6373 (N_6373,N_2414,N_1116);
nand U6374 (N_6374,N_574,N_630);
or U6375 (N_6375,N_2467,N_3640);
nor U6376 (N_6376,N_2643,N_849);
or U6377 (N_6377,N_2545,N_926);
or U6378 (N_6378,N_4375,N_4341);
and U6379 (N_6379,N_3423,N_841);
and U6380 (N_6380,N_490,N_3327);
and U6381 (N_6381,N_2351,N_4930);
and U6382 (N_6382,N_3140,N_2150);
nand U6383 (N_6383,N_3682,N_3101);
nor U6384 (N_6384,N_12,N_4952);
nor U6385 (N_6385,N_3265,N_4039);
and U6386 (N_6386,N_4514,N_3842);
or U6387 (N_6387,N_3206,N_1270);
or U6388 (N_6388,N_2325,N_1695);
xnor U6389 (N_6389,N_3399,N_2404);
nand U6390 (N_6390,N_3689,N_106);
xor U6391 (N_6391,N_476,N_773);
and U6392 (N_6392,N_720,N_1605);
nor U6393 (N_6393,N_3401,N_3788);
nor U6394 (N_6394,N_1003,N_3570);
and U6395 (N_6395,N_1863,N_3515);
nand U6396 (N_6396,N_2209,N_1434);
nand U6397 (N_6397,N_3512,N_3995);
and U6398 (N_6398,N_1378,N_3382);
and U6399 (N_6399,N_393,N_1202);
nor U6400 (N_6400,N_359,N_1152);
nand U6401 (N_6401,N_1799,N_2485);
nand U6402 (N_6402,N_4329,N_2452);
or U6403 (N_6403,N_4622,N_455);
xnor U6404 (N_6404,N_887,N_210);
nand U6405 (N_6405,N_4869,N_1746);
or U6406 (N_6406,N_4887,N_3575);
and U6407 (N_6407,N_1735,N_1538);
xor U6408 (N_6408,N_3760,N_2475);
and U6409 (N_6409,N_2657,N_4641);
nor U6410 (N_6410,N_4521,N_444);
nand U6411 (N_6411,N_3930,N_1917);
xnor U6412 (N_6412,N_1096,N_3435);
xnor U6413 (N_6413,N_3137,N_1272);
and U6414 (N_6414,N_365,N_1205);
and U6415 (N_6415,N_844,N_4984);
nand U6416 (N_6416,N_1930,N_3119);
or U6417 (N_6417,N_2177,N_1629);
nand U6418 (N_6418,N_777,N_2350);
and U6419 (N_6419,N_2642,N_1927);
nor U6420 (N_6420,N_3081,N_1244);
xor U6421 (N_6421,N_4576,N_4969);
xor U6422 (N_6422,N_370,N_3005);
nand U6423 (N_6423,N_1720,N_4983);
or U6424 (N_6424,N_3602,N_1234);
and U6425 (N_6425,N_2022,N_3283);
nand U6426 (N_6426,N_3422,N_1329);
nor U6427 (N_6427,N_2633,N_2889);
and U6428 (N_6428,N_1362,N_4712);
xor U6429 (N_6429,N_1627,N_1793);
and U6430 (N_6430,N_411,N_1176);
xnor U6431 (N_6431,N_149,N_610);
or U6432 (N_6432,N_4883,N_306);
xnor U6433 (N_6433,N_3068,N_3409);
nand U6434 (N_6434,N_3981,N_864);
xnor U6435 (N_6435,N_3562,N_3183);
or U6436 (N_6436,N_1679,N_1425);
xnor U6437 (N_6437,N_1327,N_3644);
nor U6438 (N_6438,N_1586,N_467);
nor U6439 (N_6439,N_4558,N_3843);
nor U6440 (N_6440,N_2226,N_4013);
xnor U6441 (N_6441,N_3335,N_4851);
or U6442 (N_6442,N_4225,N_2613);
or U6443 (N_6443,N_72,N_1809);
nand U6444 (N_6444,N_3095,N_2819);
nor U6445 (N_6445,N_2398,N_2388);
nor U6446 (N_6446,N_4660,N_1184);
and U6447 (N_6447,N_641,N_1724);
and U6448 (N_6448,N_1518,N_2605);
and U6449 (N_6449,N_4985,N_3698);
nand U6450 (N_6450,N_2555,N_1028);
and U6451 (N_6451,N_1513,N_2344);
nor U6452 (N_6452,N_4638,N_3458);
nand U6453 (N_6453,N_37,N_3895);
nor U6454 (N_6454,N_1960,N_4689);
or U6455 (N_6455,N_1782,N_4582);
xnor U6456 (N_6456,N_929,N_3841);
nor U6457 (N_6457,N_3700,N_1776);
and U6458 (N_6458,N_2737,N_585);
nor U6459 (N_6459,N_4787,N_3175);
nor U6460 (N_6460,N_4333,N_3768);
and U6461 (N_6461,N_2504,N_1725);
xnor U6462 (N_6462,N_2708,N_3009);
and U6463 (N_6463,N_3816,N_2828);
or U6464 (N_6464,N_4159,N_751);
and U6465 (N_6465,N_2071,N_4708);
and U6466 (N_6466,N_2043,N_1328);
nand U6467 (N_6467,N_3257,N_1693);
nor U6468 (N_6468,N_1572,N_2802);
or U6469 (N_6469,N_4360,N_799);
or U6470 (N_6470,N_2730,N_1182);
nand U6471 (N_6471,N_4575,N_2032);
xor U6472 (N_6472,N_3871,N_4846);
or U6473 (N_6473,N_2830,N_2262);
or U6474 (N_6474,N_1045,N_493);
or U6475 (N_6475,N_3668,N_525);
xor U6476 (N_6476,N_1166,N_3713);
xnor U6477 (N_6477,N_2460,N_4758);
nor U6478 (N_6478,N_2725,N_1145);
xnor U6479 (N_6479,N_2566,N_454);
or U6480 (N_6480,N_276,N_4997);
nor U6481 (N_6481,N_4903,N_3326);
or U6482 (N_6482,N_2971,N_1818);
nand U6483 (N_6483,N_163,N_2280);
or U6484 (N_6484,N_2477,N_2656);
or U6485 (N_6485,N_2824,N_2322);
nand U6486 (N_6486,N_4811,N_4139);
xnor U6487 (N_6487,N_3970,N_3762);
nor U6488 (N_6488,N_2029,N_3279);
xor U6489 (N_6489,N_1525,N_3984);
xor U6490 (N_6490,N_1030,N_2580);
or U6491 (N_6491,N_1056,N_2674);
and U6492 (N_6492,N_2455,N_700);
xor U6493 (N_6493,N_51,N_3662);
nor U6494 (N_6494,N_3425,N_4424);
xnor U6495 (N_6495,N_2500,N_992);
xor U6496 (N_6496,N_1457,N_989);
nand U6497 (N_6497,N_3599,N_4165);
nand U6498 (N_6498,N_627,N_4768);
xor U6499 (N_6499,N_2706,N_3136);
or U6500 (N_6500,N_709,N_3663);
nor U6501 (N_6501,N_3509,N_1342);
xor U6502 (N_6502,N_3528,N_4801);
or U6503 (N_6503,N_4567,N_2315);
nand U6504 (N_6504,N_2324,N_2223);
and U6505 (N_6505,N_315,N_4388);
nor U6506 (N_6506,N_948,N_4989);
and U6507 (N_6507,N_2553,N_3791);
nor U6508 (N_6508,N_1905,N_531);
nand U6509 (N_6509,N_2008,N_4453);
nand U6510 (N_6510,N_331,N_3933);
nand U6511 (N_6511,N_2732,N_4819);
or U6512 (N_6512,N_2921,N_288);
nand U6513 (N_6513,N_4934,N_1544);
or U6514 (N_6514,N_2765,N_4702);
or U6515 (N_6515,N_1463,N_489);
nor U6516 (N_6516,N_216,N_986);
or U6517 (N_6517,N_2328,N_4384);
or U6518 (N_6518,N_1044,N_4534);
nor U6519 (N_6519,N_2559,N_944);
xnor U6520 (N_6520,N_4222,N_1800);
or U6521 (N_6521,N_1269,N_1090);
xor U6522 (N_6522,N_4395,N_2079);
and U6523 (N_6523,N_762,N_609);
nor U6524 (N_6524,N_3785,N_2053);
nor U6525 (N_6525,N_2479,N_1977);
nor U6526 (N_6526,N_4674,N_1188);
or U6527 (N_6527,N_2251,N_4348);
and U6528 (N_6528,N_1158,N_3162);
nand U6529 (N_6529,N_19,N_4017);
nor U6530 (N_6530,N_321,N_217);
xor U6531 (N_6531,N_4790,N_4184);
or U6532 (N_6532,N_3354,N_1487);
nand U6533 (N_6533,N_2926,N_724);
nor U6534 (N_6534,N_225,N_735);
nand U6535 (N_6535,N_2697,N_4221);
nor U6536 (N_6536,N_945,N_3783);
or U6537 (N_6537,N_4312,N_1549);
xor U6538 (N_6538,N_1123,N_2283);
nor U6539 (N_6539,N_15,N_1599);
xnor U6540 (N_6540,N_3330,N_2791);
nor U6541 (N_6541,N_2610,N_4434);
nand U6542 (N_6542,N_4240,N_3209);
and U6543 (N_6543,N_3315,N_374);
xor U6544 (N_6544,N_2377,N_2814);
or U6545 (N_6545,N_1758,N_2365);
and U6546 (N_6546,N_702,N_1852);
or U6547 (N_6547,N_2473,N_2454);
or U6548 (N_6548,N_2860,N_3019);
and U6549 (N_6549,N_2214,N_2135);
and U6550 (N_6550,N_3456,N_1670);
nand U6551 (N_6551,N_4640,N_2984);
and U6552 (N_6552,N_3879,N_1231);
nor U6553 (N_6553,N_1744,N_2640);
nand U6554 (N_6554,N_423,N_638);
nand U6555 (N_6555,N_4152,N_3514);
nor U6556 (N_6556,N_1093,N_4260);
nand U6557 (N_6557,N_4091,N_910);
and U6558 (N_6558,N_3352,N_4581);
nor U6559 (N_6559,N_3346,N_895);
and U6560 (N_6560,N_1554,N_3138);
or U6561 (N_6561,N_4878,N_4667);
and U6562 (N_6562,N_404,N_30);
nand U6563 (N_6563,N_4501,N_3376);
xor U6564 (N_6564,N_2941,N_1664);
and U6565 (N_6565,N_603,N_4203);
and U6566 (N_6566,N_2385,N_4191);
nand U6567 (N_6567,N_3980,N_4426);
and U6568 (N_6568,N_1859,N_260);
nor U6569 (N_6569,N_2153,N_2242);
xor U6570 (N_6570,N_3038,N_970);
and U6571 (N_6571,N_2612,N_2578);
or U6572 (N_6572,N_828,N_1830);
nand U6573 (N_6573,N_3294,N_2628);
and U6574 (N_6574,N_6,N_335);
xnor U6575 (N_6575,N_4451,N_2788);
nand U6576 (N_6576,N_3902,N_1851);
nand U6577 (N_6577,N_4533,N_1479);
nor U6578 (N_6578,N_142,N_1739);
nor U6579 (N_6579,N_1305,N_2911);
nand U6580 (N_6580,N_3237,N_1472);
nor U6581 (N_6581,N_1383,N_2440);
or U6582 (N_6582,N_1973,N_4532);
and U6583 (N_6583,N_201,N_4528);
xnor U6584 (N_6584,N_3426,N_1541);
and U6585 (N_6585,N_1994,N_1421);
or U6586 (N_6586,N_2994,N_1986);
xnor U6587 (N_6587,N_4271,N_2821);
or U6588 (N_6588,N_1115,N_4909);
and U6589 (N_6589,N_1650,N_268);
or U6590 (N_6590,N_1084,N_2011);
and U6591 (N_6591,N_1786,N_4270);
or U6592 (N_6592,N_2317,N_1989);
and U6593 (N_6593,N_2938,N_3888);
or U6594 (N_6594,N_726,N_2426);
xor U6595 (N_6595,N_3181,N_1192);
or U6596 (N_6596,N_619,N_2241);
nor U6597 (N_6597,N_2729,N_3049);
nand U6598 (N_6598,N_1662,N_274);
nand U6599 (N_6599,N_4071,N_1772);
xor U6600 (N_6600,N_4145,N_4015);
nor U6601 (N_6601,N_852,N_793);
and U6602 (N_6602,N_1326,N_4657);
nand U6603 (N_6603,N_4325,N_4552);
nor U6604 (N_6604,N_4645,N_1260);
xor U6605 (N_6605,N_4083,N_4119);
and U6606 (N_6606,N_4268,N_3011);
nand U6607 (N_6607,N_776,N_843);
nor U6608 (N_6608,N_599,N_2621);
xor U6609 (N_6609,N_865,N_84);
or U6610 (N_6610,N_3427,N_255);
and U6611 (N_6611,N_534,N_290);
nor U6612 (N_6612,N_1077,N_3358);
nor U6613 (N_6613,N_3715,N_1745);
nand U6614 (N_6614,N_1806,N_4662);
or U6615 (N_6615,N_640,N_178);
or U6616 (N_6616,N_367,N_3965);
xor U6617 (N_6617,N_3825,N_1265);
nand U6618 (N_6618,N_2331,N_3397);
nand U6619 (N_6619,N_2924,N_3943);
and U6620 (N_6620,N_1430,N_4295);
nor U6621 (N_6621,N_1533,N_4940);
or U6622 (N_6622,N_4337,N_96);
or U6623 (N_6623,N_2746,N_2086);
and U6624 (N_6624,N_1626,N_1227);
xor U6625 (N_6625,N_4155,N_4389);
and U6626 (N_6626,N_3062,N_1928);
or U6627 (N_6627,N_2771,N_2256);
or U6628 (N_6628,N_1598,N_4065);
and U6629 (N_6629,N_1729,N_1368);
or U6630 (N_6630,N_4066,N_886);
nor U6631 (N_6631,N_3418,N_3919);
nor U6632 (N_6632,N_2275,N_2090);
nor U6633 (N_6633,N_1473,N_2785);
nand U6634 (N_6634,N_57,N_2913);
and U6635 (N_6635,N_477,N_3208);
nand U6636 (N_6636,N_3150,N_2439);
nor U6637 (N_6637,N_636,N_2812);
nand U6638 (N_6638,N_1984,N_1174);
or U6639 (N_6639,N_280,N_4124);
and U6640 (N_6640,N_2589,N_775);
xnor U6641 (N_6641,N_4540,N_785);
or U6642 (N_6642,N_2021,N_3664);
nor U6643 (N_6643,N_2822,N_2048);
nand U6644 (N_6644,N_4211,N_2113);
or U6645 (N_6645,N_1937,N_2877);
or U6646 (N_6646,N_263,N_1961);
and U6647 (N_6647,N_1250,N_3345);
or U6648 (N_6648,N_1224,N_2438);
nor U6649 (N_6649,N_1236,N_505);
or U6650 (N_6650,N_1433,N_1647);
nor U6651 (N_6651,N_3516,N_3487);
nand U6652 (N_6652,N_2854,N_1461);
xor U6653 (N_6653,N_3149,N_3731);
and U6654 (N_6654,N_4193,N_1253);
and U6655 (N_6655,N_1027,N_3491);
xnor U6656 (N_6656,N_1914,N_3156);
xor U6657 (N_6657,N_1657,N_2222);
or U6658 (N_6658,N_4971,N_1153);
or U6659 (N_6659,N_4349,N_1922);
nand U6660 (N_6660,N_4442,N_4280);
or U6661 (N_6661,N_3799,N_3288);
or U6662 (N_6662,N_3765,N_1257);
and U6663 (N_6663,N_118,N_54);
or U6664 (N_6664,N_4141,N_3985);
xor U6665 (N_6665,N_1258,N_126);
or U6666 (N_6666,N_2496,N_3660);
nand U6667 (N_6667,N_360,N_2476);
or U6668 (N_6668,N_3061,N_654);
and U6669 (N_6669,N_781,N_510);
nor U6670 (N_6670,N_3779,N_2973);
or U6671 (N_6671,N_3322,N_4217);
or U6672 (N_6672,N_221,N_4042);
nand U6673 (N_6673,N_2694,N_4783);
and U6674 (N_6674,N_1886,N_1471);
nor U6675 (N_6675,N_3164,N_4524);
nor U6676 (N_6676,N_809,N_2098);
and U6677 (N_6677,N_4913,N_1847);
xnor U6678 (N_6678,N_354,N_1094);
or U6679 (N_6679,N_1671,N_4177);
xnor U6680 (N_6680,N_4749,N_1857);
nor U6681 (N_6681,N_2072,N_3186);
nand U6682 (N_6682,N_4571,N_1058);
xor U6683 (N_6683,N_3567,N_1713);
nand U6684 (N_6684,N_3596,N_2817);
nand U6685 (N_6685,N_2357,N_4283);
or U6686 (N_6686,N_2898,N_326);
or U6687 (N_6687,N_1040,N_1774);
or U6688 (N_6688,N_2230,N_1843);
nand U6689 (N_6689,N_4972,N_4037);
or U6690 (N_6690,N_3821,N_836);
nor U6691 (N_6691,N_3218,N_2138);
nor U6692 (N_6692,N_1869,N_3604);
nor U6693 (N_6693,N_2549,N_1308);
nand U6694 (N_6694,N_380,N_2080);
xor U6695 (N_6695,N_3818,N_2077);
nor U6696 (N_6696,N_2296,N_2623);
xnor U6697 (N_6697,N_3010,N_4178);
nand U6698 (N_6698,N_3060,N_3798);
or U6699 (N_6699,N_177,N_60);
nor U6700 (N_6700,N_2881,N_3998);
xnor U6701 (N_6701,N_4507,N_4854);
or U6702 (N_6702,N_806,N_29);
nand U6703 (N_6703,N_279,N_3591);
nor U6704 (N_6704,N_3801,N_3772);
xor U6705 (N_6705,N_878,N_155);
nor U6706 (N_6706,N_2883,N_3360);
xor U6707 (N_6707,N_1048,N_1684);
nor U6708 (N_6708,N_3612,N_2128);
xor U6709 (N_6709,N_1854,N_794);
or U6710 (N_6710,N_3568,N_4723);
nand U6711 (N_6711,N_197,N_447);
and U6712 (N_6712,N_4735,N_3770);
and U6713 (N_6713,N_2453,N_3249);
xnor U6714 (N_6714,N_2042,N_387);
nand U6715 (N_6715,N_2618,N_2403);
nand U6716 (N_6716,N_4928,N_3959);
or U6717 (N_6717,N_3145,N_3356);
xnor U6718 (N_6718,N_3868,N_3833);
and U6719 (N_6719,N_4088,N_2916);
or U6720 (N_6720,N_4234,N_3851);
nor U6721 (N_6721,N_897,N_3319);
xnor U6722 (N_6722,N_2093,N_4265);
and U6723 (N_6723,N_338,N_1228);
and U6724 (N_6724,N_1547,N_133);
or U6725 (N_6725,N_3819,N_1012);
nor U6726 (N_6726,N_3073,N_2923);
and U6727 (N_6727,N_1010,N_146);
nor U6728 (N_6728,N_3215,N_4616);
and U6729 (N_6729,N_3594,N_372);
and U6730 (N_6730,N_3481,N_3473);
or U6731 (N_6731,N_3479,N_4503);
xor U6732 (N_6732,N_626,N_622);
and U6733 (N_6733,N_935,N_547);
nand U6734 (N_6734,N_3907,N_4825);
nor U6735 (N_6735,N_1187,N_3386);
or U6736 (N_6736,N_4100,N_1568);
nor U6737 (N_6737,N_2111,N_573);
nand U6738 (N_6738,N_1885,N_2742);
or U6739 (N_6739,N_4778,N_4885);
nor U6740 (N_6740,N_3536,N_3990);
nand U6741 (N_6741,N_3974,N_541);
and U6742 (N_6742,N_3691,N_4806);
and U6743 (N_6743,N_495,N_3546);
or U6744 (N_6744,N_3307,N_3949);
xor U6745 (N_6745,N_898,N_2604);
nand U6746 (N_6746,N_3657,N_437);
nor U6747 (N_6747,N_760,N_3222);
nor U6748 (N_6748,N_2498,N_954);
nand U6749 (N_6749,N_4374,N_2413);
nor U6750 (N_6750,N_192,N_314);
or U6751 (N_6751,N_884,N_4879);
nand U6752 (N_6752,N_2070,N_3524);
or U6753 (N_6753,N_729,N_174);
or U6754 (N_6754,N_1805,N_2155);
nand U6755 (N_6755,N_3406,N_1427);
xor U6756 (N_6756,N_469,N_3986);
and U6757 (N_6757,N_3296,N_1451);
or U6758 (N_6758,N_2972,N_2436);
nand U6759 (N_6759,N_3631,N_4135);
xnor U6760 (N_6760,N_4003,N_407);
or U6761 (N_6761,N_4153,N_909);
or U6762 (N_6762,N_4021,N_4276);
nand U6763 (N_6763,N_1601,N_608);
and U6764 (N_6764,N_4589,N_218);
nor U6765 (N_6765,N_1159,N_2920);
or U6766 (N_6766,N_4132,N_1286);
xnor U6767 (N_6767,N_2159,N_3784);
or U6768 (N_6768,N_3710,N_243);
nor U6769 (N_6769,N_693,N_4482);
or U6770 (N_6770,N_2225,N_4686);
xor U6771 (N_6771,N_3378,N_2195);
nor U6772 (N_6772,N_1636,N_3751);
or U6773 (N_6773,N_1454,N_4588);
nor U6774 (N_6774,N_1148,N_4580);
nor U6775 (N_6775,N_2579,N_2885);
and U6776 (N_6776,N_1752,N_2362);
and U6777 (N_6777,N_451,N_1575);
xnor U6778 (N_6778,N_4792,N_1140);
or U6779 (N_6779,N_4130,N_1682);
nand U6780 (N_6780,N_748,N_3999);
xor U6781 (N_6781,N_2287,N_4975);
or U6782 (N_6782,N_4491,N_435);
nand U6783 (N_6783,N_977,N_358);
nand U6784 (N_6784,N_3486,N_3342);
xor U6785 (N_6785,N_2597,N_4951);
and U6786 (N_6786,N_4598,N_1395);
nand U6787 (N_6787,N_2866,N_1255);
or U6788 (N_6788,N_4069,N_1249);
nand U6789 (N_6789,N_1825,N_4852);
or U6790 (N_6790,N_1521,N_1408);
or U6791 (N_6791,N_116,N_4051);
nand U6792 (N_6792,N_1059,N_1794);
and U6793 (N_6793,N_3008,N_2142);
and U6794 (N_6794,N_2215,N_1025);
or U6795 (N_6795,N_968,N_1501);
nor U6796 (N_6796,N_4664,N_2833);
nor U6797 (N_6797,N_1783,N_2074);
xor U6798 (N_6798,N_2078,N_4336);
xor U6799 (N_6799,N_2837,N_2571);
nor U6800 (N_6800,N_4035,N_3633);
and U6801 (N_6801,N_1151,N_2741);
nand U6802 (N_6802,N_2699,N_2887);
nand U6803 (N_6803,N_2904,N_687);
and U6804 (N_6804,N_1666,N_4381);
xor U6805 (N_6805,N_4569,N_2347);
and U6806 (N_6806,N_769,N_1838);
or U6807 (N_6807,N_1894,N_2840);
nor U6808 (N_6808,N_698,N_494);
and U6809 (N_6809,N_4692,N_500);
nor U6810 (N_6810,N_1138,N_2999);
and U6811 (N_6811,N_4857,N_3961);
or U6812 (N_6812,N_4390,N_1306);
and U6813 (N_6813,N_2320,N_804);
nor U6814 (N_6814,N_137,N_3840);
nand U6815 (N_6815,N_2505,N_1637);
nor U6816 (N_6816,N_4429,N_623);
and U6817 (N_6817,N_1920,N_66);
and U6818 (N_6818,N_4095,N_1005);
nand U6819 (N_6819,N_254,N_4919);
or U6820 (N_6820,N_4961,N_4583);
and U6821 (N_6821,N_1620,N_1162);
or U6822 (N_6822,N_4856,N_2790);
or U6823 (N_6823,N_1309,N_3440);
nor U6824 (N_6824,N_3236,N_2761);
and U6825 (N_6825,N_465,N_417);
nand U6826 (N_6826,N_956,N_2083);
and U6827 (N_6827,N_1870,N_784);
nand U6828 (N_6828,N_1559,N_1066);
xor U6829 (N_6829,N_2123,N_3776);
xnor U6830 (N_6830,N_4369,N_4872);
nor U6831 (N_6831,N_4099,N_1929);
xnor U6832 (N_6832,N_3255,N_4882);
nor U6833 (N_6833,N_5,N_4495);
xnor U6834 (N_6834,N_1673,N_2655);
xnor U6835 (N_6835,N_3324,N_139);
nand U6836 (N_6836,N_851,N_934);
and U6837 (N_6837,N_2268,N_4830);
nand U6838 (N_6838,N_2066,N_4833);
and U6839 (N_6839,N_2980,N_1591);
nand U6840 (N_6840,N_4073,N_347);
nand U6841 (N_6841,N_3103,N_4045);
nand U6842 (N_6842,N_4126,N_2547);
or U6843 (N_6843,N_1715,N_4996);
nor U6844 (N_6844,N_3143,N_120);
nand U6845 (N_6845,N_1444,N_563);
nand U6846 (N_6846,N_4542,N_3523);
xnor U6847 (N_6847,N_4117,N_4650);
nand U6848 (N_6848,N_2378,N_4210);
xnor U6849 (N_6849,N_2363,N_3558);
nand U6850 (N_6850,N_361,N_2672);
nor U6851 (N_6851,N_3437,N_4420);
xnor U6852 (N_6852,N_4522,N_4009);
nor U6853 (N_6853,N_2169,N_984);
xnor U6854 (N_6854,N_2340,N_248);
or U6855 (N_6855,N_3958,N_1792);
nand U6856 (N_6856,N_3989,N_879);
nand U6857 (N_6857,N_842,N_2899);
xor U6858 (N_6858,N_432,N_4054);
xnor U6859 (N_6859,N_3605,N_1069);
nor U6860 (N_6860,N_1526,N_3166);
nor U6861 (N_6861,N_4428,N_3015);
or U6862 (N_6862,N_1125,N_3380);
xnor U6863 (N_6863,N_4350,N_2635);
or U6864 (N_6864,N_1871,N_2129);
xnor U6865 (N_6865,N_1137,N_234);
or U6866 (N_6866,N_3229,N_4929);
nand U6867 (N_6867,N_1414,N_2291);
nand U6868 (N_6868,N_4237,N_156);
nand U6869 (N_6869,N_2484,N_4242);
nand U6870 (N_6870,N_3293,N_860);
xor U6871 (N_6871,N_2314,N_4036);
or U6872 (N_6872,N_4960,N_2145);
nor U6873 (N_6873,N_4603,N_3925);
and U6874 (N_6874,N_1971,N_3834);
and U6875 (N_6875,N_4956,N_295);
nor U6876 (N_6876,N_4804,N_462);
nor U6877 (N_6877,N_3099,N_3264);
xor U6878 (N_6878,N_4246,N_2012);
nand U6879 (N_6879,N_4461,N_4056);
or U6880 (N_6880,N_333,N_3205);
nor U6881 (N_6881,N_2849,N_1211);
nand U6882 (N_6882,N_521,N_4599);
or U6883 (N_6883,N_2092,N_3622);
nor U6884 (N_6884,N_1958,N_182);
nor U6885 (N_6885,N_2735,N_1196);
and U6886 (N_6886,N_758,N_4058);
or U6887 (N_6887,N_2606,N_2216);
or U6888 (N_6888,N_2122,N_3982);
nor U6889 (N_6889,N_4147,N_148);
nor U6890 (N_6890,N_369,N_4332);
nand U6891 (N_6891,N_3085,N_4973);
nand U6892 (N_6892,N_3151,N_1452);
xnor U6893 (N_6893,N_2934,N_939);
nand U6894 (N_6894,N_3320,N_4346);
nor U6895 (N_6895,N_4033,N_2947);
nand U6896 (N_6896,N_958,N_35);
xor U6897 (N_6897,N_870,N_2535);
xnor U6898 (N_6898,N_1733,N_4468);
or U6899 (N_6899,N_4752,N_4076);
or U6900 (N_6900,N_4537,N_3086);
nand U6901 (N_6901,N_2110,N_1910);
or U6902 (N_6902,N_220,N_2076);
nor U6903 (N_6903,N_1691,N_4957);
nor U6904 (N_6904,N_2068,N_4863);
or U6905 (N_6905,N_727,N_2562);
or U6906 (N_6906,N_1766,N_737);
nor U6907 (N_6907,N_4843,N_1223);
xnor U6908 (N_6908,N_615,N_503);
xnor U6909 (N_6909,N_1619,N_1569);
nand U6910 (N_6910,N_812,N_2793);
and U6911 (N_6911,N_602,N_4681);
xor U6912 (N_6912,N_591,N_2590);
xnor U6913 (N_6913,N_77,N_58);
or U6914 (N_6914,N_3621,N_1201);
or U6915 (N_6915,N_410,N_1206);
nor U6916 (N_6916,N_379,N_3471);
xnor U6917 (N_6917,N_2034,N_4556);
nor U6918 (N_6918,N_570,N_1563);
xnor U6919 (N_6919,N_1240,N_3122);
nor U6920 (N_6920,N_3364,N_3414);
xnor U6921 (N_6921,N_4195,N_2680);
or U6922 (N_6922,N_71,N_4498);
nand U6923 (N_6923,N_3295,N_982);
nand U6924 (N_6924,N_4602,N_1593);
or U6925 (N_6925,N_692,N_1523);
or U6926 (N_6926,N_2781,N_2588);
nor U6927 (N_6927,N_233,N_4256);
or U6928 (N_6928,N_4214,N_3525);
and U6929 (N_6929,N_213,N_1952);
nand U6930 (N_6930,N_1186,N_1437);
and U6931 (N_6931,N_532,N_2124);
nand U6932 (N_6932,N_278,N_2519);
nor U6933 (N_6933,N_2407,N_3276);
nor U6934 (N_6934,N_733,N_1318);
and U6935 (N_6935,N_14,N_4316);
and U6936 (N_6936,N_919,N_526);
or U6937 (N_6937,N_3203,N_97);
or U6938 (N_6938,N_2179,N_2886);
nor U6939 (N_6939,N_4192,N_3752);
nand U6940 (N_6940,N_3432,N_4931);
xor U6941 (N_6941,N_2641,N_3996);
or U6942 (N_6942,N_663,N_4617);
xor U6943 (N_6943,N_2067,N_858);
nor U6944 (N_6944,N_2132,N_3272);
nor U6945 (N_6945,N_540,N_4029);
xnor U6946 (N_6946,N_4803,N_4865);
and U6947 (N_6947,N_4508,N_4649);
xnor U6948 (N_6948,N_1263,N_3291);
xor U6949 (N_6949,N_2019,N_3650);
nor U6950 (N_6950,N_3976,N_4387);
and U6951 (N_6951,N_11,N_61);
nand U6952 (N_6952,N_1603,N_2893);
or U6953 (N_6953,N_2301,N_2276);
nand U6954 (N_6954,N_1144,N_406);
and U6955 (N_6955,N_41,N_488);
or U6956 (N_6956,N_4510,N_2798);
or U6957 (N_6957,N_763,N_270);
and U6958 (N_6958,N_833,N_613);
xnor U6959 (N_6959,N_4464,N_4367);
xnor U6960 (N_6960,N_2200,N_3160);
xnor U6961 (N_6961,N_4323,N_2292);
nor U6962 (N_6962,N_33,N_2992);
nor U6963 (N_6963,N_3259,N_4823);
nor U6964 (N_6964,N_3736,N_4639);
and U6965 (N_6965,N_1718,N_4609);
nand U6966 (N_6966,N_2593,N_3493);
and U6967 (N_6967,N_2928,N_3336);
nand U6968 (N_6968,N_4815,N_1400);
xor U6969 (N_6969,N_717,N_4835);
or U6970 (N_6970,N_807,N_124);
nor U6971 (N_6971,N_3359,N_482);
or U6972 (N_6972,N_2338,N_3074);
nand U6973 (N_6973,N_3942,N_1588);
or U6974 (N_6974,N_3313,N_2731);
and U6975 (N_6975,N_4912,N_275);
or U6976 (N_6976,N_4171,N_634);
nor U6977 (N_6977,N_1740,N_2486);
or U6978 (N_6978,N_4307,N_528);
xnor U6979 (N_6979,N_673,N_3674);
or U6980 (N_6980,N_4317,N_2461);
xnor U6981 (N_6981,N_4632,N_4994);
or U6982 (N_6982,N_3954,N_891);
or U6983 (N_6983,N_3171,N_2679);
nand U6984 (N_6984,N_3993,N_3632);
and U6985 (N_6985,N_3634,N_3012);
xor U6986 (N_6986,N_394,N_2238);
and U6987 (N_6987,N_552,N_859);
or U6988 (N_6988,N_2651,N_491);
and U6989 (N_6989,N_3187,N_551);
and U6990 (N_6990,N_863,N_3771);
xor U6991 (N_6991,N_1302,N_4027);
and U6992 (N_6992,N_4231,N_2639);
nand U6993 (N_6993,N_3120,N_1163);
nor U6994 (N_6994,N_2293,N_685);
nor U6995 (N_6995,N_2146,N_4807);
or U6996 (N_6996,N_1428,N_3297);
nor U6997 (N_6997,N_4512,N_2733);
xor U6998 (N_6998,N_1264,N_4515);
or U6999 (N_6999,N_889,N_3232);
and U7000 (N_7000,N_2103,N_4497);
or U7001 (N_7001,N_1741,N_449);
or U7002 (N_7002,N_2198,N_3531);
xor U7003 (N_7003,N_282,N_4123);
nor U7004 (N_7004,N_4055,N_3687);
and U7005 (N_7005,N_1097,N_2515);
nand U7006 (N_7006,N_2190,N_4149);
and U7007 (N_7007,N_4699,N_1901);
or U7008 (N_7008,N_40,N_1916);
nand U7009 (N_7009,N_3882,N_3131);
xnor U7010 (N_7010,N_1172,N_3658);
and U7011 (N_7011,N_4810,N_1828);
or U7012 (N_7012,N_2969,N_3170);
nor U7013 (N_7013,N_1837,N_3268);
nand U7014 (N_7014,N_4642,N_2332);
nor U7015 (N_7015,N_4773,N_1714);
xnor U7016 (N_7016,N_4243,N_1936);
xor U7017 (N_7017,N_2826,N_1476);
or U7018 (N_7018,N_512,N_1915);
and U7019 (N_7019,N_4425,N_3475);
or U7020 (N_7020,N_3251,N_3220);
or U7021 (N_7021,N_4352,N_2003);
or U7022 (N_7022,N_4138,N_1483);
xor U7023 (N_7023,N_1891,N_3070);
nand U7024 (N_7024,N_660,N_3075);
nand U7025 (N_7025,N_4566,N_3105);
nor U7026 (N_7026,N_3937,N_4643);
and U7027 (N_7027,N_4950,N_1589);
xnor U7028 (N_7028,N_4979,N_1445);
nand U7029 (N_7029,N_3781,N_3022);
nor U7030 (N_7030,N_3667,N_1814);
and U7031 (N_7031,N_3155,N_1950);
nand U7032 (N_7032,N_2489,N_2100);
nand U7033 (N_7033,N_1278,N_4207);
nor U7034 (N_7034,N_4772,N_3132);
xor U7035 (N_7035,N_3951,N_3245);
nor U7036 (N_7036,N_1,N_4067);
xor U7037 (N_7037,N_2786,N_284);
or U7038 (N_7038,N_2720,N_3178);
nand U7039 (N_7039,N_1420,N_4591);
and U7040 (N_7040,N_560,N_1968);
and U7041 (N_7041,N_266,N_3973);
and U7042 (N_7042,N_719,N_1555);
or U7043 (N_7043,N_1527,N_339);
and U7044 (N_7044,N_1866,N_2097);
nor U7045 (N_7045,N_586,N_1815);
and U7046 (N_7046,N_381,N_2894);
and U7047 (N_7047,N_676,N_1207);
or U7048 (N_7048,N_1844,N_1271);
and U7049 (N_7049,N_4386,N_1143);
nand U7050 (N_7050,N_4606,N_2313);
nand U7051 (N_7051,N_2859,N_1293);
nand U7052 (N_7052,N_4627,N_3286);
and U7053 (N_7053,N_839,N_4549);
and U7054 (N_7054,N_1208,N_774);
or U7055 (N_7055,N_716,N_2796);
and U7056 (N_7056,N_672,N_1455);
nor U7057 (N_7057,N_2139,N_2339);
nor U7058 (N_7058,N_2197,N_2037);
and U7059 (N_7059,N_3340,N_3306);
and U7060 (N_7060,N_4456,N_2065);
nor U7061 (N_7061,N_3446,N_2265);
or U7062 (N_7062,N_872,N_20);
xor U7063 (N_7063,N_4266,N_99);
xor U7064 (N_7064,N_677,N_3539);
nor U7065 (N_7065,N_1459,N_4492);
nor U7066 (N_7066,N_2531,N_1610);
nor U7067 (N_7067,N_2808,N_1431);
and U7068 (N_7068,N_4244,N_4340);
nand U7069 (N_7069,N_770,N_1548);
nand U7070 (N_7070,N_223,N_725);
and U7071 (N_7071,N_2237,N_4910);
or U7072 (N_7072,N_987,N_1456);
xor U7073 (N_7073,N_938,N_409);
nand U7074 (N_7074,N_2152,N_4874);
and U7075 (N_7075,N_2944,N_3542);
or U7076 (N_7076,N_562,N_199);
nand U7077 (N_7077,N_1665,N_1811);
nor U7078 (N_7078,N_4137,N_2162);
nand U7079 (N_7079,N_530,N_1098);
nor U7080 (N_7080,N_1982,N_1900);
nand U7081 (N_7081,N_319,N_1130);
nor U7082 (N_7082,N_4877,N_237);
nor U7083 (N_7083,N_3679,N_170);
xnor U7084 (N_7084,N_487,N_2288);
nor U7085 (N_7085,N_3944,N_2677);
xor U7086 (N_7086,N_2902,N_1015);
nor U7087 (N_7087,N_3560,N_1394);
nand U7088 (N_7088,N_3517,N_4070);
and U7089 (N_7089,N_2499,N_389);
nand U7090 (N_7090,N_1191,N_976);
nand U7091 (N_7091,N_188,N_1060);
nor U7092 (N_7092,N_4590,N_3732);
and U7093 (N_7093,N_3769,N_3462);
nand U7094 (N_7094,N_1332,N_1248);
or U7095 (N_7095,N_1275,N_4286);
or U7096 (N_7096,N_1279,N_2355);
xor U7097 (N_7097,N_419,N_2141);
and U7098 (N_7098,N_4229,N_3507);
and U7099 (N_7099,N_4732,N_1323);
xor U7100 (N_7100,N_348,N_3447);
and U7101 (N_7101,N_4328,N_2986);
xor U7102 (N_7102,N_2059,N_1831);
and U7103 (N_7103,N_257,N_837);
or U7104 (N_7104,N_193,N_2007);
nor U7105 (N_7105,N_2570,N_4959);
or U7106 (N_7106,N_1867,N_1608);
nand U7107 (N_7107,N_300,N_3541);
nand U7108 (N_7108,N_251,N_4729);
xor U7109 (N_7109,N_3859,N_1001);
or U7110 (N_7110,N_4049,N_355);
nand U7111 (N_7111,N_2513,N_3001);
or U7112 (N_7112,N_2687,N_23);
or U7113 (N_7113,N_3697,N_1631);
and U7114 (N_7114,N_4871,N_1369);
nand U7115 (N_7115,N_1061,N_2457);
nand U7116 (N_7116,N_3831,N_4077);
and U7117 (N_7117,N_4751,N_4624);
nand U7118 (N_7118,N_1316,N_4813);
xor U7119 (N_7119,N_1583,N_3185);
xor U7120 (N_7120,N_3852,N_2646);
or U7121 (N_7121,N_704,N_363);
and U7122 (N_7122,N_2041,N_316);
and U7123 (N_7123,N_4460,N_3039);
xnor U7124 (N_7124,N_478,N_4726);
nand U7125 (N_7125,N_607,N_4288);
xnor U7126 (N_7126,N_1737,N_3375);
nor U7127 (N_7127,N_2492,N_4447);
nand U7128 (N_7128,N_4467,N_1661);
nor U7129 (N_7129,N_4281,N_375);
nor U7130 (N_7130,N_788,N_3572);
and U7131 (N_7131,N_1100,N_4096);
and U7132 (N_7132,N_1450,N_1785);
nand U7133 (N_7133,N_1711,N_1653);
nand U7134 (N_7134,N_1621,N_85);
or U7135 (N_7135,N_1874,N_4449);
xnor U7136 (N_7136,N_4194,N_2939);
xor U7137 (N_7137,N_1401,N_4829);
xor U7138 (N_7138,N_231,N_3726);
and U7139 (N_7139,N_4899,N_4764);
nor U7140 (N_7140,N_2966,N_4072);
nor U7141 (N_7141,N_2723,N_3498);
nor U7142 (N_7142,N_2243,N_4761);
xnor U7143 (N_7143,N_3738,N_2922);
or U7144 (N_7144,N_356,N_3735);
or U7145 (N_7145,N_4506,N_4547);
or U7146 (N_7146,N_3952,N_1379);
xor U7147 (N_7147,N_1424,N_2165);
xor U7148 (N_7148,N_3045,N_950);
xor U7149 (N_7149,N_1354,N_2520);
and U7150 (N_7150,N_4140,N_3389);
nor U7151 (N_7151,N_3247,N_3918);
or U7152 (N_7152,N_3836,N_4143);
or U7153 (N_7153,N_1364,N_684);
nor U7154 (N_7154,N_1888,N_1835);
xnor U7155 (N_7155,N_4943,N_1924);
nor U7156 (N_7156,N_4326,N_222);
nand U7157 (N_7157,N_1520,N_4678);
xor U7158 (N_7158,N_3740,N_1304);
or U7159 (N_7159,N_343,N_1890);
nor U7160 (N_7160,N_4038,N_2990);
and U7161 (N_7161,N_390,N_3620);
or U7162 (N_7162,N_2342,N_537);
nor U7163 (N_7163,N_4324,N_2036);
or U7164 (N_7164,N_2666,N_4430);
and U7165 (N_7165,N_4555,N_2088);
nor U7166 (N_7166,N_4255,N_17);
xor U7167 (N_7167,N_557,N_4538);
or U7168 (N_7168,N_4479,N_2149);
xor U7169 (N_7169,N_1658,N_384);
or U7170 (N_7170,N_2106,N_3040);
nor U7171 (N_7171,N_4781,N_1763);
and U7172 (N_7172,N_1198,N_3887);
xnor U7173 (N_7173,N_4172,N_4721);
or U7174 (N_7174,N_594,N_3115);
xnor U7175 (N_7175,N_4041,N_1602);
nand U7176 (N_7176,N_136,N_3302);
nor U7177 (N_7177,N_1054,N_2663);
xnor U7178 (N_7178,N_1677,N_2337);
nand U7179 (N_7179,N_1993,N_4064);
and U7180 (N_7180,N_606,N_308);
nand U7181 (N_7181,N_1909,N_4291);
xor U7182 (N_7182,N_4080,N_908);
and U7183 (N_7183,N_4010,N_3134);
or U7184 (N_7184,N_56,N_4739);
nor U7185 (N_7185,N_4915,N_1251);
xor U7186 (N_7186,N_2912,N_1403);
and U7187 (N_7187,N_2010,N_4935);
nand U7188 (N_7188,N_4675,N_4298);
nor U7189 (N_7189,N_4821,N_2977);
nand U7190 (N_7190,N_548,N_4916);
xnor U7191 (N_7191,N_75,N_443);
and U7192 (N_7192,N_3948,N_4385);
or U7193 (N_7193,N_1282,N_690);
and U7194 (N_7194,N_4378,N_2429);
xnor U7195 (N_7195,N_1484,N_4967);
xnor U7196 (N_7196,N_1399,N_1183);
nor U7197 (N_7197,N_1988,N_1943);
xnor U7198 (N_7198,N_2466,N_4000);
or U7199 (N_7199,N_324,N_1678);
xnor U7200 (N_7200,N_2692,N_3477);
and U7201 (N_7201,N_4895,N_2853);
nor U7202 (N_7202,N_1949,N_1812);
and U7203 (N_7203,N_4530,N_3526);
nand U7204 (N_7204,N_4964,N_1164);
or U7205 (N_7205,N_2745,N_3680);
nor U7206 (N_7206,N_184,N_4557);
or U7207 (N_7207,N_4098,N_2393);
or U7208 (N_7208,N_3439,N_2714);
and U7209 (N_7209,N_4226,N_4791);
and U7210 (N_7210,N_2949,N_3058);
nand U7211 (N_7211,N_3393,N_670);
and U7212 (N_7212,N_1419,N_750);
and U7213 (N_7213,N_2002,N_3204);
nor U7214 (N_7214,N_2168,N_2172);
nor U7215 (N_7215,N_1113,N_2446);
or U7216 (N_7216,N_2044,N_400);
and U7217 (N_7217,N_3934,N_2117);
nor U7218 (N_7218,N_4397,N_1507);
nand U7219 (N_7219,N_553,N_3747);
or U7220 (N_7220,N_481,N_3182);
and U7221 (N_7221,N_4383,N_3613);
xor U7222 (N_7222,N_3850,N_1349);
nand U7223 (N_7223,N_4554,N_4261);
and U7224 (N_7224,N_668,N_757);
and U7225 (N_7225,N_3533,N_445);
xor U7226 (N_7226,N_3002,N_2719);
nor U7227 (N_7227,N_2373,N_1065);
and U7228 (N_7228,N_4398,N_3400);
nor U7229 (N_7229,N_2105,N_3552);
xor U7230 (N_7230,N_2333,N_4285);
and U7231 (N_7231,N_1216,N_1076);
xor U7232 (N_7232,N_62,N_3866);
nand U7233 (N_7233,N_4565,N_4998);
or U7234 (N_7234,N_3225,N_2389);
nor U7235 (N_7235,N_2550,N_3932);
nand U7236 (N_7236,N_2514,N_4167);
nand U7237 (N_7237,N_3547,N_2607);
or U7238 (N_7238,N_1311,N_313);
xor U7239 (N_7239,N_4836,N_396);
or U7240 (N_7240,N_114,N_4128);
nor U7241 (N_7241,N_1350,N_292);
nand U7242 (N_7242,N_2544,N_3374);
xor U7243 (N_7243,N_2868,N_2411);
xor U7244 (N_7244,N_1611,N_1038);
or U7245 (N_7245,N_3802,N_3957);
nor U7246 (N_7246,N_3305,N_4902);
nor U7247 (N_7247,N_646,N_4470);
nor U7248 (N_7248,N_3017,N_791);
and U7249 (N_7249,N_2502,N_1043);
and U7250 (N_7250,N_1480,N_683);
nand U7251 (N_7251,N_689,N_4858);
and U7252 (N_7252,N_4022,N_4766);
nor U7253 (N_7253,N_3849,N_647);
nor U7254 (N_7254,N_430,N_4845);
or U7255 (N_7255,N_52,N_1291);
xnor U7256 (N_7256,N_25,N_4644);
nor U7257 (N_7257,N_398,N_3855);
and U7258 (N_7258,N_3269,N_714);
or U7259 (N_7259,N_2870,N_1194);
xnor U7260 (N_7260,N_3803,N_4315);
xor U7261 (N_7261,N_1014,N_3905);
xor U7262 (N_7262,N_1529,N_4894);
or U7263 (N_7263,N_907,N_4587);
xor U7264 (N_7264,N_1906,N_2799);
or U7265 (N_7265,N_2625,N_3025);
nor U7266 (N_7266,N_2734,N_497);
nor U7267 (N_7267,N_3125,N_795);
nand U7268 (N_7268,N_2370,N_3645);
or U7269 (N_7269,N_4052,N_3343);
xor U7270 (N_7270,N_3147,N_4047);
and U7271 (N_7271,N_4005,N_937);
nand U7272 (N_7272,N_2587,N_320);
and U7273 (N_7273,N_924,N_3139);
nand U7274 (N_7274,N_1606,N_829);
and U7275 (N_7275,N_332,N_4308);
xor U7276 (N_7276,N_4441,N_2935);
xor U7277 (N_7277,N_4016,N_3053);
or U7278 (N_7278,N_835,N_2415);
nor U7279 (N_7279,N_3318,N_1156);
xnor U7280 (N_7280,N_8,N_2380);
nand U7281 (N_7281,N_2852,N_618);
xor U7282 (N_7282,N_2126,N_1581);
nor U7283 (N_7283,N_2227,N_1754);
xnor U7284 (N_7284,N_1072,N_3082);
nor U7285 (N_7285,N_3743,N_3127);
nor U7286 (N_7286,N_990,N_2503);
nand U7287 (N_7287,N_4672,N_1361);
xnor U7288 (N_7288,N_2919,N_1633);
or U7289 (N_7289,N_4637,N_4209);
or U7290 (N_7290,N_2062,N_168);
nor U7291 (N_7291,N_2488,N_4423);
nand U7292 (N_7292,N_1726,N_1652);
nand U7293 (N_7293,N_1133,N_2574);
nor U7294 (N_7294,N_1062,N_2769);
and U7295 (N_7295,N_1789,N_715);
and U7296 (N_7296,N_1939,N_3863);
xor U7297 (N_7297,N_1903,N_1127);
or U7298 (N_7298,N_1897,N_2386);
and U7299 (N_7299,N_1976,N_1904);
nand U7300 (N_7300,N_2267,N_3729);
nor U7301 (N_7301,N_2523,N_3384);
and U7302 (N_7302,N_195,N_767);
or U7303 (N_7303,N_3699,N_4517);
xnor U7304 (N_7304,N_1985,N_2804);
nand U7305 (N_7305,N_3588,N_845);
xnor U7306 (N_7306,N_3714,N_961);
nand U7307 (N_7307,N_2171,N_4608);
and U7308 (N_7308,N_428,N_4379);
nand U7309 (N_7309,N_848,N_2753);
nor U7310 (N_7310,N_187,N_2948);
and U7311 (N_7311,N_706,N_782);
xor U7312 (N_7312,N_4754,N_4053);
nor U7313 (N_7313,N_3569,N_1991);
nand U7314 (N_7314,N_401,N_904);
and U7315 (N_7315,N_4980,N_3043);
or U7316 (N_7316,N_1534,N_4030);
and U7317 (N_7317,N_4753,N_2255);
xnor U7318 (N_7318,N_3659,N_4974);
xnor U7319 (N_7319,N_3929,N_2766);
xor U7320 (N_7320,N_3889,N_2705);
or U7321 (N_7321,N_2151,N_1376);
and U7322 (N_7322,N_764,N_4889);
nand U7323 (N_7323,N_4239,N_366);
or U7324 (N_7324,N_3344,N_3256);
nand U7325 (N_7325,N_4160,N_2601);
and U7326 (N_7326,N_3083,N_1017);
nor U7327 (N_7327,N_92,N_4864);
xnor U7328 (N_7328,N_1256,N_746);
and U7329 (N_7329,N_3088,N_1180);
nand U7330 (N_7330,N_2929,N_1839);
or U7331 (N_7331,N_1567,N_4061);
nand U7332 (N_7332,N_4944,N_3601);
and U7333 (N_7333,N_4011,N_2603);
nor U7334 (N_7334,N_3646,N_3429);
nand U7335 (N_7335,N_2527,N_2959);
and U7336 (N_7336,N_3817,N_2743);
xor U7337 (N_7337,N_2865,N_3623);
nand U7338 (N_7338,N_4818,N_269);
nand U7339 (N_7339,N_3231,N_4924);
nor U7340 (N_7340,N_1579,N_2069);
nor U7341 (N_7341,N_2956,N_963);
or U7342 (N_7342,N_285,N_3174);
xnor U7343 (N_7343,N_1396,N_2740);
nor U7344 (N_7344,N_27,N_82);
nor U7345 (N_7345,N_4319,N_3266);
nand U7346 (N_7346,N_1026,N_697);
xnor U7347 (N_7347,N_3847,N_1956);
nor U7348 (N_7348,N_2832,N_3200);
xor U7349 (N_7349,N_3808,N_1849);
and U7350 (N_7350,N_969,N_1055);
or U7351 (N_7351,N_755,N_4636);
nand U7352 (N_7352,N_433,N_1343);
and U7353 (N_7353,N_743,N_966);
nand U7354 (N_7354,N_209,N_4416);
xor U7355 (N_7355,N_2462,N_2624);
and U7356 (N_7356,N_4125,N_1035);
nand U7357 (N_7357,N_952,N_569);
xor U7358 (N_7358,N_1363,N_1300);
xnor U7359 (N_7359,N_1779,N_2428);
xnor U7360 (N_7360,N_3648,N_3595);
and U7361 (N_7361,N_3298,N_4847);
and U7362 (N_7362,N_3348,N_1290);
nand U7363 (N_7363,N_4331,N_1021);
nor U7364 (N_7364,N_731,N_3449);
and U7365 (N_7365,N_2180,N_2051);
nand U7366 (N_7366,N_1980,N_2133);
and U7367 (N_7367,N_2258,N_70);
nand U7368 (N_7368,N_1592,N_2356);
or U7369 (N_7369,N_1000,N_4812);
and U7370 (N_7370,N_1528,N_3445);
nor U7371 (N_7371,N_2712,N_2353);
nor U7372 (N_7372,N_1409,N_3609);
nor U7373 (N_7373,N_100,N_4939);
and U7374 (N_7374,N_1218,N_866);
and U7375 (N_7375,N_4190,N_203);
nor U7376 (N_7376,N_4572,N_1481);
xor U7377 (N_7377,N_1795,N_3861);
nor U7378 (N_7378,N_336,N_3472);
xor U7379 (N_7379,N_4513,N_2592);
or U7380 (N_7380,N_2176,N_1380);
and U7381 (N_7381,N_1149,N_3672);
xnor U7382 (N_7382,N_517,N_2736);
nand U7383 (N_7383,N_2253,N_2248);
and U7384 (N_7384,N_3979,N_1022);
or U7385 (N_7385,N_1721,N_2084);
or U7386 (N_7386,N_3584,N_4965);
xor U7387 (N_7387,N_3192,N_3195);
or U7388 (N_7388,N_4206,N_3189);
or U7389 (N_7389,N_575,N_3468);
or U7390 (N_7390,N_104,N_3417);
nor U7391 (N_7391,N_3202,N_2565);
or U7392 (N_7392,N_4404,N_3080);
xor U7393 (N_7393,N_138,N_1384);
nor U7394 (N_7394,N_4500,N_4489);
or U7395 (N_7395,N_4488,N_1698);
xor U7396 (N_7396,N_1466,N_198);
xor U7397 (N_7397,N_273,N_1078);
xor U7398 (N_7398,N_3975,N_1220);
and U7399 (N_7399,N_4452,N_1953);
nor U7400 (N_7400,N_351,N_1997);
and U7401 (N_7401,N_2494,N_1181);
and U7402 (N_7402,N_3885,N_3681);
and U7403 (N_7403,N_2434,N_4301);
and U7404 (N_7404,N_3299,N_4084);
or U7405 (N_7405,N_728,N_1190);
and U7406 (N_7406,N_2968,N_730);
or U7407 (N_7407,N_4106,N_173);
and U7408 (N_7408,N_4475,N_2478);
nor U7409 (N_7409,N_1821,N_4809);
nand U7410 (N_7410,N_1965,N_1325);
nor U7411 (N_7411,N_1303,N_3908);
and U7412 (N_7412,N_119,N_4202);
nor U7413 (N_7413,N_3308,N_3655);
or U7414 (N_7414,N_128,N_1913);
and U7415 (N_7415,N_4898,N_925);
or U7416 (N_7416,N_473,N_658);
or U7417 (N_7417,N_3873,N_4278);
and U7418 (N_7418,N_103,N_4941);
nand U7419 (N_7419,N_2204,N_4104);
nor U7420 (N_7420,N_3371,N_965);
nor U7421 (N_7421,N_470,N_238);
nand U7422 (N_7422,N_4081,N_1074);
nand U7423 (N_7423,N_972,N_893);
nor U7424 (N_7424,N_2390,N_1964);
nand U7425 (N_7425,N_1313,N_1699);
or U7426 (N_7426,N_4162,N_1495);
nand U7427 (N_7427,N_4313,N_4377);
nand U7428 (N_7428,N_2334,N_2463);
nor U7429 (N_7429,N_3037,N_1552);
or U7430 (N_7430,N_911,N_235);
xor U7431 (N_7431,N_458,N_572);
and U7432 (N_7432,N_2619,N_1467);
xor U7433 (N_7433,N_571,N_1945);
nor U7434 (N_7434,N_3494,N_244);
nor U7435 (N_7435,N_3270,N_2696);
nor U7436 (N_7436,N_584,N_1881);
nand U7437 (N_7437,N_3593,N_2468);
or U7438 (N_7438,N_420,N_980);
or U7439 (N_7439,N_4937,N_3978);
or U7440 (N_7440,N_3642,N_402);
nor U7441 (N_7441,N_3969,N_3865);
nor U7442 (N_7442,N_2591,N_1612);
nand U7443 (N_7443,N_2464,N_2542);
or U7444 (N_7444,N_207,N_3390);
xor U7445 (N_7445,N_4380,N_823);
or U7446 (N_7446,N_4004,N_1558);
nand U7447 (N_7447,N_287,N_1781);
or U7448 (N_7448,N_3906,N_2235);
or U7449 (N_7449,N_3117,N_4724);
or U7450 (N_7450,N_2526,N_299);
or U7451 (N_7451,N_4355,N_4927);
or U7452 (N_7452,N_2319,N_4579);
and U7453 (N_7453,N_4074,N_2311);
or U7454 (N_7454,N_2933,N_2632);
nor U7455 (N_7455,N_2143,N_3872);
xnor U7456 (N_7456,N_1536,N_151);
xor U7457 (N_7457,N_86,N_2880);
nor U7458 (N_7458,N_742,N_4048);
xnor U7459 (N_7459,N_2810,N_4594);
nor U7460 (N_7460,N_1808,N_4896);
and U7461 (N_7461,N_1639,N_2263);
nand U7462 (N_7462,N_3968,N_2371);
nor U7463 (N_7463,N_1574,N_4215);
or U7464 (N_7464,N_2095,N_1596);
or U7465 (N_7465,N_107,N_3627);
xnor U7466 (N_7466,N_1983,N_4693);
or U7467 (N_7467,N_2148,N_4188);
nand U7468 (N_7468,N_3501,N_624);
xnor U7469 (N_7469,N_2121,N_3052);
nand U7470 (N_7470,N_3431,N_805);
or U7471 (N_7471,N_2181,N_4709);
nand U7472 (N_7472,N_3543,N_1962);
xnor U7473 (N_7473,N_4635,N_1957);
or U7474 (N_7474,N_376,N_80);
and U7475 (N_7475,N_3651,N_4306);
nor U7476 (N_7476,N_2801,N_3520);
and U7477 (N_7477,N_2101,N_227);
nor U7478 (N_7478,N_3277,N_4502);
and U7479 (N_7479,N_74,N_4748);
and U7480 (N_7480,N_3903,N_3807);
nand U7481 (N_7481,N_1167,N_4322);
and U7482 (N_7482,N_2767,N_3549);
or U7483 (N_7483,N_2974,N_1489);
xnor U7484 (N_7484,N_1875,N_1546);
nand U7485 (N_7485,N_2953,N_3071);
xnor U7486 (N_7486,N_1522,N_3007);
xnor U7487 (N_7487,N_2670,N_2234);
and U7488 (N_7488,N_2784,N_4175);
xnor U7489 (N_7489,N_3098,N_3096);
and U7490 (N_7490,N_2700,N_486);
nand U7491 (N_7491,N_2054,N_3832);
or U7492 (N_7492,N_2958,N_3626);
nand U7493 (N_7493,N_4982,N_3561);
and U7494 (N_7494,N_1214,N_2186);
or U7495 (N_7495,N_4493,N_2541);
and U7496 (N_7496,N_4150,N_2594);
or U7497 (N_7497,N_1974,N_2001);
and U7498 (N_7498,N_1556,N_1595);
nand U7499 (N_7499,N_2867,N_4901);
xnor U7500 (N_7500,N_2470,N_3583);
nand U7501 (N_7501,N_4236,N_4546);
xnor U7502 (N_7502,N_1025,N_2425);
nor U7503 (N_7503,N_3780,N_2664);
xor U7504 (N_7504,N_640,N_2978);
or U7505 (N_7505,N_997,N_1044);
or U7506 (N_7506,N_4963,N_2410);
nand U7507 (N_7507,N_1748,N_4606);
nor U7508 (N_7508,N_3372,N_731);
nor U7509 (N_7509,N_3496,N_3749);
nor U7510 (N_7510,N_1663,N_3153);
nor U7511 (N_7511,N_2196,N_894);
or U7512 (N_7512,N_2283,N_2892);
nor U7513 (N_7513,N_4013,N_2612);
or U7514 (N_7514,N_2765,N_4744);
xnor U7515 (N_7515,N_2517,N_978);
nor U7516 (N_7516,N_3225,N_1355);
xor U7517 (N_7517,N_937,N_1907);
nor U7518 (N_7518,N_4232,N_1210);
and U7519 (N_7519,N_1113,N_2135);
nor U7520 (N_7520,N_1996,N_1840);
nand U7521 (N_7521,N_1235,N_4025);
or U7522 (N_7522,N_4472,N_1691);
nand U7523 (N_7523,N_4339,N_1689);
nand U7524 (N_7524,N_4499,N_1026);
nor U7525 (N_7525,N_625,N_489);
or U7526 (N_7526,N_4109,N_2449);
and U7527 (N_7527,N_2900,N_4804);
or U7528 (N_7528,N_1418,N_1920);
nor U7529 (N_7529,N_1150,N_3545);
nor U7530 (N_7530,N_885,N_2199);
xor U7531 (N_7531,N_484,N_3063);
nand U7532 (N_7532,N_1464,N_3007);
nor U7533 (N_7533,N_3674,N_2464);
nor U7534 (N_7534,N_1654,N_841);
or U7535 (N_7535,N_1906,N_4230);
and U7536 (N_7536,N_705,N_4449);
or U7537 (N_7537,N_1479,N_4350);
nor U7538 (N_7538,N_2331,N_2774);
nand U7539 (N_7539,N_2270,N_827);
nor U7540 (N_7540,N_709,N_2127);
nor U7541 (N_7541,N_4478,N_1088);
nor U7542 (N_7542,N_4830,N_3872);
nor U7543 (N_7543,N_2256,N_2299);
nand U7544 (N_7544,N_1563,N_4923);
nor U7545 (N_7545,N_2633,N_140);
or U7546 (N_7546,N_1158,N_1049);
and U7547 (N_7547,N_3766,N_467);
and U7548 (N_7548,N_286,N_601);
and U7549 (N_7549,N_1883,N_2109);
or U7550 (N_7550,N_1084,N_4902);
nand U7551 (N_7551,N_4509,N_4920);
nor U7552 (N_7552,N_740,N_546);
xor U7553 (N_7553,N_610,N_1703);
nor U7554 (N_7554,N_3491,N_1988);
xor U7555 (N_7555,N_280,N_4860);
nand U7556 (N_7556,N_1671,N_3469);
nor U7557 (N_7557,N_2048,N_2909);
xor U7558 (N_7558,N_1776,N_3492);
and U7559 (N_7559,N_1214,N_447);
nor U7560 (N_7560,N_4486,N_1547);
nor U7561 (N_7561,N_553,N_4539);
and U7562 (N_7562,N_1392,N_3331);
nor U7563 (N_7563,N_1721,N_4279);
xnor U7564 (N_7564,N_1806,N_4226);
or U7565 (N_7565,N_2089,N_1435);
nor U7566 (N_7566,N_2913,N_3891);
nand U7567 (N_7567,N_86,N_868);
and U7568 (N_7568,N_641,N_313);
nand U7569 (N_7569,N_810,N_965);
or U7570 (N_7570,N_1978,N_4304);
nand U7571 (N_7571,N_2552,N_2716);
nand U7572 (N_7572,N_3554,N_2573);
and U7573 (N_7573,N_1388,N_3358);
nor U7574 (N_7574,N_2424,N_4043);
and U7575 (N_7575,N_4263,N_3918);
nand U7576 (N_7576,N_873,N_4123);
nand U7577 (N_7577,N_2889,N_2325);
xor U7578 (N_7578,N_1701,N_4857);
nor U7579 (N_7579,N_175,N_2266);
or U7580 (N_7580,N_1115,N_4194);
xor U7581 (N_7581,N_785,N_3934);
or U7582 (N_7582,N_3677,N_667);
or U7583 (N_7583,N_1569,N_3279);
nor U7584 (N_7584,N_1815,N_3312);
or U7585 (N_7585,N_190,N_1165);
nor U7586 (N_7586,N_4716,N_1157);
xnor U7587 (N_7587,N_4161,N_2690);
nand U7588 (N_7588,N_481,N_3772);
and U7589 (N_7589,N_2398,N_1408);
and U7590 (N_7590,N_3534,N_4061);
xnor U7591 (N_7591,N_1217,N_2468);
nand U7592 (N_7592,N_1835,N_2179);
nand U7593 (N_7593,N_3064,N_1927);
nand U7594 (N_7594,N_2433,N_1999);
and U7595 (N_7595,N_757,N_45);
or U7596 (N_7596,N_144,N_3293);
or U7597 (N_7597,N_3989,N_577);
or U7598 (N_7598,N_3741,N_3949);
and U7599 (N_7599,N_552,N_4989);
and U7600 (N_7600,N_2719,N_562);
nand U7601 (N_7601,N_4808,N_720);
xnor U7602 (N_7602,N_4908,N_3225);
and U7603 (N_7603,N_4188,N_4217);
nor U7604 (N_7604,N_1412,N_2664);
nand U7605 (N_7605,N_845,N_1255);
or U7606 (N_7606,N_660,N_3767);
xnor U7607 (N_7607,N_2874,N_4699);
or U7608 (N_7608,N_723,N_4648);
and U7609 (N_7609,N_697,N_1881);
nand U7610 (N_7610,N_4086,N_1918);
and U7611 (N_7611,N_3652,N_441);
and U7612 (N_7612,N_2572,N_3436);
and U7613 (N_7613,N_618,N_3304);
xor U7614 (N_7614,N_3687,N_2546);
nand U7615 (N_7615,N_778,N_4626);
and U7616 (N_7616,N_2912,N_2645);
nor U7617 (N_7617,N_1178,N_3574);
nor U7618 (N_7618,N_4675,N_4478);
nor U7619 (N_7619,N_3879,N_4649);
and U7620 (N_7620,N_407,N_4194);
nor U7621 (N_7621,N_2398,N_1435);
xnor U7622 (N_7622,N_1728,N_2880);
or U7623 (N_7623,N_847,N_4179);
nor U7624 (N_7624,N_1153,N_506);
xnor U7625 (N_7625,N_3826,N_319);
xnor U7626 (N_7626,N_2121,N_3056);
xnor U7627 (N_7627,N_431,N_2609);
or U7628 (N_7628,N_1523,N_4285);
nor U7629 (N_7629,N_1392,N_653);
or U7630 (N_7630,N_1545,N_241);
nand U7631 (N_7631,N_4993,N_1139);
nand U7632 (N_7632,N_623,N_3730);
nor U7633 (N_7633,N_4432,N_4158);
nand U7634 (N_7634,N_2450,N_2345);
and U7635 (N_7635,N_3000,N_3324);
and U7636 (N_7636,N_3728,N_3524);
xnor U7637 (N_7637,N_2750,N_821);
or U7638 (N_7638,N_1135,N_4296);
nor U7639 (N_7639,N_1664,N_4622);
or U7640 (N_7640,N_778,N_2637);
xor U7641 (N_7641,N_4925,N_630);
nor U7642 (N_7642,N_548,N_4953);
nand U7643 (N_7643,N_1159,N_880);
nor U7644 (N_7644,N_4161,N_4273);
xor U7645 (N_7645,N_4581,N_764);
or U7646 (N_7646,N_1148,N_2765);
and U7647 (N_7647,N_1055,N_4527);
xnor U7648 (N_7648,N_2122,N_1990);
or U7649 (N_7649,N_1750,N_3840);
and U7650 (N_7650,N_453,N_3542);
nand U7651 (N_7651,N_1203,N_861);
or U7652 (N_7652,N_3388,N_3355);
and U7653 (N_7653,N_4794,N_1363);
xor U7654 (N_7654,N_1363,N_4949);
and U7655 (N_7655,N_200,N_4261);
and U7656 (N_7656,N_2422,N_3103);
or U7657 (N_7657,N_1689,N_323);
or U7658 (N_7658,N_2122,N_4877);
nand U7659 (N_7659,N_4326,N_2071);
nand U7660 (N_7660,N_826,N_4274);
and U7661 (N_7661,N_4953,N_3175);
and U7662 (N_7662,N_1887,N_4777);
nor U7663 (N_7663,N_2392,N_973);
nor U7664 (N_7664,N_940,N_4930);
xor U7665 (N_7665,N_4926,N_1100);
and U7666 (N_7666,N_2001,N_1352);
or U7667 (N_7667,N_967,N_3492);
or U7668 (N_7668,N_1543,N_555);
xor U7669 (N_7669,N_2345,N_3986);
nor U7670 (N_7670,N_1787,N_4064);
or U7671 (N_7671,N_2918,N_2946);
or U7672 (N_7672,N_4921,N_2194);
and U7673 (N_7673,N_3772,N_6);
or U7674 (N_7674,N_1291,N_4020);
and U7675 (N_7675,N_1861,N_2787);
nand U7676 (N_7676,N_3688,N_1540);
nor U7677 (N_7677,N_2648,N_226);
or U7678 (N_7678,N_1831,N_3044);
or U7679 (N_7679,N_854,N_114);
and U7680 (N_7680,N_2389,N_4321);
and U7681 (N_7681,N_1125,N_4189);
and U7682 (N_7682,N_1453,N_1858);
nor U7683 (N_7683,N_4834,N_922);
and U7684 (N_7684,N_739,N_1398);
nor U7685 (N_7685,N_2725,N_2166);
or U7686 (N_7686,N_4466,N_1726);
nor U7687 (N_7687,N_3328,N_537);
nor U7688 (N_7688,N_2194,N_4436);
xor U7689 (N_7689,N_508,N_183);
nor U7690 (N_7690,N_3304,N_4314);
and U7691 (N_7691,N_1190,N_4568);
and U7692 (N_7692,N_2376,N_3505);
or U7693 (N_7693,N_2673,N_3648);
nor U7694 (N_7694,N_1958,N_3336);
nor U7695 (N_7695,N_4416,N_2491);
and U7696 (N_7696,N_3107,N_82);
nand U7697 (N_7697,N_1813,N_1820);
nor U7698 (N_7698,N_803,N_647);
or U7699 (N_7699,N_1968,N_3036);
and U7700 (N_7700,N_2798,N_4361);
nor U7701 (N_7701,N_4173,N_3881);
nand U7702 (N_7702,N_1810,N_4747);
or U7703 (N_7703,N_1914,N_4144);
nand U7704 (N_7704,N_3412,N_4003);
nor U7705 (N_7705,N_662,N_4273);
xnor U7706 (N_7706,N_4768,N_3536);
or U7707 (N_7707,N_3208,N_2086);
and U7708 (N_7708,N_1320,N_2320);
nand U7709 (N_7709,N_4910,N_993);
xor U7710 (N_7710,N_4693,N_2530);
nor U7711 (N_7711,N_1487,N_3442);
nor U7712 (N_7712,N_4503,N_641);
or U7713 (N_7713,N_1605,N_4763);
or U7714 (N_7714,N_562,N_796);
xnor U7715 (N_7715,N_4519,N_2017);
or U7716 (N_7716,N_2540,N_3403);
or U7717 (N_7717,N_2899,N_310);
or U7718 (N_7718,N_158,N_4240);
and U7719 (N_7719,N_3872,N_3000);
and U7720 (N_7720,N_3872,N_2580);
and U7721 (N_7721,N_3634,N_4155);
and U7722 (N_7722,N_2032,N_3693);
xnor U7723 (N_7723,N_2182,N_611);
or U7724 (N_7724,N_823,N_2441);
nor U7725 (N_7725,N_4915,N_3173);
nand U7726 (N_7726,N_555,N_1851);
nor U7727 (N_7727,N_656,N_3662);
nand U7728 (N_7728,N_2755,N_3410);
nor U7729 (N_7729,N_3524,N_1829);
nand U7730 (N_7730,N_1761,N_1943);
nor U7731 (N_7731,N_2399,N_2056);
or U7732 (N_7732,N_2556,N_639);
and U7733 (N_7733,N_776,N_2773);
or U7734 (N_7734,N_1999,N_1416);
xor U7735 (N_7735,N_2699,N_4065);
or U7736 (N_7736,N_2548,N_4116);
or U7737 (N_7737,N_2266,N_3066);
or U7738 (N_7738,N_4238,N_156);
and U7739 (N_7739,N_4463,N_2137);
nand U7740 (N_7740,N_3978,N_3984);
nor U7741 (N_7741,N_744,N_2935);
nor U7742 (N_7742,N_576,N_2498);
and U7743 (N_7743,N_4873,N_1124);
xor U7744 (N_7744,N_1496,N_330);
and U7745 (N_7745,N_2467,N_284);
nand U7746 (N_7746,N_1897,N_110);
nor U7747 (N_7747,N_402,N_3149);
and U7748 (N_7748,N_4175,N_2329);
nand U7749 (N_7749,N_2825,N_1315);
nor U7750 (N_7750,N_1767,N_3672);
nand U7751 (N_7751,N_3670,N_416);
nand U7752 (N_7752,N_2413,N_485);
and U7753 (N_7753,N_419,N_3427);
nor U7754 (N_7754,N_1631,N_4353);
xnor U7755 (N_7755,N_4386,N_2430);
xnor U7756 (N_7756,N_2912,N_2126);
or U7757 (N_7757,N_3986,N_3664);
nand U7758 (N_7758,N_4684,N_1244);
xor U7759 (N_7759,N_270,N_1074);
or U7760 (N_7760,N_2984,N_4650);
and U7761 (N_7761,N_3177,N_255);
and U7762 (N_7762,N_2701,N_86);
nor U7763 (N_7763,N_2920,N_3869);
nand U7764 (N_7764,N_1434,N_4072);
and U7765 (N_7765,N_809,N_2632);
and U7766 (N_7766,N_3213,N_4476);
nor U7767 (N_7767,N_690,N_2327);
nand U7768 (N_7768,N_3123,N_3961);
nor U7769 (N_7769,N_1576,N_2885);
or U7770 (N_7770,N_1928,N_1200);
nor U7771 (N_7771,N_2421,N_4234);
xor U7772 (N_7772,N_2984,N_4700);
or U7773 (N_7773,N_2720,N_1532);
or U7774 (N_7774,N_2182,N_839);
or U7775 (N_7775,N_3765,N_1629);
xor U7776 (N_7776,N_590,N_4861);
nor U7777 (N_7777,N_3214,N_3697);
and U7778 (N_7778,N_516,N_328);
and U7779 (N_7779,N_2603,N_1733);
xor U7780 (N_7780,N_1422,N_4784);
or U7781 (N_7781,N_3895,N_3892);
nand U7782 (N_7782,N_200,N_3447);
xor U7783 (N_7783,N_1404,N_2133);
or U7784 (N_7784,N_2501,N_3572);
nor U7785 (N_7785,N_4915,N_392);
nor U7786 (N_7786,N_3528,N_4291);
and U7787 (N_7787,N_1348,N_4020);
or U7788 (N_7788,N_3166,N_491);
nand U7789 (N_7789,N_2159,N_2358);
or U7790 (N_7790,N_3103,N_1964);
or U7791 (N_7791,N_3166,N_3586);
xnor U7792 (N_7792,N_1387,N_4819);
xor U7793 (N_7793,N_3757,N_197);
nand U7794 (N_7794,N_1540,N_4439);
and U7795 (N_7795,N_2268,N_1491);
xnor U7796 (N_7796,N_4470,N_3867);
and U7797 (N_7797,N_2300,N_2182);
xor U7798 (N_7798,N_81,N_3168);
nand U7799 (N_7799,N_2552,N_2693);
nand U7800 (N_7800,N_4944,N_1849);
nand U7801 (N_7801,N_2399,N_3825);
nor U7802 (N_7802,N_2369,N_3773);
xor U7803 (N_7803,N_2165,N_3060);
nor U7804 (N_7804,N_2365,N_3629);
nand U7805 (N_7805,N_3418,N_166);
or U7806 (N_7806,N_660,N_1798);
xnor U7807 (N_7807,N_665,N_3303);
nand U7808 (N_7808,N_3807,N_1768);
xor U7809 (N_7809,N_402,N_716);
xnor U7810 (N_7810,N_3996,N_3965);
nor U7811 (N_7811,N_2175,N_3215);
and U7812 (N_7812,N_3340,N_4482);
or U7813 (N_7813,N_254,N_2876);
nand U7814 (N_7814,N_4564,N_1250);
nand U7815 (N_7815,N_2515,N_1773);
xnor U7816 (N_7816,N_1456,N_3701);
nor U7817 (N_7817,N_3638,N_977);
and U7818 (N_7818,N_24,N_2000);
nand U7819 (N_7819,N_3621,N_308);
nand U7820 (N_7820,N_3815,N_4307);
nor U7821 (N_7821,N_4056,N_436);
xor U7822 (N_7822,N_1219,N_2276);
xnor U7823 (N_7823,N_4140,N_4399);
nand U7824 (N_7824,N_1872,N_4930);
and U7825 (N_7825,N_4783,N_3370);
xor U7826 (N_7826,N_539,N_4199);
or U7827 (N_7827,N_4893,N_1321);
or U7828 (N_7828,N_2408,N_2026);
nor U7829 (N_7829,N_1401,N_3202);
and U7830 (N_7830,N_2694,N_2539);
nor U7831 (N_7831,N_824,N_1809);
nand U7832 (N_7832,N_3929,N_2308);
and U7833 (N_7833,N_3967,N_4191);
nor U7834 (N_7834,N_2458,N_1132);
xor U7835 (N_7835,N_1403,N_1628);
nand U7836 (N_7836,N_437,N_526);
or U7837 (N_7837,N_3328,N_2715);
and U7838 (N_7838,N_246,N_3282);
or U7839 (N_7839,N_3152,N_4876);
and U7840 (N_7840,N_771,N_4023);
nor U7841 (N_7841,N_59,N_1147);
nor U7842 (N_7842,N_3591,N_1174);
nand U7843 (N_7843,N_3018,N_2572);
nand U7844 (N_7844,N_1018,N_3926);
nand U7845 (N_7845,N_25,N_4020);
nand U7846 (N_7846,N_3902,N_1463);
nor U7847 (N_7847,N_4184,N_1557);
nand U7848 (N_7848,N_3801,N_4734);
and U7849 (N_7849,N_3395,N_4724);
xnor U7850 (N_7850,N_510,N_3204);
xnor U7851 (N_7851,N_4436,N_4165);
nand U7852 (N_7852,N_1210,N_1538);
or U7853 (N_7853,N_2163,N_3186);
and U7854 (N_7854,N_3339,N_487);
and U7855 (N_7855,N_3025,N_4796);
and U7856 (N_7856,N_1719,N_2308);
and U7857 (N_7857,N_4856,N_1716);
and U7858 (N_7858,N_581,N_2140);
or U7859 (N_7859,N_757,N_238);
nand U7860 (N_7860,N_1410,N_4179);
and U7861 (N_7861,N_1041,N_2867);
or U7862 (N_7862,N_2497,N_3089);
and U7863 (N_7863,N_2477,N_3439);
nor U7864 (N_7864,N_882,N_2640);
and U7865 (N_7865,N_1300,N_2567);
nand U7866 (N_7866,N_4021,N_4391);
or U7867 (N_7867,N_813,N_1573);
nand U7868 (N_7868,N_1711,N_1146);
nand U7869 (N_7869,N_3914,N_4909);
nor U7870 (N_7870,N_2982,N_97);
nand U7871 (N_7871,N_699,N_1155);
nand U7872 (N_7872,N_967,N_2940);
or U7873 (N_7873,N_3024,N_595);
and U7874 (N_7874,N_4433,N_3706);
and U7875 (N_7875,N_950,N_827);
nor U7876 (N_7876,N_1832,N_1136);
nor U7877 (N_7877,N_1648,N_4546);
or U7878 (N_7878,N_1495,N_144);
or U7879 (N_7879,N_4438,N_3027);
and U7880 (N_7880,N_764,N_1791);
nand U7881 (N_7881,N_3665,N_986);
xnor U7882 (N_7882,N_661,N_1010);
nor U7883 (N_7883,N_4612,N_3366);
and U7884 (N_7884,N_1847,N_484);
and U7885 (N_7885,N_4260,N_4751);
nor U7886 (N_7886,N_58,N_518);
and U7887 (N_7887,N_4695,N_4600);
nor U7888 (N_7888,N_1722,N_1628);
or U7889 (N_7889,N_188,N_4542);
or U7890 (N_7890,N_1769,N_3857);
xnor U7891 (N_7891,N_2057,N_2007);
nand U7892 (N_7892,N_3338,N_1149);
nand U7893 (N_7893,N_3351,N_2766);
nor U7894 (N_7894,N_3269,N_3962);
nand U7895 (N_7895,N_4513,N_4219);
and U7896 (N_7896,N_2589,N_986);
xor U7897 (N_7897,N_2106,N_3546);
and U7898 (N_7898,N_2358,N_2354);
or U7899 (N_7899,N_2296,N_160);
nor U7900 (N_7900,N_4315,N_386);
nor U7901 (N_7901,N_4079,N_2493);
or U7902 (N_7902,N_4642,N_4713);
and U7903 (N_7903,N_1214,N_2102);
and U7904 (N_7904,N_4837,N_869);
nand U7905 (N_7905,N_144,N_751);
or U7906 (N_7906,N_3517,N_208);
nand U7907 (N_7907,N_218,N_1762);
and U7908 (N_7908,N_2900,N_248);
xor U7909 (N_7909,N_908,N_1896);
or U7910 (N_7910,N_996,N_1141);
nand U7911 (N_7911,N_4930,N_4395);
or U7912 (N_7912,N_1900,N_2978);
nor U7913 (N_7913,N_4727,N_4792);
nand U7914 (N_7914,N_1144,N_4623);
xnor U7915 (N_7915,N_4797,N_4902);
xor U7916 (N_7916,N_3665,N_4967);
nor U7917 (N_7917,N_2392,N_3316);
nand U7918 (N_7918,N_832,N_3736);
nand U7919 (N_7919,N_4744,N_3974);
xnor U7920 (N_7920,N_4072,N_2261);
nor U7921 (N_7921,N_1048,N_3785);
and U7922 (N_7922,N_2684,N_388);
xor U7923 (N_7923,N_4473,N_2325);
nor U7924 (N_7924,N_4841,N_4333);
nand U7925 (N_7925,N_4184,N_4846);
nand U7926 (N_7926,N_2489,N_3865);
xor U7927 (N_7927,N_2018,N_500);
or U7928 (N_7928,N_2615,N_4734);
and U7929 (N_7929,N_2077,N_1643);
xor U7930 (N_7930,N_2048,N_3764);
and U7931 (N_7931,N_532,N_3451);
nor U7932 (N_7932,N_4225,N_780);
or U7933 (N_7933,N_3079,N_1150);
and U7934 (N_7934,N_2033,N_2254);
nor U7935 (N_7935,N_4976,N_4294);
nor U7936 (N_7936,N_4875,N_4630);
xnor U7937 (N_7937,N_2250,N_4813);
or U7938 (N_7938,N_3214,N_915);
or U7939 (N_7939,N_3984,N_4867);
or U7940 (N_7940,N_214,N_968);
nand U7941 (N_7941,N_3428,N_2779);
nand U7942 (N_7942,N_2767,N_3632);
and U7943 (N_7943,N_4608,N_280);
nor U7944 (N_7944,N_1974,N_1441);
nor U7945 (N_7945,N_3145,N_2158);
or U7946 (N_7946,N_601,N_3086);
nor U7947 (N_7947,N_1232,N_1040);
nor U7948 (N_7948,N_4022,N_4838);
xor U7949 (N_7949,N_480,N_3212);
xor U7950 (N_7950,N_4801,N_695);
and U7951 (N_7951,N_3612,N_2109);
xor U7952 (N_7952,N_2489,N_2887);
nand U7953 (N_7953,N_2719,N_4482);
xnor U7954 (N_7954,N_2021,N_344);
or U7955 (N_7955,N_1617,N_3154);
xnor U7956 (N_7956,N_1280,N_4749);
or U7957 (N_7957,N_1847,N_4931);
nand U7958 (N_7958,N_3876,N_220);
nor U7959 (N_7959,N_3010,N_3480);
or U7960 (N_7960,N_2401,N_2425);
and U7961 (N_7961,N_4535,N_3927);
xnor U7962 (N_7962,N_3376,N_1848);
nand U7963 (N_7963,N_2343,N_1063);
and U7964 (N_7964,N_1564,N_4682);
nor U7965 (N_7965,N_4201,N_4904);
and U7966 (N_7966,N_376,N_791);
xnor U7967 (N_7967,N_130,N_2349);
and U7968 (N_7968,N_1220,N_276);
nand U7969 (N_7969,N_2657,N_3792);
nand U7970 (N_7970,N_2593,N_923);
nor U7971 (N_7971,N_4780,N_932);
xnor U7972 (N_7972,N_623,N_1197);
and U7973 (N_7973,N_4307,N_3476);
or U7974 (N_7974,N_3362,N_49);
nor U7975 (N_7975,N_1692,N_3816);
nor U7976 (N_7976,N_4463,N_685);
nand U7977 (N_7977,N_1054,N_4657);
or U7978 (N_7978,N_323,N_306);
nand U7979 (N_7979,N_2450,N_2247);
xor U7980 (N_7980,N_3730,N_3560);
nor U7981 (N_7981,N_2043,N_4678);
nor U7982 (N_7982,N_2437,N_235);
or U7983 (N_7983,N_3530,N_76);
xnor U7984 (N_7984,N_4717,N_4080);
nand U7985 (N_7985,N_2523,N_2807);
nor U7986 (N_7986,N_3213,N_3341);
or U7987 (N_7987,N_2947,N_1605);
or U7988 (N_7988,N_4809,N_335);
and U7989 (N_7989,N_1536,N_2016);
nor U7990 (N_7990,N_1911,N_2921);
and U7991 (N_7991,N_1484,N_2552);
xor U7992 (N_7992,N_2355,N_643);
nor U7993 (N_7993,N_2606,N_2247);
and U7994 (N_7994,N_4204,N_1064);
nor U7995 (N_7995,N_3882,N_3165);
and U7996 (N_7996,N_3888,N_4594);
and U7997 (N_7997,N_222,N_2831);
and U7998 (N_7998,N_1403,N_4715);
and U7999 (N_7999,N_282,N_4021);
nand U8000 (N_8000,N_2539,N_3875);
xor U8001 (N_8001,N_2290,N_3585);
nor U8002 (N_8002,N_3011,N_1368);
xor U8003 (N_8003,N_2565,N_4495);
xnor U8004 (N_8004,N_3154,N_2377);
nand U8005 (N_8005,N_269,N_2919);
nor U8006 (N_8006,N_3898,N_1049);
nand U8007 (N_8007,N_3809,N_2967);
and U8008 (N_8008,N_3173,N_3878);
or U8009 (N_8009,N_2156,N_4562);
xor U8010 (N_8010,N_4590,N_2410);
nor U8011 (N_8011,N_1398,N_2638);
xor U8012 (N_8012,N_1390,N_4983);
or U8013 (N_8013,N_4929,N_197);
and U8014 (N_8014,N_254,N_2810);
nor U8015 (N_8015,N_1497,N_4076);
nand U8016 (N_8016,N_3975,N_4185);
nor U8017 (N_8017,N_2905,N_4599);
or U8018 (N_8018,N_24,N_2631);
xor U8019 (N_8019,N_1921,N_4803);
nor U8020 (N_8020,N_654,N_2015);
and U8021 (N_8021,N_2906,N_1542);
xor U8022 (N_8022,N_1614,N_1227);
nand U8023 (N_8023,N_3172,N_2461);
or U8024 (N_8024,N_4438,N_2851);
and U8025 (N_8025,N_3994,N_1176);
and U8026 (N_8026,N_975,N_1994);
and U8027 (N_8027,N_301,N_3688);
nor U8028 (N_8028,N_2725,N_1764);
nor U8029 (N_8029,N_3289,N_901);
nand U8030 (N_8030,N_3670,N_1593);
and U8031 (N_8031,N_1819,N_3420);
xnor U8032 (N_8032,N_3289,N_1583);
and U8033 (N_8033,N_435,N_4959);
and U8034 (N_8034,N_3148,N_2895);
or U8035 (N_8035,N_1923,N_3651);
and U8036 (N_8036,N_1458,N_329);
or U8037 (N_8037,N_2216,N_762);
nor U8038 (N_8038,N_3986,N_292);
and U8039 (N_8039,N_1854,N_4499);
xnor U8040 (N_8040,N_3769,N_3095);
and U8041 (N_8041,N_3133,N_837);
and U8042 (N_8042,N_3248,N_2720);
xor U8043 (N_8043,N_1940,N_4872);
xnor U8044 (N_8044,N_3739,N_2577);
xnor U8045 (N_8045,N_382,N_4203);
and U8046 (N_8046,N_2666,N_3284);
or U8047 (N_8047,N_3022,N_879);
xnor U8048 (N_8048,N_4095,N_1894);
nand U8049 (N_8049,N_4557,N_3247);
nand U8050 (N_8050,N_2818,N_2935);
and U8051 (N_8051,N_2352,N_4358);
and U8052 (N_8052,N_3833,N_711);
and U8053 (N_8053,N_3927,N_471);
nor U8054 (N_8054,N_229,N_3932);
xor U8055 (N_8055,N_551,N_67);
xor U8056 (N_8056,N_2772,N_2003);
nand U8057 (N_8057,N_83,N_1917);
nand U8058 (N_8058,N_4917,N_4360);
or U8059 (N_8059,N_2319,N_2681);
xor U8060 (N_8060,N_3045,N_4);
or U8061 (N_8061,N_4890,N_1669);
or U8062 (N_8062,N_4316,N_4028);
nor U8063 (N_8063,N_572,N_4374);
or U8064 (N_8064,N_3490,N_2482);
xnor U8065 (N_8065,N_220,N_4059);
nand U8066 (N_8066,N_910,N_104);
nand U8067 (N_8067,N_4826,N_481);
or U8068 (N_8068,N_260,N_1291);
nor U8069 (N_8069,N_3604,N_1914);
nor U8070 (N_8070,N_2948,N_1808);
or U8071 (N_8071,N_81,N_1191);
nand U8072 (N_8072,N_4984,N_4051);
nand U8073 (N_8073,N_1571,N_2963);
or U8074 (N_8074,N_2132,N_1483);
nor U8075 (N_8075,N_2292,N_329);
xnor U8076 (N_8076,N_2461,N_3568);
and U8077 (N_8077,N_2934,N_4901);
and U8078 (N_8078,N_4695,N_229);
and U8079 (N_8079,N_1441,N_553);
nand U8080 (N_8080,N_2917,N_1556);
or U8081 (N_8081,N_391,N_665);
nor U8082 (N_8082,N_3292,N_2246);
xnor U8083 (N_8083,N_4935,N_1493);
and U8084 (N_8084,N_3546,N_199);
or U8085 (N_8085,N_3536,N_3890);
or U8086 (N_8086,N_4795,N_1642);
nand U8087 (N_8087,N_1739,N_1637);
and U8088 (N_8088,N_2648,N_2018);
nand U8089 (N_8089,N_4026,N_3470);
xnor U8090 (N_8090,N_1470,N_1344);
or U8091 (N_8091,N_3198,N_4523);
xor U8092 (N_8092,N_1903,N_2634);
nand U8093 (N_8093,N_3408,N_729);
and U8094 (N_8094,N_1758,N_3641);
and U8095 (N_8095,N_4295,N_637);
xor U8096 (N_8096,N_3432,N_1800);
and U8097 (N_8097,N_1691,N_1189);
nand U8098 (N_8098,N_3014,N_477);
nor U8099 (N_8099,N_3669,N_351);
and U8100 (N_8100,N_1547,N_3568);
xor U8101 (N_8101,N_517,N_581);
xnor U8102 (N_8102,N_1125,N_4956);
nor U8103 (N_8103,N_2955,N_1489);
xnor U8104 (N_8104,N_1902,N_1403);
and U8105 (N_8105,N_3295,N_3833);
and U8106 (N_8106,N_1219,N_4686);
nor U8107 (N_8107,N_4398,N_2437);
and U8108 (N_8108,N_1292,N_3723);
and U8109 (N_8109,N_3686,N_2686);
or U8110 (N_8110,N_475,N_4164);
nor U8111 (N_8111,N_2284,N_1574);
nand U8112 (N_8112,N_2199,N_606);
or U8113 (N_8113,N_4844,N_426);
nand U8114 (N_8114,N_4434,N_3520);
xor U8115 (N_8115,N_670,N_3987);
xor U8116 (N_8116,N_1058,N_3560);
nand U8117 (N_8117,N_4079,N_2343);
nand U8118 (N_8118,N_3732,N_2741);
or U8119 (N_8119,N_4880,N_3222);
or U8120 (N_8120,N_431,N_4645);
nand U8121 (N_8121,N_699,N_4628);
nor U8122 (N_8122,N_1998,N_1212);
xor U8123 (N_8123,N_690,N_1410);
nor U8124 (N_8124,N_3215,N_3389);
or U8125 (N_8125,N_331,N_2522);
nor U8126 (N_8126,N_899,N_4994);
or U8127 (N_8127,N_2530,N_1448);
or U8128 (N_8128,N_366,N_3431);
xor U8129 (N_8129,N_3174,N_2807);
nor U8130 (N_8130,N_4248,N_1048);
xor U8131 (N_8131,N_1661,N_3172);
xor U8132 (N_8132,N_4159,N_3310);
or U8133 (N_8133,N_271,N_3522);
and U8134 (N_8134,N_1184,N_4520);
xnor U8135 (N_8135,N_4681,N_3341);
nand U8136 (N_8136,N_157,N_3726);
xnor U8137 (N_8137,N_1842,N_1039);
and U8138 (N_8138,N_4203,N_187);
and U8139 (N_8139,N_48,N_4739);
or U8140 (N_8140,N_575,N_4319);
or U8141 (N_8141,N_3088,N_3296);
nor U8142 (N_8142,N_4544,N_3610);
or U8143 (N_8143,N_4219,N_3915);
and U8144 (N_8144,N_4900,N_4711);
or U8145 (N_8145,N_1861,N_4989);
nand U8146 (N_8146,N_3629,N_170);
or U8147 (N_8147,N_4387,N_439);
or U8148 (N_8148,N_4353,N_229);
and U8149 (N_8149,N_4828,N_3815);
xnor U8150 (N_8150,N_2972,N_221);
xor U8151 (N_8151,N_2974,N_2646);
or U8152 (N_8152,N_3390,N_4762);
xnor U8153 (N_8153,N_1443,N_1495);
or U8154 (N_8154,N_333,N_1471);
and U8155 (N_8155,N_4744,N_3671);
nor U8156 (N_8156,N_3433,N_926);
or U8157 (N_8157,N_3959,N_3697);
nor U8158 (N_8158,N_2938,N_2640);
and U8159 (N_8159,N_370,N_2015);
or U8160 (N_8160,N_4049,N_4295);
and U8161 (N_8161,N_1904,N_2273);
or U8162 (N_8162,N_2850,N_1746);
xor U8163 (N_8163,N_3124,N_1795);
nand U8164 (N_8164,N_2912,N_2465);
nand U8165 (N_8165,N_3882,N_3384);
or U8166 (N_8166,N_1030,N_4087);
xnor U8167 (N_8167,N_1616,N_935);
or U8168 (N_8168,N_4939,N_254);
or U8169 (N_8169,N_4386,N_1125);
xnor U8170 (N_8170,N_723,N_4991);
xor U8171 (N_8171,N_402,N_3703);
or U8172 (N_8172,N_2720,N_2706);
nand U8173 (N_8173,N_629,N_474);
nand U8174 (N_8174,N_3882,N_854);
and U8175 (N_8175,N_1594,N_404);
and U8176 (N_8176,N_3133,N_4866);
xor U8177 (N_8177,N_2820,N_3397);
xnor U8178 (N_8178,N_3544,N_2017);
and U8179 (N_8179,N_3348,N_2526);
or U8180 (N_8180,N_4906,N_3418);
or U8181 (N_8181,N_1127,N_3589);
nand U8182 (N_8182,N_2730,N_940);
and U8183 (N_8183,N_2127,N_4884);
or U8184 (N_8184,N_717,N_3078);
and U8185 (N_8185,N_4398,N_1843);
nor U8186 (N_8186,N_4398,N_243);
nand U8187 (N_8187,N_1656,N_448);
nand U8188 (N_8188,N_1822,N_283);
nand U8189 (N_8189,N_1311,N_3883);
nand U8190 (N_8190,N_2915,N_2571);
and U8191 (N_8191,N_3945,N_3967);
nor U8192 (N_8192,N_379,N_3009);
xor U8193 (N_8193,N_2085,N_1396);
xnor U8194 (N_8194,N_623,N_3083);
xor U8195 (N_8195,N_4333,N_4322);
nor U8196 (N_8196,N_2789,N_3187);
xor U8197 (N_8197,N_4386,N_3872);
or U8198 (N_8198,N_3702,N_4219);
and U8199 (N_8199,N_1423,N_4385);
nand U8200 (N_8200,N_968,N_2103);
xor U8201 (N_8201,N_1570,N_4844);
nand U8202 (N_8202,N_1625,N_1432);
or U8203 (N_8203,N_4009,N_2148);
nor U8204 (N_8204,N_307,N_479);
nand U8205 (N_8205,N_473,N_2317);
nor U8206 (N_8206,N_1757,N_3674);
or U8207 (N_8207,N_618,N_4139);
xor U8208 (N_8208,N_1600,N_3755);
or U8209 (N_8209,N_1920,N_59);
xnor U8210 (N_8210,N_1277,N_1189);
and U8211 (N_8211,N_4494,N_2382);
and U8212 (N_8212,N_820,N_3915);
nand U8213 (N_8213,N_2559,N_2952);
nor U8214 (N_8214,N_1338,N_1162);
xnor U8215 (N_8215,N_4589,N_4700);
xor U8216 (N_8216,N_2679,N_1451);
xnor U8217 (N_8217,N_4587,N_4378);
and U8218 (N_8218,N_869,N_110);
xor U8219 (N_8219,N_3877,N_3153);
nand U8220 (N_8220,N_4102,N_4407);
xnor U8221 (N_8221,N_4444,N_2259);
or U8222 (N_8222,N_856,N_181);
or U8223 (N_8223,N_2234,N_2969);
nor U8224 (N_8224,N_4346,N_2033);
and U8225 (N_8225,N_2684,N_2457);
and U8226 (N_8226,N_4482,N_309);
and U8227 (N_8227,N_425,N_3190);
nor U8228 (N_8228,N_1220,N_1936);
or U8229 (N_8229,N_945,N_3344);
and U8230 (N_8230,N_4238,N_59);
nand U8231 (N_8231,N_1545,N_4468);
or U8232 (N_8232,N_3509,N_2686);
nand U8233 (N_8233,N_4891,N_1770);
xor U8234 (N_8234,N_1377,N_4596);
and U8235 (N_8235,N_1725,N_4968);
nand U8236 (N_8236,N_3481,N_2773);
xor U8237 (N_8237,N_621,N_3822);
or U8238 (N_8238,N_3900,N_4300);
xor U8239 (N_8239,N_4426,N_4757);
xnor U8240 (N_8240,N_737,N_2146);
or U8241 (N_8241,N_4300,N_3492);
xor U8242 (N_8242,N_1287,N_3865);
and U8243 (N_8243,N_4312,N_1792);
or U8244 (N_8244,N_629,N_537);
xor U8245 (N_8245,N_1534,N_2297);
or U8246 (N_8246,N_4007,N_836);
nand U8247 (N_8247,N_4617,N_315);
and U8248 (N_8248,N_1314,N_4126);
xor U8249 (N_8249,N_489,N_1922);
or U8250 (N_8250,N_1575,N_3179);
and U8251 (N_8251,N_1343,N_2463);
xor U8252 (N_8252,N_2075,N_602);
or U8253 (N_8253,N_1828,N_1545);
or U8254 (N_8254,N_2682,N_1958);
nand U8255 (N_8255,N_3406,N_409);
nand U8256 (N_8256,N_362,N_3807);
or U8257 (N_8257,N_2058,N_3428);
nor U8258 (N_8258,N_3941,N_1558);
xnor U8259 (N_8259,N_658,N_2359);
nand U8260 (N_8260,N_1797,N_4283);
and U8261 (N_8261,N_129,N_1129);
or U8262 (N_8262,N_3522,N_3654);
xor U8263 (N_8263,N_1646,N_712);
and U8264 (N_8264,N_905,N_4421);
or U8265 (N_8265,N_3831,N_1461);
or U8266 (N_8266,N_1526,N_2321);
nand U8267 (N_8267,N_3492,N_814);
or U8268 (N_8268,N_362,N_1468);
nor U8269 (N_8269,N_2816,N_3823);
or U8270 (N_8270,N_601,N_3375);
nor U8271 (N_8271,N_4961,N_141);
or U8272 (N_8272,N_3560,N_3054);
nand U8273 (N_8273,N_2589,N_4336);
nor U8274 (N_8274,N_194,N_4705);
nor U8275 (N_8275,N_1148,N_513);
nor U8276 (N_8276,N_226,N_3732);
and U8277 (N_8277,N_954,N_4177);
nor U8278 (N_8278,N_4347,N_2954);
nand U8279 (N_8279,N_3001,N_1061);
xor U8280 (N_8280,N_1440,N_1133);
nand U8281 (N_8281,N_18,N_2146);
nor U8282 (N_8282,N_727,N_44);
nor U8283 (N_8283,N_2220,N_604);
nor U8284 (N_8284,N_839,N_2382);
nor U8285 (N_8285,N_4285,N_1649);
nand U8286 (N_8286,N_4440,N_1042);
or U8287 (N_8287,N_1627,N_2757);
and U8288 (N_8288,N_3895,N_1129);
nor U8289 (N_8289,N_3870,N_36);
and U8290 (N_8290,N_4878,N_3844);
xor U8291 (N_8291,N_219,N_235);
or U8292 (N_8292,N_2508,N_4481);
nand U8293 (N_8293,N_3639,N_2831);
xnor U8294 (N_8294,N_3020,N_4185);
xnor U8295 (N_8295,N_2261,N_1527);
and U8296 (N_8296,N_1139,N_4555);
and U8297 (N_8297,N_2365,N_4706);
xnor U8298 (N_8298,N_2054,N_2917);
and U8299 (N_8299,N_4423,N_3038);
and U8300 (N_8300,N_1862,N_594);
nand U8301 (N_8301,N_1624,N_58);
and U8302 (N_8302,N_2864,N_848);
nor U8303 (N_8303,N_741,N_3096);
nor U8304 (N_8304,N_4838,N_1035);
or U8305 (N_8305,N_4087,N_3711);
xor U8306 (N_8306,N_537,N_1765);
and U8307 (N_8307,N_2890,N_3556);
or U8308 (N_8308,N_4690,N_1399);
xor U8309 (N_8309,N_4980,N_4963);
nor U8310 (N_8310,N_4577,N_2771);
xnor U8311 (N_8311,N_1537,N_2952);
and U8312 (N_8312,N_2540,N_521);
nand U8313 (N_8313,N_109,N_113);
or U8314 (N_8314,N_1267,N_450);
or U8315 (N_8315,N_2375,N_3494);
nor U8316 (N_8316,N_4930,N_2933);
and U8317 (N_8317,N_4645,N_2507);
nand U8318 (N_8318,N_2359,N_925);
nor U8319 (N_8319,N_68,N_4969);
xor U8320 (N_8320,N_3601,N_1861);
nor U8321 (N_8321,N_203,N_3366);
and U8322 (N_8322,N_1539,N_4868);
nand U8323 (N_8323,N_997,N_4032);
nand U8324 (N_8324,N_4960,N_3750);
nor U8325 (N_8325,N_289,N_4085);
xor U8326 (N_8326,N_2527,N_2035);
xnor U8327 (N_8327,N_1273,N_1938);
and U8328 (N_8328,N_147,N_1547);
nand U8329 (N_8329,N_2981,N_3792);
and U8330 (N_8330,N_3460,N_1782);
and U8331 (N_8331,N_3685,N_3038);
and U8332 (N_8332,N_440,N_2930);
xor U8333 (N_8333,N_3856,N_1089);
and U8334 (N_8334,N_2872,N_4525);
nand U8335 (N_8335,N_4434,N_2173);
nand U8336 (N_8336,N_793,N_1178);
nand U8337 (N_8337,N_1843,N_3200);
nor U8338 (N_8338,N_2636,N_960);
or U8339 (N_8339,N_3541,N_2702);
or U8340 (N_8340,N_776,N_4966);
xnor U8341 (N_8341,N_2697,N_4382);
or U8342 (N_8342,N_1677,N_4514);
nor U8343 (N_8343,N_2188,N_1001);
or U8344 (N_8344,N_1567,N_4297);
nor U8345 (N_8345,N_1517,N_3691);
nand U8346 (N_8346,N_1450,N_1273);
and U8347 (N_8347,N_934,N_4672);
xor U8348 (N_8348,N_2787,N_4139);
nor U8349 (N_8349,N_1201,N_2537);
or U8350 (N_8350,N_191,N_3115);
nand U8351 (N_8351,N_381,N_584);
or U8352 (N_8352,N_1015,N_1429);
or U8353 (N_8353,N_633,N_3579);
nor U8354 (N_8354,N_3026,N_197);
nand U8355 (N_8355,N_3147,N_4854);
or U8356 (N_8356,N_2099,N_2059);
xnor U8357 (N_8357,N_1044,N_1020);
and U8358 (N_8358,N_4628,N_407);
or U8359 (N_8359,N_882,N_572);
and U8360 (N_8360,N_35,N_3320);
nor U8361 (N_8361,N_2486,N_4906);
or U8362 (N_8362,N_1097,N_2474);
nor U8363 (N_8363,N_2494,N_4059);
xor U8364 (N_8364,N_675,N_4916);
nor U8365 (N_8365,N_766,N_4471);
xnor U8366 (N_8366,N_708,N_1609);
nor U8367 (N_8367,N_3513,N_2081);
nor U8368 (N_8368,N_4918,N_4);
nor U8369 (N_8369,N_1251,N_1010);
xnor U8370 (N_8370,N_144,N_3902);
xnor U8371 (N_8371,N_1453,N_1741);
nor U8372 (N_8372,N_2048,N_916);
nand U8373 (N_8373,N_1757,N_985);
or U8374 (N_8374,N_1273,N_3368);
and U8375 (N_8375,N_1995,N_459);
nor U8376 (N_8376,N_1819,N_2760);
xor U8377 (N_8377,N_4819,N_2887);
nand U8378 (N_8378,N_3997,N_441);
nand U8379 (N_8379,N_2509,N_4189);
xor U8380 (N_8380,N_1164,N_1978);
nand U8381 (N_8381,N_2174,N_251);
or U8382 (N_8382,N_4950,N_2929);
nor U8383 (N_8383,N_1823,N_2145);
nor U8384 (N_8384,N_2222,N_1512);
xor U8385 (N_8385,N_1036,N_1804);
or U8386 (N_8386,N_2342,N_3223);
nand U8387 (N_8387,N_1671,N_3588);
nor U8388 (N_8388,N_3520,N_2623);
xnor U8389 (N_8389,N_1258,N_2940);
xnor U8390 (N_8390,N_511,N_3427);
xor U8391 (N_8391,N_168,N_2150);
and U8392 (N_8392,N_4271,N_4010);
and U8393 (N_8393,N_2425,N_1495);
nand U8394 (N_8394,N_3132,N_3256);
and U8395 (N_8395,N_4754,N_2545);
nor U8396 (N_8396,N_4174,N_3125);
and U8397 (N_8397,N_1869,N_3118);
xor U8398 (N_8398,N_179,N_287);
and U8399 (N_8399,N_3750,N_3359);
and U8400 (N_8400,N_3368,N_4440);
nand U8401 (N_8401,N_1013,N_163);
xor U8402 (N_8402,N_608,N_407);
nand U8403 (N_8403,N_3647,N_3373);
nor U8404 (N_8404,N_4055,N_4362);
xor U8405 (N_8405,N_290,N_3333);
and U8406 (N_8406,N_2612,N_3385);
nand U8407 (N_8407,N_182,N_3150);
nor U8408 (N_8408,N_1850,N_122);
or U8409 (N_8409,N_354,N_4190);
and U8410 (N_8410,N_4723,N_4009);
and U8411 (N_8411,N_4338,N_390);
nand U8412 (N_8412,N_2062,N_2459);
nand U8413 (N_8413,N_2382,N_3792);
nor U8414 (N_8414,N_3592,N_2202);
and U8415 (N_8415,N_4836,N_1165);
xor U8416 (N_8416,N_2717,N_2734);
or U8417 (N_8417,N_2314,N_2453);
or U8418 (N_8418,N_2934,N_3776);
nand U8419 (N_8419,N_4993,N_2630);
xor U8420 (N_8420,N_3024,N_3727);
nand U8421 (N_8421,N_864,N_931);
nand U8422 (N_8422,N_2571,N_2759);
xnor U8423 (N_8423,N_4398,N_4502);
or U8424 (N_8424,N_1920,N_2708);
xor U8425 (N_8425,N_1210,N_1222);
and U8426 (N_8426,N_936,N_3201);
nor U8427 (N_8427,N_3396,N_4965);
xnor U8428 (N_8428,N_3100,N_4475);
and U8429 (N_8429,N_835,N_4832);
or U8430 (N_8430,N_4526,N_2878);
or U8431 (N_8431,N_1918,N_2187);
nand U8432 (N_8432,N_4032,N_961);
nor U8433 (N_8433,N_1127,N_3146);
nor U8434 (N_8434,N_4978,N_3428);
nand U8435 (N_8435,N_3264,N_4266);
xnor U8436 (N_8436,N_888,N_702);
nor U8437 (N_8437,N_4062,N_3619);
nand U8438 (N_8438,N_1094,N_1203);
nand U8439 (N_8439,N_1230,N_1745);
and U8440 (N_8440,N_4091,N_3652);
nand U8441 (N_8441,N_2724,N_3139);
xor U8442 (N_8442,N_4396,N_3580);
or U8443 (N_8443,N_215,N_541);
nor U8444 (N_8444,N_4295,N_3014);
or U8445 (N_8445,N_494,N_4220);
xnor U8446 (N_8446,N_468,N_149);
or U8447 (N_8447,N_4523,N_4307);
and U8448 (N_8448,N_117,N_1690);
and U8449 (N_8449,N_2140,N_3389);
nand U8450 (N_8450,N_4850,N_2615);
and U8451 (N_8451,N_4489,N_832);
xnor U8452 (N_8452,N_2369,N_799);
xnor U8453 (N_8453,N_225,N_3427);
xnor U8454 (N_8454,N_3196,N_2964);
nor U8455 (N_8455,N_465,N_1172);
or U8456 (N_8456,N_1999,N_316);
and U8457 (N_8457,N_4452,N_2018);
or U8458 (N_8458,N_705,N_3715);
xnor U8459 (N_8459,N_1550,N_489);
and U8460 (N_8460,N_926,N_532);
xnor U8461 (N_8461,N_1224,N_1951);
xor U8462 (N_8462,N_540,N_237);
or U8463 (N_8463,N_2645,N_4749);
nand U8464 (N_8464,N_2251,N_3841);
nand U8465 (N_8465,N_1199,N_1840);
or U8466 (N_8466,N_2659,N_276);
nor U8467 (N_8467,N_2025,N_4880);
xnor U8468 (N_8468,N_1216,N_4472);
or U8469 (N_8469,N_1895,N_12);
nor U8470 (N_8470,N_2527,N_434);
xor U8471 (N_8471,N_2298,N_4217);
or U8472 (N_8472,N_2683,N_838);
or U8473 (N_8473,N_3074,N_3556);
nor U8474 (N_8474,N_689,N_3663);
xnor U8475 (N_8475,N_4122,N_4707);
and U8476 (N_8476,N_3495,N_2017);
or U8477 (N_8477,N_741,N_262);
and U8478 (N_8478,N_2437,N_3625);
and U8479 (N_8479,N_2851,N_2221);
xor U8480 (N_8480,N_833,N_2181);
xnor U8481 (N_8481,N_3553,N_4232);
or U8482 (N_8482,N_4020,N_4855);
or U8483 (N_8483,N_873,N_1532);
and U8484 (N_8484,N_3021,N_3368);
nand U8485 (N_8485,N_3138,N_3601);
nor U8486 (N_8486,N_2368,N_4763);
nand U8487 (N_8487,N_1137,N_998);
xor U8488 (N_8488,N_1076,N_113);
or U8489 (N_8489,N_1342,N_1552);
xor U8490 (N_8490,N_1863,N_3627);
and U8491 (N_8491,N_3045,N_4199);
nor U8492 (N_8492,N_4633,N_4191);
nand U8493 (N_8493,N_41,N_4321);
or U8494 (N_8494,N_2984,N_3180);
and U8495 (N_8495,N_3856,N_4979);
nand U8496 (N_8496,N_3273,N_451);
xor U8497 (N_8497,N_4387,N_1883);
or U8498 (N_8498,N_1354,N_2298);
nand U8499 (N_8499,N_191,N_485);
xor U8500 (N_8500,N_4889,N_2208);
nand U8501 (N_8501,N_225,N_959);
xor U8502 (N_8502,N_331,N_262);
nor U8503 (N_8503,N_2848,N_3057);
or U8504 (N_8504,N_3429,N_1407);
nor U8505 (N_8505,N_3897,N_2067);
nand U8506 (N_8506,N_4901,N_3014);
nor U8507 (N_8507,N_2783,N_735);
nand U8508 (N_8508,N_4962,N_4256);
nor U8509 (N_8509,N_1359,N_4282);
xnor U8510 (N_8510,N_3634,N_3626);
and U8511 (N_8511,N_725,N_2998);
nor U8512 (N_8512,N_1861,N_3469);
and U8513 (N_8513,N_2917,N_1397);
and U8514 (N_8514,N_2427,N_4303);
xnor U8515 (N_8515,N_3822,N_2093);
or U8516 (N_8516,N_3898,N_3858);
xor U8517 (N_8517,N_4593,N_4317);
or U8518 (N_8518,N_4007,N_1402);
xor U8519 (N_8519,N_2306,N_725);
nor U8520 (N_8520,N_1735,N_329);
nor U8521 (N_8521,N_4974,N_4964);
nand U8522 (N_8522,N_709,N_3613);
or U8523 (N_8523,N_4927,N_1934);
or U8524 (N_8524,N_1276,N_603);
nand U8525 (N_8525,N_4359,N_1354);
and U8526 (N_8526,N_4207,N_1487);
nand U8527 (N_8527,N_1131,N_2970);
nand U8528 (N_8528,N_924,N_3667);
xnor U8529 (N_8529,N_2052,N_1135);
and U8530 (N_8530,N_2699,N_2175);
nor U8531 (N_8531,N_4523,N_438);
or U8532 (N_8532,N_3347,N_1329);
nand U8533 (N_8533,N_696,N_4081);
or U8534 (N_8534,N_4555,N_975);
nand U8535 (N_8535,N_4466,N_4223);
xor U8536 (N_8536,N_4334,N_876);
xnor U8537 (N_8537,N_2508,N_4647);
nor U8538 (N_8538,N_2705,N_284);
nor U8539 (N_8539,N_4677,N_1991);
and U8540 (N_8540,N_2059,N_621);
nor U8541 (N_8541,N_1996,N_3195);
nor U8542 (N_8542,N_1919,N_1367);
xnor U8543 (N_8543,N_506,N_2935);
and U8544 (N_8544,N_1647,N_1670);
xnor U8545 (N_8545,N_2128,N_1624);
and U8546 (N_8546,N_1062,N_388);
and U8547 (N_8547,N_1656,N_2608);
xor U8548 (N_8548,N_2968,N_2150);
and U8549 (N_8549,N_1679,N_809);
or U8550 (N_8550,N_193,N_2294);
nand U8551 (N_8551,N_2859,N_4027);
nand U8552 (N_8552,N_4158,N_811);
nand U8553 (N_8553,N_3820,N_3955);
nor U8554 (N_8554,N_335,N_3765);
nand U8555 (N_8555,N_360,N_4992);
and U8556 (N_8556,N_4376,N_4964);
nor U8557 (N_8557,N_4473,N_3644);
nor U8558 (N_8558,N_1550,N_3186);
or U8559 (N_8559,N_1636,N_3331);
xor U8560 (N_8560,N_2157,N_2878);
nand U8561 (N_8561,N_85,N_1244);
nand U8562 (N_8562,N_1150,N_4459);
nor U8563 (N_8563,N_1146,N_406);
and U8564 (N_8564,N_4658,N_3433);
nor U8565 (N_8565,N_2683,N_617);
nor U8566 (N_8566,N_3751,N_1365);
xnor U8567 (N_8567,N_1126,N_2236);
or U8568 (N_8568,N_630,N_730);
nor U8569 (N_8569,N_3725,N_4728);
nand U8570 (N_8570,N_3116,N_340);
and U8571 (N_8571,N_3349,N_4743);
xnor U8572 (N_8572,N_3383,N_415);
and U8573 (N_8573,N_4527,N_1194);
xnor U8574 (N_8574,N_3255,N_2833);
xnor U8575 (N_8575,N_4866,N_2956);
nor U8576 (N_8576,N_504,N_4205);
and U8577 (N_8577,N_103,N_3504);
nand U8578 (N_8578,N_259,N_2787);
or U8579 (N_8579,N_2451,N_4626);
xor U8580 (N_8580,N_148,N_67);
xnor U8581 (N_8581,N_4913,N_4427);
nor U8582 (N_8582,N_247,N_4091);
nor U8583 (N_8583,N_1918,N_4546);
xnor U8584 (N_8584,N_2253,N_3550);
nand U8585 (N_8585,N_4757,N_2698);
or U8586 (N_8586,N_3399,N_2148);
nor U8587 (N_8587,N_4959,N_2906);
and U8588 (N_8588,N_4395,N_4892);
nor U8589 (N_8589,N_2491,N_2016);
and U8590 (N_8590,N_4754,N_4602);
or U8591 (N_8591,N_1000,N_1977);
and U8592 (N_8592,N_1312,N_3344);
nor U8593 (N_8593,N_2522,N_3421);
nand U8594 (N_8594,N_1598,N_3282);
and U8595 (N_8595,N_1995,N_2635);
and U8596 (N_8596,N_1251,N_2583);
nor U8597 (N_8597,N_502,N_4051);
nand U8598 (N_8598,N_109,N_1521);
or U8599 (N_8599,N_1218,N_2579);
or U8600 (N_8600,N_1509,N_2798);
or U8601 (N_8601,N_3457,N_4223);
nand U8602 (N_8602,N_3683,N_763);
and U8603 (N_8603,N_3221,N_651);
and U8604 (N_8604,N_4373,N_3132);
nand U8605 (N_8605,N_2581,N_4599);
or U8606 (N_8606,N_3548,N_2953);
nor U8607 (N_8607,N_2168,N_2457);
and U8608 (N_8608,N_1877,N_2114);
and U8609 (N_8609,N_745,N_4407);
xor U8610 (N_8610,N_2953,N_4907);
nand U8611 (N_8611,N_1143,N_1376);
nor U8612 (N_8612,N_3066,N_1201);
nor U8613 (N_8613,N_2197,N_1173);
nand U8614 (N_8614,N_4955,N_3130);
and U8615 (N_8615,N_4327,N_319);
nor U8616 (N_8616,N_4546,N_2464);
xor U8617 (N_8617,N_1647,N_1525);
and U8618 (N_8618,N_3505,N_657);
nand U8619 (N_8619,N_191,N_370);
or U8620 (N_8620,N_3029,N_3562);
xor U8621 (N_8621,N_2208,N_3783);
nor U8622 (N_8622,N_2391,N_1126);
or U8623 (N_8623,N_2144,N_3222);
nand U8624 (N_8624,N_1079,N_3530);
and U8625 (N_8625,N_1238,N_653);
nand U8626 (N_8626,N_4679,N_1488);
xor U8627 (N_8627,N_99,N_654);
or U8628 (N_8628,N_2012,N_3816);
nand U8629 (N_8629,N_2279,N_2253);
nor U8630 (N_8630,N_2098,N_3784);
xor U8631 (N_8631,N_3501,N_269);
nor U8632 (N_8632,N_3441,N_2585);
nor U8633 (N_8633,N_877,N_2876);
or U8634 (N_8634,N_4131,N_4443);
nand U8635 (N_8635,N_249,N_4130);
nor U8636 (N_8636,N_2582,N_2535);
xnor U8637 (N_8637,N_4382,N_1133);
xor U8638 (N_8638,N_2912,N_2553);
xnor U8639 (N_8639,N_4273,N_621);
nand U8640 (N_8640,N_1656,N_132);
and U8641 (N_8641,N_2453,N_1000);
xnor U8642 (N_8642,N_184,N_4651);
nor U8643 (N_8643,N_4149,N_2789);
xor U8644 (N_8644,N_2485,N_3657);
nand U8645 (N_8645,N_546,N_1961);
nor U8646 (N_8646,N_630,N_1657);
nand U8647 (N_8647,N_548,N_2877);
nor U8648 (N_8648,N_3289,N_2487);
and U8649 (N_8649,N_3354,N_3889);
xor U8650 (N_8650,N_4525,N_4020);
nor U8651 (N_8651,N_356,N_2685);
nand U8652 (N_8652,N_3548,N_240);
or U8653 (N_8653,N_309,N_995);
nor U8654 (N_8654,N_3890,N_3729);
and U8655 (N_8655,N_3208,N_2365);
xor U8656 (N_8656,N_3754,N_4215);
or U8657 (N_8657,N_4798,N_4641);
and U8658 (N_8658,N_2079,N_1000);
xnor U8659 (N_8659,N_3793,N_2674);
or U8660 (N_8660,N_1125,N_1984);
or U8661 (N_8661,N_609,N_4593);
xor U8662 (N_8662,N_2662,N_850);
or U8663 (N_8663,N_828,N_1282);
and U8664 (N_8664,N_1339,N_4691);
nor U8665 (N_8665,N_906,N_1113);
xor U8666 (N_8666,N_4796,N_289);
nor U8667 (N_8667,N_3975,N_1918);
and U8668 (N_8668,N_4040,N_2497);
nand U8669 (N_8669,N_484,N_3454);
and U8670 (N_8670,N_4295,N_900);
nor U8671 (N_8671,N_3693,N_1414);
and U8672 (N_8672,N_1378,N_3512);
and U8673 (N_8673,N_996,N_3439);
xor U8674 (N_8674,N_600,N_1118);
xor U8675 (N_8675,N_1423,N_2167);
or U8676 (N_8676,N_2471,N_4367);
or U8677 (N_8677,N_4011,N_3100);
and U8678 (N_8678,N_4450,N_4584);
or U8679 (N_8679,N_3326,N_4017);
xor U8680 (N_8680,N_4865,N_4011);
or U8681 (N_8681,N_1334,N_3828);
nand U8682 (N_8682,N_2101,N_1951);
and U8683 (N_8683,N_4594,N_1386);
nor U8684 (N_8684,N_2260,N_1584);
nand U8685 (N_8685,N_90,N_235);
xnor U8686 (N_8686,N_1388,N_3914);
and U8687 (N_8687,N_1731,N_2792);
nand U8688 (N_8688,N_2861,N_1074);
xnor U8689 (N_8689,N_1752,N_3026);
and U8690 (N_8690,N_1919,N_4067);
or U8691 (N_8691,N_3002,N_1257);
nor U8692 (N_8692,N_1729,N_3414);
nand U8693 (N_8693,N_2211,N_2005);
xnor U8694 (N_8694,N_1209,N_4187);
nand U8695 (N_8695,N_3152,N_962);
xor U8696 (N_8696,N_1153,N_3731);
and U8697 (N_8697,N_3103,N_1648);
or U8698 (N_8698,N_4368,N_4412);
xnor U8699 (N_8699,N_177,N_1446);
and U8700 (N_8700,N_1826,N_2638);
xor U8701 (N_8701,N_1146,N_1869);
or U8702 (N_8702,N_1170,N_3843);
or U8703 (N_8703,N_108,N_4351);
xnor U8704 (N_8704,N_4593,N_3942);
or U8705 (N_8705,N_306,N_64);
and U8706 (N_8706,N_2417,N_2240);
and U8707 (N_8707,N_1236,N_2904);
or U8708 (N_8708,N_429,N_598);
nand U8709 (N_8709,N_2714,N_1204);
nor U8710 (N_8710,N_1788,N_3122);
or U8711 (N_8711,N_718,N_2684);
nor U8712 (N_8712,N_1945,N_1840);
nand U8713 (N_8713,N_3299,N_9);
or U8714 (N_8714,N_366,N_229);
nand U8715 (N_8715,N_2850,N_4296);
and U8716 (N_8716,N_2543,N_3238);
or U8717 (N_8717,N_2606,N_668);
and U8718 (N_8718,N_2501,N_1279);
and U8719 (N_8719,N_2213,N_841);
xor U8720 (N_8720,N_3222,N_1043);
nor U8721 (N_8721,N_1028,N_1041);
nand U8722 (N_8722,N_2129,N_3535);
xor U8723 (N_8723,N_3265,N_4257);
xnor U8724 (N_8724,N_2634,N_4923);
nand U8725 (N_8725,N_2998,N_16);
nand U8726 (N_8726,N_4953,N_2013);
xnor U8727 (N_8727,N_2201,N_4490);
nor U8728 (N_8728,N_3712,N_3962);
and U8729 (N_8729,N_3473,N_4331);
nand U8730 (N_8730,N_173,N_3242);
xnor U8731 (N_8731,N_2305,N_3306);
nand U8732 (N_8732,N_3126,N_640);
nand U8733 (N_8733,N_3465,N_1633);
nand U8734 (N_8734,N_4936,N_3596);
or U8735 (N_8735,N_4121,N_2456);
nor U8736 (N_8736,N_2793,N_4901);
nor U8737 (N_8737,N_1010,N_2402);
nor U8738 (N_8738,N_2530,N_1665);
or U8739 (N_8739,N_2539,N_420);
nor U8740 (N_8740,N_3706,N_4719);
nor U8741 (N_8741,N_2708,N_329);
or U8742 (N_8742,N_1574,N_4070);
nand U8743 (N_8743,N_59,N_3461);
nor U8744 (N_8744,N_604,N_3236);
or U8745 (N_8745,N_1902,N_3469);
and U8746 (N_8746,N_1604,N_1468);
xnor U8747 (N_8747,N_2857,N_1283);
xnor U8748 (N_8748,N_2401,N_4371);
nor U8749 (N_8749,N_3825,N_881);
nand U8750 (N_8750,N_3426,N_525);
xor U8751 (N_8751,N_845,N_4141);
nor U8752 (N_8752,N_4695,N_2504);
nand U8753 (N_8753,N_3868,N_2628);
or U8754 (N_8754,N_2039,N_4230);
and U8755 (N_8755,N_503,N_1447);
nand U8756 (N_8756,N_966,N_704);
xor U8757 (N_8757,N_2221,N_298);
nor U8758 (N_8758,N_833,N_4813);
or U8759 (N_8759,N_826,N_3851);
or U8760 (N_8760,N_2146,N_530);
nand U8761 (N_8761,N_3117,N_4436);
nand U8762 (N_8762,N_1498,N_4495);
nand U8763 (N_8763,N_3631,N_565);
xnor U8764 (N_8764,N_4127,N_4799);
nand U8765 (N_8765,N_1477,N_4075);
nand U8766 (N_8766,N_375,N_3206);
nor U8767 (N_8767,N_2069,N_3671);
xnor U8768 (N_8768,N_3187,N_4452);
nor U8769 (N_8769,N_3999,N_664);
nor U8770 (N_8770,N_800,N_1944);
nor U8771 (N_8771,N_739,N_1403);
nor U8772 (N_8772,N_1256,N_3971);
or U8773 (N_8773,N_4384,N_4599);
nor U8774 (N_8774,N_2255,N_602);
or U8775 (N_8775,N_1875,N_3647);
nand U8776 (N_8776,N_4003,N_3857);
nand U8777 (N_8777,N_2660,N_688);
nand U8778 (N_8778,N_4508,N_4608);
or U8779 (N_8779,N_4739,N_2133);
nand U8780 (N_8780,N_4578,N_969);
and U8781 (N_8781,N_1093,N_3315);
nor U8782 (N_8782,N_1449,N_4938);
nand U8783 (N_8783,N_3155,N_2542);
nor U8784 (N_8784,N_2853,N_4000);
xor U8785 (N_8785,N_1546,N_3904);
nor U8786 (N_8786,N_1444,N_4434);
or U8787 (N_8787,N_81,N_1935);
nand U8788 (N_8788,N_4761,N_1);
nand U8789 (N_8789,N_1301,N_895);
and U8790 (N_8790,N_339,N_272);
nor U8791 (N_8791,N_4194,N_4141);
nor U8792 (N_8792,N_279,N_4579);
nor U8793 (N_8793,N_3928,N_4387);
nand U8794 (N_8794,N_1234,N_3836);
or U8795 (N_8795,N_306,N_4279);
nand U8796 (N_8796,N_598,N_2350);
or U8797 (N_8797,N_2579,N_211);
or U8798 (N_8798,N_3236,N_2211);
or U8799 (N_8799,N_923,N_4332);
nand U8800 (N_8800,N_1445,N_1962);
and U8801 (N_8801,N_3210,N_2992);
and U8802 (N_8802,N_436,N_2823);
nand U8803 (N_8803,N_1771,N_2950);
nor U8804 (N_8804,N_2074,N_275);
and U8805 (N_8805,N_912,N_2950);
xor U8806 (N_8806,N_3237,N_4736);
nor U8807 (N_8807,N_836,N_1549);
or U8808 (N_8808,N_2183,N_4086);
nor U8809 (N_8809,N_3738,N_797);
nor U8810 (N_8810,N_1075,N_4157);
and U8811 (N_8811,N_1793,N_2844);
nor U8812 (N_8812,N_2653,N_369);
and U8813 (N_8813,N_4304,N_1826);
nand U8814 (N_8814,N_2807,N_1538);
nand U8815 (N_8815,N_4637,N_4498);
nor U8816 (N_8816,N_2907,N_3603);
and U8817 (N_8817,N_4522,N_955);
nor U8818 (N_8818,N_1737,N_2127);
nand U8819 (N_8819,N_4565,N_949);
or U8820 (N_8820,N_237,N_314);
or U8821 (N_8821,N_522,N_1289);
nand U8822 (N_8822,N_1470,N_2423);
xnor U8823 (N_8823,N_4071,N_1478);
or U8824 (N_8824,N_4560,N_4820);
and U8825 (N_8825,N_2181,N_4991);
or U8826 (N_8826,N_4632,N_2395);
xnor U8827 (N_8827,N_2662,N_2591);
and U8828 (N_8828,N_2647,N_4997);
and U8829 (N_8829,N_4315,N_4515);
nor U8830 (N_8830,N_3705,N_1573);
or U8831 (N_8831,N_272,N_2752);
or U8832 (N_8832,N_2494,N_1110);
or U8833 (N_8833,N_3974,N_536);
nor U8834 (N_8834,N_672,N_1081);
xor U8835 (N_8835,N_4111,N_4317);
or U8836 (N_8836,N_3328,N_4747);
xnor U8837 (N_8837,N_3324,N_1395);
nor U8838 (N_8838,N_4584,N_723);
nor U8839 (N_8839,N_1436,N_3759);
xor U8840 (N_8840,N_4594,N_3925);
nor U8841 (N_8841,N_2868,N_4252);
xor U8842 (N_8842,N_2179,N_924);
or U8843 (N_8843,N_857,N_4322);
nand U8844 (N_8844,N_3440,N_3732);
nor U8845 (N_8845,N_3636,N_2546);
xnor U8846 (N_8846,N_2788,N_2919);
xnor U8847 (N_8847,N_4948,N_3338);
nand U8848 (N_8848,N_550,N_754);
or U8849 (N_8849,N_3521,N_2836);
and U8850 (N_8850,N_3359,N_4416);
or U8851 (N_8851,N_829,N_4070);
xnor U8852 (N_8852,N_1242,N_4607);
nor U8853 (N_8853,N_4088,N_2455);
nand U8854 (N_8854,N_1837,N_40);
xor U8855 (N_8855,N_3822,N_229);
nor U8856 (N_8856,N_4190,N_2214);
xor U8857 (N_8857,N_2141,N_2376);
or U8858 (N_8858,N_891,N_561);
or U8859 (N_8859,N_83,N_536);
xnor U8860 (N_8860,N_2808,N_1427);
nor U8861 (N_8861,N_4579,N_2670);
nor U8862 (N_8862,N_1917,N_79);
and U8863 (N_8863,N_4771,N_207);
and U8864 (N_8864,N_4390,N_1337);
nand U8865 (N_8865,N_1257,N_4402);
nor U8866 (N_8866,N_2296,N_3536);
nand U8867 (N_8867,N_2785,N_860);
and U8868 (N_8868,N_1733,N_1699);
nor U8869 (N_8869,N_2443,N_3101);
and U8870 (N_8870,N_122,N_1032);
or U8871 (N_8871,N_3717,N_3693);
or U8872 (N_8872,N_4117,N_144);
xor U8873 (N_8873,N_2358,N_2300);
and U8874 (N_8874,N_4118,N_2409);
nand U8875 (N_8875,N_3043,N_3017);
nor U8876 (N_8876,N_3871,N_1099);
xnor U8877 (N_8877,N_711,N_1972);
xnor U8878 (N_8878,N_3329,N_1776);
and U8879 (N_8879,N_2641,N_3625);
and U8880 (N_8880,N_1121,N_1930);
nand U8881 (N_8881,N_9,N_1009);
xor U8882 (N_8882,N_2486,N_3304);
and U8883 (N_8883,N_4078,N_2426);
and U8884 (N_8884,N_939,N_4687);
and U8885 (N_8885,N_1683,N_4982);
nor U8886 (N_8886,N_1161,N_4214);
or U8887 (N_8887,N_1077,N_2819);
xnor U8888 (N_8888,N_730,N_2670);
and U8889 (N_8889,N_3171,N_1791);
or U8890 (N_8890,N_4243,N_4343);
nand U8891 (N_8891,N_4984,N_3885);
nor U8892 (N_8892,N_1941,N_3517);
or U8893 (N_8893,N_375,N_3630);
xnor U8894 (N_8894,N_4612,N_2195);
xor U8895 (N_8895,N_4959,N_906);
and U8896 (N_8896,N_4479,N_3313);
xnor U8897 (N_8897,N_4903,N_1788);
nand U8898 (N_8898,N_4742,N_3626);
xor U8899 (N_8899,N_2758,N_4055);
or U8900 (N_8900,N_2967,N_121);
nor U8901 (N_8901,N_1439,N_3764);
nor U8902 (N_8902,N_2153,N_3340);
nand U8903 (N_8903,N_831,N_4392);
or U8904 (N_8904,N_4500,N_3792);
xnor U8905 (N_8905,N_4580,N_4752);
or U8906 (N_8906,N_4084,N_4305);
xnor U8907 (N_8907,N_3479,N_291);
nor U8908 (N_8908,N_165,N_4325);
nand U8909 (N_8909,N_1887,N_4127);
nand U8910 (N_8910,N_1367,N_2618);
or U8911 (N_8911,N_4637,N_986);
nand U8912 (N_8912,N_2031,N_1040);
xor U8913 (N_8913,N_3257,N_4599);
nor U8914 (N_8914,N_2918,N_3832);
xnor U8915 (N_8915,N_2136,N_3460);
or U8916 (N_8916,N_3893,N_119);
nor U8917 (N_8917,N_2319,N_2640);
nor U8918 (N_8918,N_373,N_1516);
xnor U8919 (N_8919,N_2049,N_1857);
or U8920 (N_8920,N_3589,N_4286);
xnor U8921 (N_8921,N_4442,N_3259);
or U8922 (N_8922,N_4508,N_787);
nor U8923 (N_8923,N_970,N_1287);
nor U8924 (N_8924,N_1102,N_4828);
or U8925 (N_8925,N_918,N_2975);
nand U8926 (N_8926,N_346,N_2214);
xnor U8927 (N_8927,N_2341,N_3329);
or U8928 (N_8928,N_4546,N_1973);
nor U8929 (N_8929,N_1516,N_4379);
or U8930 (N_8930,N_4740,N_1495);
nor U8931 (N_8931,N_2729,N_858);
or U8932 (N_8932,N_2606,N_3296);
nor U8933 (N_8933,N_3157,N_563);
and U8934 (N_8934,N_959,N_997);
nor U8935 (N_8935,N_3485,N_2699);
and U8936 (N_8936,N_463,N_4702);
nand U8937 (N_8937,N_855,N_472);
xnor U8938 (N_8938,N_2268,N_2701);
xnor U8939 (N_8939,N_1825,N_733);
nor U8940 (N_8940,N_1351,N_1629);
nor U8941 (N_8941,N_2184,N_2677);
nor U8942 (N_8942,N_1732,N_3895);
nand U8943 (N_8943,N_1611,N_1588);
xnor U8944 (N_8944,N_4876,N_2749);
and U8945 (N_8945,N_1632,N_1287);
xor U8946 (N_8946,N_1354,N_2461);
and U8947 (N_8947,N_2677,N_964);
xor U8948 (N_8948,N_3215,N_1863);
or U8949 (N_8949,N_871,N_1009);
and U8950 (N_8950,N_391,N_1874);
nor U8951 (N_8951,N_2042,N_3551);
nor U8952 (N_8952,N_3467,N_3312);
or U8953 (N_8953,N_1183,N_3363);
or U8954 (N_8954,N_1533,N_2808);
xor U8955 (N_8955,N_3293,N_1052);
nor U8956 (N_8956,N_4307,N_4263);
and U8957 (N_8957,N_1041,N_1054);
xor U8958 (N_8958,N_4580,N_4837);
xnor U8959 (N_8959,N_1824,N_3164);
nand U8960 (N_8960,N_4766,N_3108);
and U8961 (N_8961,N_747,N_3077);
xor U8962 (N_8962,N_4056,N_1629);
and U8963 (N_8963,N_1855,N_4787);
and U8964 (N_8964,N_962,N_3424);
nor U8965 (N_8965,N_860,N_4170);
nand U8966 (N_8966,N_1584,N_78);
nand U8967 (N_8967,N_2373,N_4497);
nor U8968 (N_8968,N_3558,N_2347);
nor U8969 (N_8969,N_4305,N_3476);
xor U8970 (N_8970,N_4995,N_3638);
nor U8971 (N_8971,N_4726,N_1545);
xor U8972 (N_8972,N_214,N_270);
or U8973 (N_8973,N_4851,N_638);
or U8974 (N_8974,N_2041,N_3931);
nor U8975 (N_8975,N_1488,N_2741);
nand U8976 (N_8976,N_1648,N_3741);
xnor U8977 (N_8977,N_1470,N_668);
nand U8978 (N_8978,N_2962,N_720);
nor U8979 (N_8979,N_4621,N_3854);
or U8980 (N_8980,N_4935,N_3840);
and U8981 (N_8981,N_1056,N_4372);
xor U8982 (N_8982,N_1029,N_1286);
nor U8983 (N_8983,N_426,N_1959);
nand U8984 (N_8984,N_1676,N_4129);
xnor U8985 (N_8985,N_4605,N_4028);
and U8986 (N_8986,N_2653,N_2405);
nand U8987 (N_8987,N_82,N_1136);
nand U8988 (N_8988,N_2476,N_3307);
nor U8989 (N_8989,N_568,N_1055);
and U8990 (N_8990,N_2101,N_2995);
and U8991 (N_8991,N_111,N_3342);
nand U8992 (N_8992,N_1420,N_1155);
xor U8993 (N_8993,N_3174,N_2794);
and U8994 (N_8994,N_4672,N_4042);
nand U8995 (N_8995,N_4904,N_373);
and U8996 (N_8996,N_3649,N_3837);
and U8997 (N_8997,N_321,N_3638);
or U8998 (N_8998,N_4453,N_1370);
xnor U8999 (N_8999,N_711,N_3469);
or U9000 (N_9000,N_3736,N_2832);
and U9001 (N_9001,N_3544,N_1870);
and U9002 (N_9002,N_3545,N_3392);
nand U9003 (N_9003,N_294,N_3578);
xor U9004 (N_9004,N_4333,N_3585);
nand U9005 (N_9005,N_3346,N_2696);
xor U9006 (N_9006,N_4987,N_1107);
and U9007 (N_9007,N_892,N_1362);
and U9008 (N_9008,N_2270,N_3736);
or U9009 (N_9009,N_1288,N_710);
xnor U9010 (N_9010,N_4046,N_1325);
or U9011 (N_9011,N_3467,N_2599);
and U9012 (N_9012,N_3360,N_1315);
nand U9013 (N_9013,N_3338,N_2314);
xor U9014 (N_9014,N_1078,N_2828);
and U9015 (N_9015,N_2055,N_525);
xnor U9016 (N_9016,N_1214,N_3778);
xnor U9017 (N_9017,N_3235,N_3772);
xnor U9018 (N_9018,N_1041,N_3080);
and U9019 (N_9019,N_3746,N_860);
nand U9020 (N_9020,N_2310,N_757);
or U9021 (N_9021,N_2983,N_1124);
nand U9022 (N_9022,N_2440,N_2658);
nand U9023 (N_9023,N_4466,N_333);
or U9024 (N_9024,N_4178,N_1628);
nor U9025 (N_9025,N_4919,N_2068);
nand U9026 (N_9026,N_240,N_4439);
or U9027 (N_9027,N_1474,N_2079);
nor U9028 (N_9028,N_3237,N_3086);
xor U9029 (N_9029,N_4858,N_796);
or U9030 (N_9030,N_4046,N_4194);
xor U9031 (N_9031,N_1742,N_3822);
nand U9032 (N_9032,N_3505,N_3601);
or U9033 (N_9033,N_3697,N_3902);
and U9034 (N_9034,N_611,N_3688);
and U9035 (N_9035,N_1709,N_833);
nor U9036 (N_9036,N_3856,N_1233);
nor U9037 (N_9037,N_627,N_4226);
nor U9038 (N_9038,N_2979,N_2519);
or U9039 (N_9039,N_3050,N_4150);
and U9040 (N_9040,N_1158,N_3220);
and U9041 (N_9041,N_4062,N_1245);
and U9042 (N_9042,N_3345,N_32);
nor U9043 (N_9043,N_592,N_4815);
or U9044 (N_9044,N_4953,N_198);
nand U9045 (N_9045,N_4359,N_195);
nand U9046 (N_9046,N_3602,N_3612);
or U9047 (N_9047,N_1960,N_590);
and U9048 (N_9048,N_683,N_1107);
and U9049 (N_9049,N_68,N_1792);
xor U9050 (N_9050,N_4670,N_3851);
nor U9051 (N_9051,N_1710,N_794);
and U9052 (N_9052,N_4986,N_2840);
or U9053 (N_9053,N_4169,N_1153);
nor U9054 (N_9054,N_2509,N_3325);
or U9055 (N_9055,N_1126,N_997);
or U9056 (N_9056,N_725,N_2362);
nand U9057 (N_9057,N_4267,N_4551);
xnor U9058 (N_9058,N_2206,N_4217);
or U9059 (N_9059,N_4424,N_177);
nor U9060 (N_9060,N_2439,N_1685);
nor U9061 (N_9061,N_2267,N_652);
or U9062 (N_9062,N_4859,N_4590);
nor U9063 (N_9063,N_2832,N_198);
and U9064 (N_9064,N_1166,N_4111);
or U9065 (N_9065,N_4839,N_847);
nand U9066 (N_9066,N_2003,N_4473);
nand U9067 (N_9067,N_3445,N_721);
xor U9068 (N_9068,N_444,N_2255);
or U9069 (N_9069,N_4689,N_1156);
nand U9070 (N_9070,N_3851,N_3026);
xor U9071 (N_9071,N_1521,N_2825);
xor U9072 (N_9072,N_1784,N_639);
nor U9073 (N_9073,N_1175,N_3545);
nand U9074 (N_9074,N_2517,N_2275);
or U9075 (N_9075,N_3634,N_4857);
xor U9076 (N_9076,N_552,N_433);
nor U9077 (N_9077,N_2478,N_1905);
or U9078 (N_9078,N_4366,N_236);
xor U9079 (N_9079,N_3640,N_2690);
nand U9080 (N_9080,N_2599,N_643);
or U9081 (N_9081,N_4978,N_732);
or U9082 (N_9082,N_3108,N_3686);
nor U9083 (N_9083,N_3628,N_3224);
and U9084 (N_9084,N_62,N_277);
or U9085 (N_9085,N_4103,N_838);
or U9086 (N_9086,N_1852,N_765);
nand U9087 (N_9087,N_4841,N_3692);
or U9088 (N_9088,N_4408,N_1278);
nor U9089 (N_9089,N_2087,N_542);
nand U9090 (N_9090,N_1207,N_4572);
nor U9091 (N_9091,N_4933,N_325);
nor U9092 (N_9092,N_3648,N_2108);
and U9093 (N_9093,N_4180,N_2167);
nand U9094 (N_9094,N_1289,N_287);
and U9095 (N_9095,N_3340,N_4959);
xnor U9096 (N_9096,N_2810,N_1576);
nand U9097 (N_9097,N_4041,N_3497);
nor U9098 (N_9098,N_810,N_3632);
nand U9099 (N_9099,N_2256,N_1922);
xor U9100 (N_9100,N_3726,N_2604);
nand U9101 (N_9101,N_457,N_2219);
or U9102 (N_9102,N_4692,N_887);
or U9103 (N_9103,N_844,N_1847);
or U9104 (N_9104,N_1909,N_4154);
nand U9105 (N_9105,N_2906,N_3497);
or U9106 (N_9106,N_1388,N_3287);
nor U9107 (N_9107,N_127,N_4797);
nor U9108 (N_9108,N_343,N_1113);
nand U9109 (N_9109,N_471,N_2111);
nor U9110 (N_9110,N_1520,N_713);
xor U9111 (N_9111,N_3367,N_1965);
nor U9112 (N_9112,N_1694,N_23);
nor U9113 (N_9113,N_1885,N_465);
xor U9114 (N_9114,N_122,N_4078);
or U9115 (N_9115,N_3303,N_4851);
nand U9116 (N_9116,N_1392,N_2829);
nor U9117 (N_9117,N_2059,N_4806);
nand U9118 (N_9118,N_907,N_3200);
nand U9119 (N_9119,N_3153,N_2657);
or U9120 (N_9120,N_325,N_2865);
xor U9121 (N_9121,N_4150,N_36);
nor U9122 (N_9122,N_2050,N_4556);
or U9123 (N_9123,N_4858,N_226);
nand U9124 (N_9124,N_4988,N_2832);
or U9125 (N_9125,N_326,N_3131);
or U9126 (N_9126,N_3539,N_2452);
and U9127 (N_9127,N_3857,N_1989);
and U9128 (N_9128,N_3330,N_4834);
and U9129 (N_9129,N_4734,N_2884);
and U9130 (N_9130,N_649,N_4103);
and U9131 (N_9131,N_1767,N_4498);
nor U9132 (N_9132,N_4672,N_3463);
or U9133 (N_9133,N_2216,N_3043);
or U9134 (N_9134,N_1065,N_2692);
nor U9135 (N_9135,N_854,N_1096);
and U9136 (N_9136,N_1508,N_964);
or U9137 (N_9137,N_2312,N_2390);
and U9138 (N_9138,N_2021,N_3461);
nand U9139 (N_9139,N_153,N_1813);
or U9140 (N_9140,N_3711,N_568);
nand U9141 (N_9141,N_663,N_3054);
nand U9142 (N_9142,N_2706,N_4583);
and U9143 (N_9143,N_2107,N_4814);
nand U9144 (N_9144,N_4150,N_3137);
or U9145 (N_9145,N_3010,N_1893);
and U9146 (N_9146,N_3910,N_1925);
and U9147 (N_9147,N_2182,N_4000);
xnor U9148 (N_9148,N_3854,N_362);
or U9149 (N_9149,N_3102,N_2706);
nor U9150 (N_9150,N_4979,N_4817);
and U9151 (N_9151,N_1386,N_909);
nor U9152 (N_9152,N_2770,N_4713);
or U9153 (N_9153,N_3287,N_2886);
nand U9154 (N_9154,N_2569,N_4100);
or U9155 (N_9155,N_1529,N_4923);
or U9156 (N_9156,N_2664,N_3222);
and U9157 (N_9157,N_2525,N_4519);
or U9158 (N_9158,N_3187,N_4388);
xor U9159 (N_9159,N_2083,N_3102);
nor U9160 (N_9160,N_1020,N_4495);
nor U9161 (N_9161,N_260,N_1036);
nand U9162 (N_9162,N_828,N_718);
or U9163 (N_9163,N_2894,N_4021);
xor U9164 (N_9164,N_328,N_4216);
xnor U9165 (N_9165,N_4613,N_184);
xnor U9166 (N_9166,N_4797,N_4408);
or U9167 (N_9167,N_1266,N_803);
xnor U9168 (N_9168,N_4191,N_3717);
xnor U9169 (N_9169,N_1591,N_1145);
nand U9170 (N_9170,N_4857,N_1294);
nand U9171 (N_9171,N_2754,N_3992);
nand U9172 (N_9172,N_3082,N_3163);
or U9173 (N_9173,N_625,N_642);
xnor U9174 (N_9174,N_1884,N_177);
and U9175 (N_9175,N_3489,N_1757);
and U9176 (N_9176,N_3858,N_2086);
xor U9177 (N_9177,N_499,N_2301);
and U9178 (N_9178,N_1789,N_1171);
nor U9179 (N_9179,N_3137,N_4065);
and U9180 (N_9180,N_692,N_3682);
nor U9181 (N_9181,N_146,N_2827);
and U9182 (N_9182,N_3560,N_4524);
nand U9183 (N_9183,N_3757,N_527);
nor U9184 (N_9184,N_4005,N_2268);
nand U9185 (N_9185,N_4430,N_2746);
and U9186 (N_9186,N_901,N_2088);
or U9187 (N_9187,N_2665,N_2494);
xor U9188 (N_9188,N_81,N_1848);
nand U9189 (N_9189,N_4952,N_938);
nor U9190 (N_9190,N_2963,N_220);
and U9191 (N_9191,N_2875,N_4832);
nor U9192 (N_9192,N_2626,N_11);
nand U9193 (N_9193,N_777,N_54);
xnor U9194 (N_9194,N_4279,N_3889);
nor U9195 (N_9195,N_1268,N_1084);
nor U9196 (N_9196,N_3173,N_1629);
and U9197 (N_9197,N_4955,N_4669);
xor U9198 (N_9198,N_3648,N_4979);
and U9199 (N_9199,N_1105,N_3689);
nand U9200 (N_9200,N_1188,N_4612);
nand U9201 (N_9201,N_3849,N_555);
nor U9202 (N_9202,N_2637,N_661);
nand U9203 (N_9203,N_3731,N_1409);
or U9204 (N_9204,N_3158,N_3697);
or U9205 (N_9205,N_417,N_4017);
or U9206 (N_9206,N_4993,N_1301);
and U9207 (N_9207,N_453,N_4450);
xnor U9208 (N_9208,N_2137,N_4837);
nor U9209 (N_9209,N_4990,N_3021);
or U9210 (N_9210,N_2012,N_2207);
or U9211 (N_9211,N_240,N_551);
and U9212 (N_9212,N_1090,N_2940);
and U9213 (N_9213,N_3577,N_2677);
nand U9214 (N_9214,N_3075,N_3613);
and U9215 (N_9215,N_3615,N_744);
and U9216 (N_9216,N_3766,N_2924);
xnor U9217 (N_9217,N_999,N_2559);
or U9218 (N_9218,N_2446,N_3086);
and U9219 (N_9219,N_2043,N_2922);
and U9220 (N_9220,N_1064,N_1443);
xnor U9221 (N_9221,N_2380,N_1103);
xor U9222 (N_9222,N_434,N_3984);
or U9223 (N_9223,N_1466,N_508);
nand U9224 (N_9224,N_1229,N_590);
and U9225 (N_9225,N_400,N_1979);
and U9226 (N_9226,N_643,N_3081);
or U9227 (N_9227,N_3792,N_1740);
nand U9228 (N_9228,N_980,N_1446);
nand U9229 (N_9229,N_4738,N_2982);
nor U9230 (N_9230,N_3107,N_2884);
and U9231 (N_9231,N_4486,N_2626);
or U9232 (N_9232,N_653,N_2950);
xor U9233 (N_9233,N_4438,N_4282);
nor U9234 (N_9234,N_2303,N_4836);
or U9235 (N_9235,N_4567,N_976);
xnor U9236 (N_9236,N_4822,N_1432);
nand U9237 (N_9237,N_1035,N_3790);
nor U9238 (N_9238,N_168,N_1694);
nand U9239 (N_9239,N_2709,N_2334);
or U9240 (N_9240,N_3128,N_188);
or U9241 (N_9241,N_1589,N_3264);
nor U9242 (N_9242,N_2199,N_3152);
xnor U9243 (N_9243,N_1779,N_132);
nor U9244 (N_9244,N_4101,N_3447);
nand U9245 (N_9245,N_2188,N_4474);
nor U9246 (N_9246,N_4359,N_1168);
and U9247 (N_9247,N_4666,N_229);
xnor U9248 (N_9248,N_2118,N_951);
and U9249 (N_9249,N_183,N_2969);
or U9250 (N_9250,N_4914,N_2841);
nand U9251 (N_9251,N_4197,N_3208);
nor U9252 (N_9252,N_288,N_1009);
nor U9253 (N_9253,N_652,N_830);
or U9254 (N_9254,N_2384,N_3566);
nor U9255 (N_9255,N_301,N_3049);
or U9256 (N_9256,N_2768,N_1591);
and U9257 (N_9257,N_2451,N_2958);
xnor U9258 (N_9258,N_343,N_1596);
or U9259 (N_9259,N_3124,N_2199);
or U9260 (N_9260,N_3465,N_3270);
and U9261 (N_9261,N_1322,N_3454);
and U9262 (N_9262,N_2798,N_2248);
or U9263 (N_9263,N_3770,N_3064);
and U9264 (N_9264,N_2311,N_4214);
nand U9265 (N_9265,N_357,N_1449);
nor U9266 (N_9266,N_3079,N_3120);
or U9267 (N_9267,N_4336,N_1605);
xnor U9268 (N_9268,N_4587,N_4056);
nor U9269 (N_9269,N_636,N_76);
or U9270 (N_9270,N_1122,N_2188);
nand U9271 (N_9271,N_4675,N_2486);
nor U9272 (N_9272,N_4241,N_894);
nor U9273 (N_9273,N_1921,N_2218);
and U9274 (N_9274,N_2425,N_4306);
xnor U9275 (N_9275,N_4103,N_134);
and U9276 (N_9276,N_771,N_3464);
or U9277 (N_9277,N_3601,N_4067);
or U9278 (N_9278,N_4613,N_1795);
xor U9279 (N_9279,N_2470,N_4681);
or U9280 (N_9280,N_568,N_3690);
and U9281 (N_9281,N_2154,N_3070);
nor U9282 (N_9282,N_1472,N_3632);
nand U9283 (N_9283,N_2752,N_3102);
xor U9284 (N_9284,N_1374,N_1495);
and U9285 (N_9285,N_4705,N_206);
and U9286 (N_9286,N_3253,N_1318);
and U9287 (N_9287,N_1270,N_2761);
nand U9288 (N_9288,N_4203,N_1416);
nand U9289 (N_9289,N_3807,N_2774);
xnor U9290 (N_9290,N_70,N_2255);
nand U9291 (N_9291,N_3905,N_4329);
nand U9292 (N_9292,N_846,N_148);
xor U9293 (N_9293,N_4768,N_418);
or U9294 (N_9294,N_1012,N_209);
or U9295 (N_9295,N_2668,N_3828);
nor U9296 (N_9296,N_4960,N_258);
and U9297 (N_9297,N_4223,N_284);
and U9298 (N_9298,N_2914,N_2589);
nor U9299 (N_9299,N_4075,N_3973);
and U9300 (N_9300,N_3257,N_1514);
or U9301 (N_9301,N_4324,N_1143);
and U9302 (N_9302,N_3047,N_1734);
nand U9303 (N_9303,N_4823,N_3342);
nand U9304 (N_9304,N_1885,N_4367);
or U9305 (N_9305,N_76,N_3417);
nand U9306 (N_9306,N_4568,N_801);
nand U9307 (N_9307,N_3112,N_3783);
and U9308 (N_9308,N_1719,N_2228);
xor U9309 (N_9309,N_102,N_1004);
nor U9310 (N_9310,N_2685,N_4895);
nand U9311 (N_9311,N_2223,N_4338);
or U9312 (N_9312,N_535,N_4425);
or U9313 (N_9313,N_1020,N_2067);
and U9314 (N_9314,N_3342,N_1612);
xor U9315 (N_9315,N_1473,N_2862);
or U9316 (N_9316,N_769,N_2649);
nor U9317 (N_9317,N_721,N_4390);
and U9318 (N_9318,N_4711,N_623);
nand U9319 (N_9319,N_381,N_1995);
xnor U9320 (N_9320,N_287,N_2526);
nand U9321 (N_9321,N_2052,N_3549);
xor U9322 (N_9322,N_3371,N_1002);
nor U9323 (N_9323,N_932,N_3881);
nor U9324 (N_9324,N_2973,N_4426);
nand U9325 (N_9325,N_3759,N_3480);
nand U9326 (N_9326,N_933,N_1910);
xor U9327 (N_9327,N_2618,N_3350);
xnor U9328 (N_9328,N_1759,N_4184);
nand U9329 (N_9329,N_3490,N_1684);
nor U9330 (N_9330,N_2783,N_2724);
or U9331 (N_9331,N_573,N_4756);
xor U9332 (N_9332,N_2205,N_1482);
xor U9333 (N_9333,N_1311,N_2039);
nor U9334 (N_9334,N_510,N_539);
or U9335 (N_9335,N_2139,N_4524);
nor U9336 (N_9336,N_1585,N_4521);
and U9337 (N_9337,N_922,N_3183);
nor U9338 (N_9338,N_1734,N_3456);
nand U9339 (N_9339,N_2866,N_223);
xnor U9340 (N_9340,N_4685,N_3086);
nand U9341 (N_9341,N_687,N_2535);
nand U9342 (N_9342,N_1352,N_538);
xor U9343 (N_9343,N_3189,N_2721);
and U9344 (N_9344,N_444,N_3412);
or U9345 (N_9345,N_582,N_2960);
xor U9346 (N_9346,N_1605,N_1073);
or U9347 (N_9347,N_3269,N_4647);
xor U9348 (N_9348,N_1573,N_2816);
and U9349 (N_9349,N_4019,N_3498);
or U9350 (N_9350,N_2987,N_3782);
nor U9351 (N_9351,N_3325,N_3228);
nand U9352 (N_9352,N_1121,N_475);
nand U9353 (N_9353,N_2402,N_1951);
nand U9354 (N_9354,N_1241,N_3346);
nor U9355 (N_9355,N_2483,N_4076);
or U9356 (N_9356,N_1457,N_4918);
nor U9357 (N_9357,N_3029,N_4859);
nor U9358 (N_9358,N_183,N_4918);
and U9359 (N_9359,N_1615,N_1661);
and U9360 (N_9360,N_2391,N_120);
and U9361 (N_9361,N_2166,N_4605);
nor U9362 (N_9362,N_3413,N_4379);
xor U9363 (N_9363,N_2836,N_3127);
nand U9364 (N_9364,N_3584,N_1047);
and U9365 (N_9365,N_743,N_968);
xnor U9366 (N_9366,N_4405,N_4644);
nand U9367 (N_9367,N_320,N_2192);
and U9368 (N_9368,N_3719,N_4568);
xor U9369 (N_9369,N_675,N_1327);
nor U9370 (N_9370,N_1201,N_2137);
or U9371 (N_9371,N_2256,N_715);
and U9372 (N_9372,N_1197,N_2338);
xor U9373 (N_9373,N_2111,N_4187);
nand U9374 (N_9374,N_321,N_1000);
or U9375 (N_9375,N_4990,N_3642);
nand U9376 (N_9376,N_963,N_1692);
nand U9377 (N_9377,N_3363,N_1857);
or U9378 (N_9378,N_1949,N_4633);
and U9379 (N_9379,N_2858,N_4782);
xnor U9380 (N_9380,N_2014,N_2642);
or U9381 (N_9381,N_3739,N_4581);
nand U9382 (N_9382,N_1306,N_3037);
xor U9383 (N_9383,N_2207,N_4144);
xnor U9384 (N_9384,N_2124,N_2029);
nand U9385 (N_9385,N_2643,N_3512);
nor U9386 (N_9386,N_508,N_2077);
or U9387 (N_9387,N_2298,N_2096);
or U9388 (N_9388,N_3419,N_4576);
or U9389 (N_9389,N_683,N_4378);
and U9390 (N_9390,N_4666,N_4819);
nand U9391 (N_9391,N_1907,N_3602);
nor U9392 (N_9392,N_900,N_3163);
nand U9393 (N_9393,N_1895,N_1939);
nor U9394 (N_9394,N_2797,N_3376);
xnor U9395 (N_9395,N_2236,N_357);
or U9396 (N_9396,N_3135,N_4332);
and U9397 (N_9397,N_1393,N_2690);
xor U9398 (N_9398,N_3263,N_646);
nor U9399 (N_9399,N_3221,N_173);
nand U9400 (N_9400,N_866,N_1669);
nor U9401 (N_9401,N_2468,N_47);
xor U9402 (N_9402,N_1465,N_1473);
xor U9403 (N_9403,N_4716,N_2600);
nand U9404 (N_9404,N_1916,N_799);
xor U9405 (N_9405,N_1664,N_1953);
or U9406 (N_9406,N_3825,N_4516);
xor U9407 (N_9407,N_4075,N_4023);
nand U9408 (N_9408,N_3533,N_2144);
nand U9409 (N_9409,N_2988,N_4866);
or U9410 (N_9410,N_4856,N_4004);
nand U9411 (N_9411,N_4654,N_4746);
nor U9412 (N_9412,N_4014,N_1720);
xnor U9413 (N_9413,N_2570,N_4558);
xnor U9414 (N_9414,N_3488,N_2663);
xor U9415 (N_9415,N_702,N_784);
xnor U9416 (N_9416,N_3271,N_3916);
and U9417 (N_9417,N_4262,N_661);
nand U9418 (N_9418,N_3435,N_1220);
nand U9419 (N_9419,N_196,N_4472);
and U9420 (N_9420,N_315,N_1903);
nand U9421 (N_9421,N_2188,N_3118);
xor U9422 (N_9422,N_1725,N_4360);
xnor U9423 (N_9423,N_2174,N_244);
and U9424 (N_9424,N_724,N_1418);
or U9425 (N_9425,N_741,N_3958);
nor U9426 (N_9426,N_1414,N_3553);
nor U9427 (N_9427,N_4429,N_2467);
or U9428 (N_9428,N_2785,N_1480);
or U9429 (N_9429,N_1236,N_2562);
and U9430 (N_9430,N_4346,N_4143);
nand U9431 (N_9431,N_924,N_3181);
or U9432 (N_9432,N_712,N_4945);
nand U9433 (N_9433,N_4065,N_1758);
xnor U9434 (N_9434,N_3959,N_2218);
nor U9435 (N_9435,N_1238,N_535);
nor U9436 (N_9436,N_817,N_1237);
or U9437 (N_9437,N_2377,N_3192);
and U9438 (N_9438,N_2181,N_2318);
and U9439 (N_9439,N_3011,N_3529);
nor U9440 (N_9440,N_4023,N_4181);
or U9441 (N_9441,N_1969,N_2795);
xor U9442 (N_9442,N_3042,N_3500);
xor U9443 (N_9443,N_3430,N_3609);
or U9444 (N_9444,N_2673,N_1796);
nor U9445 (N_9445,N_1959,N_404);
nand U9446 (N_9446,N_3909,N_3926);
or U9447 (N_9447,N_1304,N_4208);
xor U9448 (N_9448,N_2200,N_3634);
nor U9449 (N_9449,N_4219,N_4012);
xnor U9450 (N_9450,N_3782,N_352);
xnor U9451 (N_9451,N_2413,N_3422);
or U9452 (N_9452,N_4840,N_4549);
nand U9453 (N_9453,N_4514,N_4434);
nand U9454 (N_9454,N_2239,N_4117);
nand U9455 (N_9455,N_1890,N_2641);
or U9456 (N_9456,N_3297,N_4051);
xnor U9457 (N_9457,N_3512,N_3831);
nand U9458 (N_9458,N_739,N_4938);
and U9459 (N_9459,N_4826,N_434);
nand U9460 (N_9460,N_1613,N_1166);
and U9461 (N_9461,N_2864,N_1338);
and U9462 (N_9462,N_4390,N_1474);
nand U9463 (N_9463,N_329,N_1375);
nor U9464 (N_9464,N_1137,N_2121);
and U9465 (N_9465,N_1823,N_3432);
and U9466 (N_9466,N_3765,N_1335);
or U9467 (N_9467,N_916,N_2521);
nand U9468 (N_9468,N_377,N_688);
nand U9469 (N_9469,N_4388,N_3280);
nor U9470 (N_9470,N_3524,N_2651);
nor U9471 (N_9471,N_1989,N_4216);
nor U9472 (N_9472,N_4641,N_4152);
and U9473 (N_9473,N_2546,N_4547);
or U9474 (N_9474,N_4055,N_4772);
nor U9475 (N_9475,N_2393,N_2056);
nor U9476 (N_9476,N_896,N_1812);
nor U9477 (N_9477,N_3663,N_978);
xor U9478 (N_9478,N_3689,N_1285);
xnor U9479 (N_9479,N_2098,N_1804);
and U9480 (N_9480,N_1764,N_1085);
nand U9481 (N_9481,N_2089,N_1605);
xnor U9482 (N_9482,N_3038,N_387);
xnor U9483 (N_9483,N_1148,N_1719);
or U9484 (N_9484,N_1477,N_753);
or U9485 (N_9485,N_3224,N_3269);
or U9486 (N_9486,N_4668,N_2320);
xor U9487 (N_9487,N_878,N_1329);
and U9488 (N_9488,N_445,N_4227);
or U9489 (N_9489,N_4854,N_3697);
nand U9490 (N_9490,N_3665,N_508);
or U9491 (N_9491,N_139,N_240);
and U9492 (N_9492,N_181,N_591);
or U9493 (N_9493,N_3938,N_4542);
nor U9494 (N_9494,N_1593,N_1013);
xor U9495 (N_9495,N_3354,N_878);
xor U9496 (N_9496,N_3399,N_334);
and U9497 (N_9497,N_3167,N_1847);
nor U9498 (N_9498,N_3977,N_3968);
nor U9499 (N_9499,N_2731,N_983);
nand U9500 (N_9500,N_384,N_1726);
nand U9501 (N_9501,N_1831,N_3181);
nand U9502 (N_9502,N_2854,N_26);
or U9503 (N_9503,N_1690,N_4589);
nor U9504 (N_9504,N_4458,N_77);
nor U9505 (N_9505,N_317,N_1815);
nor U9506 (N_9506,N_1529,N_278);
nand U9507 (N_9507,N_2117,N_271);
xor U9508 (N_9508,N_4898,N_1601);
nor U9509 (N_9509,N_2362,N_3265);
xor U9510 (N_9510,N_1585,N_728);
xor U9511 (N_9511,N_2905,N_3959);
and U9512 (N_9512,N_1547,N_1870);
nand U9513 (N_9513,N_4959,N_4419);
and U9514 (N_9514,N_1790,N_263);
and U9515 (N_9515,N_856,N_1141);
nand U9516 (N_9516,N_4403,N_4125);
and U9517 (N_9517,N_1178,N_1996);
xnor U9518 (N_9518,N_1405,N_453);
nand U9519 (N_9519,N_4072,N_2779);
or U9520 (N_9520,N_4918,N_3239);
or U9521 (N_9521,N_2194,N_2011);
nand U9522 (N_9522,N_611,N_411);
nor U9523 (N_9523,N_4478,N_3215);
or U9524 (N_9524,N_308,N_4466);
nor U9525 (N_9525,N_4817,N_2509);
xor U9526 (N_9526,N_1182,N_4790);
nor U9527 (N_9527,N_2885,N_2575);
or U9528 (N_9528,N_3840,N_4205);
and U9529 (N_9529,N_3436,N_4116);
or U9530 (N_9530,N_4191,N_4201);
nand U9531 (N_9531,N_3516,N_4126);
or U9532 (N_9532,N_4262,N_354);
and U9533 (N_9533,N_1919,N_504);
xnor U9534 (N_9534,N_543,N_1631);
xnor U9535 (N_9535,N_2093,N_2017);
nor U9536 (N_9536,N_4855,N_3886);
or U9537 (N_9537,N_219,N_4194);
nor U9538 (N_9538,N_2481,N_2353);
nor U9539 (N_9539,N_2374,N_1432);
and U9540 (N_9540,N_3750,N_687);
and U9541 (N_9541,N_4075,N_4140);
nand U9542 (N_9542,N_131,N_3130);
nor U9543 (N_9543,N_1515,N_1219);
xnor U9544 (N_9544,N_4985,N_901);
nor U9545 (N_9545,N_4167,N_1642);
and U9546 (N_9546,N_1906,N_2548);
nand U9547 (N_9547,N_4637,N_2351);
nor U9548 (N_9548,N_3094,N_2186);
or U9549 (N_9549,N_4760,N_3990);
nand U9550 (N_9550,N_221,N_3860);
xnor U9551 (N_9551,N_483,N_4323);
and U9552 (N_9552,N_3630,N_4914);
nand U9553 (N_9553,N_3574,N_3025);
or U9554 (N_9554,N_4359,N_3212);
xor U9555 (N_9555,N_2027,N_1318);
nand U9556 (N_9556,N_1142,N_3915);
or U9557 (N_9557,N_4726,N_588);
xnor U9558 (N_9558,N_3001,N_1024);
xnor U9559 (N_9559,N_3470,N_4019);
xnor U9560 (N_9560,N_1822,N_1680);
xnor U9561 (N_9561,N_1578,N_3982);
nor U9562 (N_9562,N_1430,N_908);
and U9563 (N_9563,N_1473,N_201);
nand U9564 (N_9564,N_2324,N_2244);
and U9565 (N_9565,N_2870,N_3368);
or U9566 (N_9566,N_113,N_10);
nand U9567 (N_9567,N_944,N_4293);
xnor U9568 (N_9568,N_219,N_1583);
nand U9569 (N_9569,N_4232,N_1877);
nand U9570 (N_9570,N_2779,N_3684);
xor U9571 (N_9571,N_1321,N_2152);
or U9572 (N_9572,N_269,N_3546);
nand U9573 (N_9573,N_4323,N_3515);
xnor U9574 (N_9574,N_4664,N_1897);
nand U9575 (N_9575,N_3477,N_958);
xnor U9576 (N_9576,N_4711,N_2536);
nand U9577 (N_9577,N_335,N_3475);
nor U9578 (N_9578,N_1530,N_4483);
nand U9579 (N_9579,N_3659,N_3047);
xnor U9580 (N_9580,N_4531,N_1517);
nor U9581 (N_9581,N_2778,N_817);
or U9582 (N_9582,N_3332,N_84);
and U9583 (N_9583,N_1267,N_2376);
or U9584 (N_9584,N_4367,N_3198);
and U9585 (N_9585,N_2122,N_4131);
nand U9586 (N_9586,N_3430,N_68);
and U9587 (N_9587,N_4279,N_3511);
and U9588 (N_9588,N_1185,N_3339);
and U9589 (N_9589,N_4577,N_2154);
xor U9590 (N_9590,N_4472,N_1480);
nor U9591 (N_9591,N_417,N_1632);
xnor U9592 (N_9592,N_2133,N_4476);
xor U9593 (N_9593,N_2385,N_4872);
and U9594 (N_9594,N_701,N_2838);
nand U9595 (N_9595,N_1728,N_3726);
or U9596 (N_9596,N_1756,N_3104);
and U9597 (N_9597,N_4856,N_2866);
nand U9598 (N_9598,N_916,N_4169);
or U9599 (N_9599,N_2489,N_4659);
and U9600 (N_9600,N_613,N_1914);
nand U9601 (N_9601,N_2178,N_2157);
xor U9602 (N_9602,N_118,N_4551);
nor U9603 (N_9603,N_2511,N_683);
and U9604 (N_9604,N_1106,N_1198);
and U9605 (N_9605,N_580,N_207);
or U9606 (N_9606,N_1219,N_620);
xor U9607 (N_9607,N_222,N_2755);
or U9608 (N_9608,N_4732,N_3509);
or U9609 (N_9609,N_607,N_3477);
or U9610 (N_9610,N_1268,N_2854);
nor U9611 (N_9611,N_3358,N_272);
and U9612 (N_9612,N_237,N_2403);
nand U9613 (N_9613,N_2029,N_3905);
nand U9614 (N_9614,N_4658,N_3140);
nand U9615 (N_9615,N_4947,N_3773);
nor U9616 (N_9616,N_310,N_2216);
nand U9617 (N_9617,N_3062,N_2252);
xor U9618 (N_9618,N_3233,N_3257);
nand U9619 (N_9619,N_1995,N_966);
nor U9620 (N_9620,N_3924,N_596);
xnor U9621 (N_9621,N_1968,N_1937);
or U9622 (N_9622,N_2570,N_3626);
nor U9623 (N_9623,N_980,N_130);
xnor U9624 (N_9624,N_1548,N_3671);
nor U9625 (N_9625,N_4152,N_1209);
or U9626 (N_9626,N_1308,N_1486);
nand U9627 (N_9627,N_1207,N_2836);
or U9628 (N_9628,N_2247,N_68);
nor U9629 (N_9629,N_2142,N_4884);
or U9630 (N_9630,N_3446,N_4133);
or U9631 (N_9631,N_929,N_1630);
or U9632 (N_9632,N_2051,N_2559);
or U9633 (N_9633,N_2754,N_4573);
and U9634 (N_9634,N_4606,N_2319);
xnor U9635 (N_9635,N_4200,N_4785);
xnor U9636 (N_9636,N_3004,N_903);
xnor U9637 (N_9637,N_4510,N_4586);
nand U9638 (N_9638,N_3458,N_4392);
xor U9639 (N_9639,N_1500,N_3131);
nor U9640 (N_9640,N_2467,N_3762);
xnor U9641 (N_9641,N_4556,N_4926);
or U9642 (N_9642,N_2043,N_1257);
and U9643 (N_9643,N_4622,N_726);
or U9644 (N_9644,N_1049,N_1299);
nor U9645 (N_9645,N_1606,N_2778);
nand U9646 (N_9646,N_1655,N_639);
or U9647 (N_9647,N_857,N_1670);
nor U9648 (N_9648,N_235,N_2662);
and U9649 (N_9649,N_4540,N_3802);
or U9650 (N_9650,N_4063,N_3904);
nor U9651 (N_9651,N_1513,N_2609);
nand U9652 (N_9652,N_549,N_168);
and U9653 (N_9653,N_938,N_2846);
nand U9654 (N_9654,N_3844,N_2850);
or U9655 (N_9655,N_2973,N_1214);
and U9656 (N_9656,N_2424,N_3487);
or U9657 (N_9657,N_3884,N_3145);
nor U9658 (N_9658,N_3717,N_3973);
nand U9659 (N_9659,N_1404,N_1041);
or U9660 (N_9660,N_2223,N_4121);
or U9661 (N_9661,N_2269,N_4401);
and U9662 (N_9662,N_2153,N_4000);
nand U9663 (N_9663,N_4299,N_1671);
xor U9664 (N_9664,N_219,N_2183);
nor U9665 (N_9665,N_3465,N_2614);
and U9666 (N_9666,N_3693,N_3466);
nor U9667 (N_9667,N_4289,N_2829);
and U9668 (N_9668,N_1335,N_4672);
and U9669 (N_9669,N_1151,N_97);
xor U9670 (N_9670,N_2206,N_663);
xnor U9671 (N_9671,N_1957,N_4461);
or U9672 (N_9672,N_1220,N_4999);
nor U9673 (N_9673,N_4636,N_1494);
nor U9674 (N_9674,N_267,N_2688);
nor U9675 (N_9675,N_2315,N_2304);
and U9676 (N_9676,N_1476,N_3434);
xor U9677 (N_9677,N_626,N_1645);
nand U9678 (N_9678,N_2397,N_2547);
xor U9679 (N_9679,N_4012,N_2166);
xnor U9680 (N_9680,N_2681,N_3358);
or U9681 (N_9681,N_1079,N_1691);
nor U9682 (N_9682,N_168,N_4014);
nand U9683 (N_9683,N_4932,N_1739);
nor U9684 (N_9684,N_4178,N_198);
and U9685 (N_9685,N_4834,N_3747);
nor U9686 (N_9686,N_4082,N_1550);
or U9687 (N_9687,N_1839,N_167);
nor U9688 (N_9688,N_1992,N_4315);
nand U9689 (N_9689,N_959,N_531);
nor U9690 (N_9690,N_318,N_2261);
xor U9691 (N_9691,N_1561,N_3689);
or U9692 (N_9692,N_2554,N_391);
and U9693 (N_9693,N_1291,N_3888);
and U9694 (N_9694,N_3915,N_1060);
nor U9695 (N_9695,N_3455,N_3996);
nand U9696 (N_9696,N_1156,N_2748);
or U9697 (N_9697,N_4497,N_4535);
nand U9698 (N_9698,N_4858,N_3055);
or U9699 (N_9699,N_2789,N_3787);
xor U9700 (N_9700,N_4987,N_1259);
nor U9701 (N_9701,N_3190,N_424);
nand U9702 (N_9702,N_651,N_2169);
nor U9703 (N_9703,N_918,N_4020);
nand U9704 (N_9704,N_1295,N_2984);
or U9705 (N_9705,N_3327,N_2777);
and U9706 (N_9706,N_752,N_947);
xor U9707 (N_9707,N_689,N_585);
and U9708 (N_9708,N_4141,N_4378);
nor U9709 (N_9709,N_104,N_24);
nand U9710 (N_9710,N_451,N_981);
or U9711 (N_9711,N_3927,N_1806);
or U9712 (N_9712,N_3728,N_4191);
nor U9713 (N_9713,N_2873,N_4068);
and U9714 (N_9714,N_892,N_3787);
and U9715 (N_9715,N_3802,N_990);
xnor U9716 (N_9716,N_4782,N_727);
or U9717 (N_9717,N_4718,N_1824);
or U9718 (N_9718,N_3252,N_754);
or U9719 (N_9719,N_1627,N_607);
nand U9720 (N_9720,N_4994,N_925);
nor U9721 (N_9721,N_4634,N_102);
nor U9722 (N_9722,N_3446,N_1959);
xnor U9723 (N_9723,N_2626,N_4462);
or U9724 (N_9724,N_3557,N_1274);
or U9725 (N_9725,N_1368,N_154);
and U9726 (N_9726,N_863,N_3260);
nand U9727 (N_9727,N_351,N_4717);
or U9728 (N_9728,N_534,N_3280);
or U9729 (N_9729,N_2029,N_4621);
nand U9730 (N_9730,N_4338,N_4573);
nor U9731 (N_9731,N_2706,N_2462);
and U9732 (N_9732,N_3849,N_2775);
nand U9733 (N_9733,N_3232,N_876);
xor U9734 (N_9734,N_4658,N_770);
xor U9735 (N_9735,N_4932,N_4915);
xor U9736 (N_9736,N_3682,N_197);
and U9737 (N_9737,N_1505,N_2931);
xnor U9738 (N_9738,N_28,N_804);
nand U9739 (N_9739,N_3410,N_2327);
nor U9740 (N_9740,N_4633,N_1020);
xor U9741 (N_9741,N_731,N_3761);
nand U9742 (N_9742,N_3958,N_3789);
and U9743 (N_9743,N_4699,N_890);
and U9744 (N_9744,N_770,N_2200);
xnor U9745 (N_9745,N_4750,N_4001);
or U9746 (N_9746,N_1187,N_3831);
xor U9747 (N_9747,N_4344,N_4418);
and U9748 (N_9748,N_4004,N_1655);
nand U9749 (N_9749,N_831,N_1773);
nor U9750 (N_9750,N_3875,N_4262);
or U9751 (N_9751,N_2971,N_4777);
and U9752 (N_9752,N_2777,N_2039);
and U9753 (N_9753,N_1296,N_1471);
nor U9754 (N_9754,N_1564,N_3066);
and U9755 (N_9755,N_2808,N_1960);
and U9756 (N_9756,N_747,N_4911);
nor U9757 (N_9757,N_2064,N_3754);
or U9758 (N_9758,N_1146,N_1489);
or U9759 (N_9759,N_3107,N_2906);
xor U9760 (N_9760,N_4709,N_709);
nor U9761 (N_9761,N_2561,N_2841);
xnor U9762 (N_9762,N_3356,N_3878);
xnor U9763 (N_9763,N_1061,N_3796);
or U9764 (N_9764,N_4658,N_3568);
xor U9765 (N_9765,N_2753,N_1541);
or U9766 (N_9766,N_2611,N_3946);
nor U9767 (N_9767,N_1994,N_216);
xnor U9768 (N_9768,N_2141,N_3457);
nand U9769 (N_9769,N_3965,N_54);
and U9770 (N_9770,N_4521,N_3629);
xnor U9771 (N_9771,N_2551,N_4507);
xnor U9772 (N_9772,N_1859,N_1439);
nand U9773 (N_9773,N_347,N_4879);
xor U9774 (N_9774,N_1692,N_4184);
nor U9775 (N_9775,N_3549,N_1034);
nor U9776 (N_9776,N_3741,N_1715);
nand U9777 (N_9777,N_2687,N_1268);
and U9778 (N_9778,N_2092,N_492);
nor U9779 (N_9779,N_3867,N_614);
or U9780 (N_9780,N_1990,N_2469);
and U9781 (N_9781,N_2099,N_1319);
xnor U9782 (N_9782,N_2849,N_3982);
and U9783 (N_9783,N_1314,N_1417);
nor U9784 (N_9784,N_1736,N_3004);
nand U9785 (N_9785,N_3227,N_4578);
nand U9786 (N_9786,N_1124,N_475);
and U9787 (N_9787,N_249,N_676);
nor U9788 (N_9788,N_269,N_2129);
nor U9789 (N_9789,N_3671,N_4921);
or U9790 (N_9790,N_3491,N_1801);
or U9791 (N_9791,N_3736,N_4489);
or U9792 (N_9792,N_4977,N_4274);
or U9793 (N_9793,N_4629,N_2223);
and U9794 (N_9794,N_2767,N_944);
xnor U9795 (N_9795,N_3917,N_3366);
nand U9796 (N_9796,N_4572,N_2893);
nand U9797 (N_9797,N_1679,N_1652);
xor U9798 (N_9798,N_589,N_3779);
nand U9799 (N_9799,N_3020,N_4899);
or U9800 (N_9800,N_1962,N_2761);
nand U9801 (N_9801,N_2565,N_3711);
xnor U9802 (N_9802,N_3099,N_1081);
and U9803 (N_9803,N_1675,N_742);
nand U9804 (N_9804,N_1558,N_3142);
or U9805 (N_9805,N_836,N_3279);
nor U9806 (N_9806,N_1207,N_2270);
nand U9807 (N_9807,N_3570,N_685);
xnor U9808 (N_9808,N_3823,N_3369);
nand U9809 (N_9809,N_2560,N_2205);
and U9810 (N_9810,N_2972,N_4825);
and U9811 (N_9811,N_527,N_11);
nand U9812 (N_9812,N_108,N_3730);
xnor U9813 (N_9813,N_3008,N_3747);
or U9814 (N_9814,N_1746,N_2976);
nand U9815 (N_9815,N_425,N_4749);
xor U9816 (N_9816,N_3341,N_3266);
nand U9817 (N_9817,N_1355,N_1991);
xnor U9818 (N_9818,N_4088,N_2580);
or U9819 (N_9819,N_4749,N_4048);
xor U9820 (N_9820,N_2631,N_2718);
nor U9821 (N_9821,N_1960,N_1987);
xor U9822 (N_9822,N_342,N_1253);
nor U9823 (N_9823,N_2855,N_3852);
and U9824 (N_9824,N_1643,N_1848);
or U9825 (N_9825,N_2434,N_2756);
or U9826 (N_9826,N_4198,N_4242);
nand U9827 (N_9827,N_4293,N_4483);
nor U9828 (N_9828,N_66,N_3773);
nor U9829 (N_9829,N_3434,N_2268);
nand U9830 (N_9830,N_4654,N_1784);
nand U9831 (N_9831,N_865,N_3131);
xnor U9832 (N_9832,N_4309,N_2883);
xnor U9833 (N_9833,N_2105,N_622);
xor U9834 (N_9834,N_4155,N_2930);
xnor U9835 (N_9835,N_1010,N_828);
nor U9836 (N_9836,N_1774,N_1178);
nor U9837 (N_9837,N_3161,N_4055);
nand U9838 (N_9838,N_251,N_1997);
or U9839 (N_9839,N_1435,N_3574);
nand U9840 (N_9840,N_4949,N_692);
nor U9841 (N_9841,N_814,N_173);
nor U9842 (N_9842,N_2907,N_2254);
nand U9843 (N_9843,N_4923,N_1870);
or U9844 (N_9844,N_2941,N_3509);
nor U9845 (N_9845,N_2150,N_581);
nor U9846 (N_9846,N_1261,N_317);
nor U9847 (N_9847,N_4923,N_3238);
or U9848 (N_9848,N_2580,N_1513);
nor U9849 (N_9849,N_1274,N_167);
or U9850 (N_9850,N_2531,N_3923);
nor U9851 (N_9851,N_4132,N_838);
xor U9852 (N_9852,N_3684,N_3460);
nor U9853 (N_9853,N_3914,N_1481);
or U9854 (N_9854,N_897,N_2705);
nor U9855 (N_9855,N_991,N_3288);
nor U9856 (N_9856,N_3265,N_1598);
xnor U9857 (N_9857,N_2531,N_3889);
nor U9858 (N_9858,N_1100,N_1968);
or U9859 (N_9859,N_4642,N_4693);
or U9860 (N_9860,N_57,N_1649);
nor U9861 (N_9861,N_1221,N_4792);
nand U9862 (N_9862,N_358,N_1711);
nor U9863 (N_9863,N_1916,N_1233);
and U9864 (N_9864,N_2824,N_3636);
and U9865 (N_9865,N_3481,N_3482);
or U9866 (N_9866,N_4788,N_597);
xor U9867 (N_9867,N_723,N_2166);
or U9868 (N_9868,N_1547,N_2966);
or U9869 (N_9869,N_3964,N_2825);
nor U9870 (N_9870,N_1085,N_2643);
or U9871 (N_9871,N_2068,N_2956);
xor U9872 (N_9872,N_527,N_2019);
or U9873 (N_9873,N_3468,N_2792);
and U9874 (N_9874,N_3966,N_804);
and U9875 (N_9875,N_4767,N_3657);
nand U9876 (N_9876,N_4000,N_2168);
and U9877 (N_9877,N_4578,N_3281);
nand U9878 (N_9878,N_634,N_3313);
xor U9879 (N_9879,N_105,N_1731);
and U9880 (N_9880,N_4615,N_401);
and U9881 (N_9881,N_448,N_3610);
xor U9882 (N_9882,N_2602,N_1553);
and U9883 (N_9883,N_104,N_2243);
and U9884 (N_9884,N_1895,N_3853);
nor U9885 (N_9885,N_806,N_984);
and U9886 (N_9886,N_2444,N_4598);
xnor U9887 (N_9887,N_2597,N_3288);
or U9888 (N_9888,N_236,N_1201);
nor U9889 (N_9889,N_1447,N_1483);
and U9890 (N_9890,N_3686,N_4348);
or U9891 (N_9891,N_2472,N_2217);
nor U9892 (N_9892,N_3506,N_1542);
nor U9893 (N_9893,N_1305,N_1928);
nand U9894 (N_9894,N_4669,N_2912);
or U9895 (N_9895,N_645,N_493);
nor U9896 (N_9896,N_2140,N_793);
nand U9897 (N_9897,N_1382,N_2374);
nand U9898 (N_9898,N_4547,N_3166);
or U9899 (N_9899,N_319,N_4502);
and U9900 (N_9900,N_1935,N_525);
and U9901 (N_9901,N_1906,N_1006);
xor U9902 (N_9902,N_4696,N_2695);
nand U9903 (N_9903,N_4043,N_3115);
or U9904 (N_9904,N_3139,N_881);
and U9905 (N_9905,N_2961,N_4689);
nor U9906 (N_9906,N_88,N_1363);
and U9907 (N_9907,N_940,N_2392);
or U9908 (N_9908,N_1209,N_318);
or U9909 (N_9909,N_1943,N_2592);
xor U9910 (N_9910,N_1990,N_2696);
and U9911 (N_9911,N_462,N_2298);
xnor U9912 (N_9912,N_2598,N_2829);
nor U9913 (N_9913,N_1426,N_3001);
xor U9914 (N_9914,N_206,N_3256);
nor U9915 (N_9915,N_4676,N_4207);
xor U9916 (N_9916,N_3553,N_1971);
nor U9917 (N_9917,N_3220,N_892);
xnor U9918 (N_9918,N_3044,N_657);
nand U9919 (N_9919,N_2319,N_711);
and U9920 (N_9920,N_4335,N_4337);
xor U9921 (N_9921,N_2166,N_669);
xor U9922 (N_9922,N_298,N_809);
xor U9923 (N_9923,N_2200,N_1769);
nor U9924 (N_9924,N_3842,N_423);
or U9925 (N_9925,N_3928,N_500);
nand U9926 (N_9926,N_2406,N_1006);
nand U9927 (N_9927,N_4766,N_259);
or U9928 (N_9928,N_3553,N_51);
xnor U9929 (N_9929,N_2220,N_1182);
and U9930 (N_9930,N_1779,N_2328);
or U9931 (N_9931,N_2802,N_4553);
xor U9932 (N_9932,N_4379,N_707);
and U9933 (N_9933,N_1604,N_4824);
xnor U9934 (N_9934,N_2054,N_3756);
nor U9935 (N_9935,N_2672,N_858);
and U9936 (N_9936,N_4394,N_914);
nand U9937 (N_9937,N_125,N_1314);
nor U9938 (N_9938,N_3431,N_2707);
nand U9939 (N_9939,N_2943,N_1316);
or U9940 (N_9940,N_3848,N_3192);
or U9941 (N_9941,N_1501,N_4808);
and U9942 (N_9942,N_864,N_816);
nand U9943 (N_9943,N_3513,N_3264);
nand U9944 (N_9944,N_1231,N_3264);
nand U9945 (N_9945,N_241,N_4778);
or U9946 (N_9946,N_2650,N_476);
and U9947 (N_9947,N_4076,N_840);
nand U9948 (N_9948,N_3924,N_2967);
xnor U9949 (N_9949,N_3427,N_732);
xor U9950 (N_9950,N_2149,N_990);
or U9951 (N_9951,N_304,N_2094);
xnor U9952 (N_9952,N_1397,N_4069);
xnor U9953 (N_9953,N_4052,N_4579);
or U9954 (N_9954,N_2051,N_3377);
and U9955 (N_9955,N_4183,N_3087);
nand U9956 (N_9956,N_2582,N_666);
nor U9957 (N_9957,N_3364,N_4677);
nand U9958 (N_9958,N_2854,N_3667);
xor U9959 (N_9959,N_3006,N_4726);
nand U9960 (N_9960,N_4451,N_3822);
nand U9961 (N_9961,N_4200,N_4373);
xnor U9962 (N_9962,N_975,N_4529);
nor U9963 (N_9963,N_1442,N_4299);
or U9964 (N_9964,N_1121,N_2103);
nand U9965 (N_9965,N_2058,N_540);
and U9966 (N_9966,N_4981,N_1088);
and U9967 (N_9967,N_3989,N_303);
xor U9968 (N_9968,N_4230,N_4463);
and U9969 (N_9969,N_2228,N_1755);
or U9970 (N_9970,N_1790,N_3097);
xnor U9971 (N_9971,N_4108,N_1242);
xnor U9972 (N_9972,N_4163,N_4154);
nor U9973 (N_9973,N_1094,N_2281);
nor U9974 (N_9974,N_3305,N_598);
xnor U9975 (N_9975,N_3475,N_1016);
nand U9976 (N_9976,N_614,N_4877);
xnor U9977 (N_9977,N_1753,N_4830);
xor U9978 (N_9978,N_2356,N_4826);
xnor U9979 (N_9979,N_3855,N_1475);
or U9980 (N_9980,N_406,N_1429);
nor U9981 (N_9981,N_4498,N_1623);
and U9982 (N_9982,N_2092,N_3900);
or U9983 (N_9983,N_429,N_146);
xnor U9984 (N_9984,N_3525,N_3181);
nand U9985 (N_9985,N_302,N_1293);
nor U9986 (N_9986,N_4044,N_4089);
or U9987 (N_9987,N_2129,N_1857);
or U9988 (N_9988,N_3020,N_2773);
or U9989 (N_9989,N_4577,N_3689);
xnor U9990 (N_9990,N_1281,N_2362);
nor U9991 (N_9991,N_4045,N_721);
nand U9992 (N_9992,N_1326,N_186);
nand U9993 (N_9993,N_1489,N_1550);
or U9994 (N_9994,N_619,N_459);
and U9995 (N_9995,N_1236,N_156);
or U9996 (N_9996,N_3035,N_1285);
nor U9997 (N_9997,N_304,N_3857);
nor U9998 (N_9998,N_206,N_3892);
xnor U9999 (N_9999,N_4065,N_4618);
nor U10000 (N_10000,N_9768,N_9317);
nand U10001 (N_10001,N_9981,N_7804);
and U10002 (N_10002,N_9180,N_6530);
and U10003 (N_10003,N_8615,N_9688);
nor U10004 (N_10004,N_6411,N_7100);
and U10005 (N_10005,N_6157,N_6707);
nand U10006 (N_10006,N_5642,N_8184);
or U10007 (N_10007,N_6531,N_9661);
xnor U10008 (N_10008,N_7914,N_8998);
or U10009 (N_10009,N_5677,N_9301);
xor U10010 (N_10010,N_5128,N_9789);
xnor U10011 (N_10011,N_5892,N_7254);
nand U10012 (N_10012,N_6621,N_7979);
xnor U10013 (N_10013,N_7536,N_5152);
nand U10014 (N_10014,N_5590,N_9266);
and U10015 (N_10015,N_8919,N_6589);
nand U10016 (N_10016,N_8338,N_5540);
xor U10017 (N_10017,N_5006,N_9860);
nor U10018 (N_10018,N_9181,N_5557);
and U10019 (N_10019,N_5685,N_8992);
nand U10020 (N_10020,N_9184,N_6058);
xnor U10021 (N_10021,N_7028,N_6034);
or U10022 (N_10022,N_8723,N_8562);
nand U10023 (N_10023,N_5635,N_8162);
nor U10024 (N_10024,N_6973,N_5888);
nor U10025 (N_10025,N_9073,N_8342);
nand U10026 (N_10026,N_6410,N_6808);
xnor U10027 (N_10027,N_9072,N_9047);
nand U10028 (N_10028,N_8747,N_6256);
nand U10029 (N_10029,N_9604,N_5388);
or U10030 (N_10030,N_7431,N_9159);
xnor U10031 (N_10031,N_5970,N_9349);
nor U10032 (N_10032,N_5855,N_9854);
nand U10033 (N_10033,N_8667,N_7751);
nor U10034 (N_10034,N_7374,N_5830);
nand U10035 (N_10035,N_5127,N_5334);
nor U10036 (N_10036,N_5779,N_6997);
xor U10037 (N_10037,N_7604,N_5533);
or U10038 (N_10038,N_9834,N_8971);
and U10039 (N_10039,N_6921,N_5694);
or U10040 (N_10040,N_7112,N_9025);
nor U10041 (N_10041,N_9203,N_7967);
xor U10042 (N_10042,N_5930,N_8076);
nand U10043 (N_10043,N_7455,N_5975);
nor U10044 (N_10044,N_8328,N_5449);
nand U10045 (N_10045,N_5714,N_6265);
xnor U10046 (N_10046,N_9412,N_5534);
nand U10047 (N_10047,N_7192,N_7872);
and U10048 (N_10048,N_7246,N_5638);
or U10049 (N_10049,N_8847,N_9482);
xnor U10050 (N_10050,N_5078,N_7720);
and U10051 (N_10051,N_6364,N_9080);
nor U10052 (N_10052,N_6243,N_7518);
or U10053 (N_10053,N_8395,N_5292);
nand U10054 (N_10054,N_5394,N_9125);
and U10055 (N_10055,N_8004,N_7625);
or U10056 (N_10056,N_7305,N_6879);
nand U10057 (N_10057,N_7996,N_5671);
and U10058 (N_10058,N_9450,N_6992);
and U10059 (N_10059,N_9322,N_5938);
or U10060 (N_10060,N_7560,N_5556);
xnor U10061 (N_10061,N_8127,N_9426);
and U10062 (N_10062,N_5310,N_6732);
and U10063 (N_10063,N_8298,N_7044);
xnor U10064 (N_10064,N_6931,N_5360);
nor U10065 (N_10065,N_7243,N_6886);
nand U10066 (N_10066,N_6587,N_8142);
nor U10067 (N_10067,N_8973,N_7787);
and U10068 (N_10068,N_5357,N_7828);
xnor U10069 (N_10069,N_8085,N_7571);
and U10070 (N_10070,N_9598,N_7497);
nand U10071 (N_10071,N_7249,N_9877);
nor U10072 (N_10072,N_9676,N_6194);
nand U10073 (N_10073,N_7792,N_5336);
nand U10074 (N_10074,N_6214,N_7393);
nand U10075 (N_10075,N_6271,N_7178);
nor U10076 (N_10076,N_5641,N_9919);
nor U10077 (N_10077,N_6618,N_5335);
and U10078 (N_10078,N_6154,N_6081);
and U10079 (N_10079,N_7170,N_6519);
nor U10080 (N_10080,N_6311,N_7578);
or U10081 (N_10081,N_8222,N_6091);
xnor U10082 (N_10082,N_8924,N_8420);
xor U10083 (N_10083,N_6090,N_6834);
or U10084 (N_10084,N_8054,N_7209);
nand U10085 (N_10085,N_9776,N_9762);
or U10086 (N_10086,N_9393,N_9878);
or U10087 (N_10087,N_5002,N_9424);
nor U10088 (N_10088,N_8185,N_5272);
xor U10089 (N_10089,N_7382,N_7826);
xnor U10090 (N_10090,N_9136,N_6987);
or U10091 (N_10091,N_7356,N_6906);
or U10092 (N_10092,N_9015,N_6959);
nand U10093 (N_10093,N_5312,N_8831);
and U10094 (N_10094,N_9248,N_5160);
nand U10095 (N_10095,N_8535,N_9351);
nand U10096 (N_10096,N_5913,N_9137);
xor U10097 (N_10097,N_6257,N_6767);
or U10098 (N_10098,N_9879,N_5765);
and U10099 (N_10099,N_7895,N_7780);
nor U10100 (N_10100,N_5601,N_6596);
or U10101 (N_10101,N_8560,N_6898);
nand U10102 (N_10102,N_6783,N_9871);
nor U10103 (N_10103,N_8801,N_9537);
xnor U10104 (N_10104,N_8122,N_7109);
xnor U10105 (N_10105,N_6466,N_8337);
nor U10106 (N_10106,N_9651,N_5353);
or U10107 (N_10107,N_9019,N_6417);
and U10108 (N_10108,N_7025,N_6447);
and U10109 (N_10109,N_5835,N_9944);
nand U10110 (N_10110,N_9416,N_7355);
or U10111 (N_10111,N_7221,N_8216);
xor U10112 (N_10112,N_9131,N_5223);
and U10113 (N_10113,N_8452,N_6473);
and U10114 (N_10114,N_5481,N_6831);
nand U10115 (N_10115,N_5964,N_8611);
xnor U10116 (N_10116,N_6538,N_8997);
xnor U10117 (N_10117,N_6747,N_6163);
nand U10118 (N_10118,N_6375,N_5675);
or U10119 (N_10119,N_9826,N_5375);
nor U10120 (N_10120,N_7897,N_7181);
nand U10121 (N_10121,N_9990,N_8379);
xnor U10122 (N_10122,N_5246,N_8412);
nor U10123 (N_10123,N_5212,N_7291);
and U10124 (N_10124,N_8273,N_9237);
nor U10125 (N_10125,N_6757,N_5242);
and U10126 (N_10126,N_9547,N_9198);
nand U10127 (N_10127,N_8920,N_8211);
and U10128 (N_10128,N_8171,N_7389);
nor U10129 (N_10129,N_9512,N_7763);
or U10130 (N_10130,N_6526,N_7615);
nand U10131 (N_10131,N_7327,N_6175);
nand U10132 (N_10132,N_9880,N_5528);
or U10133 (N_10133,N_7885,N_5281);
xnor U10134 (N_10134,N_5553,N_6843);
or U10135 (N_10135,N_9507,N_6288);
xnor U10136 (N_10136,N_6598,N_6093);
nand U10137 (N_10137,N_5185,N_9590);
and U10138 (N_10138,N_9617,N_8866);
and U10139 (N_10139,N_6019,N_9001);
xnor U10140 (N_10140,N_5796,N_5509);
and U10141 (N_10141,N_6160,N_7513);
nand U10142 (N_10142,N_8303,N_7328);
nand U10143 (N_10143,N_6405,N_5674);
nand U10144 (N_10144,N_8626,N_8652);
xor U10145 (N_10145,N_8900,N_5931);
nand U10146 (N_10146,N_5555,N_9387);
xnor U10147 (N_10147,N_6941,N_6867);
xnor U10148 (N_10148,N_9295,N_5118);
xor U10149 (N_10149,N_8887,N_5434);
or U10150 (N_10150,N_5395,N_6200);
nor U10151 (N_10151,N_8729,N_8341);
or U10152 (N_10152,N_9844,N_6728);
xor U10153 (N_10153,N_7095,N_6646);
nand U10154 (N_10154,N_8755,N_7592);
or U10155 (N_10155,N_9693,N_9551);
nand U10156 (N_10156,N_6491,N_7313);
or U10157 (N_10157,N_7941,N_6020);
nand U10158 (N_10158,N_6448,N_8218);
nor U10159 (N_10159,N_9908,N_5278);
xnor U10160 (N_10160,N_6320,N_9925);
nand U10161 (N_10161,N_8650,N_9913);
nand U10162 (N_10162,N_8225,N_8721);
nand U10163 (N_10163,N_5010,N_7739);
xor U10164 (N_10164,N_7390,N_8367);
and U10165 (N_10165,N_8763,N_6030);
or U10166 (N_10166,N_9898,N_9696);
xor U10167 (N_10167,N_7676,N_8491);
and U10168 (N_10168,N_5709,N_6292);
or U10169 (N_10169,N_7117,N_8619);
or U10170 (N_10170,N_6610,N_6450);
and U10171 (N_10171,N_8289,N_6104);
or U10172 (N_10172,N_9583,N_8479);
and U10173 (N_10173,N_6310,N_8196);
nand U10174 (N_10174,N_5700,N_7013);
or U10175 (N_10175,N_5898,N_9704);
xor U10176 (N_10176,N_5932,N_6439);
nand U10177 (N_10177,N_9397,N_9709);
and U10178 (N_10178,N_7980,N_8709);
or U10179 (N_10179,N_8457,N_5844);
nand U10180 (N_10180,N_5494,N_5114);
xnor U10181 (N_10181,N_5268,N_6655);
nor U10182 (N_10182,N_7774,N_5056);
nand U10183 (N_10183,N_6167,N_6472);
nor U10184 (N_10184,N_5724,N_6343);
or U10185 (N_10185,N_8017,N_6703);
xor U10186 (N_10186,N_6438,N_7679);
xnor U10187 (N_10187,N_6823,N_7907);
and U10188 (N_10188,N_6877,N_5754);
xor U10189 (N_10189,N_9999,N_6348);
or U10190 (N_10190,N_6952,N_6219);
and U10191 (N_10191,N_7363,N_8348);
nand U10192 (N_10192,N_8632,N_7434);
or U10193 (N_10193,N_5066,N_7075);
nor U10194 (N_10194,N_8829,N_9660);
nand U10195 (N_10195,N_7517,N_9356);
nor U10196 (N_10196,N_8025,N_5804);
nor U10197 (N_10197,N_9865,N_7285);
and U10198 (N_10198,N_5057,N_9057);
or U10199 (N_10199,N_8439,N_8096);
and U10200 (N_10200,N_6443,N_8056);
nor U10201 (N_10201,N_9020,N_9851);
nand U10202 (N_10202,N_5839,N_7801);
nor U10203 (N_10203,N_8679,N_5093);
and U10204 (N_10204,N_6100,N_9307);
and U10205 (N_10205,N_9143,N_7778);
or U10206 (N_10206,N_8346,N_6112);
and U10207 (N_10207,N_7712,N_9639);
xor U10208 (N_10208,N_5381,N_6077);
or U10209 (N_10209,N_5045,N_9765);
and U10210 (N_10210,N_5291,N_8411);
xnor U10211 (N_10211,N_5123,N_9933);
nand U10212 (N_10212,N_9366,N_6361);
nor U10213 (N_10213,N_6687,N_7407);
nand U10214 (N_10214,N_9570,N_5202);
nor U10215 (N_10215,N_6520,N_7096);
or U10216 (N_10216,N_9461,N_7334);
xor U10217 (N_10217,N_5860,N_7397);
and U10218 (N_10218,N_6553,N_9384);
xor U10219 (N_10219,N_6057,N_6558);
nand U10220 (N_10220,N_8882,N_7820);
or U10221 (N_10221,N_7522,N_5462);
or U10222 (N_10222,N_9050,N_9953);
or U10223 (N_10223,N_5595,N_8953);
nand U10224 (N_10224,N_7053,N_8767);
and U10225 (N_10225,N_5684,N_8204);
or U10226 (N_10226,N_5774,N_6678);
and U10227 (N_10227,N_9297,N_7038);
or U10228 (N_10228,N_7071,N_9697);
nor U10229 (N_10229,N_9627,N_9827);
xnor U10230 (N_10230,N_5001,N_8373);
nor U10231 (N_10231,N_7198,N_8871);
nor U10232 (N_10232,N_5717,N_8195);
and U10233 (N_10233,N_7590,N_9171);
xor U10234 (N_10234,N_5900,N_5289);
nor U10235 (N_10235,N_6393,N_7557);
xor U10236 (N_10236,N_9669,N_9973);
or U10237 (N_10237,N_7087,N_8711);
and U10238 (N_10238,N_7951,N_5872);
or U10239 (N_10239,N_9622,N_8790);
or U10240 (N_10240,N_9935,N_7311);
and U10241 (N_10241,N_9152,N_6717);
xor U10242 (N_10242,N_5654,N_7974);
nor U10243 (N_10243,N_7015,N_5859);
and U10244 (N_10244,N_9090,N_8945);
and U10245 (N_10245,N_6305,N_8212);
nor U10246 (N_10246,N_8727,N_6825);
or U10247 (N_10247,N_7594,N_7149);
nor U10248 (N_10248,N_7770,N_7846);
and U10249 (N_10249,N_7890,N_9846);
nand U10250 (N_10250,N_6430,N_5981);
or U10251 (N_10251,N_9600,N_8016);
or U10252 (N_10252,N_6000,N_8362);
nor U10253 (N_10253,N_7860,N_9138);
and U10254 (N_10254,N_9443,N_6208);
and U10255 (N_10255,N_9216,N_9040);
nor U10256 (N_10256,N_7202,N_5230);
xnor U10257 (N_10257,N_8000,N_9031);
nor U10258 (N_10258,N_9611,N_9597);
nand U10259 (N_10259,N_5258,N_8179);
or U10260 (N_10260,N_8116,N_9772);
nand U10261 (N_10261,N_8978,N_7638);
or U10262 (N_10262,N_6778,N_8365);
xor U10263 (N_10263,N_8715,N_5541);
nor U10264 (N_10264,N_7191,N_9787);
nand U10265 (N_10265,N_8297,N_6578);
xor U10266 (N_10266,N_8284,N_6171);
or U10267 (N_10267,N_6894,N_9733);
nor U10268 (N_10268,N_8778,N_7495);
and U10269 (N_10269,N_5234,N_9148);
xnor U10270 (N_10270,N_5990,N_6691);
and U10271 (N_10271,N_7000,N_9228);
and U10272 (N_10272,N_6087,N_5323);
and U10273 (N_10273,N_9529,N_6359);
and U10274 (N_10274,N_9921,N_9308);
or U10275 (N_10275,N_9417,N_5593);
nor U10276 (N_10276,N_6927,N_9304);
or U10277 (N_10277,N_7637,N_7174);
xor U10278 (N_10278,N_9711,N_9166);
xor U10279 (N_10279,N_9499,N_6713);
nor U10280 (N_10280,N_7460,N_6527);
nor U10281 (N_10281,N_5411,N_8524);
nor U10282 (N_10282,N_5708,N_5822);
and U10283 (N_10283,N_8481,N_5021);
nor U10284 (N_10284,N_9315,N_5924);
nand U10285 (N_10285,N_7268,N_7569);
and U10286 (N_10286,N_6571,N_9847);
nand U10287 (N_10287,N_7290,N_5703);
nand U10288 (N_10288,N_5226,N_5348);
nor U10289 (N_10289,N_8570,N_5618);
nand U10290 (N_10290,N_9059,N_9657);
nor U10291 (N_10291,N_6739,N_7292);
xnor U10292 (N_10292,N_9717,N_6037);
and U10293 (N_10293,N_6164,N_9608);
or U10294 (N_10294,N_6442,N_8423);
nor U10295 (N_10295,N_9823,N_9036);
nand U10296 (N_10296,N_8340,N_6561);
nor U10297 (N_10297,N_6124,N_6948);
nor U10298 (N_10298,N_6401,N_8509);
nor U10299 (N_10299,N_8386,N_5018);
and U10300 (N_10300,N_5795,N_5472);
or U10301 (N_10301,N_7107,N_8701);
nor U10302 (N_10302,N_9386,N_5178);
nand U10303 (N_10303,N_6501,N_6661);
xor U10304 (N_10304,N_9883,N_5768);
or U10305 (N_10305,N_6052,N_6696);
and U10306 (N_10306,N_7915,N_6727);
nand U10307 (N_10307,N_9543,N_7866);
or U10308 (N_10308,N_6239,N_9432);
nand U10309 (N_10309,N_8482,N_9361);
and U10310 (N_10310,N_7151,N_7725);
nor U10311 (N_10311,N_7958,N_9100);
nand U10312 (N_10312,N_6882,N_9338);
or U10313 (N_10313,N_8514,N_9261);
nor U10314 (N_10314,N_6299,N_9803);
xor U10315 (N_10315,N_5342,N_8772);
nor U10316 (N_10316,N_5393,N_5535);
nor U10317 (N_10317,N_8664,N_7534);
and U10318 (N_10318,N_9993,N_8084);
nand U10319 (N_10319,N_7591,N_8425);
nand U10320 (N_10320,N_9625,N_9016);
and U10321 (N_10321,N_5794,N_9656);
or U10322 (N_10322,N_6762,N_9235);
and U10323 (N_10323,N_9449,N_9948);
and U10324 (N_10324,N_7500,N_6435);
or U10325 (N_10325,N_7934,N_9044);
and U10326 (N_10326,N_8534,N_5518);
xnor U10327 (N_10327,N_8589,N_5364);
and U10328 (N_10328,N_8990,N_5440);
and U10329 (N_10329,N_7420,N_6666);
nand U10330 (N_10330,N_5179,N_5994);
and U10331 (N_10331,N_6805,N_5792);
xnor U10332 (N_10332,N_7027,N_5505);
xnor U10333 (N_10333,N_7546,N_9634);
or U10334 (N_10334,N_6920,N_7841);
or U10335 (N_10335,N_8832,N_8005);
xor U10336 (N_10336,N_5391,N_6204);
xor U10337 (N_10337,N_9911,N_8811);
nand U10338 (N_10338,N_5044,N_8272);
nor U10339 (N_10339,N_9623,N_7299);
nand U10340 (N_10340,N_7115,N_7396);
and U10341 (N_10341,N_8666,N_7484);
xnor U10342 (N_10342,N_6181,N_9348);
or U10343 (N_10343,N_8550,N_7066);
xor U10344 (N_10344,N_9299,N_7714);
or U10345 (N_10345,N_9952,N_5250);
or U10346 (N_10346,N_9637,N_8549);
nand U10347 (N_10347,N_6990,N_8880);
nand U10348 (N_10348,N_8132,N_6830);
xnor U10349 (N_10349,N_9609,N_5124);
xor U10350 (N_10350,N_6721,N_6695);
or U10351 (N_10351,N_5162,N_7579);
or U10352 (N_10352,N_7375,N_7671);
and U10353 (N_10353,N_7039,N_8192);
nand U10354 (N_10354,N_8969,N_6564);
xor U10355 (N_10355,N_6741,N_8818);
and U10356 (N_10356,N_9343,N_6807);
nand U10357 (N_10357,N_8639,N_6441);
xor U10358 (N_10358,N_9647,N_6001);
xor U10359 (N_10359,N_9858,N_5279);
and U10360 (N_10360,N_9177,N_9089);
nand U10361 (N_10361,N_9283,N_7807);
xnor U10362 (N_10362,N_9538,N_6746);
and U10363 (N_10363,N_7628,N_5038);
nor U10364 (N_10364,N_8935,N_9968);
nand U10365 (N_10365,N_9144,N_8143);
nor U10366 (N_10366,N_8984,N_8051);
xnor U10367 (N_10367,N_8636,N_8938);
xor U10368 (N_10368,N_9402,N_8508);
xor U10369 (N_10369,N_5565,N_8910);
nor U10370 (N_10370,N_8922,N_6337);
nand U10371 (N_10371,N_6550,N_6813);
nand U10372 (N_10372,N_7861,N_6709);
nor U10373 (N_10373,N_6437,N_5101);
nand U10374 (N_10374,N_9553,N_7364);
xor U10375 (N_10375,N_9884,N_8609);
nand U10376 (N_10376,N_6567,N_5487);
nor U10377 (N_10377,N_8513,N_8069);
xnor U10378 (N_10378,N_9404,N_9903);
xnor U10379 (N_10379,N_6766,N_8546);
nand U10380 (N_10380,N_8925,N_7554);
xnor U10381 (N_10381,N_6743,N_9197);
or U10382 (N_10382,N_6047,N_8704);
nor U10383 (N_10383,N_9747,N_8307);
and U10384 (N_10384,N_8561,N_8392);
xor U10385 (N_10385,N_7539,N_6493);
xor U10386 (N_10386,N_5524,N_7694);
and U10387 (N_10387,N_8287,N_9066);
and U10388 (N_10388,N_6115,N_5222);
and U10389 (N_10389,N_7678,N_9009);
or U10390 (N_10390,N_9629,N_5425);
xor U10391 (N_10391,N_6988,N_6017);
nand U10392 (N_10392,N_5271,N_5899);
or U10393 (N_10393,N_8898,N_8187);
or U10394 (N_10394,N_6335,N_9668);
or U10395 (N_10395,N_6933,N_9620);
or U10396 (N_10396,N_8158,N_7666);
nand U10397 (N_10397,N_7667,N_8045);
and U10398 (N_10398,N_7796,N_8417);
and U10399 (N_10399,N_9905,N_5568);
nor U10400 (N_10400,N_9749,N_6652);
or U10401 (N_10401,N_5298,N_7810);
nor U10402 (N_10402,N_6424,N_5877);
and U10403 (N_10403,N_6094,N_7506);
and U10404 (N_10404,N_5682,N_7378);
and U10405 (N_10405,N_7600,N_9396);
or U10406 (N_10406,N_7701,N_9147);
and U10407 (N_10407,N_8761,N_6366);
or U10408 (N_10408,N_7352,N_7092);
nand U10409 (N_10409,N_8011,N_5052);
nand U10410 (N_10410,N_8872,N_7783);
nand U10411 (N_10411,N_8419,N_9335);
nor U10412 (N_10412,N_6462,N_6718);
nand U10413 (N_10413,N_8435,N_8219);
or U10414 (N_10414,N_7972,N_8857);
nand U10415 (N_10415,N_8776,N_9061);
and U10416 (N_10416,N_8201,N_7805);
and U10417 (N_10417,N_9729,N_7247);
and U10418 (N_10418,N_5960,N_9459);
xor U10419 (N_10419,N_7983,N_6016);
or U10420 (N_10420,N_8932,N_5484);
and U10421 (N_10421,N_6399,N_9024);
nand U10422 (N_10422,N_7830,N_8533);
and U10423 (N_10423,N_6412,N_8853);
and U10424 (N_10424,N_5756,N_5126);
or U10425 (N_10425,N_7938,N_9435);
xnor U10426 (N_10426,N_8391,N_7135);
and U10427 (N_10427,N_7643,N_7614);
nor U10428 (N_10428,N_9423,N_9849);
or U10429 (N_10429,N_6372,N_9246);
and U10430 (N_10430,N_5463,N_5547);
xnor U10431 (N_10431,N_5752,N_9215);
and U10432 (N_10432,N_5785,N_5125);
nand U10433 (N_10433,N_9503,N_6475);
nor U10434 (N_10434,N_9521,N_6794);
nor U10435 (N_10435,N_7239,N_6929);
xnor U10436 (N_10436,N_8121,N_7128);
nand U10437 (N_10437,N_8764,N_8891);
nor U10438 (N_10438,N_6351,N_6280);
xor U10439 (N_10439,N_7521,N_5000);
and U10440 (N_10440,N_6195,N_9172);
or U10441 (N_10441,N_5581,N_8208);
nand U10442 (N_10442,N_5798,N_5766);
and U10443 (N_10443,N_7674,N_8699);
and U10444 (N_10444,N_7006,N_6029);
xnor U10445 (N_10445,N_6580,N_5221);
nor U10446 (N_10446,N_6733,N_7881);
nand U10447 (N_10447,N_8175,N_8041);
or U10448 (N_10448,N_6658,N_9243);
nor U10449 (N_10449,N_7966,N_5801);
nor U10450 (N_10450,N_7745,N_6905);
and U10451 (N_10451,N_5154,N_7704);
and U10452 (N_10452,N_6777,N_7058);
nor U10453 (N_10453,N_5492,N_6428);
or U10454 (N_10454,N_8731,N_6789);
and U10455 (N_10455,N_6541,N_7632);
nand U10456 (N_10456,N_6704,N_8985);
nor U10457 (N_10457,N_5843,N_6619);
xor U10458 (N_10458,N_7036,N_8518);
and U10459 (N_10459,N_8948,N_8689);
nor U10460 (N_10460,N_8266,N_8629);
nand U10461 (N_10461,N_6600,N_6773);
nor U10462 (N_10462,N_6407,N_9818);
xnor U10463 (N_10463,N_6607,N_9202);
or U10464 (N_10464,N_7509,N_5090);
or U10465 (N_10465,N_8282,N_9506);
nand U10466 (N_10466,N_7410,N_6021);
nand U10467 (N_10467,N_5163,N_8490);
xor U10468 (N_10468,N_5338,N_6007);
and U10469 (N_10469,N_8178,N_8565);
and U10470 (N_10470,N_9186,N_5315);
or U10471 (N_10471,N_5940,N_6268);
xnor U10472 (N_10472,N_7953,N_9900);
and U10473 (N_10473,N_8169,N_7472);
nor U10474 (N_10474,N_9170,N_6196);
xor U10475 (N_10475,N_8241,N_7411);
and U10476 (N_10476,N_5770,N_7492);
nor U10477 (N_10477,N_6919,N_5059);
nand U10478 (N_10478,N_9411,N_6820);
or U10479 (N_10479,N_9219,N_8726);
or U10480 (N_10480,N_9064,N_5005);
and U10481 (N_10481,N_7722,N_7899);
nand U10482 (N_10482,N_8724,N_8564);
nor U10483 (N_10483,N_8941,N_9855);
nor U10484 (N_10484,N_6464,N_9682);
nor U10485 (N_10485,N_8775,N_8129);
or U10486 (N_10486,N_6370,N_8955);
or U10487 (N_10487,N_9808,N_8140);
or U10488 (N_10488,N_6603,N_5365);
or U10489 (N_10489,N_5190,N_8936);
and U10490 (N_10490,N_8263,N_5749);
xnor U10491 (N_10491,N_8505,N_5946);
xor U10492 (N_10492,N_7216,N_8274);
xor U10493 (N_10493,N_6285,N_6753);
xnor U10494 (N_10494,N_7180,N_5396);
nand U10495 (N_10495,N_6858,N_6302);
nand U10496 (N_10496,N_5934,N_8083);
or U10497 (N_10497,N_6504,N_5971);
nor U10498 (N_10498,N_5367,N_7868);
and U10499 (N_10499,N_7991,N_7296);
nand U10500 (N_10500,N_8237,N_6188);
nor U10501 (N_10501,N_5718,N_7857);
nor U10502 (N_10502,N_5870,N_8962);
nand U10503 (N_10503,N_8052,N_8540);
and U10504 (N_10504,N_8112,N_9672);
xor U10505 (N_10505,N_5401,N_5606);
and U10506 (N_10506,N_7283,N_9519);
and U10507 (N_10507,N_8058,N_6189);
and U10508 (N_10508,N_9328,N_9923);
and U10509 (N_10509,N_6436,N_7345);
nand U10510 (N_10510,N_7839,N_5976);
and U10511 (N_10511,N_8261,N_6977);
and U10512 (N_10512,N_5742,N_8343);
and U10513 (N_10513,N_7954,N_7329);
nor U10514 (N_10514,N_8576,N_6011);
xor U10515 (N_10515,N_8408,N_5112);
nor U10516 (N_10516,N_9980,N_7700);
or U10517 (N_10517,N_6946,N_8015);
and U10518 (N_10518,N_6734,N_9093);
nand U10519 (N_10519,N_7888,N_6145);
xor U10520 (N_10520,N_6720,N_8257);
nor U10521 (N_10521,N_8840,N_8108);
xnor U10522 (N_10522,N_5175,N_7084);
nand U10523 (N_10523,N_5790,N_7023);
or U10524 (N_10524,N_6486,N_6455);
xnor U10525 (N_10525,N_5414,N_8447);
and U10526 (N_10526,N_6862,N_9941);
nor U10527 (N_10527,N_5259,N_6008);
xnor U10528 (N_10528,N_8047,N_6759);
nand U10529 (N_10529,N_9485,N_5390);
xor U10530 (N_10530,N_7186,N_6131);
nand U10531 (N_10531,N_7267,N_9516);
and U10532 (N_10532,N_8707,N_9954);
nand U10533 (N_10533,N_8104,N_6365);
nand U10534 (N_10534,N_7948,N_6184);
or U10535 (N_10535,N_8681,N_8319);
or U10536 (N_10536,N_6573,N_7514);
nor U10537 (N_10537,N_9117,N_8106);
and U10538 (N_10538,N_7445,N_9195);
or U10539 (N_10539,N_5072,N_9643);
nand U10540 (N_10540,N_9675,N_6075);
nand U10541 (N_10541,N_7964,N_7476);
nor U10542 (N_10542,N_6729,N_8013);
xnor U10543 (N_10543,N_6845,N_6606);
nand U10544 (N_10544,N_9010,N_5397);
or U10545 (N_10545,N_6431,N_9685);
xnor U10546 (N_10546,N_5270,N_6318);
nand U10547 (N_10547,N_8697,N_5139);
or U10548 (N_10548,N_7037,N_6765);
nand U10549 (N_10549,N_9500,N_7556);
xnor U10550 (N_10550,N_9885,N_7924);
and U10551 (N_10551,N_9875,N_5817);
and U10552 (N_10552,N_9571,N_8437);
xor U10553 (N_10553,N_8039,N_8306);
nor U10554 (N_10554,N_5490,N_7898);
or U10555 (N_10555,N_6193,N_7106);
nor U10556 (N_10556,N_8455,N_7438);
nor U10557 (N_10557,N_7611,N_5187);
xnor U10558 (N_10558,N_7633,N_5953);
nor U10559 (N_10559,N_8765,N_6601);
nor U10560 (N_10560,N_8888,N_5753);
xnor U10561 (N_10561,N_6649,N_8700);
and U10562 (N_10562,N_5110,N_7761);
and U10563 (N_10563,N_8098,N_9588);
xor U10564 (N_10564,N_5213,N_7682);
and U10565 (N_10565,N_7394,N_5084);
xnor U10566 (N_10566,N_7064,N_5485);
or U10567 (N_10567,N_5659,N_9870);
xor U10568 (N_10568,N_6056,N_7965);
nor U10569 (N_10569,N_9560,N_5514);
or U10570 (N_10570,N_6908,N_6252);
and U10571 (N_10571,N_5634,N_6489);
nor U10572 (N_10572,N_5710,N_6488);
xnor U10573 (N_10573,N_6545,N_7373);
nor U10574 (N_10574,N_6151,N_5895);
or U10575 (N_10575,N_9983,N_7185);
and U10576 (N_10576,N_6426,N_8376);
xnor U10577 (N_10577,N_5302,N_7265);
or U10578 (N_10578,N_7223,N_7046);
nor U10579 (N_10579,N_5183,N_6229);
and U10580 (N_10580,N_9906,N_8344);
or U10581 (N_10581,N_9201,N_6612);
nor U10582 (N_10582,N_7508,N_5917);
nor U10583 (N_10583,N_5444,N_8139);
nor U10584 (N_10584,N_6631,N_5379);
xnor U10585 (N_10585,N_5751,N_9873);
nor U10586 (N_10586,N_8145,N_8050);
and U10587 (N_10587,N_8165,N_6686);
nor U10588 (N_10588,N_8057,N_7850);
and U10589 (N_10589,N_8680,N_9223);
and U10590 (N_10590,N_8993,N_5074);
or U10591 (N_10591,N_6677,N_7147);
xnor U10592 (N_10592,N_8149,N_7368);
and U10593 (N_10593,N_7496,N_5207);
or U10594 (N_10594,N_7994,N_9413);
or U10595 (N_10595,N_5085,N_8913);
and U10596 (N_10596,N_7094,N_7727);
xnor U10597 (N_10597,N_6918,N_6383);
xnor U10598 (N_10598,N_7755,N_7901);
and U10599 (N_10599,N_5341,N_7498);
nand U10600 (N_10600,N_8504,N_6497);
xor U10601 (N_10601,N_7875,N_9452);
xor U10602 (N_10602,N_5297,N_9638);
and U10603 (N_10603,N_9751,N_9679);
or U10604 (N_10604,N_5103,N_7806);
and U10605 (N_10605,N_5285,N_9715);
and U10606 (N_10606,N_7813,N_5427);
nor U10607 (N_10607,N_7256,N_8231);
and U10608 (N_10608,N_9641,N_5113);
nor U10609 (N_10609,N_5430,N_5906);
or U10610 (N_10610,N_8279,N_5003);
nand U10611 (N_10611,N_5108,N_7440);
nor U10612 (N_10612,N_7098,N_9850);
or U10613 (N_10613,N_5412,N_6636);
xor U10614 (N_10614,N_9501,N_6150);
nor U10615 (N_10615,N_6590,N_5173);
xor U10616 (N_10616,N_7210,N_6764);
nand U10617 (N_10617,N_5918,N_5923);
nor U10618 (N_10618,N_8494,N_5846);
nor U10619 (N_10619,N_9213,N_6408);
nor U10620 (N_10620,N_7733,N_7136);
or U10621 (N_10621,N_7258,N_6889);
nand U10622 (N_10622,N_9326,N_8663);
xor U10623 (N_10623,N_6785,N_8506);
and U10624 (N_10624,N_5224,N_6819);
nand U10625 (N_10625,N_5215,N_9294);
or U10626 (N_10626,N_9777,N_5554);
or U10627 (N_10627,N_6585,N_5043);
or U10628 (N_10628,N_7320,N_9401);
or U10629 (N_10629,N_5382,N_5570);
nor U10630 (N_10630,N_7728,N_5466);
or U10631 (N_10631,N_6331,N_7419);
xnor U10632 (N_10632,N_9891,N_6779);
and U10633 (N_10633,N_7226,N_5061);
nor U10634 (N_10634,N_9788,N_5419);
or U10635 (N_10635,N_7681,N_9007);
nor U10636 (N_10636,N_7273,N_7260);
nand U10637 (N_10637,N_8507,N_5189);
or U10638 (N_10638,N_8965,N_7929);
or U10639 (N_10639,N_7623,N_5167);
or U10640 (N_10640,N_5197,N_6847);
nor U10641 (N_10641,N_7491,N_7781);
and U10642 (N_10642,N_9385,N_9899);
or U10643 (N_10643,N_6515,N_5973);
nand U10644 (N_10644,N_6367,N_6683);
nor U10645 (N_10645,N_6900,N_8862);
and U10646 (N_10646,N_7634,N_9610);
nor U10647 (N_10647,N_9209,N_9782);
nand U10648 (N_10648,N_9454,N_7433);
and U10649 (N_10649,N_9277,N_6199);
xnor U10650 (N_10650,N_9965,N_8323);
nand U10651 (N_10651,N_6688,N_5542);
nor U10652 (N_10652,N_7586,N_5022);
xor U10653 (N_10653,N_5275,N_8363);
nor U10654 (N_10654,N_6849,N_6025);
nand U10655 (N_10655,N_8656,N_9271);
and U10656 (N_10656,N_5713,N_7130);
and U10657 (N_10657,N_5543,N_9798);
xor U10658 (N_10658,N_6995,N_8690);
nand U10659 (N_10659,N_5020,N_6735);
xnor U10660 (N_10660,N_7910,N_6960);
and U10661 (N_10661,N_9596,N_5984);
nand U10662 (N_10662,N_8038,N_9577);
xor U10663 (N_10663,N_5455,N_8559);
xor U10664 (N_10664,N_8557,N_7886);
nor U10665 (N_10665,N_9800,N_8027);
nor U10666 (N_10666,N_8421,N_7162);
nand U10667 (N_10667,N_6312,N_7335);
xor U10668 (N_10668,N_7482,N_7403);
nor U10669 (N_10669,N_9951,N_9528);
and U10670 (N_10670,N_9947,N_7575);
and U10671 (N_10671,N_6148,N_9146);
nand U10672 (N_10672,N_7713,N_8465);
or U10673 (N_10673,N_5893,N_8023);
nor U10674 (N_10674,N_5587,N_7920);
and U10675 (N_10675,N_5823,N_8812);
or U10676 (N_10676,N_8625,N_5767);
and U10677 (N_10677,N_6176,N_5456);
nor U10678 (N_10678,N_6962,N_6485);
nand U10679 (N_10679,N_8159,N_7322);
and U10680 (N_10680,N_5992,N_5636);
or U10681 (N_10681,N_6211,N_9584);
or U10682 (N_10682,N_8428,N_6134);
or U10683 (N_10683,N_7609,N_9058);
or U10684 (N_10684,N_8695,N_7748);
and U10685 (N_10685,N_8610,N_7655);
xor U10686 (N_10686,N_8368,N_8708);
and U10687 (N_10687,N_5235,N_8033);
or U10688 (N_10688,N_7999,N_7332);
xnor U10689 (N_10689,N_5939,N_6063);
and U10690 (N_10690,N_9303,N_5157);
nor U10691 (N_10691,N_5878,N_7836);
nand U10692 (N_10692,N_7424,N_9559);
nand U10693 (N_10693,N_8865,N_9579);
nand U10694 (N_10694,N_6220,N_5443);
nor U10695 (N_10695,N_9876,N_6775);
or U10696 (N_10696,N_8809,N_7931);
nor U10697 (N_10697,N_5459,N_5837);
nand U10698 (N_10698,N_6719,N_5191);
or U10699 (N_10699,N_7159,N_7458);
and U10700 (N_10700,N_5177,N_8281);
and U10701 (N_10701,N_5529,N_7589);
nor U10702 (N_10702,N_9262,N_5603);
nor U10703 (N_10703,N_5827,N_8080);
or U10704 (N_10704,N_5783,N_9567);
and U10705 (N_10705,N_9451,N_5260);
nor U10706 (N_10706,N_9476,N_7385);
nor U10707 (N_10707,N_9801,N_7118);
xor U10708 (N_10708,N_6066,N_5182);
nor U10709 (N_10709,N_9646,N_6106);
nor U10710 (N_10710,N_7809,N_9273);
or U10711 (N_10711,N_8471,N_7963);
nand U10712 (N_10712,N_7082,N_6521);
nand U10713 (N_10713,N_6332,N_9644);
or U10714 (N_10714,N_8335,N_7222);
and U10715 (N_10715,N_6935,N_6137);
and U10716 (N_10716,N_8097,N_6110);
or U10717 (N_10717,N_6274,N_7309);
and U10718 (N_10718,N_8583,N_7636);
or U10719 (N_10719,N_9409,N_8845);
or U10720 (N_10720,N_7163,N_6236);
or U10721 (N_10721,N_5284,N_6223);
or U10722 (N_10722,N_7673,N_9909);
or U10723 (N_10723,N_8065,N_6179);
nand U10724 (N_10724,N_7703,N_8907);
and U10725 (N_10725,N_7702,N_7133);
nor U10726 (N_10726,N_6432,N_7940);
xor U10727 (N_10727,N_7050,N_8377);
or U10728 (N_10728,N_8986,N_8644);
xor U10729 (N_10729,N_8624,N_9220);
and U10730 (N_10730,N_6770,N_6290);
xnor U10731 (N_10731,N_5987,N_6357);
nor U10732 (N_10732,N_9975,N_6197);
nand U10733 (N_10733,N_5165,N_6934);
xnor U10734 (N_10734,N_8813,N_5612);
nand U10735 (N_10735,N_6963,N_7357);
xor U10736 (N_10736,N_5032,N_6287);
or U10737 (N_10737,N_8299,N_6391);
nand U10738 (N_10738,N_8008,N_8804);
nor U10739 (N_10739,N_8749,N_8905);
and U10740 (N_10740,N_8841,N_7652);
xnor U10741 (N_10741,N_5600,N_9189);
nor U10742 (N_10742,N_5115,N_7777);
and U10743 (N_10743,N_7630,N_6301);
xnor U10744 (N_10744,N_8133,N_6002);
xor U10745 (N_10745,N_9440,N_9422);
and U10746 (N_10746,N_7173,N_7797);
xor U10747 (N_10747,N_6769,N_5969);
xnor U10748 (N_10748,N_8669,N_8734);
or U10749 (N_10749,N_6062,N_7892);
nor U10750 (N_10750,N_9667,N_9406);
nor U10751 (N_10751,N_9889,N_9008);
nand U10752 (N_10752,N_9760,N_5004);
or U10753 (N_10753,N_7194,N_6989);
or U10754 (N_10754,N_9564,N_5512);
xor U10755 (N_10755,N_5399,N_7869);
or U10756 (N_10756,N_6141,N_8600);
or U10757 (N_10757,N_7388,N_6629);
xnor U10758 (N_10758,N_9939,N_6951);
xor U10759 (N_10759,N_6284,N_9241);
xor U10760 (N_10760,N_6868,N_7443);
and U10761 (N_10761,N_7879,N_9103);
nand U10762 (N_10762,N_6654,N_8259);
or U10763 (N_10763,N_7552,N_6552);
nor U10764 (N_10764,N_7852,N_8779);
xnor U10765 (N_10765,N_5013,N_7183);
nand U10766 (N_10766,N_8136,N_5404);
nand U10767 (N_10767,N_8488,N_8703);
and U10768 (N_10768,N_6048,N_6013);
nor U10769 (N_10769,N_5225,N_6912);
and U10770 (N_10770,N_7475,N_7289);
nor U10771 (N_10771,N_9244,N_6043);
or U10772 (N_10772,N_5922,N_8168);
nor U10773 (N_10773,N_7812,N_5951);
and U10774 (N_10774,N_9523,N_7212);
nor U10775 (N_10775,N_7052,N_5778);
and U10776 (N_10776,N_5428,N_6096);
or U10777 (N_10777,N_5429,N_5145);
nand U10778 (N_10778,N_7838,N_9395);
or U10779 (N_10779,N_5611,N_5623);
and U10780 (N_10780,N_8808,N_5998);
and U10781 (N_10781,N_5009,N_9522);
nand U10782 (N_10782,N_5627,N_6574);
and U10783 (N_10783,N_7610,N_7776);
xnor U10784 (N_10784,N_5324,N_5451);
xnor U10785 (N_10785,N_9724,N_8621);
or U10786 (N_10786,N_6968,N_8798);
or U10787 (N_10787,N_6270,N_9160);
nand U10788 (N_10788,N_7775,N_7504);
xor U10789 (N_10789,N_8590,N_9357);
and U10790 (N_10790,N_7867,N_9207);
xor U10791 (N_10791,N_9270,N_9280);
and U10792 (N_10792,N_6266,N_8959);
and U10793 (N_10793,N_8308,N_8618);
or U10794 (N_10794,N_6350,N_5062);
or U10795 (N_10795,N_8276,N_9014);
and U10796 (N_10796,N_7204,N_7489);
nand U10797 (N_10797,N_7297,N_7259);
or U10798 (N_10798,N_5442,N_7889);
xnor U10799 (N_10799,N_6915,N_6829);
or U10800 (N_10800,N_9323,N_9862);
nor U10801 (N_10801,N_6763,N_5218);
xor U10802 (N_10802,N_7876,N_6738);
and U10803 (N_10803,N_8381,N_6045);
and U10804 (N_10804,N_6303,N_7690);
or U10805 (N_10805,N_8574,N_9017);
nor U10806 (N_10806,N_9365,N_5937);
and U10807 (N_10807,N_8215,N_8725);
nor U10808 (N_10808,N_5024,N_5192);
nand U10809 (N_10809,N_8598,N_6040);
xor U10810 (N_10810,N_8354,N_9897);
or U10811 (N_10811,N_5136,N_9231);
nor U10812 (N_10812,N_5274,N_6662);
or U10813 (N_10813,N_7306,N_9794);
nor U10814 (N_10814,N_5482,N_9473);
nand U10815 (N_10815,N_9388,N_7631);
xor U10816 (N_10816,N_9606,N_7422);
and U10817 (N_10817,N_5863,N_8825);
xor U10818 (N_10818,N_9541,N_6283);
xor U10819 (N_10819,N_8599,N_8751);
nor U10820 (N_10820,N_5099,N_6402);
nand U10821 (N_10821,N_7142,N_5508);
or U10822 (N_10822,N_7765,N_5818);
xnor U10823 (N_10823,N_9253,N_5632);
nand U10824 (N_10824,N_5257,N_5051);
and U10825 (N_10825,N_6138,N_5858);
nand U10826 (N_10826,N_5977,N_6699);
xor U10827 (N_10827,N_7069,N_6152);
and U10828 (N_10828,N_7099,N_6863);
xnor U10829 (N_10829,N_8197,N_7894);
and U10830 (N_10830,N_6463,N_7235);
nand U10831 (N_10831,N_7278,N_8760);
nand U10832 (N_10832,N_9698,N_7161);
nor U10833 (N_10833,N_8630,N_7692);
or U10834 (N_10834,N_8819,N_5862);
or U10835 (N_10835,N_5340,N_7429);
or U10836 (N_10836,N_6705,N_8714);
xor U10837 (N_10837,N_7768,N_6714);
nand U10838 (N_10838,N_7957,N_7912);
and U10839 (N_10839,N_5354,N_5019);
or U10840 (N_10840,N_8946,N_8105);
and U10841 (N_10841,N_5688,N_9678);
or U10842 (N_10842,N_7141,N_9814);
xor U10843 (N_10843,N_9108,N_5488);
or U10844 (N_10844,N_7577,N_6522);
or U10845 (N_10845,N_8003,N_9251);
xor U10846 (N_10846,N_8816,N_9824);
nor U10847 (N_10847,N_8320,N_9525);
and U10848 (N_10848,N_9796,N_8628);
xor U10849 (N_10849,N_5491,N_9081);
nor U10850 (N_10850,N_8958,N_7333);
or U10851 (N_10851,N_6715,N_9446);
nor U10852 (N_10852,N_5732,N_9377);
or U10853 (N_10853,N_8115,N_5049);
and U10854 (N_10854,N_6306,N_9764);
xor U10855 (N_10855,N_6130,N_9659);
or U10856 (N_10856,N_9568,N_6928);
and U10857 (N_10857,N_6264,N_7817);
nand U10858 (N_10858,N_8399,N_8603);
nor U10859 (N_10859,N_6413,N_5214);
xnor U10860 (N_10860,N_7909,N_8166);
and U10861 (N_10861,N_6872,N_8596);
nand U10862 (N_10862,N_9182,N_9561);
xor U10863 (N_10863,N_5532,N_6420);
or U10864 (N_10864,N_6812,N_9352);
xnor U10865 (N_10865,N_9265,N_6523);
nor U10866 (N_10866,N_8528,N_9305);
and U10867 (N_10867,N_5889,N_9874);
xor U10868 (N_10868,N_7583,N_8009);
xnor U10869 (N_10869,N_8090,N_6861);
nand U10870 (N_10870,N_6605,N_9652);
nand U10871 (N_10871,N_6005,N_7824);
and U10872 (N_10872,N_7724,N_9421);
xnor U10873 (N_10873,N_8327,N_6827);
nor U10874 (N_10874,N_6095,N_6967);
xor U10875 (N_10875,N_9687,N_5479);
or U10876 (N_10876,N_9539,N_8785);
and U10877 (N_10877,N_7599,N_9805);
nor U10878 (N_10878,N_8092,N_7108);
nor U10879 (N_10879,N_8782,N_8743);
and U10880 (N_10880,N_9894,N_9534);
nor U10881 (N_10881,N_8238,N_6560);
nor U10882 (N_10882,N_7771,N_6397);
or U10883 (N_10883,N_5789,N_5838);
or U10884 (N_10884,N_8444,N_6185);
xor U10885 (N_10885,N_8234,N_6317);
or U10886 (N_10886,N_7772,N_7754);
and U10887 (N_10887,N_6039,N_8107);
nand U10888 (N_10888,N_7045,N_7709);
xor U10889 (N_10889,N_9991,N_6088);
nor U10890 (N_10890,N_9554,N_9272);
and U10891 (N_10891,N_6471,N_6864);
nor U10892 (N_10892,N_6132,N_8995);
xor U10893 (N_10893,N_8820,N_6498);
and U10894 (N_10894,N_8060,N_7942);
or U10895 (N_10895,N_8130,N_9267);
nor U10896 (N_10896,N_7353,N_6947);
nand U10897 (N_10897,N_6329,N_6787);
or U10898 (N_10898,N_8269,N_9940);
xor U10899 (N_10899,N_9188,N_7896);
nand U10900 (N_10900,N_7795,N_9249);
nand U10901 (N_10901,N_8332,N_8738);
xnor U10902 (N_10902,N_9312,N_7450);
nand U10903 (N_10903,N_6878,N_9839);
and U10904 (N_10904,N_9509,N_8568);
and U10905 (N_10905,N_7650,N_9628);
and U10906 (N_10906,N_8588,N_5697);
and U10907 (N_10907,N_9332,N_5513);
or U10908 (N_10908,N_8957,N_7295);
nand U10909 (N_10909,N_6140,N_5869);
xnor U10910 (N_10910,N_6233,N_9479);
nor U10911 (N_10911,N_6453,N_9792);
xor U10912 (N_10912,N_5293,N_7686);
nor U10913 (N_10913,N_6736,N_8484);
nand U10914 (N_10914,N_7131,N_8188);
nand U10915 (N_10915,N_5263,N_8890);
and U10916 (N_10916,N_5339,N_7481);
or U10917 (N_10917,N_7950,N_5716);
xnor U10918 (N_10918,N_9268,N_7959);
and U10919 (N_10919,N_8944,N_8352);
nand U10920 (N_10920,N_7960,N_6957);
xor U10921 (N_10921,N_9809,N_7488);
xor U10922 (N_10922,N_5596,N_5489);
xnor U10923 (N_10923,N_7619,N_9042);
and U10924 (N_10924,N_6118,N_7726);
nand U10925 (N_10925,N_6876,N_6282);
or U10926 (N_10926,N_9391,N_7858);
or U10927 (N_10927,N_6468,N_7325);
nand U10928 (N_10928,N_7236,N_8413);
or U10929 (N_10929,N_6496,N_6180);
nor U10930 (N_10930,N_9517,N_9971);
or U10931 (N_10931,N_6456,N_7048);
or U10932 (N_10932,N_9949,N_6832);
xor U10933 (N_10933,N_9505,N_9976);
nand U10934 (N_10934,N_9121,N_7469);
nor U10935 (N_10935,N_7662,N_8290);
nand U10936 (N_10936,N_6400,N_6076);
nand U10937 (N_10937,N_6804,N_5676);
nor U10938 (N_10938,N_9130,N_9242);
or U10939 (N_10939,N_7113,N_6213);
nand U10940 (N_10940,N_9106,N_7218);
nand U10941 (N_10941,N_9165,N_9199);
xnor U10942 (N_10942,N_8889,N_5168);
nor U10943 (N_10943,N_5407,N_7971);
nand U10944 (N_10944,N_7818,N_6556);
xnor U10945 (N_10945,N_6984,N_8543);
nand U10946 (N_10946,N_9549,N_6856);
and U10947 (N_10947,N_8321,N_5562);
and U10948 (N_10948,N_8526,N_6708);
or U10949 (N_10949,N_7308,N_8569);
and U10950 (N_10950,N_5739,N_5909);
or U10951 (N_10951,N_9964,N_5807);
nand U10952 (N_10952,N_5572,N_8587);
and U10953 (N_10953,N_5686,N_5660);
xnor U10954 (N_10954,N_9399,N_6544);
xor U10955 (N_10955,N_8539,N_7231);
xnor U10956 (N_10956,N_8554,N_7367);
nand U10957 (N_10957,N_9363,N_8933);
xor U10958 (N_10958,N_8156,N_6851);
xnor U10959 (N_10959,N_9987,N_6895);
xnor U10960 (N_10960,N_8525,N_8369);
and U10961 (N_10961,N_8181,N_5299);
nand U10962 (N_10962,N_5744,N_6866);
and U10963 (N_10963,N_8607,N_9928);
xor U10964 (N_10964,N_5614,N_7786);
nor U10965 (N_10965,N_6887,N_7143);
and U10966 (N_10966,N_5200,N_8662);
and U10967 (N_10967,N_7166,N_8402);
and U10968 (N_10968,N_8418,N_6186);
xor U10969 (N_10969,N_7961,N_7698);
or U10970 (N_10970,N_7416,N_8713);
or U10971 (N_10971,N_5417,N_8719);
nor U10972 (N_10972,N_5782,N_8601);
nor U10973 (N_10973,N_8915,N_8516);
nor U10974 (N_10974,N_9240,N_6679);
or U10975 (N_10975,N_6904,N_9133);
and U10976 (N_10976,N_7103,N_6269);
and U10977 (N_10977,N_8684,N_7391);
and U10978 (N_10978,N_9438,N_5195);
or U10979 (N_10979,N_8748,N_9836);
or U10980 (N_10980,N_7418,N_5696);
xor U10981 (N_10981,N_7863,N_7877);
or U10982 (N_10982,N_6873,N_7360);
nor U10983 (N_10983,N_9778,N_5138);
nor U10984 (N_10984,N_7878,N_6682);
nand U10985 (N_10985,N_6659,N_7925);
or U10986 (N_10986,N_5504,N_8854);
nor U10987 (N_10987,N_6726,N_8312);
xnor U10988 (N_10988,N_5616,N_9282);
or U10989 (N_10989,N_6267,N_8432);
nor U10990 (N_10990,N_5231,N_5153);
xor U10991 (N_10991,N_8788,N_8458);
or U10992 (N_10992,N_7341,N_6330);
xor U10993 (N_10993,N_5243,N_7642);
nand U10994 (N_10994,N_7284,N_7598);
and U10995 (N_10995,N_6632,N_7968);
xor U10996 (N_10996,N_6107,N_7057);
and U10997 (N_10997,N_5667,N_8326);
nor U10998 (N_10998,N_7009,N_9086);
nand U10999 (N_10999,N_9795,N_5637);
nor U11000 (N_11000,N_5669,N_7120);
xnor U11001 (N_11001,N_7398,N_7548);
and U11002 (N_11002,N_8313,N_6074);
nor U11003 (N_11003,N_5347,N_5228);
nand U11004 (N_11004,N_5236,N_5416);
nor U11005 (N_11005,N_7280,N_6802);
or U11006 (N_11006,N_9649,N_6380);
nor U11007 (N_11007,N_5811,N_5629);
nor U11008 (N_11008,N_9566,N_9918);
or U11009 (N_11009,N_8975,N_5011);
or U11010 (N_11010,N_5111,N_8930);
or U11011 (N_11011,N_7022,N_8300);
or U11012 (N_11012,N_6650,N_6404);
nand U11013 (N_11013,N_5240,N_7784);
nor U11014 (N_11014,N_8247,N_8918);
and U11015 (N_11015,N_9961,N_5692);
xor U11016 (N_11016,N_6899,N_9390);
or U11017 (N_11017,N_9204,N_8758);
or U11018 (N_11018,N_5552,N_9757);
nand U11019 (N_11019,N_6392,N_5949);
nor U11020 (N_11020,N_8430,N_6476);
xor U11021 (N_11021,N_9780,N_8330);
or U11022 (N_11022,N_7248,N_8031);
or U11023 (N_11023,N_5276,N_9557);
nor U11024 (N_11024,N_9739,N_5608);
nand U11025 (N_11025,N_7843,N_6210);
xnor U11026 (N_11026,N_6996,N_9868);
nand U11027 (N_11027,N_7670,N_7102);
and U11028 (N_11028,N_9514,N_7211);
xor U11029 (N_11029,N_9067,N_9264);
xnor U11030 (N_11030,N_6328,N_8459);
or U11031 (N_11031,N_9217,N_8850);
and U11032 (N_11032,N_9002,N_6027);
nor U11033 (N_11033,N_7408,N_9817);
nand U11034 (N_11034,N_6575,N_8378);
or U11035 (N_11035,N_8586,N_6880);
xnor U11036 (N_11036,N_9892,N_9821);
xnor U11037 (N_11037,N_6051,N_9573);
and U11038 (N_11038,N_8899,N_6698);
xnor U11039 (N_11039,N_8789,N_8649);
nor U11040 (N_11040,N_8822,N_8393);
nand U11041 (N_11041,N_5273,N_5329);
or U11042 (N_11042,N_7732,N_7448);
or U11043 (N_11043,N_9018,N_5092);
nand U11044 (N_11044,N_7926,N_7127);
nand U11045 (N_11045,N_7427,N_7381);
and U11046 (N_11046,N_5321,N_9670);
and U11047 (N_11047,N_6053,N_7620);
nor U11048 (N_11048,N_6512,N_8658);
xnor U11049 (N_11049,N_8870,N_7602);
and U11050 (N_11050,N_6414,N_9370);
nor U11051 (N_11051,N_7715,N_9236);
or U11052 (N_11052,N_8795,N_7913);
nor U11053 (N_11053,N_7132,N_7264);
nor U11054 (N_11054,N_6761,N_6103);
nand U11055 (N_11055,N_5699,N_6336);
or U11056 (N_11056,N_7040,N_7545);
and U11057 (N_11057,N_8581,N_9151);
nand U11058 (N_11058,N_7487,N_8141);
nand U11059 (N_11059,N_5216,N_5251);
xnor U11060 (N_11060,N_8593,N_5853);
and U11061 (N_11061,N_7613,N_8774);
nand U11062 (N_11062,N_9379,N_6974);
nor U11063 (N_11063,N_6126,N_6932);
and U11064 (N_11064,N_9038,N_8202);
nor U11065 (N_11065,N_7310,N_6752);
xor U11066 (N_11066,N_8291,N_7101);
nor U11067 (N_11067,N_9071,N_7413);
nand U11068 (N_11068,N_9205,N_9756);
xor U11069 (N_11069,N_7205,N_7582);
nand U11070 (N_11070,N_8796,N_6971);
xnor U11071 (N_11071,N_6253,N_8375);
nand U11072 (N_11072,N_6445,N_5094);
nand U11073 (N_11073,N_7687,N_7695);
and U11074 (N_11074,N_5301,N_8720);
xnor U11075 (N_11075,N_7904,N_5673);
and U11076 (N_11076,N_5615,N_9774);
and U11077 (N_11077,N_8495,N_5760);
nor U11078 (N_11078,N_8824,N_7286);
nand U11079 (N_11079,N_8670,N_8856);
xnor U11080 (N_11080,N_5501,N_8157);
xnor U11081 (N_11081,N_7116,N_5569);
and U11082 (N_11082,N_8044,N_7148);
nor U11083 (N_11083,N_9163,N_5622);
nor U11084 (N_11084,N_7454,N_9056);
or U11085 (N_11085,N_7316,N_8138);
or U11086 (N_11086,N_7573,N_5683);
xor U11087 (N_11087,N_6642,N_7743);
xnor U11088 (N_11088,N_6434,N_9716);
nand U11089 (N_11089,N_8088,N_9284);
nand U11090 (N_11090,N_5269,N_8843);
nand U11091 (N_11091,N_5193,N_7584);
or U11092 (N_11092,N_5330,N_6060);
nand U11093 (N_11093,N_8400,N_6535);
or U11094 (N_11094,N_7140,N_6221);
xnor U11095 (N_11095,N_8048,N_6240);
nand U11096 (N_11096,N_9960,N_6910);
xnor U11097 (N_11097,N_5319,N_5467);
and U11098 (N_11098,N_8294,N_8081);
nor U11099 (N_11099,N_9104,N_5469);
and U11100 (N_11100,N_7799,N_6218);
nand U11101 (N_11101,N_7561,N_8070);
nor U11102 (N_11102,N_5400,N_7995);
nand U11103 (N_11103,N_7018,N_8698);
nand U11104 (N_11104,N_7547,N_9587);
nand U11105 (N_11105,N_9989,N_6855);
xnor U11106 (N_11106,N_8385,N_8160);
nor U11107 (N_11107,N_5647,N_6890);
and U11108 (N_11108,N_8415,N_9748);
and U11109 (N_11109,N_9497,N_7485);
or U11110 (N_11110,N_5159,N_7663);
or U11111 (N_11111,N_8099,N_6477);
xor U11112 (N_11112,N_7446,N_6913);
or U11113 (N_11113,N_8792,N_9094);
xor U11114 (N_11114,N_5435,N_8293);
or U11115 (N_11115,N_7906,N_8722);
and U11116 (N_11116,N_6092,N_8331);
xor U11117 (N_11117,N_6551,N_6162);
and U11118 (N_11118,N_5851,N_7281);
nand U11119 (N_11119,N_9582,N_7606);
or U11120 (N_11120,N_9496,N_5812);
xor U11121 (N_11121,N_7791,N_9477);
nand U11122 (N_11122,N_6492,N_7644);
and U11123 (N_11123,N_5639,N_6232);
and U11124 (N_11124,N_8584,N_8256);
xor U11125 (N_11125,N_6251,N_5915);
nand U11126 (N_11126,N_5054,N_5887);
nand U11127 (N_11127,N_8390,N_8851);
nand U11128 (N_11128,N_8405,N_5640);
nor U11129 (N_11129,N_6395,N_9978);
or U11130 (N_11130,N_5267,N_6892);
nor U11131 (N_11131,N_7017,N_8191);
nand U11132 (N_11132,N_6237,N_9075);
or U11133 (N_11133,N_7993,N_7184);
and U11134 (N_11134,N_5447,N_9740);
nand U11135 (N_11135,N_6192,N_9972);
nand U11136 (N_11136,N_6147,N_9546);
nand U11137 (N_11137,N_5882,N_8497);
nand U11138 (N_11138,N_7708,N_7526);
and U11139 (N_11139,N_5704,N_8807);
nand U11140 (N_11140,N_5248,N_7607);
nor U11141 (N_11141,N_5219,N_6339);
and U11142 (N_11142,N_9333,N_9355);
xor U11143 (N_11143,N_6230,N_6344);
and U11144 (N_11144,N_5678,N_8863);
nand U11145 (N_11145,N_5868,N_7344);
or U11146 (N_11146,N_8787,N_6663);
xor U11147 (N_11147,N_8682,N_9498);
nor U11148 (N_11148,N_5132,N_8264);
nor U11149 (N_11149,N_9958,N_6121);
xor U11150 (N_11150,N_5266,N_9178);
and U11151 (N_11151,N_5201,N_6860);
and U11152 (N_11152,N_5962,N_9200);
xnor U11153 (N_11153,N_8203,N_6760);
nor U11154 (N_11154,N_5264,N_6640);
nand U11155 (N_11155,N_8500,N_6222);
and U11156 (N_11156,N_9400,N_7660);
xnor U11157 (N_11157,N_5493,N_9319);
nand U11158 (N_11158,N_6795,N_9750);
or U11159 (N_11159,N_8318,N_7737);
nand U11160 (N_11160,N_5071,N_7479);
xor U11161 (N_11161,N_5849,N_9076);
xnor U11162 (N_11162,N_8270,N_7893);
and U11163 (N_11163,N_9469,N_9771);
nor U11164 (N_11164,N_5331,N_9122);
or U11165 (N_11165,N_9336,N_8167);
xnor U11166 (N_11166,N_8248,N_7990);
nor U11167 (N_11167,N_6870,N_7621);
nor U11168 (N_11168,N_9313,N_9445);
nor U11169 (N_11169,N_9344,N_5280);
and U11170 (N_11170,N_5545,N_7900);
xnor U11171 (N_11171,N_9706,N_8366);
nand U11172 (N_11172,N_8737,N_7480);
nor U11173 (N_11173,N_9383,N_5176);
xor U11174 (N_11174,N_9544,N_6604);
or U11175 (N_11175,N_9096,N_8280);
or U11176 (N_11176,N_7347,N_6722);
or U11177 (N_11177,N_8022,N_7486);
or U11178 (N_11178,N_7016,N_6319);
xnor U11179 (N_11179,N_7031,N_6702);
or U11180 (N_11180,N_8867,N_5933);
xnor U11181 (N_11181,N_6966,N_7540);
nor U11182 (N_11182,N_6893,N_9705);
nand U11183 (N_11183,N_7024,N_9664);
and U11184 (N_11184,N_9193,N_7844);
nand U11185 (N_11185,N_5131,N_6891);
nand U11186 (N_11186,N_8766,N_8754);
nor U11187 (N_11187,N_7939,N_7842);
or U11188 (N_11188,N_8802,N_6291);
and U11189 (N_11189,N_9929,N_9979);
or U11190 (N_11190,N_5666,N_8311);
and U11191 (N_11191,N_9812,N_5881);
nand U11192 (N_11192,N_7474,N_9819);
nand U11193 (N_11193,N_6217,N_8794);
and U11194 (N_11194,N_5873,N_9632);
xnor U11195 (N_11195,N_5290,N_9095);
xor U11196 (N_11196,N_8642,N_9084);
nor U11197 (N_11197,N_6577,N_6263);
nand U11198 (N_11198,N_7441,N_8974);
or U11199 (N_11199,N_6626,N_7596);
xor U11200 (N_11200,N_8753,N_6202);
xor U11201 (N_11201,N_7146,N_9594);
and U11202 (N_11202,N_6358,N_9330);
or U11203 (N_11203,N_6624,N_5210);
and U11204 (N_11204,N_6125,N_7089);
or U11205 (N_11205,N_8396,N_7800);
or U11206 (N_11206,N_6791,N_5065);
and U11207 (N_11207,N_9502,N_6511);
xnor U11208 (N_11208,N_6293,N_5531);
xor U11209 (N_11209,N_7261,N_7559);
or U11210 (N_11210,N_5362,N_7085);
xnor U11211 (N_11211,N_8759,N_5734);
xnor U11212 (N_11212,N_8278,N_9613);
or U11213 (N_11213,N_8620,N_8988);
and U11214 (N_11214,N_6116,N_5773);
or U11215 (N_11215,N_7520,N_7717);
xor U11216 (N_11216,N_5475,N_6458);
and U11217 (N_11217,N_7228,N_7507);
xnor U11218 (N_11218,N_8982,N_5426);
nor U11219 (N_11219,N_6254,N_8893);
nand U11220 (N_11220,N_5371,N_5351);
nand U11221 (N_11221,N_9077,N_8360);
or U11222 (N_11222,N_9769,N_5548);
and U11223 (N_11223,N_8523,N_9309);
or U11224 (N_11224,N_7414,N_8967);
and U11225 (N_11225,N_5896,N_7207);
nor U11226 (N_11226,N_7675,N_9692);
nor U11227 (N_11227,N_8226,N_8793);
nand U11228 (N_11228,N_9187,N_7550);
and U11229 (N_11229,N_9480,N_7199);
xnor U11230 (N_11230,N_5031,N_5521);
nand U11231 (N_11231,N_6638,N_7648);
xor U11232 (N_11232,N_9119,N_5668);
xnor U11233 (N_11233,N_5861,N_9382);
or U11234 (N_11234,N_6536,N_6822);
or U11235 (N_11235,N_5650,N_8489);
nor U11236 (N_11236,N_5385,N_5820);
nor U11237 (N_11237,N_7232,N_7114);
or U11238 (N_11238,N_5736,N_5701);
and U11239 (N_11239,N_5980,N_5520);
or U11240 (N_11240,N_5564,N_9977);
nor U11241 (N_11241,N_5037,N_5726);
xor U11242 (N_11242,N_6588,N_9690);
nor U11243 (N_11243,N_7303,N_8999);
or U11244 (N_11244,N_6609,N_7555);
xnor U11245 (N_11245,N_8937,N_8827);
and U11246 (N_11246,N_6871,N_6885);
nor U11247 (N_11247,N_9784,N_8414);
xor U11248 (N_11248,N_5530,N_9252);
nor U11249 (N_11249,N_6128,N_9430);
or U11250 (N_11250,N_9286,N_8110);
and U11251 (N_11251,N_7426,N_9055);
nor U11252 (N_11252,N_7736,N_6700);
nand U11253 (N_11253,N_8828,N_8844);
nor U11254 (N_11254,N_8094,N_6625);
and U11255 (N_11255,N_7710,N_7346);
xor U11256 (N_11256,N_5117,N_8314);
xnor U11257 (N_11257,N_8786,N_7399);
xor U11258 (N_11258,N_9766,N_6467);
nand U11259 (N_11259,N_9214,N_6242);
nand U11260 (N_11260,N_9255,N_8895);
and U11261 (N_11261,N_9591,N_5916);
nor U11262 (N_11262,N_7257,N_8251);
and U11263 (N_11263,N_7430,N_6298);
nand U11264 (N_11264,N_5558,N_9695);
nand U11265 (N_11265,N_8387,N_6506);
and U11266 (N_11266,N_5538,N_6500);
xnor U11267 (N_11267,N_6035,N_5067);
nor U11268 (N_11268,N_5815,N_6750);
nand U11269 (N_11269,N_5378,N_7779);
nand U11270 (N_11270,N_5328,N_6911);
nor U11271 (N_11271,N_7477,N_6022);
xor U11272 (N_11272,N_5741,N_9468);
nand U11273 (N_11273,N_8756,N_5196);
or U11274 (N_11274,N_9943,N_6776);
xnor U11275 (N_11275,N_9287,N_5473);
xnor U11276 (N_11276,N_9694,N_5800);
or U11277 (N_11277,N_9493,N_5810);
nand U11278 (N_11278,N_5775,N_5383);
nand U11279 (N_11279,N_5363,N_5631);
xor U11280 (N_11280,N_6546,N_6874);
and U11281 (N_11281,N_9082,N_5403);
nand U11282 (N_11282,N_6394,N_8733);
and U11283 (N_11283,N_8032,N_6896);
xnor U11284 (N_11284,N_9278,N_5307);
nor U11285 (N_11285,N_5088,N_5884);
or U11286 (N_11286,N_7067,N_5826);
nand U11287 (N_11287,N_5941,N_5852);
nand U11288 (N_11288,N_8267,N_9037);
or U11289 (N_11289,N_5626,N_8803);
nand U11290 (N_11290,N_6907,N_5055);
nor U11291 (N_11291,N_8677,N_7654);
and U11292 (N_11292,N_6643,N_7563);
nand U11293 (N_11293,N_5327,N_5719);
and U11294 (N_11294,N_9232,N_6031);
nand U11295 (N_11295,N_8053,N_5963);
xnor U11296 (N_11296,N_9902,N_6660);
and U11297 (N_11297,N_7597,N_9562);
or U11298 (N_11298,N_9707,N_9852);
nor U11299 (N_11299,N_5693,N_8544);
xor U11300 (N_11300,N_7989,N_8972);
and U11301 (N_11301,N_8152,N_7757);
xor U11302 (N_11302,N_5865,N_9853);
nand U11303 (N_11303,N_7657,N_6304);
and U11304 (N_11304,N_7339,N_7529);
and U11305 (N_11305,N_6120,N_5566);
or U11306 (N_11306,N_5586,N_9937);
or U11307 (N_11307,N_9410,N_7883);
xnor U11308 (N_11308,N_8475,N_8347);
and U11309 (N_11309,N_6205,N_5589);
or U11310 (N_11310,N_8705,N_5745);
nand U11311 (N_11311,N_9996,N_9490);
nor U11312 (N_11312,N_8448,N_7197);
nand U11313 (N_11313,N_8671,N_7921);
nand U11314 (N_11314,N_8742,N_7377);
and U11315 (N_11315,N_9720,N_5438);
and U11316 (N_11316,N_7729,N_9208);
and U11317 (N_11317,N_9212,N_8858);
or U11318 (N_11318,N_6796,N_6156);
nor U11319 (N_11319,N_5252,N_5053);
and U11320 (N_11320,N_9605,N_9957);
xnor U11321 (N_11321,N_8878,N_5605);
and U11322 (N_11322,N_7917,N_5422);
and U11323 (N_11323,N_8894,N_7002);
and U11324 (N_11324,N_6346,N_6015);
and U11325 (N_11325,N_9191,N_8460);
nand U11326 (N_11326,N_7196,N_9135);
or U11327 (N_11327,N_7225,N_7121);
xnor U11328 (N_11328,N_8977,N_8991);
xor U11329 (N_11329,N_6079,N_5249);
nand U11330 (N_11330,N_6525,N_8906);
and U11331 (N_11331,N_5070,N_6371);
nor U11332 (N_11332,N_9465,N_5655);
and U11333 (N_11333,N_8001,N_7880);
or U11334 (N_11334,N_6983,N_8255);
and U11335 (N_11335,N_9427,N_6690);
xor U11336 (N_11336,N_5854,N_6352);
or U11337 (N_11337,N_7138,N_9258);
xnor U11338 (N_11338,N_7010,N_5784);
xnor U11339 (N_11339,N_5777,N_5983);
nor U11340 (N_11340,N_6023,N_7307);
nand U11341 (N_11341,N_6178,N_5689);
nor U11342 (N_11342,N_6113,N_5722);
and U11343 (N_11343,N_6547,N_8848);
nor U11344 (N_11344,N_8146,N_8409);
nor U11345 (N_11345,N_6422,N_6172);
xor U11346 (N_11346,N_7672,N_9269);
nand U11347 (N_11347,N_8093,N_6080);
or U11348 (N_11348,N_6965,N_5891);
xnor U11349 (N_11349,N_9755,N_8359);
or U11350 (N_11350,N_6068,N_5613);
or U11351 (N_11351,N_9527,N_5253);
and U11352 (N_11352,N_5325,N_5141);
nand U11353 (N_11353,N_9492,N_9097);
or U11354 (N_11354,N_6692,N_5389);
xor U11355 (N_11355,N_9601,N_8914);
nor U11356 (N_11356,N_7029,N_9540);
and U11357 (N_11357,N_5386,N_5942);
nand U11358 (N_11358,N_5203,N_9581);
or U11359 (N_11359,N_5908,N_7423);
or U11360 (N_11360,N_8114,N_8548);
xnor U11361 (N_11361,N_5787,N_8538);
and U11362 (N_11362,N_9334,N_8869);
xor U11363 (N_11363,N_7090,N_6144);
xnor U11364 (N_11364,N_6903,N_5060);
nor U11365 (N_11365,N_5993,N_5431);
nor U11366 (N_11366,N_7056,N_7635);
xor U11367 (N_11367,N_8739,N_6259);
or U11368 (N_11368,N_8467,N_9633);
or U11369 (N_11369,N_7949,N_7417);
or U11370 (N_11370,N_8361,N_9671);
and U11371 (N_11371,N_5198,N_7862);
nand U11372 (N_11372,N_5947,N_6459);
or U11373 (N_11373,N_6073,N_6465);
or U11374 (N_11374,N_8450,N_5100);
and U11375 (N_11375,N_7080,N_7252);
nand U11376 (N_11376,N_6421,N_8427);
nor U11377 (N_11377,N_7970,N_7324);
or U11378 (N_11378,N_9091,N_9068);
xnor U11379 (N_11379,N_7503,N_7696);
nand U11380 (N_11380,N_7215,N_6307);
nand U11381 (N_11381,N_7903,N_8324);
xor U11382 (N_11382,N_6235,N_8633);
nand U11383 (N_11383,N_6009,N_7735);
or U11384 (N_11384,N_8814,N_5926);
and U11385 (N_11385,N_6191,N_5705);
or U11386 (N_11386,N_9257,N_5140);
and U11387 (N_11387,N_6382,N_7206);
or U11388 (N_11388,N_5578,N_8086);
and U11389 (N_11389,N_5727,N_8647);
and U11390 (N_11390,N_9259,N_7859);
nor U11391 (N_11391,N_6206,N_8243);
or U11392 (N_11392,N_7001,N_7908);
nor U11393 (N_11393,N_6433,N_6944);
or U11394 (N_11394,N_5095,N_8095);
nand U11395 (N_11395,N_9124,N_7165);
xor U11396 (N_11396,N_7716,N_7734);
nor U11397 (N_11397,N_5262,N_5134);
or U11398 (N_11398,N_9092,N_6321);
and U11399 (N_11399,N_6853,N_8172);
or U11400 (N_11400,N_5082,N_5080);
xnor U11401 (N_11401,N_8486,N_7998);
nor U11402 (N_11402,N_8153,N_6674);
xnor U11403 (N_11403,N_7188,N_6756);
nand U11404 (N_11404,N_6884,N_5027);
nand U11405 (N_11405,N_9845,N_6044);
or U11406 (N_11406,N_5244,N_9856);
nor U11407 (N_11407,N_8464,N_9233);
and U11408 (N_11408,N_8580,N_8217);
or U11409 (N_11409,N_5625,N_9293);
nand U11410 (N_11410,N_8189,N_9722);
or U11411 (N_11411,N_8846,N_7653);
nor U11412 (N_11412,N_6554,N_8456);
or U11413 (N_11413,N_6334,N_5220);
xor U11414 (N_11414,N_8049,N_5954);
or U11415 (N_11415,N_7220,N_6681);
nor U11416 (N_11416,N_7665,N_8675);
xnor U11417 (N_11417,N_5030,N_8638);
nand U11418 (N_11418,N_5832,N_9132);
xnor U11419 (N_11419,N_7656,N_5156);
and U11420 (N_11420,N_8443,N_8665);
or U11421 (N_11421,N_5651,N_6423);
or U11422 (N_11422,N_9799,N_7825);
and U11423 (N_11423,N_9662,N_6308);
or U11424 (N_11424,N_7168,N_6032);
nor U11425 (N_11425,N_7558,N_8288);
or U11426 (N_11426,N_6668,N_7093);
or U11427 (N_11427,N_6824,N_5690);
nor U11428 (N_11428,N_5776,N_9022);
nand U11429 (N_11429,N_6012,N_7988);
or U11430 (N_11430,N_6014,N_5551);
nor U11431 (N_11431,N_7668,N_8908);
xor U11432 (N_11432,N_9615,N_8061);
nor U11433 (N_11433,N_6129,N_7987);
xor U11434 (N_11434,N_8897,N_7350);
or U11435 (N_11435,N_7054,N_8126);
and U11436 (N_11436,N_7527,N_7255);
or U11437 (N_11437,N_7337,N_9663);
or U11438 (N_11438,N_6842,N_7008);
or U11439 (N_11439,N_6540,N_6848);
nand U11440 (N_11440,N_9936,N_5519);
nor U11441 (N_11441,N_9110,N_7229);
or U11442 (N_11442,N_9088,N_8454);
nand U11443 (N_11443,N_7362,N_9790);
nor U11444 (N_11444,N_9011,N_8555);
nor U11445 (N_11445,N_6954,N_7640);
xor U11446 (N_11446,N_7241,N_7079);
or U11447 (N_11447,N_9127,N_7821);
xnor U11448 (N_11448,N_7553,N_7705);
or U11449 (N_11449,N_5015,N_5876);
and U11450 (N_11450,N_7499,N_8752);
xnor U11451 (N_11451,N_5116,N_5155);
xnor U11452 (N_11452,N_7645,N_5186);
nor U11453 (N_11453,N_7088,N_5781);
nand U11454 (N_11454,N_9041,N_5476);
or U11455 (N_11455,N_5109,N_7616);
xor U11456 (N_11456,N_6924,N_9350);
nand U11457 (N_11457,N_7275,N_6085);
and U11458 (N_11458,N_7887,N_6671);
and U11459 (N_11459,N_6142,N_5028);
nor U11460 (N_11460,N_7565,N_6591);
xnor U11461 (N_11461,N_9032,N_7059);
xor U11462 (N_11462,N_7263,N_8404);
and U11463 (N_11463,N_7245,N_5579);
nor U11464 (N_11464,N_9107,N_9924);
xor U11465 (N_11465,N_6712,N_5721);
and U11466 (N_11466,N_6922,N_5645);
nand U11467 (N_11467,N_8861,N_6262);
nand U11468 (N_11468,N_6425,N_9726);
xnor U11469 (N_11469,N_5965,N_9083);
xor U11470 (N_11470,N_8556,N_5372);
nor U11471 (N_11471,N_7936,N_5763);
or U11472 (N_11472,N_6565,N_8968);
nor U11473 (N_11473,N_9816,N_5809);
and U11474 (N_11474,N_7927,N_9945);
nand U11475 (N_11475,N_6356,N_9732);
or U11476 (N_11476,N_9619,N_8687);
nor U11477 (N_11477,N_6645,N_5437);
xor U11478 (N_11478,N_5656,N_5296);
or U11479 (N_11479,N_9730,N_9029);
nor U11480 (N_11480,N_9045,N_6781);
or U11481 (N_11481,N_8144,N_6309);
xor U11482 (N_11482,N_9475,N_5149);
and U11483 (N_11483,N_5927,N_5706);
nand U11484 (N_11484,N_5988,N_7219);
xnor U11485 (N_11485,N_8123,N_8545);
and U11486 (N_11486,N_9362,N_5408);
xnor U11487 (N_11487,N_6224,N_6583);
and U11488 (N_11488,N_6484,N_6542);
xor U11489 (N_11489,N_5537,N_5384);
xor U11490 (N_11490,N_8834,N_6386);
nand U11491 (N_11491,N_8996,N_7747);
nor U11492 (N_11492,N_5525,N_7282);
and U11493 (N_11493,N_8770,N_5048);
or U11494 (N_11494,N_8228,N_5016);
nand U11495 (N_11495,N_8515,N_7274);
nand U11496 (N_11496,N_6689,N_7365);
nand U11497 (N_11497,N_7923,N_6294);
nand U11498 (N_11498,N_7203,N_8976);
xnor U11499 (N_11499,N_5130,N_9642);
or U11500 (N_11500,N_5539,N_5255);
xor U11501 (N_11501,N_7829,N_8462);
nand U11502 (N_11502,N_8388,N_7759);
nand U11503 (N_11503,N_6231,N_6026);
or U11504 (N_11504,N_7380,N_7605);
xor U11505 (N_11505,N_7803,N_7156);
nor U11506 (N_11506,N_6828,N_6341);
nand U11507 (N_11507,N_6360,N_9783);
nor U11508 (N_11508,N_5033,N_9256);
and U11509 (N_11509,N_8492,N_7511);
nor U11510 (N_11510,N_6937,N_9491);
nand U11511 (N_11511,N_8014,N_9746);
and U11512 (N_11512,N_6099,N_8892);
nor U11513 (N_11513,N_9488,N_5366);
nand U11514 (N_11514,N_8292,N_7302);
or U11515 (N_11515,N_6811,N_5332);
nand U11516 (N_11516,N_8579,N_8077);
and U11517 (N_11517,N_6883,N_9345);
nand U11518 (N_11518,N_5064,N_8939);
or U11519 (N_11519,N_9316,N_7359);
xor U11520 (N_11520,N_6102,N_9442);
and U11521 (N_11521,N_9574,N_6385);
or U11522 (N_11522,N_7453,N_9320);
nand U11523 (N_11523,N_6633,N_8686);
nor U11524 (N_11524,N_5885,N_9098);
xor U11525 (N_11525,N_5205,N_6353);
or U11526 (N_11526,N_5630,N_5320);
nand U11527 (N_11527,N_9956,N_9721);
or U11528 (N_11528,N_5758,N_6406);
or U11529 (N_11529,N_8072,N_7651);
and U11530 (N_11530,N_7317,N_6479);
xor U11531 (N_11531,N_7371,N_8532);
and U11532 (N_11532,N_7808,N_5560);
nand U11533 (N_11533,N_6478,N_6215);
xor U11534 (N_11534,N_9190,N_5549);
xor U11535 (N_11535,N_5040,N_7819);
xnor U11536 (N_11536,N_9230,N_9291);
or U11537 (N_11537,N_9369,N_5867);
or U11538 (N_11538,N_6127,N_5617);
nor U11539 (N_11539,N_7612,N_9224);
and U11540 (N_11540,N_8478,N_6390);
or U11541 (N_11541,N_6275,N_9917);
nand U11542 (N_11542,N_8042,N_7847);
or U11543 (N_11543,N_7618,N_9229);
nor U11544 (N_11544,N_6069,N_7068);
nand U11545 (N_11545,N_9448,N_8043);
and U11546 (N_11546,N_8470,N_7340);
and U11547 (N_11547,N_6644,N_5344);
or U11548 (N_11548,N_9250,N_9758);
xnor U11549 (N_11549,N_6279,N_9735);
nor U11550 (N_11550,N_5757,N_5604);
xor U11551 (N_11551,N_6817,N_7425);
and U11552 (N_11552,N_5317,N_8821);
or U11553 (N_11553,N_6495,N_6524);
nand U11554 (N_11554,N_7134,N_9680);
nor U11555 (N_11555,N_6991,N_7435);
or U11556 (N_11556,N_8627,N_8911);
nand U11557 (N_11557,N_5592,N_6227);
xnor U11558 (N_11558,N_5510,N_9298);
nor U11559 (N_11559,N_5406,N_9453);
and U11560 (N_11560,N_6667,N_6993);
nor U11561 (N_11561,N_8956,N_5516);
xnor U11562 (N_11562,N_8403,N_7014);
or U11563 (N_11563,N_8493,N_6945);
and U11564 (N_11564,N_7318,N_9723);
or U11565 (N_11565,N_5245,N_8271);
or U11566 (N_11566,N_8718,N_9149);
or U11567 (N_11567,N_8265,N_9358);
nand U11568 (N_11568,N_5418,N_8260);
xnor U11569 (N_11569,N_9185,N_7985);
nor U11570 (N_11570,N_8594,N_9281);
xor U11571 (N_11571,N_7790,N_8572);
xor U11572 (N_11572,N_6836,N_9441);
nor U11573 (N_11573,N_9665,N_9359);
or U11574 (N_11574,N_7977,N_5958);
xor U11575 (N_11575,N_6723,N_9302);
nand U11576 (N_11576,N_6173,N_7731);
nand U11577 (N_11577,N_8310,N_6226);
xnor U11578 (N_11578,N_9158,N_6249);
or U11579 (N_11579,N_6975,N_5507);
nand U11580 (N_11580,N_7155,N_7276);
nand U11581 (N_11581,N_7767,N_7190);
nand U11582 (N_11582,N_8485,N_5679);
nor U11583 (N_11583,N_6480,N_5461);
xor U11584 (N_11584,N_9274,N_6772);
nand U11585 (N_11585,N_8177,N_5129);
and U11586 (N_11586,N_7119,N_8511);
or U11587 (N_11587,N_8150,N_6569);
nor U11588 (N_11588,N_8401,N_7749);
and U11589 (N_11589,N_8118,N_9864);
and U11590 (N_11590,N_8370,N_9703);
xor U11591 (N_11591,N_5107,N_7182);
nand U11592 (N_11592,N_9371,N_6599);
nand U11593 (N_11593,N_5423,N_6273);
and U11594 (N_11594,N_8781,N_5352);
nand U11595 (N_11595,N_7449,N_8073);
and U11596 (N_11596,N_6809,N_6248);
and U11597 (N_11597,N_7406,N_9481);
nor U11598 (N_11598,N_8155,N_8877);
xnor U11599 (N_11599,N_9691,N_5806);
nand U11600 (N_11600,N_9922,N_8244);
or U11601 (N_11601,N_7851,N_7840);
nor U11602 (N_11602,N_7171,N_5643);
nor U11603 (N_11603,N_5633,N_5583);
xor U11604 (N_11604,N_9841,N_5069);
nor U11605 (N_11605,N_7312,N_8597);
nand U11606 (N_11606,N_7756,N_6835);
and U11607 (N_11607,N_8205,N_7788);
xor U11608 (N_11608,N_5928,N_7932);
nor U11609 (N_11609,N_8522,N_9109);
nor U11610 (N_11610,N_9881,N_6611);
xnor U11611 (N_11611,N_8283,N_9456);
nand U11612 (N_11612,N_5050,N_9708);
nor U11613 (N_11613,N_5575,N_5986);
nor U11614 (N_11614,N_5377,N_5445);
nor U11615 (N_11615,N_5972,N_6446);
and U11616 (N_11616,N_9893,N_9063);
xnor U11617 (N_11617,N_5410,N_9013);
and U11618 (N_11618,N_8213,N_8902);
xnor U11619 (N_11619,N_6369,N_9314);
or U11620 (N_11620,N_5730,N_6630);
nand U11621 (N_11621,N_7468,N_8876);
xnor U11622 (N_11622,N_9078,N_6710);
xnor U11623 (N_11623,N_8424,N_5890);
nor U11624 (N_11624,N_7208,N_5358);
or U11625 (N_11625,N_7832,N_9607);
and U11626 (N_11626,N_6909,N_7217);
and U11627 (N_11627,N_5480,N_7699);
or U11628 (N_11628,N_9914,N_7608);
nor U11629 (N_11629,N_8438,N_5144);
and U11630 (N_11630,N_6788,N_9890);
nand U11631 (N_11631,N_5911,N_9113);
or U11632 (N_11632,N_6228,N_6295);
nand U11633 (N_11633,N_7387,N_8383);
or U11634 (N_11634,N_7160,N_6740);
nor U11635 (N_11635,N_6517,N_8062);
and U11636 (N_11636,N_5075,N_9254);
xor U11637 (N_11637,N_8358,N_5208);
or U11638 (N_11638,N_6119,N_8883);
nand U11639 (N_11639,N_5829,N_8917);
xor U11640 (N_11640,N_9227,N_5845);
and U11641 (N_11641,N_8059,N_5929);
or U11642 (N_11642,N_6105,N_9239);
and U11643 (N_11643,N_9192,N_5120);
xnor U11644 (N_11644,N_5563,N_7581);
and U11645 (N_11645,N_7436,N_5582);
nand U11646 (N_11646,N_6711,N_5670);
xor U11647 (N_11647,N_9327,N_8111);
or U11648 (N_11648,N_5764,N_5194);
xnor U11649 (N_11649,N_7456,N_5034);
nor U11650 (N_11650,N_6084,N_5465);
or U11651 (N_11651,N_8469,N_8732);
nand U11652 (N_11652,N_8928,N_9471);
nor U11653 (N_11653,N_7326,N_8125);
xnor U11654 (N_11654,N_7864,N_8199);
nor U11655 (N_11655,N_7947,N_8371);
and U11656 (N_11656,N_6419,N_8693);
nand U11657 (N_11657,N_8079,N_9331);
nand U11658 (N_11658,N_9701,N_9753);
nand U11659 (N_11659,N_5237,N_7452);
nor U11660 (N_11660,N_9963,N_9888);
nor U11661 (N_11661,N_8345,N_6297);
and U11662 (N_11662,N_8836,N_9062);
or U11663 (N_11663,N_7253,N_5122);
nand U11664 (N_11664,N_7730,N_7105);
nor U11665 (N_11665,N_9437,N_8660);
nor U11666 (N_11666,N_5286,N_6897);
xor U11667 (N_11667,N_6614,N_9910);
xnor U11668 (N_11668,N_6969,N_7351);
xor U11669 (N_11669,N_7535,N_6509);
nand U11670 (N_11670,N_5875,N_8659);
nor U11671 (N_11671,N_5523,N_6117);
and U11672 (N_11672,N_9226,N_5920);
nor U11673 (N_11673,N_7943,N_9162);
nand U11674 (N_11674,N_6143,N_5076);
nand U11675 (N_11675,N_5879,N_8635);
nand U11676 (N_11676,N_6109,N_7400);
and U11677 (N_11677,N_5594,N_7145);
nand U11678 (N_11678,N_5180,N_8616);
nand U11679 (N_11679,N_7593,N_5415);
and U11680 (N_11680,N_7544,N_5943);
and U11681 (N_11681,N_9603,N_9536);
or U11682 (N_11682,N_5925,N_7370);
xnor U11683 (N_11683,N_9372,N_9154);
nand U11684 (N_11684,N_7323,N_5460);
nor U11685 (N_11685,N_8036,N_8220);
xnor U11686 (N_11686,N_8245,N_8029);
or U11687 (N_11687,N_6166,N_6751);
or U11688 (N_11688,N_6487,N_8837);
xnor U11689 (N_11689,N_8302,N_6532);
xor U11690 (N_11690,N_6925,N_6656);
nor U11691 (N_11691,N_9457,N_7177);
and U11692 (N_11692,N_5121,N_8954);
nand U11693 (N_11693,N_5850,N_8431);
xnor U11694 (N_11694,N_9168,N_9101);
and U11695 (N_11695,N_8117,N_6153);
nand U11696 (N_11696,N_6950,N_8912);
nor U11697 (N_11697,N_9624,N_7383);
or U11698 (N_11698,N_8575,N_9374);
nand U11699 (N_11699,N_6114,N_9341);
and U11700 (N_11700,N_7741,N_8830);
xnor U11701 (N_11701,N_5148,N_5857);
nand U11702 (N_11702,N_7150,N_6981);
xnor U11703 (N_11703,N_9337,N_7404);
and U11704 (N_11704,N_5446,N_5073);
and U11705 (N_11705,N_5561,N_9012);
nand U11706 (N_11706,N_8180,N_8683);
nor U11707 (N_11707,N_9478,N_8087);
and U11708 (N_11708,N_8200,N_8501);
xor U11709 (N_11709,N_9221,N_9719);
nor U11710 (N_11710,N_9974,N_5424);
xnor U11711 (N_11711,N_7227,N_6748);
nand U11712 (N_11712,N_8884,N_9791);
nor U11713 (N_11713,N_8826,N_8964);
nand U11714 (N_11714,N_6584,N_7457);
or U11715 (N_11715,N_5805,N_9785);
or U11716 (N_11716,N_5580,N_6362);
nand U11717 (N_11717,N_5833,N_9006);
xnor U11718 (N_11718,N_5967,N_7992);
nor U11719 (N_11719,N_8696,N_7230);
and U11720 (N_11720,N_9763,N_9321);
or U11721 (N_11721,N_8750,N_9354);
nor U11722 (N_11722,N_5956,N_8030);
nand U11723 (N_11723,N_5720,N_9111);
nand U11724 (N_11724,N_8849,N_5387);
nand U11725 (N_11725,N_5029,N_9848);
xnor U11726 (N_11726,N_9837,N_5376);
xor U11727 (N_11727,N_8021,N_9364);
nor U11728 (N_11728,N_7815,N_6972);
and U11729 (N_11729,N_9373,N_7978);
nor U11730 (N_11730,N_5840,N_8859);
xnor U11731 (N_11731,N_9901,N_6323);
xor U11732 (N_11732,N_8246,N_9580);
xnor U11733 (N_11733,N_6799,N_9520);
and U11734 (N_11734,N_6296,N_8046);
and U11735 (N_11735,N_6942,N_6133);
nor U11736 (N_11736,N_6816,N_5041);
xnor U11737 (N_11737,N_7922,N_8440);
and U11738 (N_11738,N_9932,N_9039);
or U11739 (N_11739,N_6024,N_5755);
xor U11740 (N_11740,N_6875,N_8728);
xnor U11741 (N_11741,N_5452,N_8604);
or U11742 (N_11742,N_8137,N_8429);
nor U11743 (N_11743,N_5096,N_6255);
nor U11744 (N_11744,N_5797,N_5680);
and U11745 (N_11745,N_7693,N_6840);
nand U11746 (N_11746,N_8502,N_9904);
xor U11747 (N_11747,N_7758,N_7019);
nor U11748 (N_11748,N_7834,N_7234);
and U11749 (N_11749,N_9578,N_5077);
nand U11750 (N_11750,N_7005,N_9683);
or U11751 (N_11751,N_8529,N_5343);
or U11752 (N_11752,N_7848,N_8736);
nor U11753 (N_11753,N_9128,N_6768);
and U11754 (N_11754,N_9838,N_7464);
or U11755 (N_11755,N_8874,N_6570);
nor U11756 (N_11756,N_7955,N_6325);
xnor U11757 (N_11757,N_5502,N_9376);
xor U11758 (N_11758,N_8552,N_7753);
and U11759 (N_11759,N_6850,N_8805);
nand U11760 (N_11760,N_8477,N_5356);
or U11761 (N_11761,N_5610,N_9234);
nor U11762 (N_11762,N_9003,N_5819);
xnor U11763 (N_11763,N_5715,N_6623);
or U11764 (N_11764,N_8963,N_5322);
nor U11765 (N_11765,N_7567,N_9895);
nand U11766 (N_11766,N_7462,N_9120);
xnor U11767 (N_11767,N_5068,N_8777);
or U11768 (N_11768,N_5474,N_8446);
or U11769 (N_11769,N_7531,N_8617);
and U11770 (N_11770,N_6510,N_9339);
nor U11771 (N_11771,N_5657,N_7200);
nand U11772 (N_11772,N_8071,N_8233);
xnor U11773 (N_11773,N_8336,N_9511);
and U11774 (N_11774,N_6958,N_8040);
and U11775 (N_11775,N_6225,N_6111);
nor U11776 (N_11776,N_8190,N_8612);
xnor U11777 (N_11777,N_5910,N_6634);
nor U11778 (N_11778,N_7129,N_9407);
or U11779 (N_11779,N_9306,N_8461);
and U11780 (N_11780,N_6409,N_9759);
nand U11781 (N_11781,N_5495,N_7502);
nand U11782 (N_11782,N_8301,N_6483);
and U11783 (N_11783,N_6615,N_8643);
and U11784 (N_11784,N_5441,N_7459);
nand U11785 (N_11785,N_9026,N_9786);
nand U11786 (N_11786,N_7937,N_9532);
nand U11787 (N_11787,N_6082,N_8740);
and U11788 (N_11788,N_8221,N_8864);
and U11789 (N_11789,N_7742,N_5737);
xnor U11790 (N_11790,N_9630,N_9998);
xor U11791 (N_11791,N_7916,N_7762);
nand U11792 (N_11792,N_9245,N_8063);
nand U11793 (N_11793,N_5346,N_7238);
xnor U11794 (N_11794,N_8688,N_5814);
and U11795 (N_11795,N_8091,N_5544);
or U11796 (N_11796,N_9828,N_5968);
and U11797 (N_11797,N_8258,N_6018);
or U11798 (N_11798,N_7020,N_9175);
or U11799 (N_11799,N_9115,N_6592);
and U11800 (N_11800,N_9592,N_9419);
and U11801 (N_11801,N_6042,N_6059);
and U11802 (N_11802,N_8356,N_5164);
nor U11803 (N_11803,N_8591,N_8970);
xnor U11804 (N_11804,N_9054,N_5277);
or U11805 (N_11805,N_8353,N_5017);
nand U11806 (N_11806,N_6940,N_8349);
and U11807 (N_11807,N_6982,N_7659);
nand U11808 (N_11808,N_5591,N_8445);
nand U11809 (N_11809,N_7242,N_6449);
or U11810 (N_11810,N_9602,N_8262);
and U11811 (N_11811,N_9085,N_5996);
and U11812 (N_11812,N_8746,N_7004);
and U11813 (N_11813,N_7537,N_9431);
xnor U11814 (N_11814,N_7946,N_6568);
nand U11815 (N_11815,N_5748,N_8223);
xor U11816 (N_11816,N_9995,N_9405);
or U11817 (N_11817,N_8472,N_7658);
nor U11818 (N_11818,N_9555,N_8229);
nor U11819 (N_11819,N_8563,N_6444);
and U11820 (N_11820,N_9065,N_9126);
xnor U11821 (N_11821,N_5392,N_8842);
xnor U11822 (N_11822,N_7845,N_8163);
nor U11823 (N_11823,N_8710,N_6846);
and U11824 (N_11824,N_9857,N_9051);
and U11825 (N_11825,N_9621,N_5468);
and U11826 (N_11826,N_6187,N_5711);
or U11827 (N_11827,N_6594,N_8109);
and U11828 (N_11828,N_9545,N_5432);
and U11829 (N_11829,N_9869,N_7074);
or U11830 (N_11830,N_6158,N_9931);
or U11831 (N_11831,N_8833,N_8595);
and U11832 (N_11832,N_8154,N_7738);
xnor U11833 (N_11833,N_9565,N_5905);
nand U11834 (N_11834,N_9907,N_9745);
and U11835 (N_11835,N_7516,N_6374);
or U11836 (N_11836,N_5515,N_7576);
xnor U11837 (N_11837,N_9872,N_7680);
nor U11838 (N_11838,N_9829,N_6315);
nor U11839 (N_11839,N_7697,N_7746);
xor U11840 (N_11840,N_8901,N_9658);
xnor U11841 (N_11841,N_6190,N_6955);
and U11842 (N_11842,N_6780,N_6003);
nor U11843 (N_11843,N_5503,N_9157);
and U11844 (N_11844,N_9548,N_7288);
and U11845 (N_11845,N_6097,N_8476);
nand U11846 (N_11846,N_9556,N_6457);
nor U11847 (N_11847,N_5834,N_8102);
nand U11848 (N_11848,N_7935,N_8034);
nand U11849 (N_11849,N_6183,N_6490);
nand U11850 (N_11850,N_8673,N_9702);
and U11851 (N_11851,N_6790,N_9021);
and U11852 (N_11852,N_5652,N_9145);
xnor U11853 (N_11853,N_5089,N_6998);
nand U11854 (N_11854,N_6272,N_9982);
nor U11855 (N_11855,N_7814,N_9655);
xor U11856 (N_11856,N_5063,N_9867);
or U11857 (N_11857,N_5944,N_8678);
nor U11858 (N_11858,N_5305,N_8006);
xor U11859 (N_11859,N_9938,N_5883);
nor U11860 (N_11860,N_5536,N_7523);
nor U11861 (N_11861,N_5158,N_7617);
nor U11862 (N_11862,N_7494,N_6562);
and U11863 (N_11863,N_6754,N_9677);
xnor U11864 (N_11864,N_9599,N_9988);
xor U11865 (N_11865,N_8134,N_6247);
xor U11866 (N_11866,N_7952,N_9970);
or U11867 (N_11867,N_6461,N_9060);
or U11868 (N_11868,N_6313,N_7905);
xnor U11869 (N_11869,N_5856,N_7237);
nor U11870 (N_11870,N_7126,N_5087);
or U11871 (N_11871,N_8434,N_8916);
or U11872 (N_11872,N_7782,N_6664);
and U11873 (N_11873,N_5256,N_5402);
or U11874 (N_11874,N_5803,N_7945);
or U11875 (N_11875,N_7647,N_7012);
or U11876 (N_11876,N_6416,N_5326);
xnor U11877 (N_11877,N_5577,N_7348);
nor U11878 (N_11878,N_9533,N_6514);
nor U11879 (N_11879,N_8389,N_6833);
or U11880 (N_11880,N_5576,N_5961);
nand U11881 (N_11881,N_6041,N_5735);
and U11882 (N_11882,N_5098,N_5181);
or U11883 (N_11883,N_6201,N_8904);
nor U11884 (N_11884,N_9563,N_7769);
or U11885 (N_11885,N_9129,N_6033);
or U11886 (N_11886,N_5912,N_8651);
xor U11887 (N_11887,N_7603,N_8101);
xnor U11888 (N_11888,N_8394,N_8608);
or U11889 (N_11889,N_9340,N_9734);
or U11890 (N_11890,N_9916,N_7033);
nor U11891 (N_11891,N_6050,N_9942);
nand U11892 (N_11892,N_9447,N_6792);
or U11893 (N_11893,N_8799,N_9495);
or U11894 (N_11894,N_6976,N_5448);
nor U11895 (N_11895,N_9681,N_5188);
or U11896 (N_11896,N_7984,N_5477);
or U11897 (N_11897,N_7189,N_9699);
xor U11898 (N_11898,N_7065,N_6651);
and U11899 (N_11899,N_9458,N_5746);
nand U11900 (N_11900,N_7944,N_9194);
nor U11901 (N_11901,N_9414,N_8730);
nor U11902 (N_11902,N_8835,N_9626);
or U11903 (N_11903,N_6064,N_6377);
and U11904 (N_11904,N_8566,N_9367);
xnor U11905 (N_11905,N_6061,N_7882);
and U11906 (N_11906,N_6731,N_9462);
and U11907 (N_11907,N_8176,N_7711);
nor U11908 (N_11908,N_8952,N_8860);
xor U11909 (N_11909,N_6537,N_7409);
nor U11910 (N_11910,N_9118,N_9552);
nand U11911 (N_11911,N_5609,N_8551);
nor U11912 (N_11912,N_7076,N_5133);
xor U11913 (N_11913,N_6159,N_8527);
nand U11914 (N_11914,N_9167,N_5762);
and U11915 (N_11915,N_5824,N_8124);
and U11916 (N_11916,N_7515,N_7369);
xnor U11917 (N_11917,N_6065,N_5151);
nand U11918 (N_11918,N_6774,N_6841);
nor U11919 (N_11919,N_7510,N_8135);
and U11920 (N_11920,N_6182,N_5184);
or U11921 (N_11921,N_5086,N_6730);
nor U11922 (N_11922,N_5454,N_6316);
xor U11923 (N_11923,N_9053,N_9842);
nor U11924 (N_11924,N_9329,N_7483);
xor U11925 (N_11925,N_8161,N_8605);
nand U11926 (N_11926,N_7175,N_7689);
nor U11927 (N_11927,N_5602,N_5288);
or U11928 (N_11928,N_5825,N_7240);
and U11929 (N_11929,N_8510,N_6949);
or U11930 (N_11930,N_8309,N_7789);
and U11931 (N_11931,N_9139,N_8487);
xnor U11932 (N_11932,N_7111,N_5227);
nand U11933 (N_11933,N_9134,N_7139);
nor U11934 (N_11934,N_6639,N_9636);
nand U11935 (N_11935,N_7338,N_6207);
and U11936 (N_11936,N_7549,N_7855);
nand U11937 (N_11937,N_9775,N_7251);
nand U11938 (N_11938,N_7519,N_7760);
xor U11939 (N_11939,N_6980,N_5420);
nand U11940 (N_11940,N_9684,N_6469);
nor U11941 (N_11941,N_9392,N_5966);
or U11942 (N_11942,N_9585,N_8815);
and U11943 (N_11943,N_7366,N_8453);
and U11944 (N_11944,N_5409,N_6198);
nand U11945 (N_11945,N_5046,N_6071);
nand U11946 (N_11946,N_5649,N_5936);
nor U11947 (N_11947,N_6936,N_7402);
xor U11948 (N_11948,N_6798,N_5369);
nand U11949 (N_11949,N_9575,N_6245);
xor U11950 (N_11950,N_7060,N_7562);
nor U11951 (N_11951,N_8119,N_8285);
nand U11952 (N_11952,N_9389,N_9815);
or U11953 (N_11953,N_9802,N_7649);
nand U11954 (N_11954,N_6481,N_9811);
nand U11955 (N_11955,N_9863,N_9439);
xnor U11956 (N_11956,N_5959,N_7641);
nor U11957 (N_11957,N_8026,N_5458);
xnor U11958 (N_11958,N_7439,N_8239);
nor U11959 (N_11959,N_8449,N_5405);
and U11960 (N_11960,N_8692,N_8582);
nor U11961 (N_11961,N_8940,N_9324);
nand U11962 (N_11962,N_5047,N_9731);
nand U11963 (N_11963,N_7224,N_6926);
nor U11964 (N_11964,N_9955,N_6725);
xnor U11965 (N_11965,N_5142,N_9290);
and U11966 (N_11966,N_7811,N_6914);
and U11967 (N_11967,N_5104,N_8934);
xor U11968 (N_11968,N_5621,N_6595);
nor U11969 (N_11969,N_6617,N_8531);
nor U11970 (N_11970,N_8519,N_5311);
xor U11971 (N_11971,N_8852,N_8170);
and U11972 (N_11972,N_7962,N_6338);
and U11973 (N_11973,N_6697,N_5733);
nand U11974 (N_11974,N_8542,N_9738);
or U11975 (N_11975,N_7467,N_8295);
xnor U11976 (N_11976,N_8236,N_9310);
nor U11977 (N_11977,N_5398,N_8214);
or U11978 (N_11978,N_7833,N_7933);
or U11979 (N_11979,N_9813,N_9380);
xnor U11980 (N_11980,N_5161,N_7201);
or U11981 (N_11981,N_5517,N_5871);
and U11982 (N_11982,N_5646,N_9737);
and U11983 (N_11983,N_9030,N_8317);
and U11984 (N_11984,N_6549,N_5848);
or U11985 (N_11985,N_6388,N_5306);
nand U11986 (N_11986,N_6647,N_6216);
nand U11987 (N_11987,N_7061,N_5135);
or U11988 (N_11988,N_8640,N_7214);
nand U11989 (N_11989,N_9754,N_7386);
xnor U11990 (N_11990,N_6693,N_5874);
and U11991 (N_11991,N_5836,N_8182);
or U11992 (N_11992,N_8961,N_6363);
nand U11993 (N_11993,N_7279,N_9825);
nand U11994 (N_11994,N_5439,N_8380);
nor U11995 (N_11995,N_5974,N_7837);
nand U11996 (N_11996,N_6324,N_9470);
or U11997 (N_11997,N_6177,N_6212);
nand U11998 (N_11998,N_9985,N_6566);
or U11999 (N_11999,N_5303,N_7873);
nor U12000 (N_12000,N_6673,N_6635);
and U12001 (N_12001,N_7585,N_8981);
nand U12002 (N_12002,N_5866,N_8020);
nor U12003 (N_12003,N_9969,N_7358);
nand U12004 (N_12004,N_7319,N_6123);
nand U12005 (N_12005,N_5599,N_8468);
nand U12006 (N_12006,N_9686,N_5008);
xnor U12007 (N_12007,N_5628,N_7379);
and U12008 (N_12008,N_9612,N_7158);
and U12009 (N_12009,N_7451,N_6653);
nand U12010 (N_12010,N_8517,N_9631);
xnor U12011 (N_12011,N_7269,N_8334);
or U12012 (N_12012,N_7691,N_9986);
xnor U12013 (N_12013,N_9123,N_9840);
nor U12014 (N_12014,N_7342,N_9342);
or U12015 (N_12015,N_5247,N_8227);
nor U12016 (N_12016,N_5137,N_8654);
nand U12017 (N_12017,N_5106,N_9218);
or U12018 (N_12018,N_9489,N_7541);
or U12019 (N_12019,N_7007,N_7685);
or U12020 (N_12020,N_5747,N_9428);
or U12021 (N_12021,N_6579,N_8078);
nand U12022 (N_12022,N_5217,N_8655);
or U12023 (N_12023,N_6168,N_9114);
xor U12024 (N_12024,N_7822,N_6529);
or U12025 (N_12025,N_7669,N_7361);
and U12026 (N_12026,N_9728,N_9474);
nand U12027 (N_12027,N_7871,N_9028);
nor U12028 (N_12028,N_6349,N_8929);
or U12029 (N_12029,N_9070,N_6586);
nor U12030 (N_12030,N_5567,N_7026);
xnor U12031 (N_12031,N_8757,N_7744);
nor U12032 (N_12032,N_7764,N_5511);
xor U12033 (N_12033,N_9263,N_5105);
nor U12034 (N_12034,N_6737,N_6004);
and U12035 (N_12035,N_8235,N_7911);
nand U12036 (N_12036,N_8103,N_9984);
or U12037 (N_12037,N_7793,N_5991);
nor U12038 (N_12038,N_8921,N_6616);
xor U12039 (N_12039,N_5036,N_6685);
xor U12040 (N_12040,N_9434,N_7051);
or U12041 (N_12041,N_9650,N_9052);
and U12042 (N_12042,N_7930,N_5368);
and U12043 (N_12043,N_6078,N_7030);
and U12044 (N_12044,N_8164,N_5522);
and U12045 (N_12045,N_7588,N_7551);
nor U12046 (N_12046,N_9275,N_8886);
nand U12047 (N_12047,N_6376,N_7447);
xnor U12048 (N_12048,N_7684,N_5361);
and U12049 (N_12049,N_6070,N_5287);
and U12050 (N_12050,N_9518,N_9176);
and U12051 (N_12051,N_5743,N_6814);
or U12052 (N_12052,N_9460,N_7574);
nand U12053 (N_12053,N_7405,N_6749);
or U12054 (N_12054,N_8355,N_6675);
or U12055 (N_12055,N_6810,N_9896);
and U12056 (N_12056,N_7595,N_7294);
and U12057 (N_12057,N_5150,N_6355);
nand U12058 (N_12058,N_9806,N_5728);
nor U12059 (N_12059,N_5672,N_8329);
xnor U12060 (N_12060,N_9378,N_9420);
xnor U12061 (N_12061,N_9530,N_8623);
or U12062 (N_12062,N_7172,N_8433);
or U12063 (N_12063,N_7478,N_6403);
or U12064 (N_12064,N_9048,N_5206);
nor U12065 (N_12065,N_8442,N_9648);
or U12066 (N_12066,N_9035,N_8480);
nand U12067 (N_12067,N_6620,N_5664);
xor U12068 (N_12068,N_9472,N_8949);
or U12069 (N_12069,N_8979,N_7003);
or U12070 (N_12070,N_5828,N_5314);
xnor U12071 (N_12071,N_9966,N_5663);
nor U12072 (N_12072,N_8672,N_8075);
and U12073 (N_12073,N_5955,N_8066);
or U12074 (N_12074,N_6881,N_9425);
xor U12075 (N_12075,N_5921,N_6745);
nand U12076 (N_12076,N_8254,N_8547);
nand U12077 (N_12077,N_8614,N_7471);
or U12078 (N_12078,N_9635,N_9992);
nand U12079 (N_12079,N_5023,N_9079);
nand U12080 (N_12080,N_5498,N_7270);
and U12081 (N_12081,N_8209,N_9689);
nand U12082 (N_12082,N_6628,N_7856);
nand U12083 (N_12083,N_8646,N_8661);
xor U12084 (N_12084,N_6139,N_8571);
or U12085 (N_12085,N_7835,N_7975);
nor U12086 (N_12086,N_6648,N_6507);
and U12087 (N_12087,N_6241,N_9494);
nor U12088 (N_12088,N_7902,N_7176);
nand U12089 (N_12089,N_7870,N_7505);
nand U12090 (N_12090,N_9099,N_5058);
nor U12091 (N_12091,N_6627,N_9558);
nand U12092 (N_12092,N_7041,N_7624);
nor U12093 (N_12093,N_5995,N_7055);
and U12094 (N_12094,N_8463,N_7493);
nor U12095 (N_12095,N_9866,N_9542);
or U12096 (N_12096,N_8909,N_8496);
nor U12097 (N_12097,N_8602,N_5695);
or U12098 (N_12098,N_5619,N_5506);
nand U12099 (N_12099,N_5241,N_6939);
and U12100 (N_12100,N_7627,N_8018);
or U12101 (N_12101,N_7853,N_5574);
and U12102 (N_12102,N_7524,N_6379);
nor U12103 (N_12103,N_6758,N_7213);
xnor U12104 (N_12104,N_9004,N_7629);
nand U12105 (N_12105,N_5083,N_7432);
nand U12106 (N_12106,N_8210,N_7542);
and U12107 (N_12107,N_9743,N_8989);
or U12108 (N_12108,N_9727,N_6373);
or U12109 (N_12109,N_5232,N_6452);
and U12110 (N_12110,N_9835,N_9586);
or U12111 (N_12111,N_7157,N_9934);
nand U12112 (N_12112,N_7081,N_5759);
xnor U12113 (N_12113,N_8012,N_9962);
xor U12114 (N_12114,N_7034,N_7802);
and U12115 (N_12115,N_6174,N_5842);
nand U12116 (N_12116,N_8357,N_6502);
nor U12117 (N_12117,N_7153,N_9174);
nor U12118 (N_12118,N_9666,N_5453);
nor U12119 (N_12119,N_8521,N_8791);
nand U12120 (N_12120,N_8881,N_8410);
and U12121 (N_12121,N_9742,N_5486);
xor U12122 (N_12122,N_8304,N_8019);
and U12123 (N_12123,N_5471,N_7664);
xor U12124 (N_12124,N_5283,N_8903);
nand U12125 (N_12125,N_7354,N_7718);
nor U12126 (N_12126,N_7465,N_7973);
or U12127 (N_12127,N_8634,N_5791);
and U12128 (N_12128,N_7428,N_9105);
nand U12129 (N_12129,N_7473,N_8926);
nor U12130 (N_12130,N_5816,N_8873);
xor U12131 (N_12131,N_8483,N_9142);
xor U12132 (N_12132,N_8024,N_8592);
nand U12133 (N_12133,N_9116,N_5204);
nor U12134 (N_12134,N_5464,N_6276);
or U12135 (N_12135,N_6161,N_5081);
and U12136 (N_12136,N_5982,N_9043);
or U12137 (N_12137,N_5662,N_5620);
nor U12138 (N_12138,N_9368,N_6680);
or U12139 (N_12139,N_6803,N_6289);
nor U12140 (N_12140,N_6784,N_9027);
nor U12141 (N_12141,N_8694,N_6398);
or U12142 (N_12142,N_9589,N_8942);
nor U12143 (N_12143,N_6234,N_6901);
nand U12144 (N_12144,N_7512,N_5211);
xnor U12145 (N_12145,N_9464,N_9674);
and U12146 (N_12146,N_5349,N_7601);
nand U12147 (N_12147,N_5526,N_5333);
nand U12148 (N_12148,N_8207,N_7122);
nor U12149 (N_12149,N_5902,N_9279);
nor U12150 (N_12150,N_7538,N_7021);
nand U12151 (N_12151,N_9415,N_5624);
xor U12152 (N_12152,N_5847,N_8868);
and U12153 (N_12153,N_5014,N_7587);
or U12154 (N_12154,N_5831,N_9761);
nand U12155 (N_12155,N_9403,N_5661);
or U12156 (N_12156,N_9033,N_9736);
or U12157 (N_12157,N_5738,N_8296);
nand U12158 (N_12158,N_9206,N_8631);
or U12159 (N_12159,N_8762,N_5282);
nand U12160 (N_12160,N_8668,N_5897);
xnor U12161 (N_12161,N_5380,N_9486);
or U12162 (N_12162,N_5681,N_6800);
xnor U12163 (N_12163,N_9531,N_6839);
xnor U12164 (N_12164,N_9886,N_7884);
xor U12165 (N_12165,N_7144,N_6852);
nand U12166 (N_12166,N_8252,N_8339);
nor U12167 (N_12167,N_5585,N_5239);
nor U12168 (N_12168,N_5169,N_9074);
xnor U12169 (N_12169,N_9713,N_6429);
nor U12170 (N_12170,N_6136,N_7421);
or U12171 (N_12171,N_9381,N_6793);
and U12172 (N_12172,N_7262,N_6838);
nand U12173 (N_12173,N_5799,N_7626);
and U12174 (N_12174,N_8230,N_7287);
and U12175 (N_12175,N_8641,N_6054);
nand U12176 (N_12176,N_7125,N_7798);
or U12177 (N_12177,N_7300,N_5904);
nor U12178 (N_12178,N_5978,N_8372);
xnor U12179 (N_12179,N_5359,N_5500);
or U12180 (N_12180,N_6821,N_8147);
xnor U12181 (N_12181,N_6494,N_6503);
xor U12182 (N_12182,N_9550,N_7543);
or U12183 (N_12183,N_6953,N_8249);
and U12184 (N_12184,N_5413,N_7688);
xor U12185 (N_12185,N_8035,N_8268);
nand U12186 (N_12186,N_6072,N_5355);
and U12187 (N_12187,N_9211,N_8839);
or U12188 (N_12188,N_9000,N_7891);
nor U12189 (N_12189,N_5665,N_7490);
xor U12190 (N_12190,N_7042,N_8980);
nand U12191 (N_12191,N_7043,N_8744);
or U12192 (N_12192,N_8541,N_8148);
and U12193 (N_12193,N_7564,N_9161);
nand U12194 (N_12194,N_9833,N_8875);
nand U12195 (N_12195,N_7865,N_5550);
nand U12196 (N_12196,N_8398,N_6440);
nand U12197 (N_12197,N_7083,N_8520);
or U12198 (N_12198,N_6286,N_5821);
nand U12199 (N_12199,N_7568,N_7401);
and U12200 (N_12200,N_5374,N_8983);
nand U12201 (N_12201,N_9861,N_7266);
nor U12202 (N_12202,N_5919,N_9156);
nand U12203 (N_12203,N_8068,N_7154);
nand U12204 (N_12204,N_5945,N_5102);
xnor U12205 (N_12205,N_5607,N_5707);
nand U12206 (N_12206,N_6528,N_9718);
nor U12207 (N_12207,N_8943,N_6518);
xnor U12208 (N_12208,N_8951,N_9618);
xor U12209 (N_12209,N_5950,N_9912);
nand U12210 (N_12210,N_9595,N_9744);
or U12211 (N_12211,N_7011,N_7164);
or U12212 (N_12212,N_8987,N_7580);
nand U12213 (N_12213,N_8305,N_8374);
nor U12214 (N_12214,N_8466,N_8128);
nor U12215 (N_12215,N_5496,N_6368);
and U12216 (N_12216,N_7343,N_5771);
and U12217 (N_12217,N_6427,N_6278);
or U12218 (N_12218,N_8810,N_7528);
or U12219 (N_12219,N_5597,N_7740);
xor U12220 (N_12220,N_5042,N_5731);
nor U12221 (N_12221,N_6978,N_8530);
nor U12222 (N_12222,N_8741,N_8577);
nor U12223 (N_12223,N_5433,N_5265);
nand U12224 (N_12224,N_7104,N_9346);
nand U12225 (N_12225,N_7750,N_9455);
and U12226 (N_12226,N_9773,N_9140);
and U12227 (N_12227,N_6083,N_6389);
nor U12228 (N_12228,N_9183,N_5952);
nor U12229 (N_12229,N_8768,N_9959);
and U12230 (N_12230,N_8074,N_6837);
and U12231 (N_12231,N_9179,N_9238);
and U12232 (N_12232,N_6333,N_7997);
nor U12233 (N_12233,N_5318,N_8503);
and U12234 (N_12234,N_8277,N_5788);
nand U12235 (N_12235,N_5935,N_8325);
nor U12236 (N_12236,N_6672,N_9436);
xor U12237 (N_12237,N_9311,N_6539);
and U12238 (N_12238,N_5174,N_8089);
nor U12239 (N_12239,N_7639,N_8950);
nand U12240 (N_12240,N_6869,N_8441);
and U12241 (N_12241,N_7532,N_6250);
nand U12242 (N_12242,N_9153,N_6557);
and U12243 (N_12243,N_9276,N_7321);
and U12244 (N_12244,N_6999,N_6676);
nor U12245 (N_12245,N_9463,N_5199);
nor U12246 (N_12246,N_6396,N_9087);
and U12247 (N_12247,N_9741,N_5780);
nand U12248 (N_12248,N_6938,N_5171);
xnor U12249 (N_12249,N_7572,N_5483);
nand U12250 (N_12250,N_8499,N_7376);
nor U12251 (N_12251,N_6782,N_6665);
xor U12252 (N_12252,N_5644,N_6724);
nor U12253 (N_12253,N_9654,N_5712);
nor U12254 (N_12254,N_7570,N_6576);
xnor U12255 (N_12255,N_8382,N_8206);
nor U12256 (N_12256,N_6378,N_6961);
or U12257 (N_12257,N_6797,N_7063);
nand U12258 (N_12258,N_9408,N_5316);
nand U12259 (N_12259,N_9920,N_8406);
nand U12260 (N_12260,N_6755,N_6246);
and U12261 (N_12261,N_6742,N_6155);
xor U12262 (N_12262,N_8783,N_9535);
and U12263 (N_12263,N_6098,N_5985);
xor U12264 (N_12264,N_6122,N_6985);
nand U12265 (N_12265,N_5769,N_5894);
nor U12266 (N_12266,N_9141,N_5571);
or U12267 (N_12267,N_7233,N_7706);
or U12268 (N_12268,N_7982,N_9831);
nand U12269 (N_12269,N_9797,N_5294);
or U12270 (N_12270,N_9793,N_8422);
nand U12271 (N_12271,N_8648,N_8067);
xor U12272 (N_12272,N_8706,N_6381);
nor U12273 (N_12273,N_5421,N_9653);
or U12274 (N_12274,N_5957,N_7816);
xnor U12275 (N_12275,N_9353,N_9807);
or U12276 (N_12276,N_5499,N_6563);
and U12277 (N_12277,N_7661,N_8275);
or U12278 (N_12278,N_8896,N_7124);
nand U12279 (N_12279,N_7315,N_6505);
xnor U12280 (N_12280,N_7372,N_9289);
nor U12281 (N_12281,N_8823,N_9926);
and U12282 (N_12282,N_9398,N_7062);
or U12283 (N_12283,N_6923,N_6460);
or U12284 (N_12284,N_8426,N_6049);
and U12285 (N_12285,N_7854,N_8240);
xnor U12286 (N_12286,N_8735,N_8780);
nor U12287 (N_12287,N_9102,N_5864);
xor U12288 (N_12288,N_6165,N_5450);
and U12289 (N_12289,N_5687,N_5091);
and U12290 (N_12290,N_9484,N_9859);
xnor U12291 (N_12291,N_7073,N_7752);
or U12292 (N_12292,N_5261,N_9930);
or U12293 (N_12293,N_8322,N_8567);
nor U12294 (N_12294,N_8653,N_9700);
nand U12295 (N_12295,N_6347,N_5648);
nand U12296 (N_12296,N_5729,N_9524);
xnor U12297 (N_12297,N_6046,N_5772);
xor U12298 (N_12298,N_6010,N_6859);
or U12299 (N_12299,N_6170,N_8364);
nor U12300 (N_12300,N_8242,N_8253);
xor U12301 (N_12301,N_5559,N_7277);
nand U12302 (N_12302,N_7566,N_7078);
and U12303 (N_12303,N_7193,N_6854);
or U12304 (N_12304,N_5304,N_5146);
nor U12305 (N_12305,N_8585,N_9069);
and U12306 (N_12306,N_5079,N_6888);
or U12307 (N_12307,N_8512,N_9418);
nor U12308 (N_12308,N_6451,N_5880);
and U12309 (N_12309,N_8578,N_6340);
nor U12310 (N_12310,N_7091,N_5907);
and U12311 (N_12311,N_7444,N_5598);
and U12312 (N_12312,N_9360,N_5345);
or U12313 (N_12313,N_5761,N_8806);
and U12314 (N_12314,N_7719,N_8994);
xor U12315 (N_12315,N_7167,N_9433);
and U12316 (N_12316,N_7773,N_9300);
nor U12317 (N_12317,N_8879,N_8558);
and U12318 (N_12318,N_5172,N_9034);
and U12319 (N_12319,N_6917,N_6387);
nand U12320 (N_12320,N_5914,N_7272);
and U12321 (N_12321,N_8250,N_7785);
nand U12322 (N_12322,N_5989,N_8885);
nand U12323 (N_12323,N_8131,N_9843);
xor U12324 (N_12324,N_6669,N_6470);
or U12325 (N_12325,N_9394,N_9285);
nor U12326 (N_12326,N_8553,N_5588);
and U12327 (N_12327,N_9725,N_5470);
nor U12328 (N_12328,N_6613,N_9967);
nor U12329 (N_12329,N_8416,N_5691);
or U12330 (N_12330,N_7470,N_5350);
nand U12331 (N_12331,N_6322,N_6277);
nand U12332 (N_12332,N_8384,N_5497);
xnor U12333 (N_12333,N_6771,N_9318);
nor U12334 (N_12334,N_9640,N_8055);
nand U12335 (N_12335,N_5786,N_6806);
nand U12336 (N_12336,N_5841,N_6637);
and U12337 (N_12337,N_6036,N_8037);
nand U12338 (N_12338,N_9645,N_7827);
nor U12339 (N_12339,N_6986,N_5573);
or U12340 (N_12340,N_9781,N_7622);
nand U12341 (N_12341,N_6657,N_8931);
xor U12342 (N_12342,N_8002,N_9225);
xnor U12343 (N_12343,N_5119,N_8286);
or U12344 (N_12344,N_9169,N_8473);
and U12345 (N_12345,N_9887,N_8855);
xnor U12346 (N_12346,N_9112,N_5337);
nand U12347 (N_12347,N_8716,N_6670);
or U12348 (N_12348,N_5373,N_9164);
nand U12349 (N_12349,N_8685,N_9714);
nor U12350 (N_12350,N_7072,N_8771);
and U12351 (N_12351,N_5698,N_6694);
nor U12352 (N_12352,N_5012,N_8232);
or U12353 (N_12353,N_7301,N_7137);
nand U12354 (N_12354,N_6701,N_7525);
nand U12355 (N_12355,N_6086,N_7336);
xnor U12356 (N_12356,N_6314,N_7086);
nor U12357 (N_12357,N_5166,N_5170);
nor U12358 (N_12358,N_7986,N_8674);
and U12359 (N_12359,N_7849,N_7683);
and U12360 (N_12360,N_6602,N_9946);
nand U12361 (N_12361,N_8960,N_7442);
or U12362 (N_12362,N_5039,N_6572);
nor U12363 (N_12363,N_6979,N_8183);
or U12364 (N_12364,N_6384,N_9023);
and U12365 (N_12365,N_7298,N_8573);
nor U12366 (N_12366,N_6865,N_5233);
xnor U12367 (N_12367,N_6684,N_5309);
nor U12368 (N_12368,N_7415,N_7466);
xnor U12369 (N_12369,N_7384,N_9994);
nor U12370 (N_12370,N_5658,N_6994);
nor U12371 (N_12371,N_6354,N_8745);
nand U12372 (N_12372,N_7293,N_8151);
nand U12373 (N_12373,N_5808,N_7169);
nand U12374 (N_12374,N_6943,N_7969);
nand U12375 (N_12375,N_7049,N_8224);
nand U12376 (N_12376,N_7097,N_7070);
nand U12377 (N_12377,N_9779,N_6454);
xor U12378 (N_12378,N_7437,N_6543);
and U12379 (N_12379,N_8923,N_6258);
nand U12380 (N_12380,N_6101,N_9593);
or U12381 (N_12381,N_8613,N_9832);
or U12382 (N_12382,N_7179,N_9804);
nand U12383 (N_12383,N_9927,N_8947);
nand U12384 (N_12384,N_9569,N_8498);
and U12385 (N_12385,N_6716,N_9997);
nor U12386 (N_12386,N_5025,N_9508);
and U12387 (N_12387,N_9526,N_6006);
nand U12388 (N_12388,N_7956,N_7461);
and U12389 (N_12389,N_5147,N_6028);
xor U12390 (N_12390,N_8174,N_8451);
xor U12391 (N_12391,N_9820,N_8838);
nor U12392 (N_12392,N_6582,N_9483);
and U12393 (N_12393,N_9752,N_8800);
and U12394 (N_12394,N_8537,N_6916);
xnor U12395 (N_12395,N_9770,N_5740);
and U12396 (N_12396,N_6641,N_8333);
and U12397 (N_12397,N_5308,N_8194);
xor U12398 (N_12398,N_9673,N_7331);
or U12399 (N_12399,N_7823,N_7032);
xor U12400 (N_12400,N_6169,N_9444);
nand U12401 (N_12401,N_6744,N_7349);
nor U12402 (N_12402,N_5457,N_6548);
nor U12403 (N_12403,N_9882,N_6326);
and U12404 (N_12404,N_5478,N_9155);
nand U12405 (N_12405,N_5948,N_8198);
nand U12406 (N_12406,N_6706,N_7646);
xor U12407 (N_12407,N_8010,N_9487);
xor U12408 (N_12408,N_9150,N_8702);
or U12409 (N_12409,N_9822,N_7035);
and U12410 (N_12410,N_7919,N_7152);
nand U12411 (N_12411,N_6555,N_6608);
nand U12412 (N_12412,N_9915,N_6089);
xnor U12413 (N_12413,N_6559,N_8007);
xnor U12414 (N_12414,N_8351,N_9513);
nor U12415 (N_12415,N_5436,N_5238);
and U12416 (N_12416,N_8100,N_9288);
or U12417 (N_12417,N_8769,N_6581);
or U12418 (N_12418,N_7928,N_7304);
and U12419 (N_12419,N_7110,N_6418);
and U12420 (N_12420,N_7412,N_5750);
nand U12421 (N_12421,N_8691,N_9950);
xnor U12422 (N_12422,N_9830,N_7392);
and U12423 (N_12423,N_8316,N_6327);
and U12424 (N_12424,N_7981,N_5229);
nand U12425 (N_12425,N_5295,N_5702);
xor U12426 (N_12426,N_6135,N_9576);
nand U12427 (N_12427,N_8120,N_8173);
nand U12428 (N_12428,N_8315,N_8606);
or U12429 (N_12429,N_8676,N_5999);
or U12430 (N_12430,N_6474,N_9049);
or U12431 (N_12431,N_9325,N_9260);
and U12432 (N_12432,N_6622,N_7271);
xnor U12433 (N_12433,N_6534,N_6108);
nand U12434 (N_12434,N_9614,N_5802);
xor U12435 (N_12435,N_6146,N_6508);
and U12436 (N_12436,N_9046,N_6149);
nor U12437 (N_12437,N_6300,N_8717);
nor U12438 (N_12438,N_5143,N_8082);
or U12439 (N_12439,N_7831,N_8797);
or U12440 (N_12440,N_7723,N_7244);
nor U12441 (N_12441,N_7721,N_9767);
nand U12442 (N_12442,N_5370,N_6970);
nand U12443 (N_12443,N_8193,N_9292);
or U12444 (N_12444,N_8657,N_6038);
and U12445 (N_12445,N_5979,N_9504);
xor U12446 (N_12446,N_7463,N_6597);
or U12447 (N_12447,N_6342,N_9710);
xnor U12448 (N_12448,N_9467,N_6964);
nand U12449 (N_12449,N_8113,N_7187);
xnor U12450 (N_12450,N_9616,N_5793);
nor U12451 (N_12451,N_6818,N_9810);
nand U12452 (N_12452,N_8966,N_7677);
and U12453 (N_12453,N_8397,N_5901);
and U12454 (N_12454,N_5903,N_6281);
nand U12455 (N_12455,N_9222,N_9247);
and U12456 (N_12456,N_9347,N_6203);
nand U12457 (N_12457,N_5209,N_9429);
nor U12458 (N_12458,N_6345,N_7077);
and U12459 (N_12459,N_6533,N_8622);
nand U12460 (N_12460,N_9572,N_8927);
nor U12461 (N_12461,N_8064,N_8028);
and U12462 (N_12462,N_6415,N_9296);
or U12463 (N_12463,N_7395,N_7530);
or U12464 (N_12464,N_8407,N_8350);
or U12465 (N_12465,N_7501,N_8784);
or U12466 (N_12466,N_5546,N_5035);
xor U12467 (N_12467,N_6930,N_9515);
or U12468 (N_12468,N_5584,N_6260);
nor U12469 (N_12469,N_9005,N_6815);
nor U12470 (N_12470,N_7330,N_7874);
nor U12471 (N_12471,N_5527,N_6844);
and U12472 (N_12472,N_9510,N_6261);
xor U12473 (N_12473,N_9173,N_7047);
xor U12474 (N_12474,N_8817,N_6786);
xor U12475 (N_12475,N_7123,N_8637);
nor U12476 (N_12476,N_6244,N_5997);
xor U12477 (N_12477,N_5254,N_6801);
nor U12478 (N_12478,N_6209,N_9196);
nor U12479 (N_12479,N_7976,N_7707);
nor U12480 (N_12480,N_7918,N_6499);
xnor U12481 (N_12481,N_9375,N_5723);
and U12482 (N_12482,N_7250,N_6826);
or U12483 (N_12483,N_5026,N_6482);
nand U12484 (N_12484,N_6516,N_6067);
and U12485 (N_12485,N_6593,N_9466);
nand U12486 (N_12486,N_6857,N_5886);
and U12487 (N_12487,N_7195,N_9712);
and U12488 (N_12488,N_7794,N_6238);
and U12489 (N_12489,N_8536,N_5813);
xnor U12490 (N_12490,N_6956,N_7766);
and U12491 (N_12491,N_5007,N_5313);
xnor U12492 (N_12492,N_9210,N_6902);
xor U12493 (N_12493,N_8712,N_8773);
and U12494 (N_12494,N_7314,N_5653);
and U12495 (N_12495,N_6055,N_8474);
and U12496 (N_12496,N_7533,N_8645);
and U12497 (N_12497,N_5097,N_8186);
nand U12498 (N_12498,N_6513,N_5725);
or U12499 (N_12499,N_8436,N_5300);
and U12500 (N_12500,N_6022,N_8284);
or U12501 (N_12501,N_7912,N_5995);
nand U12502 (N_12502,N_9646,N_8597);
or U12503 (N_12503,N_6030,N_9337);
and U12504 (N_12504,N_8369,N_9417);
or U12505 (N_12505,N_6044,N_7930);
xnor U12506 (N_12506,N_5781,N_6979);
nor U12507 (N_12507,N_7462,N_8255);
or U12508 (N_12508,N_5036,N_9166);
nor U12509 (N_12509,N_5691,N_6949);
or U12510 (N_12510,N_6783,N_5027);
or U12511 (N_12511,N_8216,N_5145);
nor U12512 (N_12512,N_8428,N_5705);
nor U12513 (N_12513,N_9237,N_9541);
and U12514 (N_12514,N_8895,N_5941);
nand U12515 (N_12515,N_5713,N_8517);
nor U12516 (N_12516,N_8670,N_5314);
nand U12517 (N_12517,N_8126,N_9016);
nand U12518 (N_12518,N_9925,N_5361);
or U12519 (N_12519,N_6280,N_9136);
nand U12520 (N_12520,N_9756,N_6380);
xnor U12521 (N_12521,N_7048,N_7437);
nand U12522 (N_12522,N_5657,N_7228);
nand U12523 (N_12523,N_8306,N_7688);
nor U12524 (N_12524,N_9552,N_9844);
or U12525 (N_12525,N_6618,N_9118);
xnor U12526 (N_12526,N_5214,N_5428);
nand U12527 (N_12527,N_6727,N_6061);
nand U12528 (N_12528,N_5012,N_5863);
nand U12529 (N_12529,N_9949,N_5276);
xnor U12530 (N_12530,N_5453,N_7753);
nand U12531 (N_12531,N_9130,N_9849);
and U12532 (N_12532,N_7747,N_5873);
nor U12533 (N_12533,N_9079,N_7084);
or U12534 (N_12534,N_8264,N_8309);
or U12535 (N_12535,N_5301,N_6747);
xor U12536 (N_12536,N_6300,N_9763);
nor U12537 (N_12537,N_9543,N_7502);
xnor U12538 (N_12538,N_7643,N_9579);
nor U12539 (N_12539,N_9352,N_6644);
or U12540 (N_12540,N_9763,N_5307);
nor U12541 (N_12541,N_9304,N_8419);
and U12542 (N_12542,N_5478,N_9051);
nand U12543 (N_12543,N_8217,N_9890);
nand U12544 (N_12544,N_5392,N_8643);
xor U12545 (N_12545,N_8986,N_8335);
nand U12546 (N_12546,N_8622,N_8370);
or U12547 (N_12547,N_6050,N_5786);
and U12548 (N_12548,N_5019,N_7774);
nor U12549 (N_12549,N_7389,N_6339);
nor U12550 (N_12550,N_7110,N_8261);
xor U12551 (N_12551,N_8786,N_7476);
nand U12552 (N_12552,N_9902,N_6910);
and U12553 (N_12553,N_7335,N_6281);
nand U12554 (N_12554,N_6998,N_9779);
nand U12555 (N_12555,N_6999,N_8054);
xor U12556 (N_12556,N_5474,N_6219);
nand U12557 (N_12557,N_9953,N_8059);
xor U12558 (N_12558,N_6575,N_8749);
or U12559 (N_12559,N_8359,N_7216);
nand U12560 (N_12560,N_5676,N_6967);
nor U12561 (N_12561,N_8291,N_9700);
and U12562 (N_12562,N_7781,N_8743);
or U12563 (N_12563,N_5808,N_9912);
and U12564 (N_12564,N_8666,N_8072);
and U12565 (N_12565,N_8648,N_7941);
nor U12566 (N_12566,N_6869,N_7947);
or U12567 (N_12567,N_9272,N_9585);
xnor U12568 (N_12568,N_5266,N_6355);
xor U12569 (N_12569,N_5662,N_9989);
xnor U12570 (N_12570,N_8398,N_6622);
nor U12571 (N_12571,N_9573,N_7290);
nand U12572 (N_12572,N_9110,N_7285);
nand U12573 (N_12573,N_9401,N_7765);
or U12574 (N_12574,N_5406,N_5504);
and U12575 (N_12575,N_6825,N_9403);
or U12576 (N_12576,N_6942,N_9990);
xnor U12577 (N_12577,N_5039,N_6819);
nand U12578 (N_12578,N_7287,N_6952);
nor U12579 (N_12579,N_8121,N_5604);
xor U12580 (N_12580,N_8330,N_9615);
xor U12581 (N_12581,N_7635,N_9810);
and U12582 (N_12582,N_5801,N_9837);
or U12583 (N_12583,N_6319,N_6820);
nand U12584 (N_12584,N_5833,N_7821);
nand U12585 (N_12585,N_8946,N_5695);
xnor U12586 (N_12586,N_8571,N_9214);
nand U12587 (N_12587,N_5376,N_6635);
xnor U12588 (N_12588,N_9948,N_5248);
or U12589 (N_12589,N_7873,N_6830);
nand U12590 (N_12590,N_9664,N_9179);
nor U12591 (N_12591,N_9998,N_6627);
or U12592 (N_12592,N_9257,N_5637);
and U12593 (N_12593,N_7471,N_5111);
and U12594 (N_12594,N_8996,N_8404);
and U12595 (N_12595,N_5468,N_8608);
or U12596 (N_12596,N_7646,N_8978);
nor U12597 (N_12597,N_8154,N_6010);
or U12598 (N_12598,N_8377,N_7429);
nor U12599 (N_12599,N_8070,N_8196);
nand U12600 (N_12600,N_6804,N_5640);
xnor U12601 (N_12601,N_6871,N_8849);
or U12602 (N_12602,N_8075,N_7737);
or U12603 (N_12603,N_9875,N_6773);
nor U12604 (N_12604,N_7861,N_6977);
or U12605 (N_12605,N_8849,N_5230);
or U12606 (N_12606,N_5653,N_5445);
or U12607 (N_12607,N_6811,N_8647);
xor U12608 (N_12608,N_7986,N_7310);
or U12609 (N_12609,N_6418,N_7159);
nand U12610 (N_12610,N_9391,N_6203);
nor U12611 (N_12611,N_5538,N_7217);
or U12612 (N_12612,N_9824,N_8460);
nand U12613 (N_12613,N_9580,N_6602);
nor U12614 (N_12614,N_9146,N_7048);
nor U12615 (N_12615,N_7789,N_7577);
or U12616 (N_12616,N_8356,N_7930);
or U12617 (N_12617,N_9164,N_7338);
xor U12618 (N_12618,N_7643,N_9878);
or U12619 (N_12619,N_7690,N_8632);
or U12620 (N_12620,N_7237,N_8242);
nor U12621 (N_12621,N_7440,N_6301);
xor U12622 (N_12622,N_7558,N_6488);
xnor U12623 (N_12623,N_8972,N_9609);
xnor U12624 (N_12624,N_5386,N_6906);
or U12625 (N_12625,N_7645,N_6125);
or U12626 (N_12626,N_9451,N_6552);
and U12627 (N_12627,N_5286,N_5848);
and U12628 (N_12628,N_9466,N_7279);
xnor U12629 (N_12629,N_7729,N_5516);
and U12630 (N_12630,N_9690,N_5758);
nor U12631 (N_12631,N_7039,N_8877);
xnor U12632 (N_12632,N_5178,N_9923);
nand U12633 (N_12633,N_7127,N_8278);
xor U12634 (N_12634,N_8616,N_7908);
xnor U12635 (N_12635,N_5588,N_9108);
and U12636 (N_12636,N_9484,N_9732);
and U12637 (N_12637,N_9892,N_5617);
nor U12638 (N_12638,N_5392,N_8761);
or U12639 (N_12639,N_5139,N_6324);
nand U12640 (N_12640,N_7254,N_6954);
nand U12641 (N_12641,N_7718,N_5665);
and U12642 (N_12642,N_7804,N_8249);
xor U12643 (N_12643,N_9514,N_8659);
or U12644 (N_12644,N_5455,N_5453);
nor U12645 (N_12645,N_6596,N_8071);
nand U12646 (N_12646,N_6228,N_6256);
nor U12647 (N_12647,N_5835,N_8041);
nand U12648 (N_12648,N_7682,N_7047);
and U12649 (N_12649,N_9243,N_6161);
nor U12650 (N_12650,N_7255,N_5589);
and U12651 (N_12651,N_6420,N_9929);
and U12652 (N_12652,N_8455,N_5413);
nand U12653 (N_12653,N_6706,N_6682);
xnor U12654 (N_12654,N_6219,N_5125);
and U12655 (N_12655,N_6978,N_8841);
xnor U12656 (N_12656,N_6817,N_6277);
nor U12657 (N_12657,N_9854,N_5905);
and U12658 (N_12658,N_6294,N_7513);
xnor U12659 (N_12659,N_6283,N_8938);
or U12660 (N_12660,N_5301,N_5831);
or U12661 (N_12661,N_5732,N_9445);
nor U12662 (N_12662,N_6491,N_5912);
or U12663 (N_12663,N_9307,N_5282);
or U12664 (N_12664,N_9836,N_6936);
nand U12665 (N_12665,N_5110,N_7974);
or U12666 (N_12666,N_6044,N_6108);
nor U12667 (N_12667,N_6891,N_6128);
nand U12668 (N_12668,N_9020,N_8645);
xnor U12669 (N_12669,N_8508,N_6878);
nor U12670 (N_12670,N_6812,N_6064);
xnor U12671 (N_12671,N_7010,N_6581);
xor U12672 (N_12672,N_5410,N_5645);
nand U12673 (N_12673,N_6677,N_8728);
nand U12674 (N_12674,N_5044,N_7550);
and U12675 (N_12675,N_5286,N_9028);
nor U12676 (N_12676,N_8040,N_7568);
and U12677 (N_12677,N_5350,N_8465);
and U12678 (N_12678,N_5096,N_5546);
xor U12679 (N_12679,N_9595,N_9167);
and U12680 (N_12680,N_6929,N_6740);
xnor U12681 (N_12681,N_6429,N_5728);
nand U12682 (N_12682,N_8714,N_7214);
nand U12683 (N_12683,N_9489,N_9193);
and U12684 (N_12684,N_7746,N_5810);
nor U12685 (N_12685,N_5335,N_6248);
nand U12686 (N_12686,N_6206,N_7021);
nand U12687 (N_12687,N_9463,N_9842);
and U12688 (N_12688,N_9327,N_9902);
nor U12689 (N_12689,N_9446,N_6709);
nor U12690 (N_12690,N_8791,N_6202);
nand U12691 (N_12691,N_6544,N_7066);
nor U12692 (N_12692,N_6905,N_9428);
and U12693 (N_12693,N_8787,N_5183);
or U12694 (N_12694,N_6831,N_7903);
or U12695 (N_12695,N_6733,N_7820);
nor U12696 (N_12696,N_5804,N_5293);
and U12697 (N_12697,N_6257,N_8978);
xor U12698 (N_12698,N_8672,N_5222);
nand U12699 (N_12699,N_7344,N_5365);
nand U12700 (N_12700,N_7793,N_6280);
xnor U12701 (N_12701,N_9397,N_7462);
nand U12702 (N_12702,N_9627,N_9846);
and U12703 (N_12703,N_7798,N_8286);
nor U12704 (N_12704,N_9130,N_8416);
nor U12705 (N_12705,N_8847,N_8417);
xor U12706 (N_12706,N_9030,N_5355);
and U12707 (N_12707,N_5478,N_9036);
nor U12708 (N_12708,N_7954,N_7314);
or U12709 (N_12709,N_9295,N_6928);
nor U12710 (N_12710,N_8272,N_9450);
nor U12711 (N_12711,N_5504,N_7950);
or U12712 (N_12712,N_8582,N_7681);
nor U12713 (N_12713,N_7403,N_7677);
or U12714 (N_12714,N_5049,N_5245);
or U12715 (N_12715,N_9898,N_7553);
nor U12716 (N_12716,N_6352,N_6361);
or U12717 (N_12717,N_7601,N_7738);
nor U12718 (N_12718,N_8571,N_5189);
or U12719 (N_12719,N_9007,N_9232);
xor U12720 (N_12720,N_8599,N_8826);
and U12721 (N_12721,N_9955,N_9064);
nor U12722 (N_12722,N_5656,N_7681);
and U12723 (N_12723,N_8652,N_9936);
nand U12724 (N_12724,N_9579,N_8179);
and U12725 (N_12725,N_7465,N_5505);
nand U12726 (N_12726,N_6825,N_8985);
nand U12727 (N_12727,N_8482,N_5646);
nor U12728 (N_12728,N_5116,N_8738);
or U12729 (N_12729,N_5641,N_7640);
and U12730 (N_12730,N_7773,N_6306);
xor U12731 (N_12731,N_6737,N_8168);
and U12732 (N_12732,N_5184,N_9729);
and U12733 (N_12733,N_9735,N_7367);
and U12734 (N_12734,N_6353,N_5103);
nand U12735 (N_12735,N_7573,N_8582);
nor U12736 (N_12736,N_9925,N_5111);
or U12737 (N_12737,N_6388,N_8463);
xnor U12738 (N_12738,N_8614,N_6615);
xnor U12739 (N_12739,N_5044,N_7849);
nand U12740 (N_12740,N_8100,N_9884);
nor U12741 (N_12741,N_7096,N_8116);
xor U12742 (N_12742,N_6207,N_9320);
xor U12743 (N_12743,N_9511,N_8934);
nand U12744 (N_12744,N_5883,N_8155);
xnor U12745 (N_12745,N_6626,N_6220);
nand U12746 (N_12746,N_5210,N_7551);
and U12747 (N_12747,N_6339,N_9144);
nand U12748 (N_12748,N_5125,N_8224);
xor U12749 (N_12749,N_5785,N_9745);
nor U12750 (N_12750,N_6041,N_9433);
nor U12751 (N_12751,N_7983,N_6507);
nand U12752 (N_12752,N_5216,N_9954);
or U12753 (N_12753,N_5029,N_8615);
and U12754 (N_12754,N_8060,N_6628);
and U12755 (N_12755,N_6801,N_6282);
nor U12756 (N_12756,N_9392,N_7155);
nor U12757 (N_12757,N_5907,N_6950);
xor U12758 (N_12758,N_9050,N_6439);
or U12759 (N_12759,N_5795,N_5790);
nand U12760 (N_12760,N_5311,N_7332);
or U12761 (N_12761,N_8132,N_6902);
xor U12762 (N_12762,N_6475,N_6386);
or U12763 (N_12763,N_7883,N_7501);
nor U12764 (N_12764,N_7975,N_5451);
and U12765 (N_12765,N_7867,N_8566);
xnor U12766 (N_12766,N_6581,N_9265);
or U12767 (N_12767,N_7134,N_7040);
or U12768 (N_12768,N_8522,N_7983);
xnor U12769 (N_12769,N_6303,N_7398);
and U12770 (N_12770,N_8234,N_6244);
xor U12771 (N_12771,N_6137,N_9511);
nor U12772 (N_12772,N_6998,N_5788);
nand U12773 (N_12773,N_5723,N_8940);
or U12774 (N_12774,N_8765,N_9994);
nand U12775 (N_12775,N_6751,N_9764);
and U12776 (N_12776,N_8703,N_7197);
or U12777 (N_12777,N_7121,N_5613);
nand U12778 (N_12778,N_7447,N_7653);
and U12779 (N_12779,N_8406,N_7449);
nand U12780 (N_12780,N_8519,N_9245);
nor U12781 (N_12781,N_6567,N_9891);
and U12782 (N_12782,N_9836,N_8727);
nand U12783 (N_12783,N_9906,N_8642);
or U12784 (N_12784,N_5909,N_9145);
or U12785 (N_12785,N_6954,N_5314);
nor U12786 (N_12786,N_6726,N_8229);
or U12787 (N_12787,N_7869,N_7042);
xor U12788 (N_12788,N_7058,N_5826);
nor U12789 (N_12789,N_6944,N_7690);
xor U12790 (N_12790,N_8947,N_8834);
or U12791 (N_12791,N_7473,N_6083);
and U12792 (N_12792,N_5533,N_7590);
or U12793 (N_12793,N_7556,N_8970);
xor U12794 (N_12794,N_5623,N_9880);
and U12795 (N_12795,N_6814,N_7793);
or U12796 (N_12796,N_6208,N_7389);
nor U12797 (N_12797,N_5371,N_7243);
or U12798 (N_12798,N_5350,N_7267);
xnor U12799 (N_12799,N_5626,N_8032);
and U12800 (N_12800,N_8207,N_6467);
nand U12801 (N_12801,N_5156,N_6167);
nor U12802 (N_12802,N_8027,N_5774);
nand U12803 (N_12803,N_7239,N_6460);
nand U12804 (N_12804,N_8366,N_7939);
or U12805 (N_12805,N_6180,N_5462);
nor U12806 (N_12806,N_9590,N_6158);
or U12807 (N_12807,N_7506,N_5362);
and U12808 (N_12808,N_7003,N_9728);
and U12809 (N_12809,N_9156,N_9953);
xnor U12810 (N_12810,N_8988,N_6946);
and U12811 (N_12811,N_5317,N_5648);
nand U12812 (N_12812,N_8169,N_8741);
nand U12813 (N_12813,N_5388,N_7279);
xor U12814 (N_12814,N_6242,N_9903);
and U12815 (N_12815,N_5555,N_6471);
nand U12816 (N_12816,N_9363,N_7241);
nand U12817 (N_12817,N_6593,N_7617);
or U12818 (N_12818,N_6298,N_8578);
nor U12819 (N_12819,N_5627,N_5769);
xnor U12820 (N_12820,N_8450,N_9667);
nand U12821 (N_12821,N_5875,N_5558);
or U12822 (N_12822,N_7279,N_6240);
nor U12823 (N_12823,N_9270,N_9746);
and U12824 (N_12824,N_8878,N_9565);
xnor U12825 (N_12825,N_9712,N_8523);
and U12826 (N_12826,N_8630,N_8364);
nor U12827 (N_12827,N_8979,N_6735);
or U12828 (N_12828,N_8857,N_9143);
nor U12829 (N_12829,N_9570,N_7812);
or U12830 (N_12830,N_8675,N_7113);
and U12831 (N_12831,N_9906,N_5049);
xnor U12832 (N_12832,N_8314,N_9146);
xor U12833 (N_12833,N_6462,N_5146);
or U12834 (N_12834,N_8709,N_5153);
or U12835 (N_12835,N_5126,N_9590);
or U12836 (N_12836,N_6802,N_7390);
or U12837 (N_12837,N_6690,N_9070);
or U12838 (N_12838,N_6596,N_5654);
xnor U12839 (N_12839,N_7932,N_9299);
nand U12840 (N_12840,N_5791,N_6387);
and U12841 (N_12841,N_7858,N_6716);
nor U12842 (N_12842,N_5785,N_7614);
nand U12843 (N_12843,N_7710,N_5145);
or U12844 (N_12844,N_6974,N_8444);
nand U12845 (N_12845,N_8289,N_9977);
nand U12846 (N_12846,N_7203,N_7121);
nand U12847 (N_12847,N_8551,N_7704);
and U12848 (N_12848,N_7842,N_5005);
nand U12849 (N_12849,N_6008,N_9442);
nor U12850 (N_12850,N_9384,N_5110);
nand U12851 (N_12851,N_8050,N_6926);
nor U12852 (N_12852,N_6374,N_7293);
nor U12853 (N_12853,N_7850,N_8534);
or U12854 (N_12854,N_7868,N_8360);
nand U12855 (N_12855,N_5699,N_5575);
and U12856 (N_12856,N_8387,N_9879);
or U12857 (N_12857,N_7398,N_6322);
and U12858 (N_12858,N_7609,N_6558);
nor U12859 (N_12859,N_5249,N_7942);
or U12860 (N_12860,N_6874,N_6742);
xor U12861 (N_12861,N_8105,N_9174);
and U12862 (N_12862,N_7585,N_9048);
nor U12863 (N_12863,N_7298,N_6897);
and U12864 (N_12864,N_8073,N_9432);
nor U12865 (N_12865,N_6094,N_9326);
nor U12866 (N_12866,N_5296,N_7012);
and U12867 (N_12867,N_6446,N_8342);
and U12868 (N_12868,N_5162,N_7222);
or U12869 (N_12869,N_9127,N_8611);
xnor U12870 (N_12870,N_6359,N_7749);
nor U12871 (N_12871,N_5273,N_7944);
nor U12872 (N_12872,N_7420,N_5017);
nor U12873 (N_12873,N_8321,N_6066);
and U12874 (N_12874,N_8299,N_8549);
xnor U12875 (N_12875,N_6626,N_6753);
nor U12876 (N_12876,N_9463,N_5461);
nand U12877 (N_12877,N_9366,N_9158);
nand U12878 (N_12878,N_7406,N_6383);
and U12879 (N_12879,N_6291,N_5252);
nand U12880 (N_12880,N_8371,N_9800);
or U12881 (N_12881,N_7687,N_7164);
nor U12882 (N_12882,N_7455,N_9013);
and U12883 (N_12883,N_5131,N_5909);
or U12884 (N_12884,N_7857,N_8023);
nand U12885 (N_12885,N_6339,N_9941);
nor U12886 (N_12886,N_6497,N_8663);
or U12887 (N_12887,N_9313,N_8193);
nor U12888 (N_12888,N_9882,N_8853);
xnor U12889 (N_12889,N_7918,N_6064);
and U12890 (N_12890,N_7588,N_7468);
and U12891 (N_12891,N_6144,N_5798);
or U12892 (N_12892,N_5529,N_9709);
xnor U12893 (N_12893,N_6699,N_8972);
nand U12894 (N_12894,N_5579,N_7352);
and U12895 (N_12895,N_9148,N_7521);
xor U12896 (N_12896,N_8759,N_7882);
and U12897 (N_12897,N_7261,N_6604);
and U12898 (N_12898,N_7405,N_9408);
xor U12899 (N_12899,N_6584,N_7835);
nor U12900 (N_12900,N_8943,N_7262);
xor U12901 (N_12901,N_9633,N_8124);
nor U12902 (N_12902,N_7212,N_8643);
or U12903 (N_12903,N_5894,N_5119);
xnor U12904 (N_12904,N_9963,N_9691);
or U12905 (N_12905,N_6679,N_6312);
or U12906 (N_12906,N_8877,N_5139);
nand U12907 (N_12907,N_6241,N_5185);
and U12908 (N_12908,N_9011,N_6193);
xor U12909 (N_12909,N_9242,N_6045);
xnor U12910 (N_12910,N_7114,N_7792);
nand U12911 (N_12911,N_7419,N_9409);
and U12912 (N_12912,N_8497,N_6826);
nand U12913 (N_12913,N_8080,N_5759);
nand U12914 (N_12914,N_9521,N_6434);
nor U12915 (N_12915,N_6100,N_6505);
nand U12916 (N_12916,N_5937,N_8342);
nor U12917 (N_12917,N_9239,N_9482);
and U12918 (N_12918,N_7609,N_6191);
nor U12919 (N_12919,N_7811,N_6145);
or U12920 (N_12920,N_9041,N_6023);
xor U12921 (N_12921,N_8762,N_8297);
nand U12922 (N_12922,N_6875,N_8166);
nor U12923 (N_12923,N_7553,N_9336);
xnor U12924 (N_12924,N_9227,N_8058);
or U12925 (N_12925,N_9524,N_7065);
nor U12926 (N_12926,N_8605,N_7497);
xor U12927 (N_12927,N_7636,N_5045);
nand U12928 (N_12928,N_5120,N_7980);
xnor U12929 (N_12929,N_6405,N_9246);
xnor U12930 (N_12930,N_9849,N_5984);
nor U12931 (N_12931,N_5667,N_5374);
or U12932 (N_12932,N_9528,N_7481);
and U12933 (N_12933,N_9598,N_7893);
and U12934 (N_12934,N_9789,N_9180);
and U12935 (N_12935,N_7458,N_5654);
and U12936 (N_12936,N_5606,N_8029);
nor U12937 (N_12937,N_8274,N_9299);
xor U12938 (N_12938,N_5589,N_8231);
or U12939 (N_12939,N_8946,N_9110);
nor U12940 (N_12940,N_6419,N_9528);
xor U12941 (N_12941,N_5242,N_7584);
and U12942 (N_12942,N_8557,N_8224);
nor U12943 (N_12943,N_6152,N_5469);
xnor U12944 (N_12944,N_9292,N_7734);
or U12945 (N_12945,N_7970,N_5679);
and U12946 (N_12946,N_7663,N_8520);
xnor U12947 (N_12947,N_8889,N_8577);
xnor U12948 (N_12948,N_5048,N_6300);
nor U12949 (N_12949,N_7878,N_8410);
nand U12950 (N_12950,N_5690,N_5970);
or U12951 (N_12951,N_6558,N_7323);
nand U12952 (N_12952,N_8491,N_7372);
nor U12953 (N_12953,N_8506,N_5081);
xor U12954 (N_12954,N_7773,N_8591);
or U12955 (N_12955,N_6872,N_9525);
and U12956 (N_12956,N_5300,N_8122);
or U12957 (N_12957,N_8017,N_9606);
nor U12958 (N_12958,N_7658,N_8568);
xor U12959 (N_12959,N_7486,N_7174);
and U12960 (N_12960,N_6429,N_9342);
nand U12961 (N_12961,N_6239,N_9426);
nor U12962 (N_12962,N_8084,N_6131);
or U12963 (N_12963,N_8554,N_9830);
or U12964 (N_12964,N_7198,N_7835);
or U12965 (N_12965,N_8821,N_6075);
or U12966 (N_12966,N_7762,N_7689);
or U12967 (N_12967,N_8795,N_7002);
nor U12968 (N_12968,N_7664,N_8536);
nand U12969 (N_12969,N_8858,N_8906);
and U12970 (N_12970,N_6019,N_8807);
and U12971 (N_12971,N_6808,N_6206);
or U12972 (N_12972,N_9184,N_7244);
nor U12973 (N_12973,N_8849,N_5904);
or U12974 (N_12974,N_8218,N_7026);
and U12975 (N_12975,N_5213,N_5977);
and U12976 (N_12976,N_8105,N_7444);
nand U12977 (N_12977,N_7454,N_8735);
nor U12978 (N_12978,N_8337,N_9957);
or U12979 (N_12979,N_6326,N_7964);
xnor U12980 (N_12980,N_7776,N_9553);
and U12981 (N_12981,N_8700,N_9551);
nand U12982 (N_12982,N_7893,N_8893);
nor U12983 (N_12983,N_7794,N_9202);
nor U12984 (N_12984,N_9371,N_8449);
xnor U12985 (N_12985,N_5178,N_8432);
or U12986 (N_12986,N_9466,N_8594);
xnor U12987 (N_12987,N_6827,N_8293);
or U12988 (N_12988,N_6296,N_7113);
nor U12989 (N_12989,N_7577,N_8101);
xor U12990 (N_12990,N_6368,N_5936);
nor U12991 (N_12991,N_7310,N_6842);
xnor U12992 (N_12992,N_5604,N_6237);
or U12993 (N_12993,N_8788,N_6068);
nand U12994 (N_12994,N_9936,N_6641);
nor U12995 (N_12995,N_6094,N_5556);
nand U12996 (N_12996,N_8254,N_9805);
or U12997 (N_12997,N_6113,N_6450);
nand U12998 (N_12998,N_7960,N_9715);
xnor U12999 (N_12999,N_7184,N_6592);
nand U13000 (N_13000,N_8553,N_8149);
or U13001 (N_13001,N_7223,N_5437);
xnor U13002 (N_13002,N_6950,N_9743);
nand U13003 (N_13003,N_8272,N_5039);
xor U13004 (N_13004,N_6328,N_8782);
xnor U13005 (N_13005,N_8000,N_5263);
xor U13006 (N_13006,N_9022,N_6356);
nand U13007 (N_13007,N_9437,N_7676);
or U13008 (N_13008,N_5720,N_8286);
xnor U13009 (N_13009,N_8456,N_9640);
and U13010 (N_13010,N_7744,N_6158);
nor U13011 (N_13011,N_7143,N_9136);
nor U13012 (N_13012,N_9153,N_5632);
xor U13013 (N_13013,N_6979,N_5668);
nand U13014 (N_13014,N_7026,N_5737);
nor U13015 (N_13015,N_5530,N_7045);
nand U13016 (N_13016,N_5234,N_6605);
xnor U13017 (N_13017,N_7015,N_7333);
and U13018 (N_13018,N_8241,N_5373);
nor U13019 (N_13019,N_6894,N_9753);
xnor U13020 (N_13020,N_9435,N_6453);
nor U13021 (N_13021,N_5246,N_5826);
nand U13022 (N_13022,N_8216,N_5153);
nor U13023 (N_13023,N_5885,N_9773);
or U13024 (N_13024,N_7893,N_5092);
or U13025 (N_13025,N_7094,N_7578);
and U13026 (N_13026,N_7238,N_7275);
nor U13027 (N_13027,N_6100,N_5968);
and U13028 (N_13028,N_9265,N_7056);
and U13029 (N_13029,N_5239,N_5102);
xnor U13030 (N_13030,N_7453,N_9473);
and U13031 (N_13031,N_6365,N_7491);
xor U13032 (N_13032,N_5368,N_7015);
and U13033 (N_13033,N_7607,N_8739);
nand U13034 (N_13034,N_8203,N_7311);
and U13035 (N_13035,N_6982,N_8792);
and U13036 (N_13036,N_5537,N_8464);
and U13037 (N_13037,N_8596,N_9751);
nor U13038 (N_13038,N_6269,N_9821);
and U13039 (N_13039,N_9086,N_9712);
nand U13040 (N_13040,N_8799,N_9996);
xor U13041 (N_13041,N_7008,N_5206);
xor U13042 (N_13042,N_5917,N_9538);
nor U13043 (N_13043,N_6500,N_9874);
nor U13044 (N_13044,N_8675,N_8929);
and U13045 (N_13045,N_7337,N_5296);
nor U13046 (N_13046,N_8747,N_9096);
or U13047 (N_13047,N_7262,N_7512);
xor U13048 (N_13048,N_7972,N_7567);
or U13049 (N_13049,N_6912,N_6220);
nand U13050 (N_13050,N_8107,N_5332);
nand U13051 (N_13051,N_5476,N_7413);
xnor U13052 (N_13052,N_6582,N_5590);
nand U13053 (N_13053,N_7746,N_5430);
nor U13054 (N_13054,N_9607,N_5878);
or U13055 (N_13055,N_7836,N_5392);
or U13056 (N_13056,N_7499,N_7666);
nand U13057 (N_13057,N_5502,N_8221);
or U13058 (N_13058,N_5808,N_9991);
and U13059 (N_13059,N_6902,N_7419);
xnor U13060 (N_13060,N_5848,N_6460);
or U13061 (N_13061,N_6745,N_5482);
nor U13062 (N_13062,N_6144,N_6848);
xnor U13063 (N_13063,N_7553,N_7291);
and U13064 (N_13064,N_6848,N_8332);
xnor U13065 (N_13065,N_5897,N_8667);
xor U13066 (N_13066,N_9977,N_7833);
nand U13067 (N_13067,N_8808,N_6253);
nor U13068 (N_13068,N_6646,N_8845);
nor U13069 (N_13069,N_7626,N_8728);
nor U13070 (N_13070,N_7574,N_7059);
and U13071 (N_13071,N_7519,N_7662);
nor U13072 (N_13072,N_8897,N_9908);
nor U13073 (N_13073,N_8520,N_5570);
xnor U13074 (N_13074,N_6727,N_7475);
or U13075 (N_13075,N_8316,N_5164);
and U13076 (N_13076,N_5587,N_6819);
and U13077 (N_13077,N_7096,N_9688);
nor U13078 (N_13078,N_8125,N_9725);
or U13079 (N_13079,N_6941,N_9257);
and U13080 (N_13080,N_8993,N_8138);
nand U13081 (N_13081,N_7344,N_5356);
nor U13082 (N_13082,N_8795,N_9573);
nand U13083 (N_13083,N_5769,N_9565);
nand U13084 (N_13084,N_9572,N_7695);
or U13085 (N_13085,N_5595,N_8587);
xor U13086 (N_13086,N_9025,N_5908);
xor U13087 (N_13087,N_8139,N_8524);
or U13088 (N_13088,N_8683,N_9233);
nor U13089 (N_13089,N_5163,N_6897);
nor U13090 (N_13090,N_6593,N_9301);
xnor U13091 (N_13091,N_9432,N_5236);
xnor U13092 (N_13092,N_8770,N_5568);
nand U13093 (N_13093,N_7604,N_6169);
and U13094 (N_13094,N_6402,N_9115);
or U13095 (N_13095,N_9832,N_6039);
and U13096 (N_13096,N_7100,N_7831);
and U13097 (N_13097,N_5111,N_6397);
and U13098 (N_13098,N_6513,N_6926);
and U13099 (N_13099,N_9244,N_9974);
nor U13100 (N_13100,N_5767,N_9512);
xnor U13101 (N_13101,N_7058,N_6277);
xor U13102 (N_13102,N_9736,N_9284);
and U13103 (N_13103,N_7807,N_8179);
nor U13104 (N_13104,N_9734,N_6500);
nor U13105 (N_13105,N_9840,N_6290);
nor U13106 (N_13106,N_6477,N_9340);
xnor U13107 (N_13107,N_9629,N_5658);
nand U13108 (N_13108,N_6617,N_6052);
and U13109 (N_13109,N_5801,N_7408);
nor U13110 (N_13110,N_6799,N_9404);
xnor U13111 (N_13111,N_8931,N_9300);
and U13112 (N_13112,N_8362,N_7884);
and U13113 (N_13113,N_7292,N_9595);
and U13114 (N_13114,N_8428,N_8946);
nand U13115 (N_13115,N_7975,N_8073);
nor U13116 (N_13116,N_6083,N_6311);
xnor U13117 (N_13117,N_7420,N_9419);
xor U13118 (N_13118,N_6064,N_9987);
xor U13119 (N_13119,N_5484,N_9523);
or U13120 (N_13120,N_8377,N_7178);
and U13121 (N_13121,N_5684,N_8589);
or U13122 (N_13122,N_6410,N_6994);
xnor U13123 (N_13123,N_6448,N_9904);
nand U13124 (N_13124,N_6418,N_6156);
and U13125 (N_13125,N_9853,N_8943);
or U13126 (N_13126,N_6870,N_8202);
nor U13127 (N_13127,N_9551,N_5785);
or U13128 (N_13128,N_8847,N_9799);
xnor U13129 (N_13129,N_5979,N_7036);
and U13130 (N_13130,N_6292,N_5824);
nor U13131 (N_13131,N_9165,N_6520);
or U13132 (N_13132,N_6777,N_5622);
and U13133 (N_13133,N_9628,N_5795);
xor U13134 (N_13134,N_6636,N_5141);
xor U13135 (N_13135,N_5361,N_7869);
xor U13136 (N_13136,N_7602,N_6625);
nor U13137 (N_13137,N_9560,N_7424);
and U13138 (N_13138,N_7975,N_5979);
nor U13139 (N_13139,N_7799,N_8756);
xnor U13140 (N_13140,N_7553,N_8266);
nor U13141 (N_13141,N_7589,N_7205);
nand U13142 (N_13142,N_9506,N_6530);
nor U13143 (N_13143,N_8794,N_6033);
nand U13144 (N_13144,N_7674,N_8506);
or U13145 (N_13145,N_9333,N_8097);
and U13146 (N_13146,N_7095,N_5861);
nand U13147 (N_13147,N_7863,N_9065);
nand U13148 (N_13148,N_6065,N_7407);
and U13149 (N_13149,N_9074,N_7870);
and U13150 (N_13150,N_6027,N_7639);
nand U13151 (N_13151,N_5888,N_7107);
nor U13152 (N_13152,N_7538,N_6162);
or U13153 (N_13153,N_9601,N_8901);
or U13154 (N_13154,N_9855,N_5468);
nand U13155 (N_13155,N_6251,N_7371);
nand U13156 (N_13156,N_7722,N_9736);
nand U13157 (N_13157,N_5844,N_9664);
or U13158 (N_13158,N_8992,N_8414);
xor U13159 (N_13159,N_5784,N_8207);
xnor U13160 (N_13160,N_6267,N_8971);
nand U13161 (N_13161,N_9391,N_7274);
and U13162 (N_13162,N_7967,N_8292);
nor U13163 (N_13163,N_5293,N_5236);
and U13164 (N_13164,N_8224,N_5623);
or U13165 (N_13165,N_8977,N_7204);
xnor U13166 (N_13166,N_8590,N_6859);
or U13167 (N_13167,N_9642,N_8671);
and U13168 (N_13168,N_7793,N_9047);
or U13169 (N_13169,N_6696,N_9077);
xor U13170 (N_13170,N_8077,N_6418);
nor U13171 (N_13171,N_6933,N_5094);
xnor U13172 (N_13172,N_5829,N_9582);
nor U13173 (N_13173,N_8297,N_7604);
nor U13174 (N_13174,N_7877,N_8070);
nand U13175 (N_13175,N_7066,N_8443);
and U13176 (N_13176,N_5327,N_5654);
nor U13177 (N_13177,N_8655,N_7350);
xnor U13178 (N_13178,N_9179,N_5967);
nor U13179 (N_13179,N_6968,N_8353);
and U13180 (N_13180,N_9598,N_7618);
nor U13181 (N_13181,N_8155,N_5887);
xor U13182 (N_13182,N_7615,N_6423);
and U13183 (N_13183,N_9191,N_9969);
nor U13184 (N_13184,N_6451,N_7668);
nor U13185 (N_13185,N_8031,N_8026);
and U13186 (N_13186,N_7030,N_8943);
nor U13187 (N_13187,N_5566,N_6191);
and U13188 (N_13188,N_9390,N_8605);
xnor U13189 (N_13189,N_8355,N_8966);
or U13190 (N_13190,N_6543,N_5154);
and U13191 (N_13191,N_5612,N_5864);
and U13192 (N_13192,N_5132,N_6520);
and U13193 (N_13193,N_5273,N_9559);
nand U13194 (N_13194,N_7636,N_9888);
or U13195 (N_13195,N_5444,N_6754);
and U13196 (N_13196,N_9430,N_8791);
xnor U13197 (N_13197,N_6095,N_7355);
nand U13198 (N_13198,N_9106,N_6826);
nand U13199 (N_13199,N_9979,N_5450);
nand U13200 (N_13200,N_8027,N_9261);
nor U13201 (N_13201,N_9199,N_8890);
nor U13202 (N_13202,N_7502,N_5225);
xor U13203 (N_13203,N_5130,N_7511);
nand U13204 (N_13204,N_8888,N_6877);
nor U13205 (N_13205,N_7353,N_5992);
or U13206 (N_13206,N_8638,N_8984);
xnor U13207 (N_13207,N_8198,N_5053);
or U13208 (N_13208,N_5382,N_7690);
or U13209 (N_13209,N_9146,N_9429);
xor U13210 (N_13210,N_5563,N_9978);
nor U13211 (N_13211,N_7401,N_6466);
or U13212 (N_13212,N_8862,N_7139);
or U13213 (N_13213,N_7808,N_7734);
nor U13214 (N_13214,N_9883,N_8358);
or U13215 (N_13215,N_6408,N_8260);
and U13216 (N_13216,N_8028,N_6493);
nor U13217 (N_13217,N_7898,N_8039);
and U13218 (N_13218,N_6537,N_9498);
or U13219 (N_13219,N_5693,N_8698);
nand U13220 (N_13220,N_6579,N_6199);
nand U13221 (N_13221,N_5206,N_6874);
and U13222 (N_13222,N_7628,N_9335);
and U13223 (N_13223,N_7044,N_9584);
nand U13224 (N_13224,N_7716,N_9081);
or U13225 (N_13225,N_7914,N_9157);
and U13226 (N_13226,N_8945,N_7819);
or U13227 (N_13227,N_9634,N_6826);
and U13228 (N_13228,N_6431,N_6638);
nor U13229 (N_13229,N_7194,N_5673);
xor U13230 (N_13230,N_9456,N_8841);
nand U13231 (N_13231,N_7228,N_5855);
xor U13232 (N_13232,N_9065,N_7144);
nor U13233 (N_13233,N_9126,N_9816);
nor U13234 (N_13234,N_6427,N_9871);
nor U13235 (N_13235,N_5068,N_8806);
or U13236 (N_13236,N_6942,N_9642);
nand U13237 (N_13237,N_9750,N_5754);
nor U13238 (N_13238,N_6841,N_8638);
xnor U13239 (N_13239,N_6974,N_8212);
nand U13240 (N_13240,N_8609,N_9134);
xnor U13241 (N_13241,N_8836,N_7084);
xor U13242 (N_13242,N_5570,N_5739);
nand U13243 (N_13243,N_7803,N_9902);
xnor U13244 (N_13244,N_7264,N_5450);
or U13245 (N_13245,N_7832,N_9502);
or U13246 (N_13246,N_6709,N_8903);
and U13247 (N_13247,N_5111,N_6497);
nor U13248 (N_13248,N_7974,N_7446);
or U13249 (N_13249,N_8029,N_7750);
xnor U13250 (N_13250,N_8169,N_5901);
nand U13251 (N_13251,N_9741,N_6297);
xnor U13252 (N_13252,N_5857,N_9321);
nor U13253 (N_13253,N_7013,N_5946);
nor U13254 (N_13254,N_7379,N_5459);
nand U13255 (N_13255,N_9930,N_8659);
or U13256 (N_13256,N_9183,N_9209);
nand U13257 (N_13257,N_5745,N_7153);
and U13258 (N_13258,N_5348,N_9560);
nand U13259 (N_13259,N_7988,N_8461);
xor U13260 (N_13260,N_6092,N_5411);
and U13261 (N_13261,N_7609,N_5125);
nor U13262 (N_13262,N_9490,N_8858);
and U13263 (N_13263,N_7004,N_9468);
nand U13264 (N_13264,N_7268,N_9004);
xnor U13265 (N_13265,N_5529,N_7967);
or U13266 (N_13266,N_5058,N_7540);
nor U13267 (N_13267,N_6079,N_9180);
or U13268 (N_13268,N_6137,N_8041);
xor U13269 (N_13269,N_5258,N_6714);
or U13270 (N_13270,N_6197,N_7958);
and U13271 (N_13271,N_9531,N_5882);
or U13272 (N_13272,N_6786,N_5517);
nor U13273 (N_13273,N_8109,N_6423);
nor U13274 (N_13274,N_9396,N_6057);
or U13275 (N_13275,N_8358,N_8133);
or U13276 (N_13276,N_5687,N_9673);
or U13277 (N_13277,N_6763,N_6483);
nand U13278 (N_13278,N_5818,N_9631);
or U13279 (N_13279,N_5382,N_7388);
nor U13280 (N_13280,N_7619,N_6299);
xnor U13281 (N_13281,N_9640,N_7561);
and U13282 (N_13282,N_9249,N_8805);
or U13283 (N_13283,N_8189,N_6300);
nand U13284 (N_13284,N_9346,N_6051);
and U13285 (N_13285,N_8484,N_6934);
nor U13286 (N_13286,N_8333,N_9062);
and U13287 (N_13287,N_6060,N_6858);
xnor U13288 (N_13288,N_9127,N_7264);
nor U13289 (N_13289,N_5673,N_6456);
and U13290 (N_13290,N_6866,N_8054);
xor U13291 (N_13291,N_9774,N_7386);
or U13292 (N_13292,N_6182,N_5276);
xnor U13293 (N_13293,N_7703,N_6998);
or U13294 (N_13294,N_8774,N_7703);
nand U13295 (N_13295,N_5236,N_6966);
xor U13296 (N_13296,N_8181,N_8743);
or U13297 (N_13297,N_6563,N_8267);
or U13298 (N_13298,N_5060,N_6817);
xnor U13299 (N_13299,N_6600,N_9665);
nor U13300 (N_13300,N_7734,N_8819);
xor U13301 (N_13301,N_6809,N_8329);
nand U13302 (N_13302,N_6613,N_8717);
or U13303 (N_13303,N_5619,N_7727);
nand U13304 (N_13304,N_9178,N_8001);
or U13305 (N_13305,N_5624,N_5488);
xnor U13306 (N_13306,N_9092,N_6774);
nand U13307 (N_13307,N_8222,N_6445);
nand U13308 (N_13308,N_6859,N_6730);
nand U13309 (N_13309,N_7088,N_7189);
nand U13310 (N_13310,N_7548,N_9641);
and U13311 (N_13311,N_8436,N_6795);
and U13312 (N_13312,N_7235,N_8593);
xor U13313 (N_13313,N_6063,N_6600);
or U13314 (N_13314,N_9141,N_8546);
or U13315 (N_13315,N_5518,N_9753);
nor U13316 (N_13316,N_6529,N_5911);
nand U13317 (N_13317,N_8856,N_6974);
nand U13318 (N_13318,N_8613,N_7255);
nand U13319 (N_13319,N_8884,N_9067);
xnor U13320 (N_13320,N_5846,N_7647);
or U13321 (N_13321,N_9486,N_8570);
nand U13322 (N_13322,N_6382,N_8054);
or U13323 (N_13323,N_9522,N_5531);
nor U13324 (N_13324,N_5730,N_7779);
nor U13325 (N_13325,N_9098,N_9882);
and U13326 (N_13326,N_8138,N_6853);
or U13327 (N_13327,N_6650,N_7456);
nand U13328 (N_13328,N_9587,N_5855);
nand U13329 (N_13329,N_9330,N_5357);
xnor U13330 (N_13330,N_9652,N_8423);
nand U13331 (N_13331,N_9626,N_7046);
nand U13332 (N_13332,N_6405,N_5248);
nor U13333 (N_13333,N_8278,N_7584);
nor U13334 (N_13334,N_6322,N_9531);
nand U13335 (N_13335,N_5518,N_7771);
or U13336 (N_13336,N_7711,N_6261);
and U13337 (N_13337,N_8540,N_5401);
or U13338 (N_13338,N_5587,N_5267);
nand U13339 (N_13339,N_9447,N_6584);
and U13340 (N_13340,N_6979,N_7685);
and U13341 (N_13341,N_7276,N_9657);
xnor U13342 (N_13342,N_8974,N_9798);
nor U13343 (N_13343,N_5102,N_7957);
xnor U13344 (N_13344,N_7421,N_9553);
or U13345 (N_13345,N_6454,N_5697);
nand U13346 (N_13346,N_7122,N_6750);
xnor U13347 (N_13347,N_5207,N_6156);
and U13348 (N_13348,N_6804,N_9151);
or U13349 (N_13349,N_5099,N_6191);
and U13350 (N_13350,N_9297,N_9071);
nand U13351 (N_13351,N_7230,N_6046);
or U13352 (N_13352,N_5809,N_7370);
nor U13353 (N_13353,N_5476,N_5250);
nand U13354 (N_13354,N_9466,N_7355);
xnor U13355 (N_13355,N_5281,N_7569);
and U13356 (N_13356,N_8818,N_6885);
nand U13357 (N_13357,N_6271,N_5895);
nor U13358 (N_13358,N_5616,N_6351);
nand U13359 (N_13359,N_6183,N_7027);
nand U13360 (N_13360,N_9991,N_7381);
and U13361 (N_13361,N_9772,N_5033);
nand U13362 (N_13362,N_7667,N_5883);
or U13363 (N_13363,N_7371,N_9177);
or U13364 (N_13364,N_6782,N_5830);
xnor U13365 (N_13365,N_6774,N_9887);
nand U13366 (N_13366,N_7525,N_7693);
or U13367 (N_13367,N_6256,N_8532);
xor U13368 (N_13368,N_6488,N_5488);
nor U13369 (N_13369,N_6928,N_9051);
or U13370 (N_13370,N_8866,N_5003);
or U13371 (N_13371,N_5212,N_5437);
and U13372 (N_13372,N_5723,N_5933);
nor U13373 (N_13373,N_8704,N_8778);
or U13374 (N_13374,N_7469,N_5409);
and U13375 (N_13375,N_9356,N_6410);
and U13376 (N_13376,N_7873,N_8576);
or U13377 (N_13377,N_6959,N_9452);
xnor U13378 (N_13378,N_9898,N_7521);
and U13379 (N_13379,N_8141,N_6089);
and U13380 (N_13380,N_8720,N_5007);
or U13381 (N_13381,N_6085,N_8418);
or U13382 (N_13382,N_5311,N_9628);
or U13383 (N_13383,N_5083,N_5160);
nand U13384 (N_13384,N_7977,N_7312);
or U13385 (N_13385,N_8453,N_6169);
and U13386 (N_13386,N_9532,N_6560);
xnor U13387 (N_13387,N_5470,N_7973);
and U13388 (N_13388,N_5734,N_6698);
and U13389 (N_13389,N_8775,N_6167);
xor U13390 (N_13390,N_5312,N_8976);
and U13391 (N_13391,N_9508,N_9245);
nor U13392 (N_13392,N_9493,N_9360);
xor U13393 (N_13393,N_5840,N_5166);
and U13394 (N_13394,N_5019,N_5128);
nand U13395 (N_13395,N_8093,N_5825);
nand U13396 (N_13396,N_7725,N_5310);
or U13397 (N_13397,N_8882,N_6624);
xnor U13398 (N_13398,N_9686,N_9372);
xnor U13399 (N_13399,N_8437,N_6052);
or U13400 (N_13400,N_7750,N_5177);
xor U13401 (N_13401,N_7002,N_7220);
nor U13402 (N_13402,N_7547,N_7973);
nor U13403 (N_13403,N_5507,N_7466);
or U13404 (N_13404,N_5535,N_6461);
xnor U13405 (N_13405,N_9226,N_8846);
or U13406 (N_13406,N_5549,N_9682);
and U13407 (N_13407,N_5721,N_9831);
nor U13408 (N_13408,N_7136,N_8011);
nand U13409 (N_13409,N_8739,N_9357);
or U13410 (N_13410,N_5182,N_9986);
and U13411 (N_13411,N_9180,N_9693);
nor U13412 (N_13412,N_7783,N_5850);
and U13413 (N_13413,N_9551,N_6976);
nor U13414 (N_13414,N_8895,N_5971);
nor U13415 (N_13415,N_5581,N_8855);
nand U13416 (N_13416,N_9619,N_8195);
xor U13417 (N_13417,N_9469,N_5416);
or U13418 (N_13418,N_9202,N_8456);
and U13419 (N_13419,N_9364,N_7007);
and U13420 (N_13420,N_8560,N_8046);
nor U13421 (N_13421,N_8558,N_5822);
nand U13422 (N_13422,N_9201,N_5642);
nand U13423 (N_13423,N_8118,N_9039);
and U13424 (N_13424,N_6441,N_9229);
and U13425 (N_13425,N_9972,N_8795);
or U13426 (N_13426,N_5741,N_5397);
or U13427 (N_13427,N_7468,N_6456);
and U13428 (N_13428,N_6940,N_9893);
xor U13429 (N_13429,N_7853,N_6134);
or U13430 (N_13430,N_9206,N_5941);
xor U13431 (N_13431,N_5049,N_5916);
xor U13432 (N_13432,N_5066,N_6603);
nand U13433 (N_13433,N_6770,N_8627);
xor U13434 (N_13434,N_6828,N_5836);
nand U13435 (N_13435,N_5184,N_5235);
nor U13436 (N_13436,N_8771,N_6165);
or U13437 (N_13437,N_5617,N_8016);
nand U13438 (N_13438,N_8164,N_8550);
and U13439 (N_13439,N_6735,N_7002);
or U13440 (N_13440,N_9535,N_6332);
nor U13441 (N_13441,N_8208,N_8399);
nand U13442 (N_13442,N_7081,N_7239);
nor U13443 (N_13443,N_8719,N_8355);
xnor U13444 (N_13444,N_6184,N_6476);
nor U13445 (N_13445,N_5384,N_5240);
or U13446 (N_13446,N_7017,N_5665);
and U13447 (N_13447,N_9115,N_7316);
xnor U13448 (N_13448,N_6378,N_8570);
nand U13449 (N_13449,N_7970,N_5592);
nor U13450 (N_13450,N_9974,N_8826);
or U13451 (N_13451,N_8916,N_5320);
nor U13452 (N_13452,N_6627,N_8449);
xor U13453 (N_13453,N_7196,N_7684);
or U13454 (N_13454,N_8372,N_7200);
xor U13455 (N_13455,N_6379,N_5211);
nor U13456 (N_13456,N_8094,N_9587);
xnor U13457 (N_13457,N_8703,N_6087);
xnor U13458 (N_13458,N_7376,N_6699);
nor U13459 (N_13459,N_6490,N_7743);
nor U13460 (N_13460,N_7815,N_9401);
or U13461 (N_13461,N_5713,N_6183);
nand U13462 (N_13462,N_5353,N_7665);
or U13463 (N_13463,N_6616,N_9587);
or U13464 (N_13464,N_9600,N_7355);
nor U13465 (N_13465,N_8596,N_7700);
and U13466 (N_13466,N_8215,N_8468);
nand U13467 (N_13467,N_5064,N_5839);
or U13468 (N_13468,N_8342,N_5545);
nand U13469 (N_13469,N_5369,N_7923);
and U13470 (N_13470,N_6701,N_7738);
nor U13471 (N_13471,N_8454,N_7582);
nand U13472 (N_13472,N_5668,N_5520);
or U13473 (N_13473,N_5060,N_5697);
xor U13474 (N_13474,N_9309,N_8878);
or U13475 (N_13475,N_9723,N_8759);
or U13476 (N_13476,N_7448,N_7560);
nand U13477 (N_13477,N_7098,N_9867);
or U13478 (N_13478,N_9649,N_5123);
or U13479 (N_13479,N_9096,N_6441);
and U13480 (N_13480,N_5899,N_6123);
nor U13481 (N_13481,N_9692,N_7768);
nor U13482 (N_13482,N_9313,N_8887);
and U13483 (N_13483,N_9412,N_5511);
xor U13484 (N_13484,N_6819,N_6864);
nor U13485 (N_13485,N_9903,N_8300);
nor U13486 (N_13486,N_5431,N_7547);
nand U13487 (N_13487,N_5158,N_8874);
nand U13488 (N_13488,N_7852,N_7940);
xor U13489 (N_13489,N_7395,N_8034);
or U13490 (N_13490,N_5238,N_9059);
or U13491 (N_13491,N_6985,N_9340);
or U13492 (N_13492,N_6012,N_9448);
and U13493 (N_13493,N_5983,N_7078);
nand U13494 (N_13494,N_7397,N_7459);
or U13495 (N_13495,N_6591,N_9282);
xnor U13496 (N_13496,N_9468,N_7508);
nand U13497 (N_13497,N_8410,N_8229);
xnor U13498 (N_13498,N_6709,N_8340);
xnor U13499 (N_13499,N_6986,N_6943);
and U13500 (N_13500,N_7733,N_7049);
xor U13501 (N_13501,N_5658,N_6037);
xor U13502 (N_13502,N_8336,N_6573);
nor U13503 (N_13503,N_7162,N_7645);
nor U13504 (N_13504,N_7999,N_8165);
xnor U13505 (N_13505,N_5982,N_6373);
and U13506 (N_13506,N_9561,N_6455);
and U13507 (N_13507,N_6708,N_8124);
and U13508 (N_13508,N_9370,N_9420);
nand U13509 (N_13509,N_6744,N_5731);
and U13510 (N_13510,N_8847,N_6468);
and U13511 (N_13511,N_7054,N_5202);
and U13512 (N_13512,N_9612,N_6193);
nor U13513 (N_13513,N_6476,N_8361);
nor U13514 (N_13514,N_7210,N_5509);
or U13515 (N_13515,N_7629,N_8063);
xor U13516 (N_13516,N_5528,N_7066);
xor U13517 (N_13517,N_9911,N_6648);
nor U13518 (N_13518,N_8223,N_6341);
nand U13519 (N_13519,N_7563,N_6664);
xor U13520 (N_13520,N_9007,N_9310);
nor U13521 (N_13521,N_9027,N_7773);
xnor U13522 (N_13522,N_8521,N_5742);
nand U13523 (N_13523,N_8954,N_5063);
xor U13524 (N_13524,N_7210,N_6486);
xnor U13525 (N_13525,N_6796,N_8099);
nand U13526 (N_13526,N_7378,N_7798);
nor U13527 (N_13527,N_5692,N_6899);
xnor U13528 (N_13528,N_7749,N_7400);
nand U13529 (N_13529,N_6139,N_5440);
nor U13530 (N_13530,N_7229,N_6242);
or U13531 (N_13531,N_7477,N_7659);
or U13532 (N_13532,N_7992,N_5693);
nand U13533 (N_13533,N_9209,N_5267);
xnor U13534 (N_13534,N_8774,N_8850);
nor U13535 (N_13535,N_9326,N_8859);
nand U13536 (N_13536,N_6919,N_6233);
nand U13537 (N_13537,N_7667,N_5299);
or U13538 (N_13538,N_8456,N_7211);
or U13539 (N_13539,N_5876,N_5698);
or U13540 (N_13540,N_9833,N_5340);
and U13541 (N_13541,N_9204,N_5501);
and U13542 (N_13542,N_7414,N_6619);
nor U13543 (N_13543,N_5266,N_6055);
xnor U13544 (N_13544,N_8529,N_5950);
xor U13545 (N_13545,N_9339,N_6390);
nand U13546 (N_13546,N_5795,N_5616);
nand U13547 (N_13547,N_8472,N_7037);
or U13548 (N_13548,N_7237,N_7092);
nor U13549 (N_13549,N_7707,N_8456);
and U13550 (N_13550,N_7489,N_9255);
xnor U13551 (N_13551,N_6733,N_6918);
or U13552 (N_13552,N_5922,N_5930);
or U13553 (N_13553,N_8711,N_9992);
xnor U13554 (N_13554,N_5868,N_8286);
nand U13555 (N_13555,N_6555,N_7899);
nor U13556 (N_13556,N_6120,N_9744);
and U13557 (N_13557,N_5210,N_5043);
and U13558 (N_13558,N_7706,N_5515);
nor U13559 (N_13559,N_5419,N_9639);
nor U13560 (N_13560,N_6405,N_7647);
and U13561 (N_13561,N_6654,N_7593);
nand U13562 (N_13562,N_7083,N_7750);
and U13563 (N_13563,N_5970,N_7506);
nor U13564 (N_13564,N_6316,N_5865);
xnor U13565 (N_13565,N_8453,N_7320);
or U13566 (N_13566,N_9914,N_9640);
and U13567 (N_13567,N_5913,N_5692);
and U13568 (N_13568,N_8440,N_6875);
nand U13569 (N_13569,N_8654,N_8230);
and U13570 (N_13570,N_7551,N_6076);
nand U13571 (N_13571,N_8637,N_8241);
or U13572 (N_13572,N_6362,N_8934);
nand U13573 (N_13573,N_9845,N_7616);
nor U13574 (N_13574,N_7889,N_6256);
and U13575 (N_13575,N_9285,N_8651);
and U13576 (N_13576,N_9776,N_7239);
nor U13577 (N_13577,N_7550,N_6089);
or U13578 (N_13578,N_8744,N_9104);
nand U13579 (N_13579,N_8681,N_6383);
or U13580 (N_13580,N_7648,N_9128);
nand U13581 (N_13581,N_5947,N_9052);
nor U13582 (N_13582,N_6480,N_9283);
xor U13583 (N_13583,N_5243,N_5633);
or U13584 (N_13584,N_6687,N_6235);
and U13585 (N_13585,N_7159,N_7377);
nand U13586 (N_13586,N_7241,N_6699);
and U13587 (N_13587,N_5415,N_6767);
or U13588 (N_13588,N_6424,N_7818);
xnor U13589 (N_13589,N_6412,N_5566);
xor U13590 (N_13590,N_6936,N_6596);
or U13591 (N_13591,N_5227,N_8822);
and U13592 (N_13592,N_9779,N_7418);
nand U13593 (N_13593,N_7117,N_9619);
or U13594 (N_13594,N_5908,N_7320);
or U13595 (N_13595,N_7217,N_6228);
xnor U13596 (N_13596,N_8753,N_9074);
nand U13597 (N_13597,N_5483,N_6903);
nor U13598 (N_13598,N_5637,N_9580);
nor U13599 (N_13599,N_7334,N_5663);
xor U13600 (N_13600,N_5136,N_8773);
nand U13601 (N_13601,N_6797,N_5035);
or U13602 (N_13602,N_5077,N_7827);
and U13603 (N_13603,N_6903,N_9455);
xnor U13604 (N_13604,N_5671,N_9085);
xnor U13605 (N_13605,N_7715,N_7958);
xor U13606 (N_13606,N_9054,N_5685);
xnor U13607 (N_13607,N_6306,N_6574);
xor U13608 (N_13608,N_7472,N_5068);
nand U13609 (N_13609,N_7588,N_8750);
xor U13610 (N_13610,N_9367,N_6125);
nor U13611 (N_13611,N_5179,N_8138);
or U13612 (N_13612,N_6879,N_7733);
and U13613 (N_13613,N_6805,N_6484);
nand U13614 (N_13614,N_7391,N_9876);
xnor U13615 (N_13615,N_9874,N_7938);
nand U13616 (N_13616,N_7197,N_9361);
and U13617 (N_13617,N_7662,N_7062);
nand U13618 (N_13618,N_6581,N_5896);
nand U13619 (N_13619,N_9942,N_6807);
and U13620 (N_13620,N_6912,N_6663);
and U13621 (N_13621,N_7762,N_7282);
nor U13622 (N_13622,N_8292,N_9658);
and U13623 (N_13623,N_8190,N_9970);
and U13624 (N_13624,N_5647,N_7421);
and U13625 (N_13625,N_6161,N_7643);
nand U13626 (N_13626,N_5813,N_6481);
or U13627 (N_13627,N_7662,N_8105);
nor U13628 (N_13628,N_5551,N_5014);
and U13629 (N_13629,N_6288,N_7147);
xor U13630 (N_13630,N_7791,N_7029);
and U13631 (N_13631,N_6771,N_6303);
nand U13632 (N_13632,N_9436,N_7760);
nor U13633 (N_13633,N_5737,N_5347);
nand U13634 (N_13634,N_6493,N_7661);
or U13635 (N_13635,N_9460,N_6498);
nor U13636 (N_13636,N_7495,N_9475);
and U13637 (N_13637,N_9036,N_6544);
or U13638 (N_13638,N_8641,N_5444);
nor U13639 (N_13639,N_7502,N_7802);
nand U13640 (N_13640,N_7639,N_6430);
and U13641 (N_13641,N_7290,N_5540);
xnor U13642 (N_13642,N_7140,N_7764);
xnor U13643 (N_13643,N_9905,N_5464);
nand U13644 (N_13644,N_6975,N_8590);
nand U13645 (N_13645,N_8279,N_8095);
xnor U13646 (N_13646,N_9216,N_6340);
nand U13647 (N_13647,N_5558,N_5219);
and U13648 (N_13648,N_8502,N_6173);
nor U13649 (N_13649,N_9716,N_7704);
nand U13650 (N_13650,N_9391,N_8461);
nor U13651 (N_13651,N_9573,N_7957);
nor U13652 (N_13652,N_5719,N_6615);
nor U13653 (N_13653,N_7096,N_5166);
or U13654 (N_13654,N_8607,N_8673);
nor U13655 (N_13655,N_9155,N_7804);
xor U13656 (N_13656,N_7648,N_7393);
nand U13657 (N_13657,N_5232,N_5586);
and U13658 (N_13658,N_6717,N_9056);
xor U13659 (N_13659,N_6516,N_6949);
nand U13660 (N_13660,N_9368,N_8770);
or U13661 (N_13661,N_8184,N_6747);
nor U13662 (N_13662,N_8430,N_6127);
nand U13663 (N_13663,N_7017,N_9401);
or U13664 (N_13664,N_6704,N_9830);
xnor U13665 (N_13665,N_7679,N_6521);
nor U13666 (N_13666,N_5536,N_8566);
nor U13667 (N_13667,N_6622,N_5457);
xor U13668 (N_13668,N_7419,N_7555);
and U13669 (N_13669,N_9157,N_9227);
and U13670 (N_13670,N_8390,N_8344);
or U13671 (N_13671,N_9931,N_5525);
nand U13672 (N_13672,N_5545,N_9276);
and U13673 (N_13673,N_8503,N_9489);
xor U13674 (N_13674,N_5905,N_5145);
and U13675 (N_13675,N_5200,N_5605);
nor U13676 (N_13676,N_5989,N_7736);
or U13677 (N_13677,N_7477,N_7042);
or U13678 (N_13678,N_9220,N_8761);
or U13679 (N_13679,N_8025,N_7085);
or U13680 (N_13680,N_9579,N_7531);
nor U13681 (N_13681,N_6838,N_9318);
xnor U13682 (N_13682,N_8966,N_9008);
and U13683 (N_13683,N_6577,N_6725);
nand U13684 (N_13684,N_8300,N_5962);
and U13685 (N_13685,N_5417,N_5576);
xor U13686 (N_13686,N_9188,N_5032);
xnor U13687 (N_13687,N_5843,N_8352);
xor U13688 (N_13688,N_6786,N_7970);
or U13689 (N_13689,N_6458,N_7041);
and U13690 (N_13690,N_5583,N_7327);
nand U13691 (N_13691,N_7675,N_9236);
or U13692 (N_13692,N_9684,N_6050);
and U13693 (N_13693,N_6481,N_6550);
nand U13694 (N_13694,N_8448,N_7770);
xnor U13695 (N_13695,N_5638,N_7767);
and U13696 (N_13696,N_9950,N_8401);
or U13697 (N_13697,N_7906,N_7719);
nor U13698 (N_13698,N_6790,N_7912);
or U13699 (N_13699,N_5570,N_8943);
and U13700 (N_13700,N_5416,N_9787);
nand U13701 (N_13701,N_5181,N_9242);
and U13702 (N_13702,N_8388,N_8105);
nand U13703 (N_13703,N_7776,N_7203);
nor U13704 (N_13704,N_7541,N_7280);
and U13705 (N_13705,N_6061,N_5087);
nand U13706 (N_13706,N_5230,N_8509);
xor U13707 (N_13707,N_5425,N_8337);
or U13708 (N_13708,N_5841,N_5531);
and U13709 (N_13709,N_7278,N_8823);
nor U13710 (N_13710,N_8725,N_8167);
or U13711 (N_13711,N_9438,N_5388);
nor U13712 (N_13712,N_5021,N_5882);
nand U13713 (N_13713,N_7654,N_8341);
xor U13714 (N_13714,N_6889,N_7732);
xnor U13715 (N_13715,N_7939,N_5370);
or U13716 (N_13716,N_7007,N_7797);
xor U13717 (N_13717,N_5407,N_9708);
and U13718 (N_13718,N_9437,N_5642);
or U13719 (N_13719,N_7126,N_8783);
or U13720 (N_13720,N_6290,N_5737);
nor U13721 (N_13721,N_6920,N_7534);
nand U13722 (N_13722,N_8805,N_5762);
xnor U13723 (N_13723,N_7965,N_5743);
and U13724 (N_13724,N_9912,N_8840);
xor U13725 (N_13725,N_9469,N_9472);
nor U13726 (N_13726,N_6205,N_5753);
nor U13727 (N_13727,N_8651,N_6199);
nor U13728 (N_13728,N_9790,N_7090);
nand U13729 (N_13729,N_6841,N_9903);
nand U13730 (N_13730,N_8386,N_6453);
and U13731 (N_13731,N_6945,N_5599);
nor U13732 (N_13732,N_8515,N_7979);
nor U13733 (N_13733,N_5344,N_9239);
or U13734 (N_13734,N_5303,N_6118);
nor U13735 (N_13735,N_9941,N_8505);
nand U13736 (N_13736,N_5951,N_6331);
xor U13737 (N_13737,N_6720,N_8900);
nand U13738 (N_13738,N_6885,N_5892);
nand U13739 (N_13739,N_9925,N_5231);
and U13740 (N_13740,N_7144,N_5963);
nand U13741 (N_13741,N_6661,N_5254);
or U13742 (N_13742,N_7002,N_8258);
xor U13743 (N_13743,N_5719,N_9875);
or U13744 (N_13744,N_6747,N_8366);
xnor U13745 (N_13745,N_5190,N_6965);
and U13746 (N_13746,N_6693,N_9996);
and U13747 (N_13747,N_6447,N_7923);
or U13748 (N_13748,N_8545,N_6039);
nor U13749 (N_13749,N_9155,N_6565);
nor U13750 (N_13750,N_9903,N_8122);
and U13751 (N_13751,N_8669,N_6583);
and U13752 (N_13752,N_7027,N_7329);
and U13753 (N_13753,N_7912,N_6563);
nor U13754 (N_13754,N_6438,N_5220);
xnor U13755 (N_13755,N_7734,N_9772);
nand U13756 (N_13756,N_6374,N_8308);
or U13757 (N_13757,N_7522,N_9383);
or U13758 (N_13758,N_5008,N_5994);
and U13759 (N_13759,N_9868,N_8463);
xnor U13760 (N_13760,N_5486,N_8213);
or U13761 (N_13761,N_6297,N_6533);
or U13762 (N_13762,N_5959,N_7193);
and U13763 (N_13763,N_5241,N_6728);
nor U13764 (N_13764,N_7152,N_9540);
nor U13765 (N_13765,N_9065,N_6065);
or U13766 (N_13766,N_7499,N_7198);
nor U13767 (N_13767,N_6588,N_9427);
xor U13768 (N_13768,N_8466,N_5998);
or U13769 (N_13769,N_7624,N_6214);
or U13770 (N_13770,N_9556,N_6770);
or U13771 (N_13771,N_5928,N_8356);
or U13772 (N_13772,N_8948,N_8818);
nand U13773 (N_13773,N_5097,N_6261);
nor U13774 (N_13774,N_7455,N_5191);
xnor U13775 (N_13775,N_7538,N_9359);
nor U13776 (N_13776,N_7316,N_9324);
nor U13777 (N_13777,N_5188,N_6054);
and U13778 (N_13778,N_5137,N_9798);
nor U13779 (N_13779,N_9180,N_5316);
and U13780 (N_13780,N_9636,N_6027);
nor U13781 (N_13781,N_5478,N_5382);
and U13782 (N_13782,N_9387,N_8158);
or U13783 (N_13783,N_9852,N_8394);
nor U13784 (N_13784,N_9579,N_9582);
xnor U13785 (N_13785,N_5275,N_8766);
nand U13786 (N_13786,N_8199,N_9045);
and U13787 (N_13787,N_7895,N_8756);
xnor U13788 (N_13788,N_6982,N_5879);
or U13789 (N_13789,N_6944,N_8970);
xor U13790 (N_13790,N_8675,N_6479);
xor U13791 (N_13791,N_7083,N_9238);
nor U13792 (N_13792,N_6089,N_8186);
nor U13793 (N_13793,N_7546,N_7590);
and U13794 (N_13794,N_7901,N_7239);
xnor U13795 (N_13795,N_6857,N_7067);
nor U13796 (N_13796,N_6284,N_7914);
and U13797 (N_13797,N_5151,N_5190);
and U13798 (N_13798,N_5294,N_8293);
nor U13799 (N_13799,N_6073,N_5892);
or U13800 (N_13800,N_7752,N_7773);
or U13801 (N_13801,N_7776,N_9657);
xor U13802 (N_13802,N_7984,N_6806);
nor U13803 (N_13803,N_7011,N_7746);
or U13804 (N_13804,N_5465,N_7672);
and U13805 (N_13805,N_7859,N_5972);
xnor U13806 (N_13806,N_5155,N_7375);
or U13807 (N_13807,N_8800,N_9319);
xnor U13808 (N_13808,N_6892,N_5068);
and U13809 (N_13809,N_8999,N_7780);
and U13810 (N_13810,N_9603,N_7785);
or U13811 (N_13811,N_8075,N_6053);
and U13812 (N_13812,N_6057,N_8812);
and U13813 (N_13813,N_5318,N_7512);
nor U13814 (N_13814,N_6510,N_9065);
nor U13815 (N_13815,N_8927,N_7153);
or U13816 (N_13816,N_7600,N_8697);
nor U13817 (N_13817,N_8355,N_5201);
or U13818 (N_13818,N_8563,N_7523);
nor U13819 (N_13819,N_7044,N_7942);
nand U13820 (N_13820,N_8671,N_6614);
or U13821 (N_13821,N_5167,N_9945);
or U13822 (N_13822,N_7431,N_8219);
and U13823 (N_13823,N_7435,N_8824);
and U13824 (N_13824,N_7965,N_5348);
or U13825 (N_13825,N_9321,N_7637);
nor U13826 (N_13826,N_6039,N_6427);
xor U13827 (N_13827,N_6235,N_6290);
and U13828 (N_13828,N_7873,N_7692);
xnor U13829 (N_13829,N_7870,N_8439);
and U13830 (N_13830,N_7462,N_8001);
xor U13831 (N_13831,N_9065,N_9396);
nand U13832 (N_13832,N_9148,N_7719);
nor U13833 (N_13833,N_9287,N_6875);
and U13834 (N_13834,N_5930,N_6378);
nor U13835 (N_13835,N_6229,N_6890);
nor U13836 (N_13836,N_8297,N_6135);
nor U13837 (N_13837,N_7830,N_5476);
and U13838 (N_13838,N_7638,N_7128);
or U13839 (N_13839,N_5529,N_6803);
nand U13840 (N_13840,N_8220,N_5976);
nor U13841 (N_13841,N_7412,N_5646);
or U13842 (N_13842,N_7554,N_5320);
xor U13843 (N_13843,N_8074,N_9268);
or U13844 (N_13844,N_7046,N_9462);
nor U13845 (N_13845,N_8233,N_5410);
or U13846 (N_13846,N_6880,N_6820);
nand U13847 (N_13847,N_7456,N_6289);
xnor U13848 (N_13848,N_6830,N_7546);
xnor U13849 (N_13849,N_8549,N_9090);
and U13850 (N_13850,N_7732,N_8156);
xnor U13851 (N_13851,N_9562,N_8138);
or U13852 (N_13852,N_6865,N_8224);
and U13853 (N_13853,N_6429,N_7499);
xor U13854 (N_13854,N_8532,N_8089);
xor U13855 (N_13855,N_6304,N_6760);
nand U13856 (N_13856,N_5955,N_5799);
and U13857 (N_13857,N_5102,N_6682);
xnor U13858 (N_13858,N_7637,N_7722);
and U13859 (N_13859,N_9646,N_5878);
or U13860 (N_13860,N_5770,N_6234);
nand U13861 (N_13861,N_8883,N_5655);
nor U13862 (N_13862,N_8263,N_8608);
nand U13863 (N_13863,N_5690,N_5682);
or U13864 (N_13864,N_7477,N_9182);
and U13865 (N_13865,N_8558,N_7638);
nand U13866 (N_13866,N_6048,N_7688);
and U13867 (N_13867,N_5210,N_8858);
or U13868 (N_13868,N_7950,N_8205);
nand U13869 (N_13869,N_7291,N_5793);
and U13870 (N_13870,N_7131,N_7327);
xnor U13871 (N_13871,N_8191,N_9156);
or U13872 (N_13872,N_7350,N_5057);
nand U13873 (N_13873,N_5395,N_5051);
xnor U13874 (N_13874,N_6643,N_7025);
xnor U13875 (N_13875,N_8314,N_7838);
nand U13876 (N_13876,N_6711,N_7655);
xnor U13877 (N_13877,N_9760,N_7705);
nand U13878 (N_13878,N_7333,N_9986);
xor U13879 (N_13879,N_7666,N_6027);
or U13880 (N_13880,N_9041,N_6284);
nor U13881 (N_13881,N_8822,N_7248);
nor U13882 (N_13882,N_9480,N_9708);
nand U13883 (N_13883,N_6863,N_9423);
and U13884 (N_13884,N_7121,N_7647);
xor U13885 (N_13885,N_9946,N_6130);
nor U13886 (N_13886,N_5590,N_9228);
or U13887 (N_13887,N_6397,N_9818);
and U13888 (N_13888,N_7458,N_8298);
xnor U13889 (N_13889,N_6066,N_7804);
xor U13890 (N_13890,N_6359,N_8550);
or U13891 (N_13891,N_6179,N_7152);
and U13892 (N_13892,N_6175,N_6617);
and U13893 (N_13893,N_5596,N_8286);
or U13894 (N_13894,N_8388,N_5083);
nor U13895 (N_13895,N_9576,N_7191);
nor U13896 (N_13896,N_7867,N_6872);
and U13897 (N_13897,N_6210,N_9573);
nand U13898 (N_13898,N_9456,N_9686);
nor U13899 (N_13899,N_5394,N_5160);
or U13900 (N_13900,N_6822,N_6976);
or U13901 (N_13901,N_6268,N_8048);
nor U13902 (N_13902,N_7438,N_6087);
nand U13903 (N_13903,N_9000,N_6451);
xnor U13904 (N_13904,N_7044,N_7240);
or U13905 (N_13905,N_6723,N_8832);
or U13906 (N_13906,N_8231,N_9473);
xor U13907 (N_13907,N_5976,N_7718);
or U13908 (N_13908,N_8216,N_9625);
or U13909 (N_13909,N_6528,N_6698);
nor U13910 (N_13910,N_6897,N_8516);
nand U13911 (N_13911,N_9026,N_9502);
xnor U13912 (N_13912,N_8650,N_7314);
nand U13913 (N_13913,N_7968,N_9123);
and U13914 (N_13914,N_5585,N_5802);
or U13915 (N_13915,N_7516,N_9512);
xnor U13916 (N_13916,N_7765,N_8260);
nand U13917 (N_13917,N_9425,N_6325);
nor U13918 (N_13918,N_6872,N_7406);
nor U13919 (N_13919,N_8570,N_7061);
or U13920 (N_13920,N_7060,N_7262);
or U13921 (N_13921,N_5675,N_5590);
nand U13922 (N_13922,N_6200,N_7965);
nand U13923 (N_13923,N_6366,N_7301);
nand U13924 (N_13924,N_9297,N_6370);
and U13925 (N_13925,N_8318,N_5176);
nand U13926 (N_13926,N_5058,N_5520);
or U13927 (N_13927,N_7013,N_5672);
xnor U13928 (N_13928,N_5131,N_7933);
nand U13929 (N_13929,N_5832,N_6759);
or U13930 (N_13930,N_9031,N_7370);
xnor U13931 (N_13931,N_5541,N_5572);
or U13932 (N_13932,N_9749,N_8209);
nor U13933 (N_13933,N_6469,N_7769);
nand U13934 (N_13934,N_9319,N_5896);
xnor U13935 (N_13935,N_5358,N_7134);
xnor U13936 (N_13936,N_9471,N_6556);
xor U13937 (N_13937,N_6547,N_6050);
nor U13938 (N_13938,N_9388,N_8827);
xnor U13939 (N_13939,N_9744,N_5644);
nor U13940 (N_13940,N_6953,N_7291);
or U13941 (N_13941,N_5940,N_9877);
nor U13942 (N_13942,N_6734,N_5825);
nand U13943 (N_13943,N_8754,N_9550);
nand U13944 (N_13944,N_8535,N_5606);
or U13945 (N_13945,N_5314,N_9674);
nor U13946 (N_13946,N_5837,N_5858);
nor U13947 (N_13947,N_9296,N_7547);
and U13948 (N_13948,N_7187,N_6498);
nor U13949 (N_13949,N_6737,N_7228);
or U13950 (N_13950,N_6465,N_5376);
nor U13951 (N_13951,N_9799,N_5276);
nand U13952 (N_13952,N_7022,N_8404);
nor U13953 (N_13953,N_6702,N_8379);
or U13954 (N_13954,N_8903,N_5149);
and U13955 (N_13955,N_9172,N_8911);
xor U13956 (N_13956,N_5455,N_5170);
and U13957 (N_13957,N_9452,N_9166);
and U13958 (N_13958,N_9069,N_6249);
nor U13959 (N_13959,N_9118,N_9326);
and U13960 (N_13960,N_8672,N_8747);
or U13961 (N_13961,N_5052,N_6303);
or U13962 (N_13962,N_9451,N_5859);
or U13963 (N_13963,N_6272,N_7269);
xnor U13964 (N_13964,N_5986,N_5072);
xnor U13965 (N_13965,N_8824,N_5425);
and U13966 (N_13966,N_7605,N_6161);
and U13967 (N_13967,N_9596,N_9273);
or U13968 (N_13968,N_7513,N_6139);
nand U13969 (N_13969,N_8288,N_8969);
and U13970 (N_13970,N_6461,N_7574);
or U13971 (N_13971,N_7658,N_7736);
nor U13972 (N_13972,N_7646,N_9237);
or U13973 (N_13973,N_6289,N_6272);
and U13974 (N_13974,N_5731,N_9697);
and U13975 (N_13975,N_7300,N_7134);
nand U13976 (N_13976,N_6359,N_7543);
nand U13977 (N_13977,N_5932,N_7746);
xor U13978 (N_13978,N_6147,N_7684);
and U13979 (N_13979,N_7419,N_9072);
xor U13980 (N_13980,N_5059,N_9208);
nor U13981 (N_13981,N_9848,N_7638);
and U13982 (N_13982,N_7748,N_7364);
xor U13983 (N_13983,N_8681,N_8195);
nand U13984 (N_13984,N_5999,N_7771);
xor U13985 (N_13985,N_7231,N_8924);
or U13986 (N_13986,N_6419,N_9573);
or U13987 (N_13987,N_9572,N_8886);
and U13988 (N_13988,N_9821,N_7825);
and U13989 (N_13989,N_6423,N_7535);
nand U13990 (N_13990,N_8955,N_5900);
nand U13991 (N_13991,N_6001,N_6481);
nand U13992 (N_13992,N_9410,N_9123);
nor U13993 (N_13993,N_7776,N_6003);
nand U13994 (N_13994,N_5422,N_5838);
or U13995 (N_13995,N_7378,N_7444);
xnor U13996 (N_13996,N_9879,N_8878);
or U13997 (N_13997,N_6288,N_7031);
nor U13998 (N_13998,N_8264,N_7518);
nand U13999 (N_13999,N_9409,N_8356);
nand U14000 (N_14000,N_7960,N_6938);
nor U14001 (N_14001,N_5199,N_7459);
and U14002 (N_14002,N_7837,N_6821);
nand U14003 (N_14003,N_8366,N_8867);
nor U14004 (N_14004,N_9019,N_9522);
xor U14005 (N_14005,N_9374,N_7849);
or U14006 (N_14006,N_5638,N_5720);
nand U14007 (N_14007,N_9941,N_9162);
and U14008 (N_14008,N_6872,N_8892);
xnor U14009 (N_14009,N_9826,N_7208);
nand U14010 (N_14010,N_8115,N_7893);
and U14011 (N_14011,N_7695,N_9943);
or U14012 (N_14012,N_8332,N_7631);
xnor U14013 (N_14013,N_5080,N_5376);
nand U14014 (N_14014,N_6037,N_7142);
xor U14015 (N_14015,N_8213,N_5611);
xor U14016 (N_14016,N_6029,N_9378);
nand U14017 (N_14017,N_9398,N_8054);
xnor U14018 (N_14018,N_9446,N_5649);
or U14019 (N_14019,N_9204,N_8005);
nand U14020 (N_14020,N_6705,N_8758);
xnor U14021 (N_14021,N_9645,N_9728);
nand U14022 (N_14022,N_5301,N_7795);
and U14023 (N_14023,N_5203,N_8501);
and U14024 (N_14024,N_8615,N_6699);
or U14025 (N_14025,N_6541,N_6523);
nor U14026 (N_14026,N_8143,N_5032);
nor U14027 (N_14027,N_6914,N_8168);
nor U14028 (N_14028,N_6876,N_7260);
nand U14029 (N_14029,N_5895,N_7734);
nand U14030 (N_14030,N_9945,N_7300);
and U14031 (N_14031,N_7668,N_7380);
and U14032 (N_14032,N_9607,N_9938);
nor U14033 (N_14033,N_7494,N_5634);
nor U14034 (N_14034,N_8043,N_8711);
or U14035 (N_14035,N_9902,N_6935);
nor U14036 (N_14036,N_6288,N_6072);
nor U14037 (N_14037,N_6956,N_6087);
nor U14038 (N_14038,N_5859,N_5251);
nand U14039 (N_14039,N_8402,N_8766);
xnor U14040 (N_14040,N_5051,N_8974);
xor U14041 (N_14041,N_5090,N_8759);
nand U14042 (N_14042,N_5907,N_9005);
nor U14043 (N_14043,N_7983,N_9578);
nand U14044 (N_14044,N_7973,N_5286);
and U14045 (N_14045,N_7051,N_5181);
and U14046 (N_14046,N_9985,N_7504);
and U14047 (N_14047,N_7219,N_8543);
nand U14048 (N_14048,N_7911,N_9703);
nand U14049 (N_14049,N_5704,N_7439);
xnor U14050 (N_14050,N_8045,N_9155);
or U14051 (N_14051,N_9889,N_5438);
or U14052 (N_14052,N_5127,N_5015);
nor U14053 (N_14053,N_6388,N_6107);
xnor U14054 (N_14054,N_6759,N_8668);
or U14055 (N_14055,N_7347,N_7231);
and U14056 (N_14056,N_8632,N_6846);
and U14057 (N_14057,N_7836,N_8362);
xnor U14058 (N_14058,N_9104,N_5355);
or U14059 (N_14059,N_5509,N_9105);
or U14060 (N_14060,N_8730,N_9197);
nand U14061 (N_14061,N_7188,N_9511);
nand U14062 (N_14062,N_7530,N_9466);
nand U14063 (N_14063,N_6873,N_9586);
and U14064 (N_14064,N_5586,N_8922);
nor U14065 (N_14065,N_7127,N_7927);
or U14066 (N_14066,N_6135,N_6141);
and U14067 (N_14067,N_6539,N_9714);
or U14068 (N_14068,N_5094,N_5296);
xnor U14069 (N_14069,N_8933,N_7242);
xnor U14070 (N_14070,N_7461,N_5979);
xor U14071 (N_14071,N_9145,N_8384);
nand U14072 (N_14072,N_8348,N_6534);
and U14073 (N_14073,N_9932,N_6897);
or U14074 (N_14074,N_5057,N_8870);
nor U14075 (N_14075,N_8701,N_9287);
nor U14076 (N_14076,N_7557,N_9930);
and U14077 (N_14077,N_6613,N_9797);
and U14078 (N_14078,N_9985,N_6196);
or U14079 (N_14079,N_6276,N_6564);
or U14080 (N_14080,N_5898,N_8382);
nor U14081 (N_14081,N_6036,N_5056);
xor U14082 (N_14082,N_6236,N_7126);
nand U14083 (N_14083,N_5594,N_6157);
nor U14084 (N_14084,N_9883,N_7667);
nor U14085 (N_14085,N_7256,N_6057);
nor U14086 (N_14086,N_9153,N_7283);
xnor U14087 (N_14087,N_7766,N_7663);
xnor U14088 (N_14088,N_9128,N_7003);
or U14089 (N_14089,N_9524,N_8808);
or U14090 (N_14090,N_7977,N_8972);
and U14091 (N_14091,N_8935,N_8014);
and U14092 (N_14092,N_7291,N_5291);
or U14093 (N_14093,N_7401,N_8232);
xnor U14094 (N_14094,N_8277,N_5314);
xor U14095 (N_14095,N_6549,N_8464);
or U14096 (N_14096,N_8895,N_8725);
nand U14097 (N_14097,N_7342,N_8207);
or U14098 (N_14098,N_6542,N_5547);
nor U14099 (N_14099,N_8752,N_9500);
or U14100 (N_14100,N_8150,N_6787);
nand U14101 (N_14101,N_6637,N_6054);
and U14102 (N_14102,N_5357,N_8324);
or U14103 (N_14103,N_7852,N_5160);
xnor U14104 (N_14104,N_6843,N_8429);
nand U14105 (N_14105,N_9692,N_8210);
nand U14106 (N_14106,N_8247,N_7129);
nand U14107 (N_14107,N_5399,N_5950);
nand U14108 (N_14108,N_5921,N_8796);
and U14109 (N_14109,N_6792,N_9676);
nor U14110 (N_14110,N_5270,N_5812);
nand U14111 (N_14111,N_6733,N_7038);
or U14112 (N_14112,N_8906,N_6874);
and U14113 (N_14113,N_9863,N_9337);
xor U14114 (N_14114,N_5253,N_7390);
and U14115 (N_14115,N_6460,N_8053);
nor U14116 (N_14116,N_5746,N_5713);
or U14117 (N_14117,N_5331,N_6246);
nor U14118 (N_14118,N_9431,N_9458);
nor U14119 (N_14119,N_7181,N_9152);
xnor U14120 (N_14120,N_8814,N_6088);
xnor U14121 (N_14121,N_8758,N_9707);
nand U14122 (N_14122,N_6704,N_6145);
nand U14123 (N_14123,N_8330,N_7369);
xnor U14124 (N_14124,N_7086,N_7191);
nor U14125 (N_14125,N_5226,N_7693);
or U14126 (N_14126,N_8869,N_7145);
nand U14127 (N_14127,N_5532,N_9258);
or U14128 (N_14128,N_5817,N_9233);
nand U14129 (N_14129,N_8064,N_8697);
and U14130 (N_14130,N_7329,N_7000);
or U14131 (N_14131,N_9952,N_6347);
nor U14132 (N_14132,N_9032,N_6687);
xnor U14133 (N_14133,N_7643,N_5279);
nand U14134 (N_14134,N_6136,N_7631);
nor U14135 (N_14135,N_8662,N_9741);
or U14136 (N_14136,N_9087,N_8088);
nand U14137 (N_14137,N_9649,N_6478);
xnor U14138 (N_14138,N_7821,N_5233);
or U14139 (N_14139,N_5177,N_6263);
nand U14140 (N_14140,N_8857,N_8867);
nor U14141 (N_14141,N_8392,N_7387);
or U14142 (N_14142,N_8118,N_9453);
or U14143 (N_14143,N_8191,N_9896);
and U14144 (N_14144,N_7610,N_5141);
xnor U14145 (N_14145,N_5229,N_6350);
nor U14146 (N_14146,N_9848,N_7865);
and U14147 (N_14147,N_6535,N_5401);
nand U14148 (N_14148,N_5740,N_9394);
nor U14149 (N_14149,N_7708,N_8893);
xnor U14150 (N_14150,N_6341,N_9461);
or U14151 (N_14151,N_8528,N_9313);
xor U14152 (N_14152,N_7969,N_9865);
xnor U14153 (N_14153,N_6998,N_5940);
and U14154 (N_14154,N_7855,N_6077);
nor U14155 (N_14155,N_5148,N_9902);
or U14156 (N_14156,N_9160,N_7383);
nand U14157 (N_14157,N_7894,N_9819);
or U14158 (N_14158,N_7130,N_9953);
nand U14159 (N_14159,N_6640,N_8486);
nor U14160 (N_14160,N_5536,N_5648);
and U14161 (N_14161,N_5228,N_6248);
or U14162 (N_14162,N_5742,N_8516);
or U14163 (N_14163,N_9693,N_8045);
and U14164 (N_14164,N_9924,N_8090);
nand U14165 (N_14165,N_5872,N_7565);
xor U14166 (N_14166,N_5338,N_7752);
xor U14167 (N_14167,N_5615,N_9006);
and U14168 (N_14168,N_9364,N_7018);
or U14169 (N_14169,N_9297,N_5125);
and U14170 (N_14170,N_6320,N_8119);
nand U14171 (N_14171,N_6577,N_9479);
nand U14172 (N_14172,N_8582,N_5124);
nor U14173 (N_14173,N_7517,N_9202);
or U14174 (N_14174,N_8217,N_6101);
or U14175 (N_14175,N_7293,N_8050);
xor U14176 (N_14176,N_9033,N_5922);
and U14177 (N_14177,N_7989,N_9294);
and U14178 (N_14178,N_7602,N_6674);
nor U14179 (N_14179,N_5863,N_6679);
and U14180 (N_14180,N_9745,N_7671);
and U14181 (N_14181,N_6493,N_8457);
xnor U14182 (N_14182,N_9414,N_6331);
nand U14183 (N_14183,N_6538,N_6706);
nor U14184 (N_14184,N_6895,N_7525);
or U14185 (N_14185,N_9895,N_5488);
and U14186 (N_14186,N_5160,N_5859);
and U14187 (N_14187,N_5010,N_9270);
or U14188 (N_14188,N_6292,N_9509);
nor U14189 (N_14189,N_7668,N_5770);
xnor U14190 (N_14190,N_7759,N_5082);
nor U14191 (N_14191,N_5695,N_9212);
or U14192 (N_14192,N_5271,N_9885);
and U14193 (N_14193,N_5557,N_8777);
xor U14194 (N_14194,N_7644,N_6744);
or U14195 (N_14195,N_9545,N_5178);
or U14196 (N_14196,N_7145,N_6337);
xnor U14197 (N_14197,N_7408,N_7038);
nand U14198 (N_14198,N_7864,N_8152);
nor U14199 (N_14199,N_6676,N_5483);
or U14200 (N_14200,N_6824,N_6034);
nor U14201 (N_14201,N_7106,N_7463);
and U14202 (N_14202,N_7968,N_8561);
and U14203 (N_14203,N_8145,N_9895);
nand U14204 (N_14204,N_7019,N_8820);
nand U14205 (N_14205,N_6014,N_7071);
nor U14206 (N_14206,N_5620,N_6273);
and U14207 (N_14207,N_8868,N_5427);
nand U14208 (N_14208,N_7124,N_7567);
and U14209 (N_14209,N_6888,N_5433);
nand U14210 (N_14210,N_6235,N_5707);
xor U14211 (N_14211,N_6578,N_8093);
or U14212 (N_14212,N_8449,N_5383);
nand U14213 (N_14213,N_6689,N_5574);
nand U14214 (N_14214,N_8614,N_7199);
and U14215 (N_14215,N_9432,N_6242);
xor U14216 (N_14216,N_9959,N_8802);
nor U14217 (N_14217,N_6542,N_8266);
and U14218 (N_14218,N_5791,N_5965);
or U14219 (N_14219,N_6516,N_8162);
or U14220 (N_14220,N_7336,N_6648);
nor U14221 (N_14221,N_7990,N_7940);
nand U14222 (N_14222,N_8661,N_6814);
nor U14223 (N_14223,N_8181,N_5861);
xnor U14224 (N_14224,N_7676,N_7324);
nand U14225 (N_14225,N_5255,N_7933);
xnor U14226 (N_14226,N_6705,N_7816);
nand U14227 (N_14227,N_6572,N_9140);
or U14228 (N_14228,N_6742,N_5356);
xor U14229 (N_14229,N_9619,N_5993);
xnor U14230 (N_14230,N_9029,N_9294);
xor U14231 (N_14231,N_5656,N_7100);
nor U14232 (N_14232,N_6605,N_5124);
or U14233 (N_14233,N_6864,N_9523);
xnor U14234 (N_14234,N_9624,N_9912);
and U14235 (N_14235,N_6513,N_7949);
nor U14236 (N_14236,N_6371,N_7947);
xnor U14237 (N_14237,N_9254,N_5807);
xor U14238 (N_14238,N_6951,N_8369);
nor U14239 (N_14239,N_6134,N_9811);
and U14240 (N_14240,N_8450,N_8429);
nor U14241 (N_14241,N_6090,N_5899);
or U14242 (N_14242,N_9380,N_6691);
and U14243 (N_14243,N_7556,N_7168);
and U14244 (N_14244,N_5749,N_5183);
nor U14245 (N_14245,N_7149,N_5290);
or U14246 (N_14246,N_6921,N_5138);
nand U14247 (N_14247,N_5885,N_5651);
and U14248 (N_14248,N_9093,N_8094);
nand U14249 (N_14249,N_8887,N_9858);
or U14250 (N_14250,N_9736,N_7353);
nor U14251 (N_14251,N_5146,N_6399);
or U14252 (N_14252,N_5219,N_6885);
and U14253 (N_14253,N_6769,N_6016);
xnor U14254 (N_14254,N_7840,N_9532);
nand U14255 (N_14255,N_9376,N_9335);
or U14256 (N_14256,N_5519,N_8285);
xor U14257 (N_14257,N_7723,N_8497);
and U14258 (N_14258,N_8794,N_7650);
or U14259 (N_14259,N_5967,N_8557);
or U14260 (N_14260,N_9934,N_7504);
and U14261 (N_14261,N_5701,N_7530);
nand U14262 (N_14262,N_5128,N_6710);
and U14263 (N_14263,N_6858,N_5650);
nor U14264 (N_14264,N_5498,N_8134);
xnor U14265 (N_14265,N_6405,N_9006);
nor U14266 (N_14266,N_6526,N_7990);
nor U14267 (N_14267,N_6973,N_7282);
or U14268 (N_14268,N_5624,N_8622);
and U14269 (N_14269,N_6996,N_5112);
nand U14270 (N_14270,N_8673,N_9305);
nand U14271 (N_14271,N_5491,N_7183);
nand U14272 (N_14272,N_6012,N_5714);
nand U14273 (N_14273,N_6970,N_5091);
nor U14274 (N_14274,N_9298,N_6714);
xnor U14275 (N_14275,N_5140,N_5998);
nor U14276 (N_14276,N_9109,N_8513);
and U14277 (N_14277,N_7162,N_8587);
and U14278 (N_14278,N_9471,N_6885);
xnor U14279 (N_14279,N_5637,N_6139);
and U14280 (N_14280,N_9681,N_8789);
nand U14281 (N_14281,N_9728,N_5788);
nor U14282 (N_14282,N_6797,N_6891);
nand U14283 (N_14283,N_9783,N_9219);
or U14284 (N_14284,N_7067,N_6140);
xor U14285 (N_14285,N_7877,N_9740);
and U14286 (N_14286,N_9747,N_8630);
nand U14287 (N_14287,N_8025,N_5469);
nor U14288 (N_14288,N_5859,N_5189);
nor U14289 (N_14289,N_9440,N_5435);
nor U14290 (N_14290,N_8644,N_7508);
nor U14291 (N_14291,N_7665,N_5117);
and U14292 (N_14292,N_6009,N_5743);
nor U14293 (N_14293,N_8955,N_6590);
or U14294 (N_14294,N_8262,N_6628);
or U14295 (N_14295,N_9944,N_8773);
nand U14296 (N_14296,N_7439,N_5309);
and U14297 (N_14297,N_6209,N_5147);
and U14298 (N_14298,N_8397,N_6009);
xnor U14299 (N_14299,N_9935,N_6677);
or U14300 (N_14300,N_9657,N_6995);
and U14301 (N_14301,N_5130,N_9242);
nand U14302 (N_14302,N_8275,N_8634);
nand U14303 (N_14303,N_7496,N_9130);
xnor U14304 (N_14304,N_9930,N_6407);
nor U14305 (N_14305,N_7075,N_5958);
nor U14306 (N_14306,N_5017,N_9966);
or U14307 (N_14307,N_5465,N_7193);
xnor U14308 (N_14308,N_6975,N_9814);
nor U14309 (N_14309,N_6278,N_9423);
nor U14310 (N_14310,N_6827,N_9100);
or U14311 (N_14311,N_6825,N_5394);
nand U14312 (N_14312,N_6356,N_6086);
or U14313 (N_14313,N_6188,N_5077);
nor U14314 (N_14314,N_8856,N_6627);
nand U14315 (N_14315,N_5575,N_8573);
nand U14316 (N_14316,N_5312,N_9285);
nand U14317 (N_14317,N_5916,N_5794);
nand U14318 (N_14318,N_6770,N_8436);
nand U14319 (N_14319,N_8045,N_7958);
or U14320 (N_14320,N_7503,N_8184);
xnor U14321 (N_14321,N_9361,N_9108);
nor U14322 (N_14322,N_7122,N_5337);
and U14323 (N_14323,N_8167,N_9937);
and U14324 (N_14324,N_6478,N_6809);
xnor U14325 (N_14325,N_5775,N_9410);
nor U14326 (N_14326,N_6001,N_8403);
or U14327 (N_14327,N_6632,N_6736);
xor U14328 (N_14328,N_7705,N_5397);
and U14329 (N_14329,N_8372,N_9214);
xnor U14330 (N_14330,N_6574,N_8612);
or U14331 (N_14331,N_9652,N_8601);
or U14332 (N_14332,N_6823,N_5587);
and U14333 (N_14333,N_5583,N_5003);
nand U14334 (N_14334,N_9565,N_8280);
and U14335 (N_14335,N_6841,N_9865);
and U14336 (N_14336,N_5482,N_5384);
or U14337 (N_14337,N_5610,N_9538);
nand U14338 (N_14338,N_6796,N_8168);
nand U14339 (N_14339,N_8015,N_5593);
nor U14340 (N_14340,N_6200,N_5421);
and U14341 (N_14341,N_8317,N_9603);
and U14342 (N_14342,N_8549,N_8874);
xor U14343 (N_14343,N_7346,N_6638);
and U14344 (N_14344,N_8771,N_9701);
nand U14345 (N_14345,N_9885,N_5832);
or U14346 (N_14346,N_5282,N_6080);
xor U14347 (N_14347,N_9962,N_6182);
xor U14348 (N_14348,N_6122,N_7508);
nor U14349 (N_14349,N_5404,N_9567);
and U14350 (N_14350,N_7966,N_9000);
or U14351 (N_14351,N_5585,N_8415);
or U14352 (N_14352,N_5760,N_8049);
and U14353 (N_14353,N_5608,N_8048);
and U14354 (N_14354,N_6582,N_7856);
nand U14355 (N_14355,N_9848,N_7359);
and U14356 (N_14356,N_8677,N_5631);
xnor U14357 (N_14357,N_5131,N_9138);
and U14358 (N_14358,N_6501,N_7485);
xor U14359 (N_14359,N_7950,N_7085);
nand U14360 (N_14360,N_7413,N_7154);
and U14361 (N_14361,N_7933,N_7277);
or U14362 (N_14362,N_5456,N_9816);
or U14363 (N_14363,N_5269,N_6403);
or U14364 (N_14364,N_8256,N_6881);
nor U14365 (N_14365,N_8332,N_7763);
or U14366 (N_14366,N_5742,N_7894);
nor U14367 (N_14367,N_9017,N_5969);
and U14368 (N_14368,N_8617,N_6161);
nor U14369 (N_14369,N_9180,N_8122);
and U14370 (N_14370,N_5612,N_9398);
or U14371 (N_14371,N_5796,N_7672);
xnor U14372 (N_14372,N_8006,N_7897);
or U14373 (N_14373,N_9063,N_6116);
or U14374 (N_14374,N_6084,N_5305);
or U14375 (N_14375,N_8389,N_8177);
xor U14376 (N_14376,N_7510,N_7846);
xor U14377 (N_14377,N_8930,N_9738);
and U14378 (N_14378,N_6792,N_5532);
and U14379 (N_14379,N_5246,N_9115);
nor U14380 (N_14380,N_9943,N_8494);
and U14381 (N_14381,N_5762,N_8441);
nor U14382 (N_14382,N_7645,N_6061);
nor U14383 (N_14383,N_8805,N_8120);
nor U14384 (N_14384,N_6188,N_7966);
nand U14385 (N_14385,N_8579,N_8398);
xnor U14386 (N_14386,N_5222,N_7493);
or U14387 (N_14387,N_9570,N_5604);
and U14388 (N_14388,N_6750,N_5716);
nor U14389 (N_14389,N_9362,N_5033);
and U14390 (N_14390,N_5327,N_9926);
xnor U14391 (N_14391,N_7644,N_5238);
nor U14392 (N_14392,N_8289,N_5115);
and U14393 (N_14393,N_6161,N_8094);
nor U14394 (N_14394,N_9683,N_6401);
or U14395 (N_14395,N_6899,N_7290);
xor U14396 (N_14396,N_8919,N_6831);
xnor U14397 (N_14397,N_5760,N_7061);
and U14398 (N_14398,N_7013,N_8972);
xnor U14399 (N_14399,N_6123,N_6854);
xnor U14400 (N_14400,N_9119,N_7119);
xor U14401 (N_14401,N_6450,N_8411);
nor U14402 (N_14402,N_8347,N_8682);
nor U14403 (N_14403,N_6260,N_9585);
xnor U14404 (N_14404,N_8234,N_7511);
nand U14405 (N_14405,N_5680,N_7077);
and U14406 (N_14406,N_7879,N_9883);
and U14407 (N_14407,N_9874,N_8353);
nand U14408 (N_14408,N_5287,N_9111);
nor U14409 (N_14409,N_8626,N_9607);
nand U14410 (N_14410,N_7677,N_9596);
nand U14411 (N_14411,N_8745,N_7376);
nor U14412 (N_14412,N_8786,N_8859);
xor U14413 (N_14413,N_5531,N_6633);
xor U14414 (N_14414,N_6258,N_6293);
or U14415 (N_14415,N_6292,N_9026);
nor U14416 (N_14416,N_6898,N_9189);
xor U14417 (N_14417,N_6066,N_9899);
xor U14418 (N_14418,N_9633,N_9627);
and U14419 (N_14419,N_9932,N_7594);
and U14420 (N_14420,N_7538,N_8093);
and U14421 (N_14421,N_9868,N_8481);
and U14422 (N_14422,N_6256,N_6232);
nand U14423 (N_14423,N_5819,N_6761);
or U14424 (N_14424,N_7435,N_9159);
nor U14425 (N_14425,N_9271,N_5193);
and U14426 (N_14426,N_7704,N_6397);
xor U14427 (N_14427,N_8460,N_9736);
or U14428 (N_14428,N_8242,N_8545);
or U14429 (N_14429,N_5863,N_5852);
or U14430 (N_14430,N_8835,N_9266);
nor U14431 (N_14431,N_5319,N_8852);
nor U14432 (N_14432,N_7538,N_7494);
nor U14433 (N_14433,N_8644,N_6511);
or U14434 (N_14434,N_6383,N_5005);
or U14435 (N_14435,N_8161,N_8658);
nand U14436 (N_14436,N_6322,N_5171);
xnor U14437 (N_14437,N_6135,N_8519);
and U14438 (N_14438,N_5287,N_6775);
xnor U14439 (N_14439,N_6230,N_8464);
or U14440 (N_14440,N_9103,N_5918);
and U14441 (N_14441,N_9737,N_8737);
xnor U14442 (N_14442,N_9374,N_8196);
or U14443 (N_14443,N_6156,N_8824);
nor U14444 (N_14444,N_8151,N_8339);
nor U14445 (N_14445,N_7902,N_7864);
nand U14446 (N_14446,N_9952,N_7587);
nor U14447 (N_14447,N_9103,N_7467);
and U14448 (N_14448,N_8364,N_9741);
or U14449 (N_14449,N_8597,N_8418);
nand U14450 (N_14450,N_6474,N_7216);
nand U14451 (N_14451,N_5504,N_7376);
or U14452 (N_14452,N_8475,N_6731);
or U14453 (N_14453,N_8236,N_6626);
and U14454 (N_14454,N_6977,N_7116);
and U14455 (N_14455,N_8455,N_5173);
and U14456 (N_14456,N_7474,N_8764);
nor U14457 (N_14457,N_7229,N_7135);
and U14458 (N_14458,N_9084,N_7261);
xnor U14459 (N_14459,N_7061,N_7019);
or U14460 (N_14460,N_6179,N_8717);
nand U14461 (N_14461,N_8190,N_9892);
nand U14462 (N_14462,N_9646,N_5376);
or U14463 (N_14463,N_5934,N_9146);
or U14464 (N_14464,N_8996,N_6721);
nand U14465 (N_14465,N_9124,N_7490);
nand U14466 (N_14466,N_9072,N_5933);
nand U14467 (N_14467,N_6887,N_7802);
or U14468 (N_14468,N_9249,N_9340);
or U14469 (N_14469,N_9241,N_6741);
nor U14470 (N_14470,N_8252,N_6145);
xnor U14471 (N_14471,N_8948,N_5753);
xor U14472 (N_14472,N_8502,N_7363);
nor U14473 (N_14473,N_5605,N_6886);
and U14474 (N_14474,N_6255,N_9326);
nand U14475 (N_14475,N_5613,N_8910);
xnor U14476 (N_14476,N_6850,N_7746);
or U14477 (N_14477,N_9513,N_8375);
nor U14478 (N_14478,N_9002,N_5163);
and U14479 (N_14479,N_5068,N_6363);
and U14480 (N_14480,N_6684,N_9419);
or U14481 (N_14481,N_9075,N_8164);
or U14482 (N_14482,N_9775,N_9818);
or U14483 (N_14483,N_6049,N_6915);
nand U14484 (N_14484,N_5360,N_8099);
nand U14485 (N_14485,N_9642,N_9944);
or U14486 (N_14486,N_7078,N_7573);
and U14487 (N_14487,N_9132,N_5711);
nand U14488 (N_14488,N_5174,N_8576);
nand U14489 (N_14489,N_7211,N_8968);
nor U14490 (N_14490,N_9574,N_7965);
xor U14491 (N_14491,N_7489,N_8017);
and U14492 (N_14492,N_7803,N_9441);
or U14493 (N_14493,N_5290,N_5782);
xnor U14494 (N_14494,N_9737,N_5674);
xnor U14495 (N_14495,N_9224,N_6188);
nor U14496 (N_14496,N_9378,N_9855);
xor U14497 (N_14497,N_8694,N_6936);
xnor U14498 (N_14498,N_8492,N_8147);
xor U14499 (N_14499,N_8783,N_9236);
xor U14500 (N_14500,N_6707,N_9033);
xnor U14501 (N_14501,N_7771,N_9376);
or U14502 (N_14502,N_5779,N_8987);
xor U14503 (N_14503,N_7585,N_9130);
nand U14504 (N_14504,N_7114,N_9908);
nand U14505 (N_14505,N_6682,N_8367);
nand U14506 (N_14506,N_6501,N_5220);
nor U14507 (N_14507,N_9927,N_9318);
nand U14508 (N_14508,N_8271,N_9279);
or U14509 (N_14509,N_5867,N_9940);
xnor U14510 (N_14510,N_7181,N_8496);
nand U14511 (N_14511,N_5012,N_9234);
or U14512 (N_14512,N_5327,N_7025);
and U14513 (N_14513,N_9470,N_7573);
nor U14514 (N_14514,N_5556,N_7575);
xor U14515 (N_14515,N_7251,N_8090);
xor U14516 (N_14516,N_6945,N_6457);
nand U14517 (N_14517,N_9635,N_6516);
and U14518 (N_14518,N_5219,N_9498);
nor U14519 (N_14519,N_5381,N_5013);
nand U14520 (N_14520,N_5467,N_5310);
nand U14521 (N_14521,N_6311,N_6213);
xnor U14522 (N_14522,N_5414,N_5484);
xnor U14523 (N_14523,N_5710,N_9324);
or U14524 (N_14524,N_6572,N_5146);
nand U14525 (N_14525,N_5485,N_6385);
xnor U14526 (N_14526,N_7698,N_7063);
nand U14527 (N_14527,N_5069,N_5432);
xor U14528 (N_14528,N_8903,N_7350);
nand U14529 (N_14529,N_7738,N_9860);
nand U14530 (N_14530,N_5381,N_6674);
and U14531 (N_14531,N_8144,N_5125);
xor U14532 (N_14532,N_9144,N_7386);
and U14533 (N_14533,N_6645,N_9667);
xor U14534 (N_14534,N_7223,N_7712);
xor U14535 (N_14535,N_5493,N_7676);
nand U14536 (N_14536,N_5510,N_6702);
or U14537 (N_14537,N_8710,N_9848);
nor U14538 (N_14538,N_9411,N_5691);
nor U14539 (N_14539,N_6448,N_6563);
nor U14540 (N_14540,N_8233,N_7487);
nor U14541 (N_14541,N_6400,N_8629);
nand U14542 (N_14542,N_9687,N_5919);
or U14543 (N_14543,N_9109,N_8005);
xnor U14544 (N_14544,N_9449,N_5586);
or U14545 (N_14545,N_7167,N_7278);
nor U14546 (N_14546,N_6039,N_7908);
and U14547 (N_14547,N_8842,N_7938);
and U14548 (N_14548,N_7232,N_5054);
nand U14549 (N_14549,N_9474,N_9842);
or U14550 (N_14550,N_7122,N_7414);
xor U14551 (N_14551,N_6914,N_9617);
xor U14552 (N_14552,N_7266,N_6206);
nand U14553 (N_14553,N_9237,N_7622);
or U14554 (N_14554,N_5213,N_8584);
and U14555 (N_14555,N_6282,N_5567);
nand U14556 (N_14556,N_7381,N_5828);
xnor U14557 (N_14557,N_6876,N_7306);
xor U14558 (N_14558,N_7625,N_6117);
and U14559 (N_14559,N_5777,N_9837);
nor U14560 (N_14560,N_5498,N_6362);
nor U14561 (N_14561,N_9344,N_9621);
and U14562 (N_14562,N_8604,N_5444);
or U14563 (N_14563,N_7620,N_9999);
or U14564 (N_14564,N_9599,N_7854);
or U14565 (N_14565,N_7085,N_7368);
nand U14566 (N_14566,N_5950,N_6333);
nand U14567 (N_14567,N_9349,N_7578);
and U14568 (N_14568,N_5551,N_7009);
xnor U14569 (N_14569,N_9204,N_6554);
and U14570 (N_14570,N_5485,N_8000);
nor U14571 (N_14571,N_7023,N_5876);
and U14572 (N_14572,N_9488,N_8930);
or U14573 (N_14573,N_6834,N_8557);
xor U14574 (N_14574,N_7132,N_7526);
and U14575 (N_14575,N_7681,N_5176);
nand U14576 (N_14576,N_5310,N_9092);
xor U14577 (N_14577,N_5514,N_9533);
or U14578 (N_14578,N_8895,N_7105);
or U14579 (N_14579,N_6108,N_5535);
nor U14580 (N_14580,N_8920,N_5639);
and U14581 (N_14581,N_7680,N_6669);
nor U14582 (N_14582,N_6426,N_5215);
or U14583 (N_14583,N_5372,N_5956);
or U14584 (N_14584,N_7954,N_8493);
and U14585 (N_14585,N_9840,N_5847);
nor U14586 (N_14586,N_9620,N_9837);
nor U14587 (N_14587,N_9555,N_8122);
or U14588 (N_14588,N_5835,N_5359);
nand U14589 (N_14589,N_7850,N_8458);
or U14590 (N_14590,N_8893,N_9183);
nor U14591 (N_14591,N_8445,N_5044);
nand U14592 (N_14592,N_8288,N_8553);
and U14593 (N_14593,N_9248,N_9012);
or U14594 (N_14594,N_5593,N_5043);
xnor U14595 (N_14595,N_8138,N_9457);
nor U14596 (N_14596,N_9667,N_7359);
xor U14597 (N_14597,N_7195,N_5027);
nand U14598 (N_14598,N_5779,N_9229);
nand U14599 (N_14599,N_7606,N_8074);
and U14600 (N_14600,N_6114,N_9212);
and U14601 (N_14601,N_7716,N_8358);
or U14602 (N_14602,N_6330,N_6705);
nor U14603 (N_14603,N_9635,N_7306);
or U14604 (N_14604,N_5996,N_9227);
nand U14605 (N_14605,N_8683,N_5297);
and U14606 (N_14606,N_9640,N_8623);
and U14607 (N_14607,N_7193,N_8469);
nor U14608 (N_14608,N_6483,N_7387);
nand U14609 (N_14609,N_5364,N_6265);
xor U14610 (N_14610,N_8249,N_5674);
nor U14611 (N_14611,N_8545,N_8838);
nand U14612 (N_14612,N_8471,N_5230);
or U14613 (N_14613,N_7759,N_7275);
nor U14614 (N_14614,N_5800,N_8331);
or U14615 (N_14615,N_9743,N_5804);
and U14616 (N_14616,N_9988,N_8649);
nor U14617 (N_14617,N_6084,N_5236);
and U14618 (N_14618,N_6915,N_8383);
nand U14619 (N_14619,N_7426,N_9571);
or U14620 (N_14620,N_7536,N_7766);
nor U14621 (N_14621,N_5212,N_9656);
and U14622 (N_14622,N_6192,N_6483);
or U14623 (N_14623,N_9233,N_9259);
nor U14624 (N_14624,N_8401,N_6453);
xnor U14625 (N_14625,N_7769,N_9814);
and U14626 (N_14626,N_9090,N_6132);
nand U14627 (N_14627,N_6753,N_9393);
or U14628 (N_14628,N_6053,N_6630);
and U14629 (N_14629,N_7587,N_7121);
nor U14630 (N_14630,N_9804,N_6119);
xnor U14631 (N_14631,N_7501,N_9363);
nand U14632 (N_14632,N_9298,N_6100);
nand U14633 (N_14633,N_8328,N_7430);
xnor U14634 (N_14634,N_5576,N_5906);
and U14635 (N_14635,N_9862,N_9706);
xor U14636 (N_14636,N_6909,N_8880);
xnor U14637 (N_14637,N_7922,N_5690);
xor U14638 (N_14638,N_8627,N_8232);
or U14639 (N_14639,N_9115,N_6006);
nand U14640 (N_14640,N_8527,N_5461);
nand U14641 (N_14641,N_8117,N_7201);
nand U14642 (N_14642,N_7039,N_8027);
and U14643 (N_14643,N_9072,N_7358);
or U14644 (N_14644,N_5087,N_8645);
nand U14645 (N_14645,N_8372,N_7360);
nor U14646 (N_14646,N_7160,N_6790);
or U14647 (N_14647,N_7185,N_8834);
and U14648 (N_14648,N_6813,N_6234);
or U14649 (N_14649,N_5925,N_9975);
xor U14650 (N_14650,N_9755,N_5949);
xor U14651 (N_14651,N_7691,N_8511);
and U14652 (N_14652,N_9185,N_5854);
or U14653 (N_14653,N_8408,N_7650);
and U14654 (N_14654,N_8274,N_7839);
nor U14655 (N_14655,N_5362,N_5093);
nand U14656 (N_14656,N_7477,N_5515);
nand U14657 (N_14657,N_7428,N_9979);
nand U14658 (N_14658,N_7081,N_9787);
xnor U14659 (N_14659,N_9120,N_9465);
nand U14660 (N_14660,N_5628,N_6388);
or U14661 (N_14661,N_7857,N_6866);
xor U14662 (N_14662,N_6927,N_9236);
nand U14663 (N_14663,N_5988,N_7292);
xor U14664 (N_14664,N_9143,N_5434);
nor U14665 (N_14665,N_6969,N_8775);
or U14666 (N_14666,N_9133,N_8471);
xor U14667 (N_14667,N_6206,N_7753);
nor U14668 (N_14668,N_7427,N_6114);
or U14669 (N_14669,N_9503,N_8165);
nor U14670 (N_14670,N_8358,N_9806);
xnor U14671 (N_14671,N_9266,N_9801);
and U14672 (N_14672,N_9469,N_8049);
xnor U14673 (N_14673,N_9750,N_9568);
nor U14674 (N_14674,N_9657,N_7968);
xnor U14675 (N_14675,N_7424,N_7773);
nor U14676 (N_14676,N_9800,N_6988);
nor U14677 (N_14677,N_5957,N_7265);
or U14678 (N_14678,N_5345,N_5215);
and U14679 (N_14679,N_6071,N_6576);
or U14680 (N_14680,N_5310,N_5672);
xnor U14681 (N_14681,N_5739,N_7210);
and U14682 (N_14682,N_8003,N_8758);
or U14683 (N_14683,N_5856,N_9990);
nor U14684 (N_14684,N_5430,N_8798);
nor U14685 (N_14685,N_5641,N_7506);
or U14686 (N_14686,N_9478,N_8915);
xnor U14687 (N_14687,N_6715,N_6144);
xor U14688 (N_14688,N_6876,N_5857);
nand U14689 (N_14689,N_7464,N_8733);
or U14690 (N_14690,N_6825,N_8969);
and U14691 (N_14691,N_7127,N_5575);
nor U14692 (N_14692,N_8331,N_6702);
xor U14693 (N_14693,N_6397,N_8264);
xnor U14694 (N_14694,N_8252,N_8269);
xnor U14695 (N_14695,N_5138,N_6520);
or U14696 (N_14696,N_8895,N_8843);
and U14697 (N_14697,N_6296,N_8549);
or U14698 (N_14698,N_5285,N_6955);
or U14699 (N_14699,N_6711,N_7049);
and U14700 (N_14700,N_5414,N_8124);
or U14701 (N_14701,N_8510,N_7982);
or U14702 (N_14702,N_7325,N_5845);
nor U14703 (N_14703,N_8472,N_7355);
nor U14704 (N_14704,N_7662,N_6420);
nor U14705 (N_14705,N_8988,N_6752);
nand U14706 (N_14706,N_5614,N_7033);
or U14707 (N_14707,N_7139,N_8787);
and U14708 (N_14708,N_8042,N_8611);
and U14709 (N_14709,N_5003,N_8182);
and U14710 (N_14710,N_9226,N_5574);
or U14711 (N_14711,N_7298,N_9470);
xor U14712 (N_14712,N_9337,N_6891);
or U14713 (N_14713,N_5130,N_7499);
nor U14714 (N_14714,N_9248,N_8968);
xnor U14715 (N_14715,N_6703,N_7830);
nor U14716 (N_14716,N_9348,N_8685);
and U14717 (N_14717,N_8321,N_8327);
nand U14718 (N_14718,N_9381,N_5811);
nor U14719 (N_14719,N_8716,N_5745);
and U14720 (N_14720,N_5793,N_9264);
nor U14721 (N_14721,N_5732,N_8867);
nor U14722 (N_14722,N_7451,N_7025);
nor U14723 (N_14723,N_8987,N_5416);
nor U14724 (N_14724,N_9731,N_6035);
or U14725 (N_14725,N_7576,N_6954);
xnor U14726 (N_14726,N_7351,N_7763);
nor U14727 (N_14727,N_9391,N_9876);
nor U14728 (N_14728,N_9562,N_7783);
nand U14729 (N_14729,N_8642,N_5593);
xor U14730 (N_14730,N_7861,N_7368);
nand U14731 (N_14731,N_5446,N_8340);
nand U14732 (N_14732,N_9969,N_8283);
xnor U14733 (N_14733,N_6089,N_5223);
or U14734 (N_14734,N_6614,N_5757);
and U14735 (N_14735,N_8294,N_7979);
or U14736 (N_14736,N_9423,N_7104);
nand U14737 (N_14737,N_5536,N_9219);
xor U14738 (N_14738,N_5901,N_9080);
nand U14739 (N_14739,N_8418,N_5621);
xnor U14740 (N_14740,N_6196,N_8004);
nand U14741 (N_14741,N_8747,N_8498);
xor U14742 (N_14742,N_9600,N_9244);
or U14743 (N_14743,N_7311,N_9771);
or U14744 (N_14744,N_7650,N_8584);
xnor U14745 (N_14745,N_7850,N_6988);
or U14746 (N_14746,N_7937,N_9633);
nor U14747 (N_14747,N_6310,N_9210);
nand U14748 (N_14748,N_9139,N_6349);
nand U14749 (N_14749,N_9204,N_5132);
xnor U14750 (N_14750,N_9187,N_6660);
or U14751 (N_14751,N_6650,N_7084);
or U14752 (N_14752,N_5077,N_7485);
xor U14753 (N_14753,N_7953,N_5015);
nor U14754 (N_14754,N_9862,N_5763);
and U14755 (N_14755,N_8045,N_7170);
and U14756 (N_14756,N_7792,N_9890);
and U14757 (N_14757,N_9613,N_6683);
nor U14758 (N_14758,N_7134,N_6157);
nor U14759 (N_14759,N_8529,N_6105);
and U14760 (N_14760,N_5137,N_8198);
xnor U14761 (N_14761,N_7135,N_7647);
xnor U14762 (N_14762,N_7997,N_8130);
nand U14763 (N_14763,N_8582,N_7346);
nand U14764 (N_14764,N_5265,N_8891);
nor U14765 (N_14765,N_8791,N_7968);
and U14766 (N_14766,N_5542,N_8465);
nand U14767 (N_14767,N_7944,N_9706);
and U14768 (N_14768,N_5599,N_7582);
nand U14769 (N_14769,N_6851,N_6939);
and U14770 (N_14770,N_6565,N_7732);
xnor U14771 (N_14771,N_5462,N_5710);
nor U14772 (N_14772,N_7997,N_8159);
nand U14773 (N_14773,N_6713,N_5923);
and U14774 (N_14774,N_5126,N_6817);
xnor U14775 (N_14775,N_6579,N_8072);
nor U14776 (N_14776,N_5004,N_5215);
xnor U14777 (N_14777,N_8765,N_7327);
and U14778 (N_14778,N_6407,N_9805);
nand U14779 (N_14779,N_8201,N_6245);
and U14780 (N_14780,N_5702,N_6674);
nand U14781 (N_14781,N_5025,N_8703);
and U14782 (N_14782,N_5978,N_7376);
nand U14783 (N_14783,N_6347,N_5218);
xor U14784 (N_14784,N_9825,N_8176);
xor U14785 (N_14785,N_6384,N_8923);
nand U14786 (N_14786,N_6491,N_6110);
or U14787 (N_14787,N_5775,N_8459);
nand U14788 (N_14788,N_8718,N_7837);
or U14789 (N_14789,N_7521,N_7920);
nor U14790 (N_14790,N_7503,N_8351);
and U14791 (N_14791,N_6177,N_8671);
or U14792 (N_14792,N_7915,N_5666);
and U14793 (N_14793,N_9451,N_7077);
nor U14794 (N_14794,N_5631,N_9331);
nand U14795 (N_14795,N_6583,N_9893);
and U14796 (N_14796,N_8379,N_6733);
xnor U14797 (N_14797,N_5736,N_6648);
xnor U14798 (N_14798,N_9127,N_9435);
and U14799 (N_14799,N_8686,N_5475);
nor U14800 (N_14800,N_6748,N_7566);
nand U14801 (N_14801,N_7746,N_6645);
xnor U14802 (N_14802,N_6615,N_6765);
or U14803 (N_14803,N_9878,N_6182);
nor U14804 (N_14804,N_9181,N_7190);
nor U14805 (N_14805,N_5200,N_5203);
nand U14806 (N_14806,N_8445,N_6202);
nor U14807 (N_14807,N_8955,N_8674);
or U14808 (N_14808,N_6164,N_7569);
and U14809 (N_14809,N_7633,N_7920);
xnor U14810 (N_14810,N_8202,N_8169);
and U14811 (N_14811,N_5064,N_6295);
xnor U14812 (N_14812,N_7037,N_8807);
and U14813 (N_14813,N_7682,N_7358);
or U14814 (N_14814,N_6680,N_6604);
or U14815 (N_14815,N_8999,N_6469);
nand U14816 (N_14816,N_9066,N_6207);
xor U14817 (N_14817,N_9816,N_9538);
and U14818 (N_14818,N_8333,N_7567);
and U14819 (N_14819,N_5052,N_6848);
and U14820 (N_14820,N_5401,N_8957);
or U14821 (N_14821,N_9388,N_7959);
nand U14822 (N_14822,N_8686,N_8710);
xor U14823 (N_14823,N_5485,N_9505);
xor U14824 (N_14824,N_9397,N_9823);
and U14825 (N_14825,N_7932,N_9770);
or U14826 (N_14826,N_5571,N_8156);
nor U14827 (N_14827,N_9070,N_6704);
xnor U14828 (N_14828,N_5920,N_6805);
nor U14829 (N_14829,N_6139,N_5944);
nand U14830 (N_14830,N_6864,N_8617);
nor U14831 (N_14831,N_9641,N_5070);
nand U14832 (N_14832,N_8853,N_6354);
xnor U14833 (N_14833,N_7624,N_8060);
nand U14834 (N_14834,N_8535,N_6726);
nand U14835 (N_14835,N_8801,N_5877);
nor U14836 (N_14836,N_6061,N_7781);
xor U14837 (N_14837,N_5586,N_7985);
nand U14838 (N_14838,N_8249,N_9003);
or U14839 (N_14839,N_8980,N_7922);
xor U14840 (N_14840,N_9997,N_9386);
nor U14841 (N_14841,N_5655,N_6585);
or U14842 (N_14842,N_6968,N_5254);
and U14843 (N_14843,N_9888,N_7865);
or U14844 (N_14844,N_9584,N_7138);
or U14845 (N_14845,N_7677,N_5308);
nor U14846 (N_14846,N_7301,N_9542);
xnor U14847 (N_14847,N_6412,N_6004);
and U14848 (N_14848,N_8171,N_8411);
and U14849 (N_14849,N_7179,N_5897);
nand U14850 (N_14850,N_8913,N_8503);
xnor U14851 (N_14851,N_6330,N_7966);
xor U14852 (N_14852,N_6741,N_6263);
or U14853 (N_14853,N_8481,N_5024);
xor U14854 (N_14854,N_7092,N_5147);
and U14855 (N_14855,N_9095,N_8572);
or U14856 (N_14856,N_7262,N_5484);
nor U14857 (N_14857,N_8120,N_5165);
xor U14858 (N_14858,N_5125,N_9804);
nor U14859 (N_14859,N_6030,N_8473);
nor U14860 (N_14860,N_7011,N_6895);
nand U14861 (N_14861,N_9450,N_8530);
or U14862 (N_14862,N_9239,N_8924);
nand U14863 (N_14863,N_8926,N_9981);
or U14864 (N_14864,N_6804,N_9798);
nor U14865 (N_14865,N_9640,N_8625);
nand U14866 (N_14866,N_8413,N_9959);
xor U14867 (N_14867,N_6540,N_5628);
xor U14868 (N_14868,N_5238,N_8998);
or U14869 (N_14869,N_8997,N_7949);
xnor U14870 (N_14870,N_5125,N_8278);
nor U14871 (N_14871,N_5251,N_5333);
and U14872 (N_14872,N_7279,N_8054);
nor U14873 (N_14873,N_9738,N_6586);
nor U14874 (N_14874,N_5263,N_8058);
xor U14875 (N_14875,N_5993,N_9881);
nand U14876 (N_14876,N_7421,N_8566);
and U14877 (N_14877,N_7223,N_9649);
or U14878 (N_14878,N_6584,N_9150);
nor U14879 (N_14879,N_8675,N_6233);
nor U14880 (N_14880,N_5428,N_7318);
xor U14881 (N_14881,N_6353,N_6612);
xor U14882 (N_14882,N_5960,N_5831);
and U14883 (N_14883,N_5429,N_7383);
xor U14884 (N_14884,N_6541,N_9956);
and U14885 (N_14885,N_6453,N_9636);
nand U14886 (N_14886,N_5994,N_7149);
and U14887 (N_14887,N_9064,N_6760);
nor U14888 (N_14888,N_9840,N_7345);
or U14889 (N_14889,N_7107,N_5392);
or U14890 (N_14890,N_8097,N_8120);
and U14891 (N_14891,N_8336,N_8459);
nor U14892 (N_14892,N_6475,N_5218);
xor U14893 (N_14893,N_5280,N_6531);
and U14894 (N_14894,N_9051,N_8186);
nor U14895 (N_14895,N_7320,N_7621);
xnor U14896 (N_14896,N_8269,N_6079);
xnor U14897 (N_14897,N_5132,N_8631);
or U14898 (N_14898,N_7564,N_6259);
nand U14899 (N_14899,N_8743,N_7153);
and U14900 (N_14900,N_8470,N_7841);
xnor U14901 (N_14901,N_7735,N_5498);
nand U14902 (N_14902,N_8177,N_8597);
or U14903 (N_14903,N_6936,N_5542);
nor U14904 (N_14904,N_8320,N_8849);
or U14905 (N_14905,N_8244,N_5378);
and U14906 (N_14906,N_8514,N_7823);
and U14907 (N_14907,N_8628,N_8746);
xor U14908 (N_14908,N_8172,N_9123);
and U14909 (N_14909,N_8397,N_6767);
and U14910 (N_14910,N_7191,N_5933);
and U14911 (N_14911,N_7591,N_8659);
nand U14912 (N_14912,N_5409,N_9328);
xor U14913 (N_14913,N_6644,N_5107);
xnor U14914 (N_14914,N_9211,N_5628);
or U14915 (N_14915,N_6778,N_7837);
nand U14916 (N_14916,N_5438,N_8419);
or U14917 (N_14917,N_6687,N_8991);
xor U14918 (N_14918,N_9336,N_8419);
or U14919 (N_14919,N_6234,N_8739);
or U14920 (N_14920,N_5086,N_6851);
nor U14921 (N_14921,N_9733,N_8041);
nand U14922 (N_14922,N_6833,N_9013);
and U14923 (N_14923,N_7964,N_6643);
and U14924 (N_14924,N_9537,N_9072);
xor U14925 (N_14925,N_6700,N_5872);
nand U14926 (N_14926,N_8510,N_8788);
and U14927 (N_14927,N_5466,N_5200);
nor U14928 (N_14928,N_5056,N_6614);
or U14929 (N_14929,N_7297,N_9476);
xnor U14930 (N_14930,N_5983,N_8259);
nand U14931 (N_14931,N_6177,N_5461);
and U14932 (N_14932,N_5687,N_6458);
and U14933 (N_14933,N_9254,N_9605);
and U14934 (N_14934,N_6966,N_7441);
or U14935 (N_14935,N_9751,N_6145);
nor U14936 (N_14936,N_6151,N_6812);
or U14937 (N_14937,N_8104,N_7347);
and U14938 (N_14938,N_8442,N_9029);
xor U14939 (N_14939,N_5777,N_7610);
or U14940 (N_14940,N_8234,N_8779);
nand U14941 (N_14941,N_7271,N_6696);
and U14942 (N_14942,N_8672,N_6355);
and U14943 (N_14943,N_7555,N_5199);
or U14944 (N_14944,N_9166,N_8339);
xor U14945 (N_14945,N_8850,N_5613);
nand U14946 (N_14946,N_8450,N_7312);
or U14947 (N_14947,N_8750,N_8275);
nand U14948 (N_14948,N_8188,N_7499);
nand U14949 (N_14949,N_5408,N_7016);
xor U14950 (N_14950,N_5893,N_5016);
nand U14951 (N_14951,N_7666,N_8572);
nor U14952 (N_14952,N_5216,N_8924);
nand U14953 (N_14953,N_8116,N_7013);
xor U14954 (N_14954,N_9433,N_9547);
nor U14955 (N_14955,N_6154,N_6508);
and U14956 (N_14956,N_6614,N_9708);
xor U14957 (N_14957,N_9313,N_9587);
and U14958 (N_14958,N_6002,N_8475);
and U14959 (N_14959,N_8151,N_6325);
nand U14960 (N_14960,N_7643,N_7892);
or U14961 (N_14961,N_8819,N_8795);
nand U14962 (N_14962,N_5206,N_6355);
and U14963 (N_14963,N_6940,N_7183);
and U14964 (N_14964,N_7459,N_8176);
nor U14965 (N_14965,N_8460,N_5792);
nand U14966 (N_14966,N_7073,N_9652);
or U14967 (N_14967,N_9512,N_9330);
nor U14968 (N_14968,N_6077,N_8464);
and U14969 (N_14969,N_5333,N_9877);
nand U14970 (N_14970,N_5746,N_9733);
or U14971 (N_14971,N_8601,N_8032);
nor U14972 (N_14972,N_7310,N_5883);
or U14973 (N_14973,N_7666,N_6702);
or U14974 (N_14974,N_8884,N_5247);
or U14975 (N_14975,N_8122,N_7232);
or U14976 (N_14976,N_5828,N_9812);
nor U14977 (N_14977,N_8500,N_7040);
or U14978 (N_14978,N_6593,N_9246);
nor U14979 (N_14979,N_6175,N_5777);
and U14980 (N_14980,N_9311,N_9933);
and U14981 (N_14981,N_9358,N_5451);
nor U14982 (N_14982,N_6276,N_6713);
or U14983 (N_14983,N_7181,N_6175);
and U14984 (N_14984,N_9110,N_7300);
xor U14985 (N_14985,N_8140,N_8432);
nor U14986 (N_14986,N_9541,N_5408);
or U14987 (N_14987,N_5135,N_9213);
nand U14988 (N_14988,N_6469,N_6053);
and U14989 (N_14989,N_5772,N_8712);
nand U14990 (N_14990,N_7897,N_5102);
nor U14991 (N_14991,N_5186,N_5107);
xnor U14992 (N_14992,N_7648,N_8036);
nor U14993 (N_14993,N_7639,N_6101);
nor U14994 (N_14994,N_7537,N_8501);
nand U14995 (N_14995,N_6870,N_6664);
nand U14996 (N_14996,N_7719,N_5866);
and U14997 (N_14997,N_8143,N_5322);
xor U14998 (N_14998,N_9486,N_5699);
nand U14999 (N_14999,N_6100,N_5310);
or U15000 (N_15000,N_10104,N_11686);
xnor U15001 (N_15001,N_10077,N_13874);
xor U15002 (N_15002,N_10510,N_12746);
nand U15003 (N_15003,N_10953,N_12547);
or U15004 (N_15004,N_13541,N_10625);
nor U15005 (N_15005,N_11627,N_12026);
and U15006 (N_15006,N_13170,N_10554);
nor U15007 (N_15007,N_11073,N_13726);
or U15008 (N_15008,N_13760,N_11313);
and U15009 (N_15009,N_14058,N_11661);
and U15010 (N_15010,N_10846,N_11954);
xnor U15011 (N_15011,N_12677,N_10025);
and U15012 (N_15012,N_11936,N_11221);
xnor U15013 (N_15013,N_13941,N_13552);
nand U15014 (N_15014,N_12024,N_13278);
xor U15015 (N_15015,N_13100,N_14368);
nand U15016 (N_15016,N_14796,N_10733);
nor U15017 (N_15017,N_10518,N_12501);
nand U15018 (N_15018,N_10843,N_12496);
nand U15019 (N_15019,N_13472,N_10722);
nand U15020 (N_15020,N_12940,N_12436);
or U15021 (N_15021,N_13297,N_13818);
nor U15022 (N_15022,N_10563,N_13669);
xor U15023 (N_15023,N_10167,N_13822);
and U15024 (N_15024,N_11135,N_10052);
nor U15025 (N_15025,N_12250,N_12080);
or U15026 (N_15026,N_10443,N_14181);
or U15027 (N_15027,N_13057,N_14698);
or U15028 (N_15028,N_10979,N_12423);
and U15029 (N_15029,N_12405,N_11437);
nor U15030 (N_15030,N_10417,N_13590);
nand U15031 (N_15031,N_13881,N_11605);
xnor U15032 (N_15032,N_14697,N_13475);
or U15033 (N_15033,N_13602,N_12088);
xnor U15034 (N_15034,N_10248,N_12899);
nand U15035 (N_15035,N_12188,N_11214);
nor U15036 (N_15036,N_10924,N_12415);
and U15037 (N_15037,N_13606,N_12615);
xnor U15038 (N_15038,N_11000,N_14134);
nor U15039 (N_15039,N_14535,N_10439);
nor U15040 (N_15040,N_12360,N_14382);
xnor U15041 (N_15041,N_11930,N_10683);
and U15042 (N_15042,N_11011,N_14105);
xor U15043 (N_15043,N_14933,N_11600);
or U15044 (N_15044,N_12785,N_12097);
xnor U15045 (N_15045,N_13832,N_14706);
nand U15046 (N_15046,N_12158,N_13488);
nand U15047 (N_15047,N_13579,N_10907);
xor U15048 (N_15048,N_12947,N_14527);
xor U15049 (N_15049,N_13696,N_14829);
and U15050 (N_15050,N_10801,N_12101);
and U15051 (N_15051,N_12379,N_10111);
and U15052 (N_15052,N_14956,N_11840);
xor U15053 (N_15053,N_10365,N_12675);
or U15054 (N_15054,N_11341,N_11929);
and U15055 (N_15055,N_13289,N_11610);
nand U15056 (N_15056,N_11050,N_10824);
nand U15057 (N_15057,N_14056,N_10731);
xnor U15058 (N_15058,N_12914,N_13477);
xor U15059 (N_15059,N_12492,N_14863);
xor U15060 (N_15060,N_11459,N_13718);
xor U15061 (N_15061,N_13225,N_10705);
nor U15062 (N_15062,N_13582,N_14961);
and U15063 (N_15063,N_14051,N_14823);
xnor U15064 (N_15064,N_13308,N_10962);
xnor U15065 (N_15065,N_12511,N_10550);
or U15066 (N_15066,N_11647,N_10274);
nor U15067 (N_15067,N_13447,N_12148);
or U15068 (N_15068,N_10957,N_11898);
and U15069 (N_15069,N_11263,N_12513);
xnor U15070 (N_15070,N_14436,N_10287);
nor U15071 (N_15071,N_14252,N_12794);
and U15072 (N_15072,N_10549,N_12350);
nor U15073 (N_15073,N_13305,N_10746);
xnor U15074 (N_15074,N_11753,N_13430);
nor U15075 (N_15075,N_10454,N_10551);
nor U15076 (N_15076,N_14532,N_13844);
or U15077 (N_15077,N_10292,N_12397);
nor U15078 (N_15078,N_14544,N_12082);
and U15079 (N_15079,N_13895,N_11968);
or U15080 (N_15080,N_13827,N_13019);
nor U15081 (N_15081,N_10122,N_10372);
or U15082 (N_15082,N_12988,N_13262);
nand U15083 (N_15083,N_10301,N_11177);
nand U15084 (N_15084,N_10994,N_10164);
and U15085 (N_15085,N_10017,N_12728);
xor U15086 (N_15086,N_13834,N_10349);
and U15087 (N_15087,N_11714,N_12392);
and U15088 (N_15088,N_14695,N_10908);
nand U15089 (N_15089,N_10078,N_14007);
and U15090 (N_15090,N_14414,N_10968);
and U15091 (N_15091,N_14239,N_12506);
or U15092 (N_15092,N_14472,N_10158);
or U15093 (N_15093,N_12441,N_14700);
nor U15094 (N_15094,N_11159,N_13872);
and U15095 (N_15095,N_12731,N_11513);
or U15096 (N_15096,N_12171,N_14490);
and U15097 (N_15097,N_13087,N_12018);
and U15098 (N_15098,N_12901,N_11343);
or U15099 (N_15099,N_12775,N_13588);
or U15100 (N_15100,N_11624,N_10720);
nand U15101 (N_15101,N_14495,N_12235);
nand U15102 (N_15102,N_14144,N_12470);
or U15103 (N_15103,N_11414,N_12937);
nor U15104 (N_15104,N_11407,N_10727);
and U15105 (N_15105,N_12889,N_13415);
or U15106 (N_15106,N_14468,N_10304);
xnor U15107 (N_15107,N_14445,N_13528);
nor U15108 (N_15108,N_14627,N_13794);
or U15109 (N_15109,N_11326,N_13049);
nand U15110 (N_15110,N_10666,N_14882);
or U15111 (N_15111,N_11759,N_11470);
xor U15112 (N_15112,N_11917,N_12979);
nand U15113 (N_15113,N_10906,N_14206);
nand U15114 (N_15114,N_14210,N_12284);
and U15115 (N_15115,N_10461,N_11206);
nand U15116 (N_15116,N_14491,N_12252);
xor U15117 (N_15117,N_13843,N_13442);
nand U15118 (N_15118,N_13310,N_13445);
nand U15119 (N_15119,N_12334,N_12764);
nor U15120 (N_15120,N_14938,N_10305);
and U15121 (N_15121,N_13047,N_12231);
xor U15122 (N_15122,N_11504,N_13040);
nand U15123 (N_15123,N_13144,N_11815);
nor U15124 (N_15124,N_11888,N_12474);
nor U15125 (N_15125,N_13644,N_11473);
and U15126 (N_15126,N_11547,N_13763);
xor U15127 (N_15127,N_11290,N_10726);
or U15128 (N_15128,N_11350,N_13775);
and U15129 (N_15129,N_11429,N_14985);
xnor U15130 (N_15130,N_12568,N_10213);
or U15131 (N_15131,N_13348,N_14629);
and U15132 (N_15132,N_14519,N_14402);
xor U15133 (N_15133,N_11976,N_11531);
nand U15134 (N_15134,N_11562,N_12296);
and U15135 (N_15135,N_10343,N_10626);
nand U15136 (N_15136,N_14098,N_11544);
or U15137 (N_15137,N_12963,N_11995);
or U15138 (N_15138,N_13481,N_10141);
xnor U15139 (N_15139,N_14440,N_13373);
nand U15140 (N_15140,N_13234,N_11793);
xnor U15141 (N_15141,N_12907,N_10360);
or U15142 (N_15142,N_11446,N_13200);
and U15143 (N_15143,N_14477,N_11612);
or U15144 (N_15144,N_11814,N_13038);
nor U15145 (N_15145,N_13044,N_11994);
and U15146 (N_15146,N_11980,N_12569);
nor U15147 (N_15147,N_12434,N_12008);
and U15148 (N_15148,N_11822,N_11646);
or U15149 (N_15149,N_12555,N_11655);
nand U15150 (N_15150,N_12104,N_12461);
nand U15151 (N_15151,N_11409,N_14172);
and U15152 (N_15152,N_13386,N_10297);
and U15153 (N_15153,N_13292,N_11884);
and U15154 (N_15154,N_12773,N_14912);
and U15155 (N_15155,N_14903,N_14849);
nor U15156 (N_15156,N_10440,N_14996);
and U15157 (N_15157,N_14665,N_12673);
nor U15158 (N_15158,N_11498,N_12565);
and U15159 (N_15159,N_10136,N_10251);
nor U15160 (N_15160,N_14132,N_10790);
nor U15161 (N_15161,N_13746,N_10694);
or U15162 (N_15162,N_13111,N_14010);
or U15163 (N_15163,N_14222,N_11103);
or U15164 (N_15164,N_13615,N_11774);
xnor U15165 (N_15165,N_14501,N_11862);
nor U15166 (N_15166,N_10432,N_10816);
nor U15167 (N_15167,N_10434,N_11425);
xnor U15168 (N_15168,N_10112,N_11465);
or U15169 (N_15169,N_14958,N_12964);
nor U15170 (N_15170,N_12145,N_10307);
nand U15171 (N_15171,N_14773,N_11671);
and U15172 (N_15172,N_13989,N_13240);
or U15173 (N_15173,N_10878,N_13627);
or U15174 (N_15174,N_13565,N_12822);
and U15175 (N_15175,N_10364,N_11108);
nor U15176 (N_15176,N_14682,N_10817);
nand U15177 (N_15177,N_14974,N_14606);
and U15178 (N_15178,N_14777,N_11324);
and U15179 (N_15179,N_12955,N_14244);
or U15180 (N_15180,N_13126,N_13298);
nand U15181 (N_15181,N_13774,N_12078);
or U15182 (N_15182,N_11569,N_11376);
nand U15183 (N_15183,N_12226,N_14904);
or U15184 (N_15184,N_14536,N_10844);
and U15185 (N_15185,N_12759,N_12044);
xor U15186 (N_15186,N_13206,N_10565);
xor U15187 (N_15187,N_12227,N_12550);
nor U15188 (N_15188,N_14497,N_10330);
or U15189 (N_15189,N_10199,N_11144);
or U15190 (N_15190,N_12179,N_14167);
and U15191 (N_15191,N_12169,N_11915);
nor U15192 (N_15192,N_14048,N_11892);
nor U15193 (N_15193,N_12174,N_14135);
nor U15194 (N_15194,N_13825,N_12362);
and U15195 (N_15195,N_10665,N_13762);
xor U15196 (N_15196,N_10832,N_10766);
or U15197 (N_15197,N_14979,N_14474);
nand U15198 (N_15198,N_13016,N_12000);
nor U15199 (N_15199,N_10795,N_12049);
and U15200 (N_15200,N_12813,N_11070);
or U15201 (N_15201,N_12317,N_13913);
nor U15202 (N_15202,N_12753,N_10204);
or U15203 (N_15203,N_11743,N_14751);
or U15204 (N_15204,N_12529,N_14332);
nor U15205 (N_15205,N_13839,N_10103);
or U15206 (N_15206,N_14949,N_11101);
nor U15207 (N_15207,N_11467,N_10497);
nand U15208 (N_15208,N_12419,N_12274);
or U15209 (N_15209,N_12118,N_14290);
and U15210 (N_15210,N_12438,N_13396);
and U15211 (N_15211,N_11364,N_11777);
xnor U15212 (N_15212,N_13145,N_14537);
nor U15213 (N_15213,N_11720,N_14154);
or U15214 (N_15214,N_10948,N_12241);
or U15215 (N_15215,N_14826,N_10473);
and U15216 (N_15216,N_13227,N_13168);
and U15217 (N_15217,N_14584,N_10913);
or U15218 (N_15218,N_13522,N_12259);
and U15219 (N_15219,N_14935,N_10642);
nor U15220 (N_15220,N_14515,N_11817);
and U15221 (N_15221,N_12526,N_10211);
and U15222 (N_15222,N_10200,N_14592);
and U15223 (N_15223,N_14041,N_10259);
and U15224 (N_15224,N_14726,N_13000);
or U15225 (N_15225,N_11842,N_14412);
and U15226 (N_15226,N_11656,N_10262);
nand U15227 (N_15227,N_10714,N_13633);
nand U15228 (N_15228,N_14567,N_11054);
or U15229 (N_15229,N_12251,N_10300);
xnor U15230 (N_15230,N_11896,N_13360);
nand U15231 (N_15231,N_10560,N_13220);
xnor U15232 (N_15232,N_13248,N_11739);
or U15233 (N_15233,N_14800,N_14972);
and U15234 (N_15234,N_10427,N_13338);
and U15235 (N_15235,N_13609,N_12230);
nor U15236 (N_15236,N_10617,N_10171);
or U15237 (N_15237,N_14323,N_10866);
nand U15238 (N_15238,N_12404,N_12935);
and U15239 (N_15239,N_10992,N_11611);
nor U15240 (N_15240,N_12989,N_13328);
nor U15241 (N_15241,N_13621,N_10818);
or U15242 (N_15242,N_11044,N_14462);
or U15243 (N_15243,N_11676,N_13393);
and U15244 (N_15244,N_11440,N_13405);
or U15245 (N_15245,N_14867,N_13680);
xnor U15246 (N_15246,N_12696,N_11542);
nor U15247 (N_15247,N_11718,N_10785);
or U15248 (N_15248,N_12305,N_14464);
and U15249 (N_15249,N_10925,N_10138);
and U15250 (N_15250,N_11901,N_13083);
or U15251 (N_15251,N_13250,N_13722);
or U15252 (N_15252,N_10921,N_12195);
xnor U15253 (N_15253,N_10744,N_10387);
xor U15254 (N_15254,N_13517,N_14406);
nand U15255 (N_15255,N_12338,N_12817);
xnor U15256 (N_15256,N_10484,N_10008);
nor U15257 (N_15257,N_11525,N_14024);
xor U15258 (N_15258,N_10324,N_11348);
or U15259 (N_15259,N_10934,N_10657);
and U15260 (N_15260,N_12129,N_14730);
and U15261 (N_15261,N_14518,N_12146);
xor U15262 (N_15262,N_10511,N_11287);
nor U15263 (N_15263,N_12222,N_12875);
or U15264 (N_15264,N_12105,N_10615);
or U15265 (N_15265,N_14977,N_13189);
nand U15266 (N_15266,N_10055,N_12311);
or U15267 (N_15267,N_10202,N_12524);
and U15268 (N_15268,N_11468,N_10212);
nor U15269 (N_15269,N_13323,N_10910);
nand U15270 (N_15270,N_12545,N_12546);
nand U15271 (N_15271,N_14514,N_14159);
nand U15272 (N_15272,N_11795,N_11317);
nor U15273 (N_15273,N_10033,N_13431);
or U15274 (N_15274,N_11658,N_10827);
xnor U15275 (N_15275,N_13865,N_14469);
and U15276 (N_15276,N_11384,N_14200);
xnor U15277 (N_15277,N_11725,N_12803);
nor U15278 (N_15278,N_14423,N_14944);
nand U15279 (N_15279,N_11546,N_11450);
nor U15280 (N_15280,N_12054,N_13085);
or U15281 (N_15281,N_11941,N_10256);
nor U15282 (N_15282,N_11109,N_13318);
nand U15283 (N_15283,N_10736,N_12823);
nand U15284 (N_15284,N_13108,N_10688);
and U15285 (N_15285,N_11642,N_12318);
and U15286 (N_15286,N_14587,N_14643);
nand U15287 (N_15287,N_11204,N_10778);
xnor U15288 (N_15288,N_12688,N_10652);
or U15289 (N_15289,N_11186,N_11999);
and U15290 (N_15290,N_12059,N_12001);
nand U15291 (N_15291,N_12572,N_14272);
and U15292 (N_15292,N_11388,N_12356);
or U15293 (N_15293,N_10699,N_11367);
nand U15294 (N_15294,N_10205,N_13785);
and U15295 (N_15295,N_11768,N_12544);
and U15296 (N_15296,N_10955,N_10591);
or U15297 (N_15297,N_14182,N_13270);
nor U15298 (N_15298,N_14703,N_14088);
xnor U15299 (N_15299,N_11863,N_11675);
or U15300 (N_15300,N_14357,N_10228);
xnor U15301 (N_15301,N_13919,N_14043);
and U15302 (N_15302,N_11921,N_11758);
nand U15303 (N_15303,N_12936,N_12847);
xnor U15304 (N_15304,N_12647,N_12863);
and U15305 (N_15305,N_11229,N_13233);
or U15306 (N_15306,N_11230,N_14218);
or U15307 (N_15307,N_13909,N_14548);
nor U15308 (N_15308,N_11246,N_14451);
xor U15309 (N_15309,N_13420,N_14001);
and U15310 (N_15310,N_14969,N_11805);
nor U15311 (N_15311,N_10767,N_10054);
and U15312 (N_15312,N_13352,N_10933);
nand U15313 (N_15313,N_14114,N_13790);
and U15314 (N_15314,N_12004,N_14707);
or U15315 (N_15315,N_14008,N_10024);
and U15316 (N_15316,N_13836,N_11327);
xnor U15317 (N_15317,N_13283,N_13207);
or U15318 (N_15318,N_11620,N_10828);
and U15319 (N_15319,N_13559,N_13975);
and U15320 (N_15320,N_14087,N_14150);
or U15321 (N_15321,N_13901,N_11395);
or U15322 (N_15322,N_12225,N_11235);
nand U15323 (N_15323,N_12942,N_11811);
xnor U15324 (N_15324,N_12115,N_13162);
nor U15325 (N_15325,N_13315,N_13771);
nor U15326 (N_15326,N_12845,N_14022);
nor U15327 (N_15327,N_13056,N_10580);
and U15328 (N_15328,N_10275,N_12958);
and U15329 (N_15329,N_13698,N_12359);
or U15330 (N_15330,N_13346,N_10239);
nand U15331 (N_15331,N_10947,N_13211);
and U15332 (N_15332,N_11961,N_12483);
nand U15333 (N_15333,N_14420,N_10536);
and U15334 (N_15334,N_12207,N_10753);
or U15335 (N_15335,N_11847,N_13290);
xor U15336 (N_15336,N_10397,N_10232);
nand U15337 (N_15337,N_12915,N_10351);
or U15338 (N_15338,N_13251,N_12365);
xnor U15339 (N_15339,N_14786,N_14632);
nand U15340 (N_15340,N_13175,N_12437);
nand U15341 (N_15341,N_11571,N_10884);
nand U15342 (N_15342,N_14282,N_13706);
nand U15343 (N_15343,N_14261,N_12694);
or U15344 (N_15344,N_10875,N_11505);
and U15345 (N_15345,N_14214,N_13974);
or U15346 (N_15346,N_13084,N_14708);
or U15347 (N_15347,N_11812,N_10954);
xor U15348 (N_15348,N_10849,N_12442);
xor U15349 (N_15349,N_13473,N_14813);
or U15350 (N_15350,N_10203,N_13957);
xnor U15351 (N_15351,N_14724,N_10973);
and U15352 (N_15352,N_12194,N_11558);
nor U15353 (N_15353,N_12307,N_12690);
xnor U15354 (N_15354,N_12534,N_12751);
xor U15355 (N_15355,N_12313,N_11806);
nor U15356 (N_15356,N_13082,N_10574);
xor U15357 (N_15357,N_13092,N_13858);
and U15358 (N_15358,N_12611,N_11853);
xor U15359 (N_15359,N_12310,N_12454);
nand U15360 (N_15360,N_12142,N_13867);
nand U15361 (N_15361,N_14279,N_12765);
or U15362 (N_15362,N_11314,N_13601);
nand U15363 (N_15363,N_10247,N_13912);
xor U15364 (N_15364,N_12364,N_14669);
and U15365 (N_15365,N_13745,N_12416);
nand U15366 (N_15366,N_12384,N_10403);
or U15367 (N_15367,N_13167,N_12879);
nand U15368 (N_15368,N_12237,N_14943);
xnor U15369 (N_15369,N_10348,N_10697);
or U15370 (N_15370,N_12666,N_14783);
or U15371 (N_15371,N_10189,N_10916);
or U15372 (N_15372,N_10703,N_11088);
or U15373 (N_15373,N_14905,N_14756);
and U15374 (N_15374,N_10544,N_12363);
nand U15375 (N_15375,N_10476,N_10215);
xnor U15376 (N_15376,N_13375,N_12910);
or U15377 (N_15377,N_11706,N_10187);
nand U15378 (N_15378,N_11175,N_13112);
nor U15379 (N_15379,N_14557,N_13916);
xnor U15380 (N_15380,N_12209,N_11788);
or U15381 (N_15381,N_11514,N_12683);
nand U15382 (N_15382,N_12490,N_11443);
nor U15383 (N_15383,N_10852,N_14457);
nor U15384 (N_15384,N_12376,N_12025);
nand U15385 (N_15385,N_12370,N_12155);
and U15386 (N_15386,N_12922,N_10314);
and U15387 (N_15387,N_10378,N_10487);
nor U15388 (N_15388,N_10606,N_11248);
or U15389 (N_15389,N_14397,N_11110);
nand U15390 (N_15390,N_12090,N_13136);
nand U15391 (N_15391,N_13268,N_11277);
xnor U15392 (N_15392,N_13125,N_13221);
nor U15393 (N_15393,N_12917,N_14874);
nor U15394 (N_15394,N_10266,N_11020);
xnor U15395 (N_15395,N_14877,N_10972);
xor U15396 (N_15396,N_11259,N_12197);
nor U15397 (N_15397,N_12578,N_14338);
xnor U15398 (N_15398,N_11490,N_10963);
xor U15399 (N_15399,N_14674,N_13424);
and U15400 (N_15400,N_11267,N_13201);
or U15401 (N_15401,N_11920,N_14873);
xor U15402 (N_15402,N_13956,N_11978);
nor U15403 (N_15403,N_14269,N_10422);
and U15404 (N_15404,N_12684,N_14353);
or U15405 (N_15405,N_14216,N_10572);
and U15406 (N_15406,N_13392,N_12066);
xnor U15407 (N_15407,N_14932,N_14178);
nand U15408 (N_15408,N_11322,N_14115);
nand U15409 (N_15409,N_11712,N_13586);
nor U15410 (N_15410,N_13500,N_12238);
nand U15411 (N_15411,N_13443,N_14299);
xnor U15412 (N_15412,N_10867,N_13860);
nor U15413 (N_15413,N_14744,N_14914);
or U15414 (N_15414,N_12681,N_11986);
or U15415 (N_15415,N_12628,N_10177);
xor U15416 (N_15416,N_10649,N_12358);
nand U15417 (N_15417,N_10466,N_10858);
or U15418 (N_15418,N_10739,N_11126);
nor U15419 (N_15419,N_13725,N_11701);
and U15420 (N_15420,N_13151,N_14012);
nor U15421 (N_15421,N_14732,N_11782);
nor U15422 (N_15422,N_11055,N_12202);
or U15423 (N_15423,N_10418,N_12982);
xnor U15424 (N_15424,N_10861,N_11577);
xor U15425 (N_15425,N_12051,N_13324);
nor U15426 (N_15426,N_12626,N_10335);
nor U15427 (N_15427,N_11217,N_10964);
nor U15428 (N_15428,N_11197,N_14486);
xor U15429 (N_15429,N_10506,N_13705);
and U15430 (N_15430,N_10447,N_12554);
or U15431 (N_15431,N_14790,N_12131);
and U15432 (N_15432,N_12394,N_12399);
and U15433 (N_15433,N_12292,N_13793);
nand U15434 (N_15434,N_12232,N_13987);
nand U15435 (N_15435,N_13246,N_14550);
nor U15436 (N_15436,N_10173,N_10949);
nand U15437 (N_15437,N_10883,N_12645);
and U15438 (N_15438,N_10937,N_12872);
xor U15439 (N_15439,N_11066,N_10092);
xor U15440 (N_15440,N_13224,N_12806);
or U15441 (N_15441,N_12070,N_10429);
and U15442 (N_15442,N_13764,N_14696);
nor U15443 (N_15443,N_12272,N_13574);
xnor U15444 (N_15444,N_14298,N_14250);
and U15445 (N_15445,N_13700,N_13635);
nor U15446 (N_15446,N_10513,N_11802);
or U15447 (N_15447,N_11703,N_11825);
xnor U15448 (N_15448,N_10144,N_11821);
xnor U15449 (N_15449,N_10974,N_13026);
xnor U15450 (N_15450,N_11746,N_12596);
nor U15451 (N_15451,N_11303,N_12247);
nor U15452 (N_15452,N_12676,N_10456);
or U15453 (N_15453,N_14049,N_11633);
nand U15454 (N_15454,N_11306,N_10354);
nor U15455 (N_15455,N_12975,N_14089);
or U15456 (N_15456,N_10250,N_12289);
nand U15457 (N_15457,N_14666,N_14729);
and U15458 (N_15458,N_13469,N_12508);
nand U15459 (N_15459,N_10319,N_12199);
nor U15460 (N_15460,N_10441,N_11301);
nand U15461 (N_15461,N_10841,N_13630);
nor U15462 (N_15462,N_13846,N_10943);
or U15463 (N_15463,N_11184,N_13900);
xor U15464 (N_15464,N_12886,N_10556);
and U15465 (N_15465,N_13300,N_14163);
nor U15466 (N_15466,N_11028,N_14886);
nand U15467 (N_15467,N_11155,N_14765);
or U15468 (N_15468,N_13917,N_11724);
xnor U15469 (N_15469,N_12243,N_14547);
nand U15470 (N_15470,N_12353,N_12092);
nand U15471 (N_15471,N_14426,N_10303);
xor U15472 (N_15472,N_12750,N_10522);
nor U15473 (N_15473,N_10031,N_10263);
nand U15474 (N_15474,N_12481,N_12283);
or U15475 (N_15475,N_12099,N_10836);
nor U15476 (N_15476,N_12869,N_14915);
xnor U15477 (N_15477,N_11691,N_10600);
and U15478 (N_15478,N_10608,N_10481);
nor U15479 (N_15479,N_14395,N_13281);
nand U15480 (N_15480,N_13679,N_12498);
nor U15481 (N_15481,N_11438,N_12674);
nor U15482 (N_15482,N_10540,N_14663);
nand U15483 (N_15483,N_10107,N_12278);
nor U15484 (N_15484,N_11796,N_14066);
xnor U15485 (N_15485,N_12181,N_11697);
and U15486 (N_15486,N_14505,N_12154);
nor U15487 (N_15487,N_12956,N_13177);
nor U15488 (N_15488,N_13853,N_14750);
nand U15489 (N_15489,N_10339,N_14970);
nor U15490 (N_15490,N_12873,N_13952);
nor U15491 (N_15491,N_10759,N_14540);
nor U15492 (N_15492,N_13815,N_10571);
or U15493 (N_15493,N_12451,N_14975);
nor U15494 (N_15494,N_14122,N_13868);
nand U15495 (N_15495,N_14493,N_12968);
nor U15496 (N_15496,N_10153,N_14654);
xnor U15497 (N_15497,N_11057,N_10352);
xnor U15498 (N_15498,N_11732,N_13397);
nor U15499 (N_15499,N_12934,N_10508);
or U15500 (N_15500,N_10090,N_10186);
nor U15501 (N_15501,N_13351,N_13121);
xor U15502 (N_15502,N_10425,N_13279);
nor U15503 (N_15503,N_11756,N_14467);
or U15504 (N_15504,N_12229,N_14570);
xor U15505 (N_15505,N_11069,N_11913);
nand U15506 (N_15506,N_11269,N_14485);
nor U15507 (N_15507,N_12125,N_12014);
and U15508 (N_15508,N_10792,N_14971);
and U15509 (N_15509,N_14573,N_12699);
xnor U15510 (N_15510,N_13737,N_13271);
xor U15511 (N_15511,N_11362,N_13595);
or U15512 (N_15512,N_12439,N_11373);
nand U15513 (N_15513,N_12061,N_12168);
nand U15514 (N_15514,N_14342,N_12114);
nor U15515 (N_15515,N_10806,N_13138);
nor U15516 (N_15516,N_13479,N_11537);
xnor U15517 (N_15517,N_14901,N_10169);
nand U15518 (N_15518,N_10590,N_10175);
nand U15519 (N_15519,N_14617,N_12488);
and U15520 (N_15520,N_11310,N_12172);
nor U15521 (N_15521,N_13214,N_14856);
nor U15522 (N_15522,N_10577,N_13893);
or U15523 (N_15523,N_11064,N_11187);
or U15524 (N_15524,N_12182,N_11844);
or U15525 (N_15525,N_10022,N_12757);
and U15526 (N_15526,N_13920,N_12927);
nand U15527 (N_15527,N_11368,N_12336);
or U15528 (N_15528,N_12734,N_10881);
and U15529 (N_15529,N_11512,N_14976);
or U15530 (N_15530,N_12421,N_11342);
or U15531 (N_15531,N_11383,N_14723);
xor U15532 (N_15532,N_14631,N_14374);
nor U15533 (N_15533,N_13769,N_11990);
and U15534 (N_15534,N_12767,N_12471);
and U15535 (N_15535,N_11281,N_14145);
xor U15536 (N_15536,N_13203,N_14184);
nand U15537 (N_15537,N_12401,N_12203);
or U15538 (N_15538,N_10283,N_11022);
nor U15539 (N_15539,N_13094,N_14693);
and U15540 (N_15540,N_10401,N_12271);
xor U15541 (N_15541,N_10893,N_14075);
or U15542 (N_15542,N_13354,N_11734);
nand U15543 (N_15543,N_11635,N_14822);
or U15544 (N_15544,N_10938,N_13933);
xnor U15545 (N_15545,N_12435,N_10003);
and U15546 (N_15546,N_11018,N_13659);
nor U15547 (N_15547,N_14363,N_11889);
xnor U15548 (N_15548,N_13738,N_11565);
and U15549 (N_15549,N_13199,N_14050);
nor U15550 (N_15550,N_13123,N_10803);
xnor U15551 (N_15551,N_13810,N_10374);
and U15552 (N_15552,N_12747,N_12874);
xnor U15553 (N_15553,N_12933,N_14448);
and U15554 (N_15554,N_13589,N_13515);
and U15555 (N_15555,N_14228,N_10486);
nor U15556 (N_15556,N_13080,N_10660);
or U15557 (N_15557,N_12902,N_14590);
nor U15558 (N_15558,N_11365,N_11379);
and U15559 (N_15559,N_11711,N_14418);
xnor U15560 (N_15560,N_14266,N_12824);
nor U15561 (N_15561,N_14869,N_14568);
xor U15562 (N_15562,N_10216,N_13599);
nand U15563 (N_15563,N_11143,N_14909);
and U15564 (N_15564,N_12248,N_13039);
nand U15565 (N_15565,N_14153,N_11132);
and U15566 (N_15566,N_12037,N_12453);
nor U15567 (N_15567,N_12638,N_11588);
xor U15568 (N_15568,N_12783,N_13655);
or U15569 (N_15569,N_10745,N_11899);
or U15570 (N_15570,N_11213,N_13674);
nor U15571 (N_15571,N_12761,N_14897);
and U15572 (N_15572,N_10395,N_10246);
and U15573 (N_15573,N_11315,N_11876);
nand U15574 (N_15574,N_14265,N_13110);
nand U15575 (N_15575,N_10784,N_10168);
xnor U15576 (N_15576,N_12967,N_13452);
xnor U15577 (N_15577,N_10648,N_13657);
or U15578 (N_15578,N_10095,N_12612);
xor U15579 (N_15579,N_10416,N_12244);
xnor U15580 (N_15580,N_13611,N_13311);
xnor U15581 (N_15581,N_13930,N_10939);
and U15582 (N_15582,N_10026,N_11589);
nand U15583 (N_15583,N_10646,N_14898);
nand U15584 (N_15584,N_13878,N_13882);
and U15585 (N_15585,N_11433,N_13380);
xnor U15586 (N_15586,N_12740,N_10165);
xor U15587 (N_15587,N_12583,N_14277);
xor U15588 (N_15588,N_11049,N_14691);
and U15589 (N_15589,N_14253,N_12308);
or U15590 (N_15590,N_12352,N_12758);
or U15591 (N_15591,N_14928,N_12276);
nor U15592 (N_15592,N_12536,N_13487);
or U15593 (N_15593,N_11226,N_14094);
xnor U15594 (N_15594,N_14168,N_14188);
nand U15595 (N_15595,N_12994,N_10435);
nor U15596 (N_15596,N_14801,N_13128);
xor U15597 (N_15597,N_14437,N_10362);
or U15598 (N_15598,N_13835,N_12030);
xor U15599 (N_15599,N_14307,N_10413);
nand U15600 (N_15600,N_11062,N_13018);
nand U15601 (N_15601,N_12431,N_13772);
and U15602 (N_15602,N_10997,N_14381);
and U15603 (N_15603,N_11979,N_11183);
nand U15604 (N_15604,N_10988,N_10161);
nand U15605 (N_15605,N_13407,N_10754);
nand U15606 (N_15606,N_14967,N_14716);
xor U15607 (N_15607,N_11502,N_13526);
nand U15608 (N_15608,N_13468,N_14037);
nor U15609 (N_15609,N_10737,N_12076);
and U15610 (N_15610,N_12827,N_14992);
and U15611 (N_15611,N_12033,N_10363);
and U15612 (N_15612,N_10333,N_12156);
xor U15613 (N_15613,N_11030,N_14137);
and U15614 (N_15614,N_10316,N_12629);
nand U15615 (N_15615,N_11974,N_12480);
or U15616 (N_15616,N_14546,N_14704);
xor U15617 (N_15617,N_10010,N_10850);
nor U15618 (N_15618,N_12882,N_14787);
and U15619 (N_15619,N_11196,N_12689);
or U15620 (N_15620,N_11865,N_11606);
nand U15621 (N_15621,N_12135,N_11515);
nor U15622 (N_15622,N_10446,N_11860);
and U15623 (N_15623,N_14878,N_11232);
nand U15624 (N_15624,N_13573,N_11219);
xnor U15625 (N_15625,N_10281,N_12864);
or U15626 (N_15626,N_11621,N_11394);
and U15627 (N_15627,N_10890,N_14347);
nand U15628 (N_15628,N_11823,N_12446);
nor U15629 (N_15629,N_12159,N_10928);
nor U15630 (N_15630,N_10347,N_11244);
xnor U15631 (N_15631,N_10480,N_11192);
or U15632 (N_15632,N_14620,N_13051);
xor U15633 (N_15633,N_13977,N_13720);
nor U15634 (N_15634,N_12991,N_13403);
xor U15635 (N_15635,N_10227,N_10249);
nor U15636 (N_15636,N_11981,N_10982);
and U15637 (N_15637,N_12669,N_14375);
nand U15638 (N_15638,N_13159,N_12609);
nor U15639 (N_15639,N_13927,N_10990);
nand U15640 (N_15640,N_10477,N_14400);
nand U15641 (N_15641,N_14552,N_10588);
nand U15642 (N_15642,N_14838,N_13999);
or U15643 (N_15643,N_14694,N_10618);
nand U15644 (N_15644,N_11471,N_13652);
or U15645 (N_15645,N_12925,N_11489);
nand U15646 (N_15646,N_11906,N_12287);
xor U15647 (N_15647,N_12161,N_13748);
nor U15648 (N_15648,N_14641,N_10576);
and U15649 (N_15649,N_13583,N_10797);
nand U15650 (N_15650,N_11730,N_11090);
xor U15651 (N_15651,N_11114,N_10623);
nand U15652 (N_15652,N_11225,N_14415);
nand U15653 (N_15653,N_14482,N_12075);
xor U15654 (N_15654,N_14259,N_14162);
and U15655 (N_15655,N_13464,N_10075);
nor U15656 (N_15656,N_13581,N_11789);
xnor U15657 (N_15657,N_10667,N_10864);
xor U15658 (N_15658,N_10880,N_12640);
nor U15659 (N_15659,N_14799,N_12022);
xor U15660 (N_15660,N_11039,N_11462);
and U15661 (N_15661,N_13499,N_10479);
and U15662 (N_15662,N_10686,N_13538);
nor U15663 (N_15663,N_11903,N_10750);
or U15664 (N_15664,N_14320,N_10942);
or U15665 (N_15665,N_14411,N_14059);
xor U15666 (N_15666,N_14409,N_13640);
or U15667 (N_15667,N_11179,N_13222);
and U15668 (N_15668,N_12713,N_13587);
nand U15669 (N_15669,N_12990,N_14782);
xnor U15670 (N_15670,N_11136,N_14591);
nor U15671 (N_15671,N_14755,N_14585);
nand U15672 (N_15672,N_13950,N_14367);
or U15673 (N_15673,N_13502,N_12793);
xor U15674 (N_15674,N_14776,N_14757);
nand U15675 (N_15675,N_12263,N_10616);
nor U15676 (N_15676,N_12851,N_14577);
or U15677 (N_15677,N_13367,N_10789);
nor U15678 (N_15678,N_14312,N_14425);
and U15679 (N_15679,N_13752,N_14494);
and U15680 (N_15680,N_12723,N_12557);
xnor U15681 (N_15681,N_10218,N_13898);
nand U15682 (N_15682,N_11027,N_11923);
and U15683 (N_15683,N_13438,N_13507);
nor U15684 (N_15684,N_11122,N_13571);
or U15685 (N_15685,N_12620,N_10073);
or U15686 (N_15686,N_11168,N_14854);
nor U15687 (N_15687,N_12820,N_14255);
nor U15688 (N_15688,N_14021,N_14686);
nor U15689 (N_15689,N_14345,N_12301);
and U15690 (N_15690,N_12726,N_12390);
xor U15691 (N_15691,N_12671,N_13015);
xor U15692 (N_15692,N_13188,N_11386);
nor U15693 (N_15693,N_12661,N_10448);
or U15694 (N_15694,N_11461,N_10711);
nand U15695 (N_15695,N_14737,N_14223);
or U15696 (N_15696,N_13524,N_11526);
nor U15697 (N_15697,N_14171,N_11258);
nor U15698 (N_15698,N_13513,N_10555);
nand U15699 (N_15699,N_14980,N_10496);
or U15700 (N_15700,N_11165,N_11665);
xnor U15701 (N_15701,N_13282,N_11189);
nor U15702 (N_15702,N_11272,N_12462);
xor U15703 (N_15703,N_10041,N_13299);
nor U15704 (N_15704,N_13117,N_14774);
and U15705 (N_15705,N_11792,N_11548);
xor U15706 (N_15706,N_14942,N_11151);
and U15707 (N_15707,N_10837,N_12006);
xor U15708 (N_15708,N_10695,N_10701);
nand U15709 (N_15709,N_13017,N_13649);
nor U15710 (N_15710,N_14852,N_12881);
nand U15711 (N_15711,N_10971,N_10687);
nand U15712 (N_15712,N_10285,N_14890);
nand U15713 (N_15713,N_12837,N_14512);
nand U15714 (N_15714,N_13306,N_14816);
nor U15715 (N_15715,N_11067,N_13996);
nor U15716 (N_15716,N_14435,N_11836);
or U15717 (N_15717,N_13939,N_14834);
nand U15718 (N_15718,N_10079,N_14845);
and U15719 (N_15719,N_11951,N_12602);
nor U15720 (N_15720,N_12919,N_12987);
nand U15721 (N_15721,N_12655,N_12123);
xnor U15722 (N_15722,N_14531,N_13422);
or U15723 (N_15723,N_11463,N_10013);
or U15724 (N_15724,N_14189,N_11215);
and U15725 (N_15725,N_11664,N_11237);
xor U15726 (N_15726,N_14764,N_12619);
nand U15727 (N_15727,N_13456,N_12884);
xnor U15728 (N_15728,N_11933,N_14023);
xor U15729 (N_15729,N_10627,N_11199);
or U15730 (N_15730,N_12959,N_14990);
xor U15731 (N_15731,N_10082,N_14989);
or U15732 (N_15732,N_12433,N_10960);
nand U15733 (N_15733,N_12715,N_14575);
or U15734 (N_15734,N_10604,N_13915);
nor U15735 (N_15735,N_13413,N_14504);
or U15736 (N_15736,N_14489,N_10007);
nor U15737 (N_15737,N_11401,N_14902);
nand U15738 (N_15738,N_12053,N_13963);
xor U15739 (N_15739,N_14602,N_14104);
xor U15740 (N_15740,N_12996,N_13782);
and U15741 (N_15741,N_13228,N_11270);
nor U15742 (N_15742,N_13364,N_11366);
or U15743 (N_15743,N_14770,N_13059);
xnor U15744 (N_15744,N_12041,N_11532);
nand U15745 (N_15745,N_14175,N_10146);
and U15746 (N_15746,N_14559,N_11140);
or U15747 (N_15747,N_13149,N_11312);
nor U15748 (N_15748,N_14925,N_11162);
nor U15749 (N_15749,N_10238,N_12253);
nand U15750 (N_15750,N_14780,N_14407);
xor U15751 (N_15751,N_12584,N_14806);
xor U15752 (N_15752,N_10857,N_12932);
nor U15753 (N_15753,N_14610,N_12772);
xor U15754 (N_15754,N_12782,N_12543);
nor U15755 (N_15755,N_11009,N_14638);
nor U15756 (N_15756,N_10286,N_11094);
and U15757 (N_15757,N_10517,N_11113);
xnor U15758 (N_15758,N_13847,N_10707);
nand U15759 (N_15759,N_12657,N_13029);
nor U15760 (N_15760,N_11950,N_11946);
or U15761 (N_15761,N_14177,N_14683);
or U15762 (N_15762,N_12826,N_14047);
nor U15763 (N_15763,N_10080,N_12491);
or U15764 (N_15764,N_13542,N_10278);
nor U15765 (N_15765,N_11715,N_11966);
and U15766 (N_15766,N_13968,N_11550);
xor U15767 (N_15767,N_12805,N_11046);
or U15768 (N_15768,N_14798,N_12412);
and U15769 (N_15769,N_13454,N_14076);
nand U15770 (N_15770,N_13231,N_12293);
nor U15771 (N_15771,N_14681,N_13381);
nor U15772 (N_15772,N_14858,N_14352);
nand U15773 (N_15773,N_14335,N_11349);
nand U15774 (N_15774,N_10501,N_13792);
xnor U15775 (N_15775,N_13959,N_14067);
xnor U15776 (N_15776,N_11516,N_10894);
nor U15777 (N_15777,N_12876,N_13344);
and U15778 (N_15778,N_10233,N_14649);
nor U15779 (N_15779,N_10299,N_14880);
nand U15780 (N_15780,N_14111,N_10991);
nor U15781 (N_15781,N_10682,N_13229);
xnor U15782 (N_15782,N_14866,N_10489);
nand U15783 (N_15783,N_10094,N_13618);
nor U15784 (N_15784,N_14771,N_11733);
nor U15785 (N_15785,N_11227,N_10892);
or U15786 (N_15786,N_13178,N_12371);
or U15787 (N_15787,N_14446,N_13101);
nand U15788 (N_15788,N_11883,N_11975);
and U15789 (N_15789,N_14201,N_13483);
xnor U15790 (N_15790,N_10149,N_13462);
nand U15791 (N_15791,N_11308,N_12329);
and U15792 (N_15792,N_13455,N_14983);
nor U15793 (N_15793,N_11500,N_14158);
nor U15794 (N_15794,N_11160,N_13797);
nor U15795 (N_15795,N_11517,N_11188);
nand U15796 (N_15796,N_12570,N_11337);
nor U15797 (N_15797,N_13164,N_12650);
or U15798 (N_15798,N_14597,N_11723);
xor U15799 (N_15799,N_14198,N_14870);
nand U15800 (N_15800,N_10860,N_14046);
nor U15801 (N_15801,N_13702,N_12838);
xor U15802 (N_15802,N_11250,N_11166);
nor U15803 (N_15803,N_12303,N_11563);
or U15804 (N_15804,N_11827,N_13166);
or U15805 (N_15805,N_13350,N_13223);
nor U15806 (N_15806,N_10587,N_13174);
nand U15807 (N_15807,N_11444,N_13905);
nor U15808 (N_15808,N_13476,N_10147);
and U15809 (N_15809,N_12610,N_13607);
and U15810 (N_15810,N_14143,N_12372);
nor U15811 (N_15811,N_13814,N_10421);
and U15812 (N_15812,N_13492,N_12685);
nor U15813 (N_15813,N_10176,N_11681);
and U15814 (N_15814,N_14509,N_14562);
or U15815 (N_15815,N_13757,N_11587);
or U15816 (N_15816,N_12880,N_12643);
nand U15817 (N_15817,N_10582,N_14480);
and U15818 (N_15818,N_10909,N_10624);
xor U15819 (N_15819,N_14121,N_10188);
nand U15820 (N_15820,N_12102,N_12034);
xor U15821 (N_15821,N_12409,N_13525);
and U15822 (N_15822,N_14640,N_10672);
xor U15823 (N_15823,N_14351,N_13910);
xor U15824 (N_15824,N_10260,N_11442);
nand U15825 (N_15825,N_14921,N_12314);
and U15826 (N_15826,N_12541,N_10449);
and U15827 (N_15827,N_13063,N_10426);
and U15828 (N_15828,N_12587,N_10032);
xor U15829 (N_15829,N_10819,N_12768);
and U15830 (N_15830,N_14442,N_11059);
nand U15831 (N_15831,N_11289,N_14805);
or U15832 (N_15832,N_11195,N_11784);
nand U15833 (N_15833,N_13741,N_14292);
and U15834 (N_15834,N_10640,N_12795);
nand U15835 (N_15835,N_13436,N_13925);
nor U15836 (N_15836,N_12885,N_14701);
nor U15837 (N_15837,N_11257,N_10800);
nand U15838 (N_15838,N_11455,N_10012);
or U15839 (N_15839,N_13273,N_12651);
nor U15840 (N_15840,N_14850,N_14506);
nor U15841 (N_15841,N_12617,N_10748);
nand U15842 (N_15842,N_12732,N_12201);
or U15843 (N_15843,N_14526,N_12717);
xor U15844 (N_15844,N_14044,N_14174);
or U15845 (N_15845,N_14560,N_13389);
nand U15846 (N_15846,N_11363,N_14721);
or U15847 (N_15847,N_13802,N_11652);
xnor U15848 (N_15848,N_14100,N_10779);
or U15849 (N_15849,N_10952,N_12426);
and U15850 (N_15850,N_12100,N_10120);
or U15851 (N_15851,N_10367,N_14164);
nand U15852 (N_15852,N_11484,N_13378);
xor U15853 (N_15853,N_14667,N_13796);
and U15854 (N_15854,N_13384,N_10313);
xnor U15855 (N_15855,N_13267,N_10529);
nor U15856 (N_15856,N_12642,N_13717);
nand U15857 (N_15857,N_13682,N_10195);
xnor U15858 (N_15858,N_11153,N_13150);
nor U15859 (N_15859,N_10231,N_11578);
nand U15860 (N_15860,N_12593,N_10129);
or U15861 (N_15861,N_13013,N_11855);
or U15862 (N_15862,N_10773,N_10807);
nor U15863 (N_15863,N_11885,N_11451);
nand U15864 (N_15864,N_11288,N_10870);
xor U15865 (N_15865,N_10539,N_14660);
nor U15866 (N_15866,N_10408,N_10856);
xnor U15867 (N_15867,N_12447,N_13239);
nor U15868 (N_15868,N_13861,N_14687);
and U15869 (N_15869,N_12269,N_14644);
nor U15870 (N_15870,N_12973,N_12450);
and U15871 (N_15871,N_14593,N_13966);
nor U15872 (N_15872,N_11292,N_10108);
or U15873 (N_15873,N_10718,N_14148);
nor U15874 (N_15874,N_14302,N_10059);
or U15875 (N_15875,N_14017,N_13871);
and U15876 (N_15876,N_11038,N_14093);
and U15877 (N_15877,N_14227,N_11211);
nor U15878 (N_15878,N_14195,N_13991);
nor U15879 (N_15879,N_12871,N_10578);
nand U15880 (N_15880,N_12147,N_13172);
or U15881 (N_15881,N_10093,N_13598);
and U15882 (N_15882,N_12019,N_14441);
or U15883 (N_15883,N_12160,N_10139);
xnor U15884 (N_15884,N_11831,N_14460);
or U15885 (N_15885,N_12265,N_12810);
or U15886 (N_15886,N_11794,N_13181);
nor U15887 (N_15887,N_14794,N_12786);
nand U15888 (N_15888,N_13732,N_14948);
and U15889 (N_15889,N_10160,N_12708);
nor U15890 (N_15890,N_12064,N_11738);
nor U15891 (N_15891,N_10098,N_10369);
nand U15892 (N_15892,N_13813,N_11191);
nand U15893 (N_15893,N_12849,N_12769);
and U15894 (N_15894,N_10088,N_13805);
xor U15895 (N_15895,N_13428,N_12582);
nand U15896 (N_15896,N_13809,N_14936);
xnor U15897 (N_15897,N_13127,N_14952);
nor U15898 (N_15898,N_14978,N_11040);
xor U15899 (N_15899,N_13314,N_11634);
and U15900 (N_15900,N_10751,N_12533);
nor U15901 (N_15901,N_12711,N_13689);
or U15902 (N_15902,N_10058,N_11029);
xnor U15903 (N_15903,N_11554,N_14393);
nor U15904 (N_15904,N_11016,N_10848);
and U15905 (N_15905,N_14369,N_11048);
or U15906 (N_15906,N_10879,N_10774);
or U15907 (N_15907,N_13561,N_10756);
and U15908 (N_15908,N_11527,N_10581);
or U15909 (N_15909,N_13758,N_14802);
and U15910 (N_15910,N_10148,N_10636);
xor U15911 (N_15911,N_11735,N_10531);
or U15912 (N_15912,N_14120,N_10038);
xnor U15913 (N_15913,N_10815,N_11830);
and U15914 (N_15914,N_14241,N_10802);
xnor U15915 (N_15915,N_13943,N_10808);
nor U15916 (N_15916,N_13759,N_11494);
nand U15917 (N_15917,N_10236,N_14618);
and U15918 (N_15918,N_13302,N_12343);
or U15919 (N_15919,N_11278,N_10325);
nor U15920 (N_15920,N_11010,N_11085);
nand U15921 (N_15921,N_11210,N_10681);
and U15922 (N_15922,N_10048,N_13131);
xor U15923 (N_15923,N_11130,N_11856);
nor U15924 (N_15924,N_11116,N_13829);
or U15925 (N_15925,N_10804,N_14128);
and U15926 (N_15926,N_10791,N_10777);
nor U15927 (N_15927,N_10946,N_12648);
nor U15928 (N_15928,N_10277,N_13981);
nand U15929 (N_15929,N_10532,N_11841);
nor U15930 (N_15930,N_13990,N_10170);
xnor U15931 (N_15931,N_14719,N_14456);
and U15932 (N_15932,N_14205,N_14187);
and U15933 (N_15933,N_12531,N_12339);
nor U15934 (N_15934,N_14399,N_11032);
nor U15935 (N_15935,N_10315,N_14015);
nor U15936 (N_15936,N_13667,N_10614);
and U15937 (N_15937,N_12800,N_13628);
or U15938 (N_15938,N_14679,N_13739);
xor U15939 (N_15939,N_10293,N_11033);
xnor U15940 (N_15940,N_14965,N_10502);
nand U15941 (N_15941,N_10985,N_13347);
nor U15942 (N_15942,N_11965,N_11839);
nor U15943 (N_15943,N_10355,N_11861);
nand U15944 (N_15944,N_13449,N_13340);
and U15945 (N_15945,N_12622,N_12672);
xnor U15946 (N_15946,N_13632,N_10872);
xnor U15947 (N_15947,N_13859,N_14988);
nor U15948 (N_15948,N_10151,N_11698);
and U15949 (N_15949,N_13626,N_13093);
or U15950 (N_15950,N_14025,N_13931);
nand U15951 (N_15951,N_10128,N_12130);
or U15952 (N_15952,N_13004,N_11207);
or U15953 (N_15953,N_11075,N_13527);
and U15954 (N_15954,N_13374,N_11481);
xnor U15955 (N_15955,N_12279,N_13972);
and U15956 (N_15956,N_12068,N_11275);
nor U15957 (N_15957,N_11807,N_12972);
nor U15958 (N_15958,N_12736,N_11370);
nor U15959 (N_15959,N_13252,N_13816);
nor U15960 (N_15960,N_12150,N_14117);
and U15961 (N_15961,N_10781,N_13060);
nand U15962 (N_15962,N_10067,N_12414);
nand U15963 (N_15963,N_14300,N_13095);
or U15964 (N_15964,N_11931,N_12606);
or U15965 (N_15965,N_11757,N_11902);
nand U15966 (N_15966,N_12361,N_13052);
nor U15967 (N_15967,N_11392,N_11025);
or U15968 (N_15968,N_10191,N_12071);
nor U15969 (N_15969,N_14859,N_12067);
and U15970 (N_15970,N_10162,N_10690);
nor U15971 (N_15971,N_12776,N_10541);
nand U15972 (N_15972,N_13980,N_13743);
and U15973 (N_15973,N_10130,N_14918);
xor U15974 (N_15974,N_10632,N_12698);
nor U15975 (N_15975,N_11945,N_13140);
nor U15976 (N_15976,N_11559,N_11609);
nand U15977 (N_15977,N_11193,N_11557);
or U15978 (N_15978,N_14131,N_10102);
xor U15979 (N_15979,N_13254,N_11828);
and U15980 (N_15980,N_14835,N_13642);
nor U15981 (N_15981,N_12564,N_11754);
nor U15982 (N_15982,N_11346,N_13366);
nor U15983 (N_15983,N_13091,N_13245);
nor U15984 (N_15984,N_14247,N_10859);
or U15985 (N_15985,N_10491,N_12485);
xor U15986 (N_15986,N_13891,N_10575);
and U15987 (N_15987,N_12290,N_13781);
nand U15988 (N_15988,N_12106,N_13550);
xor U15989 (N_15989,N_14754,N_11700);
xor U15990 (N_15990,N_14444,N_10983);
and U15991 (N_15991,N_14986,N_12944);
xnor U15992 (N_15992,N_11218,N_13568);
xnor U15993 (N_15993,N_13383,N_12220);
or U15994 (N_15994,N_10868,N_11586);
nand U15995 (N_15995,N_12678,N_13119);
nor U15996 (N_15996,N_14534,N_11086);
nor U15997 (N_15997,N_14006,N_14258);
nor U15998 (N_15998,N_12087,N_11553);
nor U15999 (N_15999,N_14127,N_13471);
or U16000 (N_16000,N_11745,N_12378);
or U16001 (N_16001,N_12389,N_12766);
xor U16002 (N_16002,N_14027,N_14524);
nor U16003 (N_16003,N_10224,N_11003);
nor U16004 (N_16004,N_11200,N_14149);
nand U16005 (N_16005,N_13699,N_14677);
and U16006 (N_16006,N_12079,N_10118);
nor U16007 (N_16007,N_13744,N_14226);
nor U16008 (N_16008,N_12887,N_13210);
and U16009 (N_16009,N_14377,N_13553);
and U16010 (N_16010,N_13280,N_11773);
or U16011 (N_16011,N_13817,N_14888);
and U16012 (N_16012,N_13106,N_12812);
nor U16013 (N_16013,N_10535,N_13622);
or U16014 (N_16014,N_13723,N_12614);
nand U16015 (N_16015,N_11878,N_12576);
nand U16016 (N_16016,N_10243,N_12852);
and U16017 (N_16017,N_10004,N_11496);
or U16018 (N_16018,N_10932,N_10980);
and U16019 (N_16019,N_14843,N_12992);
xor U16020 (N_16020,N_13856,N_11551);
nand U16021 (N_16021,N_13580,N_14224);
xnor U16022 (N_16022,N_13205,N_14303);
nor U16023 (N_16023,N_12288,N_12332);
or U16024 (N_16024,N_13272,N_11835);
nor U16025 (N_16025,N_14630,N_11653);
xnor U16026 (N_16026,N_11452,N_11096);
nand U16027 (N_16027,N_10719,N_14274);
or U16028 (N_16028,N_11708,N_11037);
or U16029 (N_16029,N_10226,N_11164);
nor U16030 (N_16030,N_14808,N_13520);
and U16031 (N_16031,N_13577,N_12208);
nand U16032 (N_16032,N_13421,N_10899);
and U16033 (N_16033,N_10523,N_14380);
and U16034 (N_16034,N_12424,N_10126);
or U16035 (N_16035,N_13337,N_10273);
xnor U16036 (N_16036,N_11176,N_13512);
nor U16037 (N_16037,N_14475,N_12535);
nor U16038 (N_16038,N_10734,N_10356);
and U16039 (N_16039,N_14853,N_13255);
xor U16040 (N_16040,N_13543,N_13402);
and U16041 (N_16041,N_10524,N_12633);
nor U16042 (N_16042,N_14275,N_12829);
and U16043 (N_16043,N_11091,N_11372);
xor U16044 (N_16044,N_12113,N_10179);
xor U16045 (N_16045,N_10840,N_11726);
and U16046 (N_16046,N_12003,N_12083);
nand U16047 (N_16047,N_13215,N_11926);
nand U16048 (N_16048,N_13883,N_13077);
and U16049 (N_16049,N_10040,N_12321);
and U16050 (N_16050,N_13531,N_14572);
or U16051 (N_16051,N_13336,N_13287);
xor U16052 (N_16052,N_14141,N_12395);
or U16053 (N_16053,N_14063,N_11334);
nor U16054 (N_16054,N_11629,N_11458);
nand U16055 (N_16055,N_10490,N_11472);
nand U16056 (N_16056,N_12382,N_12178);
nor U16057 (N_16057,N_10294,N_12563);
nor U16058 (N_16058,N_13423,N_12561);
and U16059 (N_16059,N_13333,N_10647);
and U16060 (N_16060,N_11619,N_10412);
nand U16061 (N_16061,N_13335,N_14403);
and U16062 (N_16062,N_13877,N_11479);
and U16063 (N_16063,N_14349,N_12842);
nor U16064 (N_16064,N_14919,N_14533);
and U16065 (N_16065,N_12183,N_14492);
xnor U16066 (N_16066,N_11262,N_12970);
or U16067 (N_16067,N_10668,N_13516);
nand U16068 (N_16068,N_13532,N_12277);
nor U16069 (N_16069,N_11987,N_12449);
nor U16070 (N_16070,N_10409,N_10914);
nand U16071 (N_16071,N_14251,N_13412);
nand U16072 (N_16072,N_13851,N_12132);
or U16073 (N_16073,N_10965,N_13425);
nand U16074 (N_16074,N_10742,N_13938);
and U16075 (N_16075,N_13368,N_11763);
xnor U16076 (N_16076,N_11107,N_14238);
nor U16077 (N_16077,N_13730,N_11904);
and U16078 (N_16078,N_10871,N_14516);
or U16079 (N_16079,N_14688,N_10110);
nor U16080 (N_16080,N_13510,N_14458);
nor U16081 (N_16081,N_14138,N_12327);
and U16082 (N_16082,N_12151,N_12477);
and U16083 (N_16083,N_12831,N_10996);
xor U16084 (N_16084,N_12560,N_10220);
and U16085 (N_16085,N_10675,N_10855);
xor U16086 (N_16086,N_10725,N_12631);
xor U16087 (N_16087,N_13567,N_14689);
nand U16088 (N_16088,N_14438,N_10569);
and U16089 (N_16089,N_11141,N_13238);
xor U16090 (N_16090,N_13453,N_13470);
xor U16091 (N_16091,N_11752,N_14125);
and U16092 (N_16092,N_14297,N_13842);
nor U16093 (N_16093,N_11399,N_12913);
nor U16094 (N_16094,N_11019,N_13065);
or U16095 (N_16095,N_14615,N_10436);
nand U16096 (N_16096,N_13037,N_11838);
or U16097 (N_16097,N_12840,N_14452);
nor U16098 (N_16098,N_12381,N_14993);
nor U16099 (N_16099,N_12406,N_10509);
nor U16100 (N_16100,N_12931,N_12299);
nor U16101 (N_16101,N_11416,N_13716);
or U16102 (N_16102,N_12993,N_10334);
nor U16103 (N_16103,N_13320,N_12217);
nand U16104 (N_16104,N_12357,N_14410);
and U16105 (N_16105,N_12983,N_14634);
nor U16106 (N_16106,N_13556,N_10047);
and U16107 (N_16107,N_11567,N_10822);
xnor U16108 (N_16108,N_10786,N_13766);
xnor U16109 (N_16109,N_14071,N_11228);
nor U16110 (N_16110,N_14069,N_10344);
xnor U16111 (N_16111,N_13264,N_11881);
xor U16112 (N_16112,N_11405,N_13432);
nor U16113 (N_16113,N_14271,N_12403);
nand U16114 (N_16114,N_10641,N_10016);
or U16115 (N_16115,N_13465,N_13770);
or U16116 (N_16116,N_14847,N_14004);
nand U16117 (N_16117,N_11637,N_13171);
xor U16118 (N_16118,N_13971,N_10455);
and U16119 (N_16119,N_11293,N_13934);
or U16120 (N_16120,N_14728,N_13474);
or U16121 (N_16121,N_12456,N_13088);
nor U16122 (N_16122,N_13906,N_14496);
nand U16123 (N_16123,N_12601,N_13710);
and U16124 (N_16124,N_11021,N_10805);
or U16125 (N_16125,N_12185,N_13219);
nor U16126 (N_16126,N_13023,N_13703);
or U16127 (N_16127,N_10241,N_11970);
or U16128 (N_16128,N_11868,N_10463);
nand U16129 (N_16129,N_10814,N_11943);
and U16130 (N_16130,N_12219,N_12870);
nor U16131 (N_16131,N_14155,N_11285);
xor U16132 (N_16132,N_11683,N_12704);
nand U16133 (N_16133,N_13661,N_10042);
and U16134 (N_16134,N_10833,N_13173);
and U16135 (N_16135,N_12120,N_11922);
or U16136 (N_16136,N_14287,N_12938);
and U16137 (N_16137,N_10691,N_11918);
or U16138 (N_16138,N_12930,N_11787);
or U16139 (N_16139,N_14609,N_13158);
nand U16140 (N_16140,N_13285,N_10966);
xnor U16141 (N_16141,N_10995,N_13995);
xnor U16142 (N_16142,N_10474,N_13671);
or U16143 (N_16143,N_14743,N_14328);
and U16144 (N_16144,N_10366,N_11540);
nand U16145 (N_16145,N_13461,N_12236);
nor U16146 (N_16146,N_14717,N_13154);
or U16147 (N_16147,N_12962,N_14327);
nor U16148 (N_16148,N_10208,N_14781);
and U16149 (N_16149,N_14331,N_11335);
and U16150 (N_16150,N_10638,N_11869);
or U16151 (N_16151,N_11687,N_12112);
or U16152 (N_16152,N_13007,N_11408);
and U16153 (N_16153,N_10331,N_12733);
xnor U16154 (N_16154,N_10198,N_13986);
xor U16155 (N_16155,N_14851,N_11001);
nor U16156 (N_16156,N_13727,N_12939);
nor U16157 (N_16157,N_12375,N_11294);
nor U16158 (N_16158,N_13631,N_13656);
nand U16159 (N_16159,N_14123,N_10898);
nand U16160 (N_16160,N_14817,N_12953);
xnor U16161 (N_16161,N_13288,N_13001);
nor U16162 (N_16162,N_10712,N_10014);
and U16163 (N_16163,N_10896,N_14003);
xor U16164 (N_16164,N_11427,N_13020);
nand U16165 (N_16165,N_12478,N_10620);
nor U16166 (N_16166,N_11707,N_14102);
xnor U16167 (N_16167,N_10903,N_13331);
and U16168 (N_16168,N_10975,N_12916);
or U16169 (N_16169,N_13491,N_13509);
nor U16170 (N_16170,N_10302,N_11036);
nand U16171 (N_16171,N_10710,N_10630);
nor U16172 (N_16172,N_14147,N_10811);
nor U16173 (N_16173,N_12286,N_12388);
nor U16174 (N_16174,N_12868,N_11680);
nand U16175 (N_16175,N_14525,N_10545);
xor U16176 (N_16176,N_11118,N_14365);
xnor U16177 (N_16177,N_12430,N_10920);
xor U16178 (N_16178,N_10288,N_14837);
or U16179 (N_16179,N_14741,N_10650);
nor U16180 (N_16180,N_13303,N_10897);
nand U16181 (N_16181,N_10398,N_11282);
nor U16182 (N_16182,N_11776,N_14336);
nand U16183 (N_16183,N_14103,N_13357);
nand U16184 (N_16184,N_10002,N_14068);
nor U16185 (N_16185,N_14057,N_10206);
xnor U16186 (N_16186,N_14647,N_11145);
nor U16187 (N_16187,N_13707,N_13685);
and U16188 (N_16188,N_14722,N_13616);
xor U16189 (N_16189,N_10280,N_13033);
nor U16190 (N_16190,N_11742,N_13828);
or U16191 (N_16191,N_12322,N_12828);
xnor U16192 (N_16192,N_14659,N_11234);
nor U16193 (N_16193,N_13683,N_10678);
or U16194 (N_16194,N_14065,N_11956);
and U16195 (N_16195,N_12032,N_13780);
and U16196 (N_16196,N_14924,N_10519);
or U16197 (N_16197,N_14917,N_14821);
nand U16198 (N_16198,N_10772,N_12866);
nand U16199 (N_16199,N_11992,N_13275);
nor U16200 (N_16200,N_10245,N_13819);
and U16201 (N_16201,N_11239,N_10584);
nand U16202 (N_16202,N_10659,N_14242);
xor U16203 (N_16203,N_14371,N_14392);
xnor U16204 (N_16204,N_13612,N_10553);
or U16205 (N_16205,N_11599,N_12562);
and U16206 (N_16206,N_10820,N_13795);
or U16207 (N_16207,N_12211,N_10375);
and U16208 (N_16208,N_11659,N_10613);
nor U16209 (N_16209,N_14459,N_10599);
and U16210 (N_16210,N_12010,N_14084);
or U16211 (N_16211,N_14404,N_14657);
nor U16212 (N_16212,N_10684,N_12500);
and U16213 (N_16213,N_13003,N_10676);
nor U16214 (N_16214,N_12928,N_14236);
nand U16215 (N_16215,N_10611,N_12193);
and U16216 (N_16216,N_13908,N_11460);
xor U16217 (N_16217,N_12326,N_13183);
nor U16218 (N_16218,N_13301,N_10384);
and U16219 (N_16219,N_13837,N_11466);
or U16220 (N_16220,N_13676,N_13401);
and U16221 (N_16221,N_12221,N_12216);
and U16222 (N_16222,N_13286,N_13904);
or U16223 (N_16223,N_10021,N_12941);
nand U16224 (N_16224,N_11623,N_10257);
and U16225 (N_16225,N_11916,N_14040);
nand U16226 (N_16226,N_10740,N_14832);
and U16227 (N_16227,N_14819,N_13197);
xnor U16228 (N_16228,N_14285,N_10628);
nand U16229 (N_16229,N_11695,N_14016);
nand U16230 (N_16230,N_14315,N_12966);
nor U16231 (N_16231,N_14390,N_13277);
nor U16232 (N_16232,N_11078,N_10037);
or U16233 (N_16233,N_11361,N_13976);
and U16234 (N_16234,N_14656,N_12687);
nand U16235 (N_16235,N_12978,N_10635);
nor U16236 (N_16236,N_14883,N_10414);
nor U16237 (N_16237,N_11331,N_12585);
or U16238 (N_16238,N_13503,N_10831);
and U16239 (N_16239,N_13410,N_11845);
or U16240 (N_16240,N_13478,N_11900);
nor U16241 (N_16241,N_10724,N_10244);
and U16242 (N_16242,N_11877,N_13390);
nor U16243 (N_16243,N_13889,N_12906);
or U16244 (N_16244,N_14763,N_13196);
nor U16245 (N_16245,N_14389,N_14284);
and U16246 (N_16246,N_12600,N_11249);
nor U16247 (N_16247,N_12532,N_13998);
nand U16248 (N_16248,N_13369,N_12467);
nand U16249 (N_16249,N_12981,N_12797);
or U16250 (N_16250,N_11648,N_14308);
or U16251 (N_16251,N_14318,N_10629);
xor U16252 (N_16252,N_14714,N_13947);
and U16253 (N_16253,N_13496,N_11803);
nor U16254 (N_16254,N_13572,N_10664);
nor U16255 (N_16255,N_10680,N_11820);
nor U16256 (N_16256,N_13115,N_11309);
xnor U16257 (N_16257,N_10100,N_11380);
or U16258 (N_16258,N_12472,N_11099);
nor U16259 (N_16259,N_13993,N_12126);
nor U16260 (N_16260,N_13823,N_10451);
or U16261 (N_16261,N_10500,N_10716);
nor U16262 (N_16262,N_14795,N_14733);
nand U16263 (N_16263,N_11824,N_14672);
nor U16264 (N_16264,N_10956,N_12730);
and U16265 (N_16265,N_13824,N_11296);
xnor U16266 (N_16266,N_14891,N_11102);
and U16267 (N_16267,N_12089,N_13755);
xnor U16268 (N_16268,N_13362,N_10598);
xor U16269 (N_16269,N_10072,N_10053);
nand U16270 (N_16270,N_14240,N_13539);
and U16271 (N_16271,N_11297,N_11566);
and U16272 (N_16272,N_12859,N_11280);
or U16273 (N_16273,N_10542,N_10543);
nor U16274 (N_16274,N_11060,N_12855);
nand U16275 (N_16275,N_14231,N_10096);
xor U16276 (N_16276,N_12841,N_10034);
nand U16277 (N_16277,N_12005,N_13193);
xnor U16278 (N_16278,N_11809,N_14032);
xnor U16279 (N_16279,N_13547,N_10066);
xnor U16280 (N_16280,N_14405,N_12367);
xnor U16281 (N_16281,N_10887,N_12275);
xor U16282 (N_16282,N_13322,N_12377);
nor U16283 (N_16283,N_13969,N_12512);
xnor U16284 (N_16284,N_13179,N_13942);
or U16285 (N_16285,N_12951,N_10989);
xor U16286 (N_16286,N_14885,N_12028);
nor U16287 (N_16287,N_10838,N_10662);
xor U16288 (N_16288,N_11104,N_11454);
nand U16289 (N_16289,N_10087,N_11487);
and U16290 (N_16290,N_14311,N_10839);
and U16291 (N_16291,N_13854,N_13480);
xnor U16292 (N_16292,N_10810,N_14884);
or U16293 (N_16293,N_11744,N_14230);
xnor U16294 (N_16294,N_14604,N_13845);
nand U16295 (N_16295,N_12121,N_12065);
nand U16296 (N_16296,N_13592,N_10320);
nor U16297 (N_16297,N_11654,N_14428);
and U16298 (N_16298,N_14803,N_13575);
or U16299 (N_16299,N_12518,N_12214);
or U16300 (N_16300,N_10589,N_12589);
or U16301 (N_16301,N_12530,N_11846);
nand U16302 (N_16302,N_10214,N_12658);
xnor U16303 (N_16303,N_10340,N_13873);
or U16304 (N_16304,N_13377,N_14035);
or U16305 (N_16305,N_14019,N_12366);
or U16306 (N_16306,N_10562,N_11387);
nand U16307 (N_16307,N_10609,N_13961);
or U16308 (N_16308,N_11972,N_14498);
xnor U16309 (N_16309,N_11340,N_11031);
nand U16310 (N_16310,N_10747,N_12200);
or U16311 (N_16311,N_11529,N_14887);
nand U16312 (N_16312,N_12799,N_11014);
xnor U16313 (N_16313,N_12796,N_10869);
nand U16314 (N_16314,N_13928,N_11034);
xor U16315 (N_16315,N_13198,N_12507);
nor U16316 (N_16316,N_10671,N_14746);
and U16317 (N_16317,N_14582,N_14280);
nand U16318 (N_16318,N_12074,N_11352);
nand U16319 (N_16319,N_10882,N_12985);
nand U16320 (N_16320,N_10308,N_12324);
or U16321 (N_16321,N_11485,N_12094);
nor U16322 (N_16322,N_14920,N_12579);
or U16323 (N_16323,N_12165,N_12368);
nor U16324 (N_16324,N_12929,N_12411);
xnor U16325 (N_16325,N_13894,N_11360);
nor U16326 (N_16326,N_11989,N_11082);
nor U16327 (N_16327,N_12455,N_12141);
or U16328 (N_16328,N_11713,N_13497);
nand U16329 (N_16329,N_12522,N_11666);
or U16330 (N_16330,N_13426,N_13964);
or U16331 (N_16331,N_14692,N_13434);
or U16332 (N_16332,N_14848,N_11967);
nand U16333 (N_16333,N_13345,N_11436);
nor U16334 (N_16334,N_14099,N_12255);
or U16335 (N_16335,N_11543,N_11333);
and U16336 (N_16336,N_10679,N_13157);
nand U16337 (N_16337,N_12599,N_14220);
nor U16338 (N_16338,N_11727,N_13459);
or U16339 (N_16339,N_10074,N_13332);
xor U16340 (N_16340,N_10537,N_10410);
nand U16341 (N_16341,N_14879,N_12282);
xnor U16342 (N_16342,N_14014,N_13715);
and U16343 (N_16343,N_11147,N_11618);
nor U16344 (N_16344,N_13417,N_12804);
or U16345 (N_16345,N_11755,N_10585);
xnor U16346 (N_16346,N_11319,N_10172);
nand U16347 (N_16347,N_10601,N_14635);
or U16348 (N_16348,N_14054,N_10261);
or U16349 (N_16349,N_14896,N_14507);
or U16350 (N_16350,N_11194,N_10196);
and U16351 (N_16351,N_11311,N_12152);
and U16352 (N_16352,N_10951,N_14337);
or U16353 (N_16353,N_14994,N_11625);
xor U16354 (N_16354,N_11499,N_14831);
and U16355 (N_16355,N_11216,N_13068);
xnor U16356 (N_16356,N_11614,N_14624);
nand U16357 (N_16357,N_10847,N_12457);
xnor U16358 (N_16358,N_11800,N_10342);
or U16359 (N_16359,N_14797,N_11837);
and U16360 (N_16360,N_13006,N_10065);
or U16361 (N_16361,N_13783,N_13130);
nand U16362 (N_16362,N_14192,N_14096);
or U16363 (N_16363,N_10230,N_10987);
and U16364 (N_16364,N_10469,N_10876);
xor U16365 (N_16365,N_12494,N_13923);
and U16366 (N_16366,N_13852,N_13949);
nand U16367 (N_16367,N_14655,N_11575);
and U16368 (N_16368,N_11167,N_11400);
and U16369 (N_16369,N_13142,N_12801);
xnor U16370 (N_16370,N_10194,N_13668);
nand U16371 (N_16371,N_10407,N_11682);
xor U16372 (N_16372,N_12632,N_10464);
nor U16373 (N_16373,N_10853,N_11766);
or U16374 (N_16374,N_14070,N_13169);
and U16375 (N_16375,N_14678,N_12460);
nand U16376 (N_16376,N_14578,N_14510);
nand U16377 (N_16377,N_10673,N_14343);
and U16378 (N_16378,N_13742,N_13243);
nand U16379 (N_16379,N_11674,N_10154);
xnor U16380 (N_16380,N_12523,N_13557);
nand U16381 (N_16381,N_13359,N_11942);
nor U16382 (N_16382,N_10046,N_13658);
and U16383 (N_16383,N_14950,N_13064);
nand U16384 (N_16384,N_13192,N_14740);
or U16385 (N_16385,N_10124,N_12110);
xor U16386 (N_16386,N_11255,N_14957);
and U16387 (N_16387,N_14387,N_14268);
xnor U16388 (N_16388,N_12905,N_11740);
nand U16389 (N_16389,N_11518,N_12618);
xor U16390 (N_16390,N_10670,N_10530);
and U16391 (N_16391,N_12443,N_10959);
xor U16392 (N_16392,N_11080,N_12206);
nand U16393 (N_16393,N_14364,N_11305);
or U16394 (N_16394,N_11185,N_10081);
or U16395 (N_16395,N_10312,N_13439);
and U16396 (N_16396,N_11596,N_12763);
and U16397 (N_16397,N_14160,N_11667);
or U16398 (N_16398,N_13672,N_13921);
nor U16399 (N_16399,N_10326,N_13569);
or U16400 (N_16400,N_11072,N_13010);
nor U16401 (N_16401,N_14520,N_12897);
nand U16402 (N_16402,N_14812,N_12999);
or U16403 (N_16403,N_14146,N_11105);
nor U16404 (N_16404,N_11702,N_13005);
nand U16405 (N_16405,N_10264,N_14264);
and U16406 (N_16406,N_12595,N_12525);
xnor U16407 (N_16407,N_11299,N_13232);
xnor U16408 (N_16408,N_12825,N_13105);
or U16409 (N_16409,N_10166,N_13399);
and U16410 (N_16410,N_12262,N_10133);
nor U16411 (N_16411,N_11142,N_10253);
nand U16412 (N_16412,N_12396,N_12175);
nor U16413 (N_16413,N_13646,N_13241);
nand U16414 (N_16414,N_12516,N_13641);
nor U16415 (N_16415,N_14517,N_12537);
or U16416 (N_16416,N_14133,N_14731);
nand U16417 (N_16417,N_14539,N_10958);
or U16418 (N_16418,N_13293,N_14705);
nor U16419 (N_16419,N_11432,N_13504);
xor U16420 (N_16420,N_11710,N_13593);
or U16421 (N_16421,N_10270,N_12893);
or U16422 (N_16422,N_11202,N_14945);
nor U16423 (N_16423,N_11534,N_10902);
nor U16424 (N_16424,N_11864,N_12960);
and U16425 (N_16425,N_13176,N_12215);
or U16426 (N_16426,N_14881,N_13099);
nand U16427 (N_16427,N_11519,N_13316);
nand U16428 (N_16428,N_14142,N_12035);
xor U16429 (N_16429,N_14739,N_10430);
nand U16430 (N_16430,N_13821,N_14119);
and U16431 (N_16431,N_14471,N_13750);
nor U16432 (N_16432,N_11247,N_14561);
and U16433 (N_16433,N_14839,N_12860);
and U16434 (N_16434,N_12239,N_14372);
nor U16435 (N_16435,N_13263,N_12625);
nand U16436 (N_16436,N_12752,N_10912);
xnor U16437 (N_16437,N_14028,N_10911);
nand U16438 (N_16438,N_10507,N_11236);
nand U16439 (N_16439,N_14246,N_13549);
or U16440 (N_16440,N_12821,N_10018);
xor U16441 (N_16441,N_10612,N_12042);
and U16442 (N_16442,N_13684,N_14784);
xor U16443 (N_16443,N_11491,N_14810);
or U16444 (N_16444,N_12718,N_14611);
and U16445 (N_16445,N_12552,N_11065);
nand U16446 (N_16446,N_10050,N_14775);
xor U16447 (N_16447,N_10656,N_11993);
or U16448 (N_16448,N_11866,N_11699);
or U16449 (N_16449,N_10242,N_12328);
and U16450 (N_16450,N_14824,N_13876);
or U16451 (N_16451,N_10877,N_12624);
or U16452 (N_16452,N_14170,N_11241);
nor U16453 (N_16453,N_10000,N_13768);
and U16454 (N_16454,N_13495,N_14963);
and U16455 (N_16455,N_13103,N_10603);
nand U16456 (N_16456,N_10945,N_12890);
xor U16457 (N_16457,N_14447,N_13365);
nor U16458 (N_16458,N_12634,N_10485);
and U16459 (N_16459,N_12836,N_12495);
nor U16460 (N_16460,N_10235,N_10438);
or U16461 (N_16461,N_14166,N_10225);
xor U16462 (N_16462,N_12298,N_10011);
or U16463 (N_16463,N_12774,N_10637);
xnor U16464 (N_16464,N_10472,N_14747);
xnor U16465 (N_16465,N_12198,N_10036);
nand U16466 (N_16466,N_11445,N_10109);
nand U16467 (N_16467,N_12538,N_14911);
nand U16468 (N_16468,N_12224,N_12210);
and U16469 (N_16469,N_11198,N_10917);
nand U16470 (N_16470,N_14432,N_12218);
nor U16471 (N_16471,N_12482,N_12420);
xor U16472 (N_16472,N_10723,N_12023);
or U16473 (N_16473,N_11870,N_12058);
and U16474 (N_16474,N_12233,N_13544);
nor U16475 (N_16475,N_13566,N_11071);
nand U16476 (N_16476,N_14862,N_12011);
nor U16477 (N_16477,N_12081,N_11748);
xor U16478 (N_16478,N_10181,N_10605);
nand U16479 (N_16479,N_13787,N_14229);
nor U16480 (N_16480,N_10276,N_14661);
or U16481 (N_16481,N_11613,N_11651);
and U16482 (N_16482,N_12950,N_11649);
and U16483 (N_16483,N_10592,N_11015);
nor U16484 (N_16484,N_11300,N_12904);
xor U16485 (N_16485,N_13028,N_12047);
nand U16486 (N_16486,N_13032,N_11593);
nor U16487 (N_16487,N_11556,N_12012);
nand U16488 (N_16488,N_11816,N_11778);
xor U16489 (N_16489,N_10713,N_10704);
and U16490 (N_16490,N_11834,N_13009);
xor U16491 (N_16491,N_10845,N_13074);
nor U16492 (N_16492,N_13341,N_10143);
nand U16493 (N_16493,N_13932,N_12909);
xor U16494 (N_16494,N_14598,N_14995);
nor U16495 (N_16495,N_12891,N_11910);
or U16496 (N_16496,N_11536,N_12693);
nand U16497 (N_16497,N_14569,N_12700);
and U16498 (N_16498,N_11138,N_14053);
nor U16499 (N_16499,N_11506,N_13441);
nand U16500 (N_16500,N_12691,N_12998);
nor U16501 (N_16501,N_10125,N_14738);
nor U16502 (N_16502,N_13584,N_13185);
nand U16503 (N_16503,N_11749,N_11488);
nand U16504 (N_16504,N_13799,N_14116);
or U16505 (N_16505,N_12139,N_10498);
or U16506 (N_16506,N_14758,N_10442);
nor U16507 (N_16507,N_10771,N_14314);
and U16508 (N_16508,N_14194,N_13761);
nand U16509 (N_16509,N_11448,N_13650);
and U16510 (N_16510,N_12738,N_10468);
and U16511 (N_16511,N_13729,N_11638);
nor U16512 (N_16512,N_13673,N_12567);
and U16513 (N_16513,N_11403,N_11449);
xnor U16514 (N_16514,N_11223,N_11406);
and U16515 (N_16515,N_12091,N_11670);
nand U16516 (N_16516,N_11737,N_11154);
xor U16517 (N_16517,N_13585,N_14551);
nor U16518 (N_16518,N_10729,N_12727);
nand U16519 (N_16519,N_11641,N_11190);
nor U16520 (N_16520,N_11208,N_11907);
and U16521 (N_16521,N_12497,N_14959);
xnor U16522 (N_16522,N_11751,N_12748);
nand U16523 (N_16523,N_12575,N_11770);
or U16524 (N_16524,N_12444,N_12440);
nor U16525 (N_16525,N_13576,N_10393);
nand U16526 (N_16526,N_13701,N_13807);
nor U16527 (N_16527,N_12345,N_12116);
nor U16528 (N_16528,N_14060,N_11875);
xnor U16529 (N_16529,N_10918,N_11477);
xor U16530 (N_16530,N_11077,N_10919);
and U16531 (N_16531,N_11764,N_12551);
or U16532 (N_16532,N_11478,N_13398);
nor U16533 (N_16533,N_11222,N_11530);
nand U16534 (N_16534,N_10931,N_13202);
or U16535 (N_16535,N_13244,N_14443);
nor U16536 (N_16536,N_14267,N_14180);
or U16537 (N_16537,N_12918,N_11591);
or U16538 (N_16538,N_12714,N_11439);
nand U16539 (N_16539,N_13494,N_11511);
nor U16540 (N_16540,N_11393,N_12077);
or U16541 (N_16541,N_13754,N_13637);
nor U16542 (N_16542,N_11431,N_13713);
nand U16543 (N_16543,N_11507,N_10085);
and U16544 (N_16544,N_13055,N_12302);
or U16545 (N_16545,N_10131,N_14408);
or U16546 (N_16546,N_12479,N_11344);
xnor U16547 (N_16547,N_13749,N_14384);
xor U16548 (N_16548,N_10057,N_13506);
nand U16549 (N_16549,N_11630,N_13617);
xor U16550 (N_16550,N_12566,N_14036);
nand U16551 (N_16551,N_14416,N_10063);
nor U16552 (N_16552,N_11895,N_14354);
nand U16553 (N_16553,N_14894,N_13102);
nor U16554 (N_16554,N_13619,N_10999);
nand U16555 (N_16555,N_12038,N_14836);
and U16556 (N_16556,N_10229,N_10291);
nand U16557 (N_16557,N_11522,N_10512);
and U16558 (N_16558,N_11911,N_13194);
nand U16559 (N_16559,N_11808,N_13237);
xnor U16560 (N_16560,N_13356,N_12892);
or U16561 (N_16561,N_11959,N_13256);
or U16562 (N_16562,N_10715,N_13831);
xor U16563 (N_16563,N_14419,N_13490);
or U16564 (N_16564,N_14020,N_14579);
nand U16565 (N_16565,N_12119,N_13258);
or U16566 (N_16566,N_12046,N_12297);
nor U16567 (N_16567,N_12422,N_10405);
and U16568 (N_16568,N_13418,N_13530);
nor U16569 (N_16569,N_11761,N_12499);
or U16570 (N_16570,N_13918,N_12559);
xnor U16571 (N_16571,N_10217,N_11797);
and U16572 (N_16572,N_11058,N_10020);
and U16573 (N_16573,N_12281,N_14753);
and U16574 (N_16574,N_13079,N_13545);
or U16575 (N_16575,N_11415,N_11852);
nor U16576 (N_16576,N_13457,N_14653);
nor U16577 (N_16577,N_14596,N_11345);
or U16578 (N_16578,N_12834,N_13935);
xor U16579 (N_16579,N_14097,N_11321);
nand U16580 (N_16580,N_14249,N_13997);
nand U16581 (N_16581,N_14276,N_14769);
xor U16582 (N_16582,N_10515,N_11552);
or U16583 (N_16583,N_14761,N_11944);
and U16584 (N_16584,N_13113,N_14156);
or U16585 (N_16585,N_13035,N_11912);
or U16586 (N_16586,N_12133,N_10370);
xor U16587 (N_16587,N_12176,N_10926);
nand U16588 (N_16588,N_12045,N_10526);
and U16589 (N_16589,N_10396,N_11171);
nor U16590 (N_16590,N_14555,N_14190);
nor U16591 (N_16591,N_10424,N_12098);
and U16592 (N_16592,N_11128,N_12706);
and U16593 (N_16593,N_10295,N_13636);
nor U16594 (N_16594,N_13864,N_13325);
nor U16595 (N_16595,N_13887,N_11205);
or U16596 (N_16596,N_11358,N_10045);
nor U16597 (N_16597,N_10460,N_14846);
and U16598 (N_16598,N_11302,N_13022);
and U16599 (N_16599,N_13886,N_13066);
and U16600 (N_16600,N_10760,N_11382);
xnor U16601 (N_16601,N_10595,N_14664);
nand U16602 (N_16602,N_10505,N_10028);
or U16603 (N_16603,N_12707,N_12300);
nand U16604 (N_16604,N_14662,N_10488);
and U16605 (N_16605,N_10123,N_11139);
nor U16606 (N_16606,N_13134,N_10594);
or U16607 (N_16607,N_12315,N_14398);
nand U16608 (N_16608,N_14401,N_10798);
xnor U16609 (N_16609,N_11008,N_14316);
nand U16610 (N_16610,N_10525,N_10961);
and U16611 (N_16611,N_12060,N_11672);
xnor U16612 (N_16612,N_12167,N_12138);
and U16613 (N_16613,N_12295,N_14607);
nand U16614 (N_16614,N_14768,N_12652);
or U16615 (N_16615,N_14906,N_14680);
and U16616 (N_16616,N_12853,N_12965);
nor U16617 (N_16617,N_12163,N_10121);
nor U16618 (N_16618,N_11182,N_12354);
nor U16619 (N_16619,N_12459,N_13767);
and U16620 (N_16620,N_10583,N_14073);
or U16621 (N_16621,N_11220,N_12103);
or U16622 (N_16622,N_10762,N_10115);
nand U16623 (N_16623,N_11765,N_10674);
nor U16624 (N_16624,N_12487,N_14601);
nor U16625 (N_16625,N_11328,N_10528);
and U16626 (N_16626,N_11882,N_10977);
xnor U16627 (N_16627,N_11172,N_14454);
xnor U16628 (N_16628,N_10516,N_12815);
nor U16629 (N_16629,N_13450,N_14833);
or U16630 (N_16630,N_11371,N_12027);
or U16631 (N_16631,N_12463,N_14356);
xor U16632 (N_16632,N_12402,N_10775);
nand U16633 (N_16633,N_11909,N_12724);
xor U16634 (N_16634,N_10944,N_11538);
xor U16635 (N_16635,N_11535,N_14702);
or U16636 (N_16636,N_12835,N_14827);
or U16637 (N_16637,N_14818,N_14623);
xor U16638 (N_16638,N_10382,N_10696);
nand U16639 (N_16639,N_13327,N_13907);
nand U16640 (N_16640,N_11626,N_13866);
xor U16641 (N_16641,N_14955,N_11129);
nor U16642 (N_16642,N_13342,N_11084);
xnor U16643 (N_16643,N_13536,N_13960);
nor U16644 (N_16644,N_12721,N_11169);
and U16645 (N_16645,N_11283,N_13155);
or U16646 (N_16646,N_10223,N_10183);
and U16647 (N_16647,N_12486,N_10174);
or U16648 (N_16648,N_10068,N_13236);
nor U16649 (N_16649,N_10328,N_14861);
nand U16650 (N_16650,N_11663,N_11265);
and U16651 (N_16651,N_13409,N_10101);
or U16652 (N_16652,N_14711,N_10346);
or U16653 (N_16653,N_11932,N_11079);
and U16654 (N_16654,N_11692,N_10377);
and U16655 (N_16655,N_14478,N_10499);
xor U16656 (N_16656,N_10269,N_11560);
xor U16657 (N_16657,N_14842,N_13411);
or U16658 (N_16658,N_12926,N_14233);
and U16659 (N_16659,N_14605,N_13440);
and U16660 (N_16660,N_11434,N_10373);
and U16661 (N_16661,N_14907,N_11174);
and U16662 (N_16662,N_11152,N_13045);
xnor U16663 (N_16663,N_13751,N_10406);
nand U16664 (N_16664,N_12514,N_13662);
nor U16665 (N_16665,N_10863,N_11810);
nor U16666 (N_16666,N_12320,N_12997);
and U16667 (N_16667,N_12323,N_12249);
xnor U16668 (N_16668,N_14129,N_13427);
and U16669 (N_16669,N_10097,N_14388);
or U16670 (N_16670,N_13803,N_10142);
xor U16671 (N_16671,N_14987,N_14639);
nand U16672 (N_16672,N_12553,N_11963);
xor U16673 (N_16673,N_10390,N_14946);
nor U16674 (N_16674,N_13994,N_13535);
xnor U16675 (N_16675,N_11212,N_11464);
nand U16676 (N_16676,N_14927,N_14034);
nor U16677 (N_16677,N_14840,N_11493);
nor U16678 (N_16678,N_13212,N_13266);
nand U16679 (N_16679,N_11291,N_10755);
or U16680 (N_16680,N_14652,N_13848);
or U16681 (N_16681,N_11545,N_10823);
nor U16682 (N_16682,N_14791,N_10341);
and U16683 (N_16683,N_12351,N_13046);
xnor U16684 (N_16684,N_10559,N_14736);
nor U16685 (N_16685,N_10645,N_11580);
xor U16686 (N_16686,N_13031,N_13862);
nand U16687 (N_16687,N_11997,N_10357);
or U16688 (N_16688,N_10557,N_13002);
or U16689 (N_16689,N_13012,N_14009);
xor U16690 (N_16690,N_10043,N_10930);
nor U16691 (N_16691,N_12861,N_11644);
nand U16692 (N_16692,N_13624,N_11595);
xnor U16693 (N_16693,N_10904,N_11410);
or U16694 (N_16694,N_13786,N_13678);
or U16695 (N_16695,N_12735,N_14213);
xor U16696 (N_16696,N_12604,N_14185);
and U16697 (N_16697,N_10267,N_14235);
nand U16698 (N_16698,N_12789,N_13408);
and U16699 (N_16699,N_13664,N_14658);
nor U16700 (N_16700,N_14391,N_13951);
or U16701 (N_16701,N_10935,N_10970);
nor U16702 (N_16702,N_13806,N_11323);
or U16703 (N_16703,N_14072,N_10895);
or U16704 (N_16704,N_14899,N_10658);
or U16705 (N_16705,N_11041,N_14542);
and U16706 (N_16706,N_12924,N_12391);
and U16707 (N_16707,N_11938,N_10185);
nor U16708 (N_16708,N_13319,N_13451);
nand U16709 (N_16709,N_13709,N_10520);
and U16710 (N_16710,N_10450,N_11083);
or U16711 (N_16711,N_14197,N_14586);
nand U16712 (N_16712,N_12374,N_12667);
or U16713 (N_16713,N_11677,N_11304);
or U16714 (N_16714,N_12448,N_13879);
xnor U16715 (N_16715,N_13958,N_14521);
xor U16716 (N_16716,N_13603,N_13922);
xnor U16717 (N_16717,N_10338,N_11273);
and U16718 (N_16718,N_12974,N_11339);
nor U16719 (N_16719,N_11061,N_13489);
or U16720 (N_16720,N_14900,N_14082);
or U16721 (N_16721,N_14203,N_10163);
xnor U16722 (N_16722,N_13249,N_14085);
nand U16723 (N_16723,N_13724,N_14511);
or U16724 (N_16724,N_14690,N_11786);
or U16725 (N_16725,N_10950,N_10558);
nand U16726 (N_16726,N_12013,N_14502);
and U16727 (N_16727,N_11780,N_14283);
xor U16728 (N_16728,N_14453,N_12153);
nand U16729 (N_16729,N_11722,N_14309);
nor U16730 (N_16730,N_12280,N_11056);
or U16731 (N_16731,N_14871,N_13330);
nand U16732 (N_16732,N_11679,N_12294);
nor U16733 (N_16733,N_13361,N_13027);
and U16734 (N_16734,N_12373,N_13153);
xor U16735 (N_16735,N_14325,N_11998);
and U16736 (N_16736,N_12333,N_11564);
nor U16737 (N_16737,N_12539,N_12134);
xor U16738 (N_16738,N_14161,N_11274);
and U16739 (N_16739,N_12240,N_14636);
nand U16740 (N_16740,N_11495,N_11396);
nand U16741 (N_16741,N_10969,N_11684);
or U16742 (N_16742,N_14614,N_10566);
or U16743 (N_16743,N_14476,N_13523);
or U16744 (N_16744,N_14619,N_13370);
nor U16745 (N_16745,N_13147,N_13109);
and U16746 (N_16746,N_12986,N_11404);
nand U16747 (N_16747,N_11398,N_12429);
or U16748 (N_16748,N_13983,N_14508);
and U16749 (N_16749,N_14083,N_13382);
nor U16750 (N_16750,N_13226,N_11476);
and U16751 (N_16751,N_14483,N_12325);
or U16752 (N_16752,N_10327,N_14350);
or U16753 (N_16753,N_10117,N_14293);
nand U16754 (N_16754,N_11148,N_14074);
nand U16755 (N_16755,N_13519,N_13765);
and U16756 (N_16756,N_11879,N_13945);
or U16757 (N_16757,N_12057,N_14951);
or U16758 (N_16758,N_14417,N_12745);
xnor U16759 (N_16759,N_13533,N_12256);
and U16760 (N_16760,N_14566,N_11503);
nor U16761 (N_16761,N_10180,N_11914);
nand U16762 (N_16762,N_10548,N_13460);
nor U16763 (N_16763,N_11426,N_11960);
nor U16764 (N_16764,N_11092,N_11120);
nand U16765 (N_16765,N_13953,N_13433);
or U16766 (N_16766,N_12393,N_10116);
nand U16767 (N_16767,N_14973,N_12921);
or U16768 (N_16768,N_11347,N_12712);
nor U16769 (N_16769,N_10685,N_13184);
and U16770 (N_16770,N_11483,N_10361);
xnor U16771 (N_16771,N_14982,N_11051);
xor U16772 (N_16772,N_13663,N_12137);
nand U16773 (N_16773,N_12807,N_10271);
or U16774 (N_16774,N_14600,N_11035);
nand U16775 (N_16775,N_12663,N_11640);
and U16776 (N_16776,N_14212,N_11002);
or U16777 (N_16777,N_10459,N_12149);
nand U16778 (N_16778,N_11851,N_12542);
xor U16779 (N_16779,N_12484,N_13182);
nor U16780 (N_16780,N_10568,N_13604);
nor U16781 (N_16781,N_10091,N_12212);
nor U16782 (N_16782,N_13312,N_12659);
nor U16783 (N_16783,N_14379,N_11201);
nor U16784 (N_16784,N_12413,N_10689);
and U16785 (N_16785,N_12270,N_11539);
nand U16786 (N_16786,N_11937,N_12784);
xnor U16787 (N_16787,N_14960,N_13139);
or U16788 (N_16788,N_13152,N_14237);
nand U16789 (N_16789,N_13394,N_10420);
or U16790 (N_16790,N_13484,N_11829);
nand U16791 (N_16791,N_11004,N_11023);
nor U16792 (N_16792,N_10336,N_11617);
or U16793 (N_16793,N_10311,N_11233);
xnor U16794 (N_16794,N_13695,N_12464);
xor U16795 (N_16795,N_11615,N_11261);
or U16796 (N_16796,N_10265,N_12954);
nor U16797 (N_16797,N_12695,N_10345);
nor U16798 (N_16798,N_13069,N_14281);
nor U16799 (N_16799,N_14378,N_11411);
xor U16800 (N_16800,N_10764,N_14650);
or U16801 (N_16801,N_10415,N_13870);
nor U16802 (N_16802,N_10359,N_11849);
or U16803 (N_16803,N_10873,N_12641);
or U16804 (N_16804,N_13596,N_12355);
or U16805 (N_16805,N_14109,N_13830);
nand U16806 (N_16806,N_12722,N_13962);
and U16807 (N_16807,N_11353,N_14433);
or U16808 (N_16808,N_14637,N_10437);
nor U16809 (N_16809,N_14207,N_12592);
xor U16810 (N_16810,N_10561,N_12716);
and U16811 (N_16811,N_13363,N_14348);
or U16812 (N_16812,N_11093,N_11374);
nor U16813 (N_16813,N_14778,N_13902);
nor U16814 (N_16814,N_13141,N_13446);
or U16815 (N_16815,N_10769,N_12052);
xnor U16816 (N_16816,N_14538,N_11582);
xor U16817 (N_16817,N_12418,N_13660);
and U16818 (N_16818,N_12086,N_11017);
xor U16819 (N_16819,N_13058,N_14341);
and U16820 (N_16820,N_12605,N_13735);
or U16821 (N_16821,N_10639,N_13204);
or U16822 (N_16822,N_14466,N_10812);
nor U16823 (N_16823,N_12558,N_11123);
xor U16824 (N_16824,N_10654,N_10380);
and U16825 (N_16825,N_12952,N_13025);
xor U16826 (N_16826,N_14628,N_13560);
or U16827 (N_16827,N_14086,N_10106);
nor U16828 (N_16828,N_14934,N_13620);
and U16829 (N_16829,N_10462,N_13613);
nand U16830 (N_16830,N_12309,N_14556);
nor U16831 (N_16831,N_10321,N_11924);
xor U16832 (N_16832,N_14725,N_14429);
xnor U16833 (N_16833,N_14245,N_14789);
or U16834 (N_16834,N_13892,N_14968);
nand U16835 (N_16835,N_13756,N_11843);
nor U16836 (N_16836,N_11685,N_11775);
nor U16837 (N_16837,N_11521,N_13163);
xor U16838 (N_16838,N_13097,N_10927);
and U16839 (N_16839,N_14439,N_10219);
nand U16840 (N_16840,N_13811,N_10693);
or U16841 (N_16841,N_10564,N_12017);
or U16842 (N_16842,N_13050,N_10702);
or U16843 (N_16843,N_11355,N_12636);
and U16844 (N_16844,N_14113,N_10622);
or U16845 (N_16845,N_12878,N_11719);
and U16846 (N_16846,N_12109,N_12190);
nor U16847 (N_16847,N_11982,N_14612);
nand U16848 (N_16848,N_13880,N_14668);
xor U16849 (N_16849,N_14339,N_12948);
xor U16850 (N_16850,N_13992,N_12254);
xnor U16851 (N_16851,N_14889,N_13444);
nor U16852 (N_16852,N_12597,N_11253);
xor U16853 (N_16853,N_11880,N_13804);
and U16854 (N_16854,N_14340,N_12660);
and U16855 (N_16855,N_11850,N_10619);
xnor U16856 (N_16856,N_11385,N_10738);
and U16857 (N_16857,N_11354,N_13970);
and U16858 (N_16858,N_11662,N_10813);
xor U16859 (N_16859,N_11859,N_10901);
or U16860 (N_16860,N_10735,N_12521);
and U16861 (N_16861,N_11243,N_13850);
and U16862 (N_16862,N_11486,N_11245);
and U16863 (N_16863,N_10284,N_14286);
and U16864 (N_16864,N_10538,N_14500);
nor U16865 (N_16865,N_13353,N_14118);
xor U16866 (N_16866,N_14090,N_10782);
xor U16867 (N_16867,N_13265,N_12192);
xnor U16868 (N_16868,N_13313,N_11729);
nor U16869 (N_16869,N_12319,N_14713);
nor U16870 (N_16870,N_13634,N_10889);
and U16871 (N_16871,N_14396,N_12020);
nand U16872 (N_16872,N_12850,N_13329);
and U16873 (N_16873,N_13148,N_14038);
nor U16874 (N_16874,N_11897,N_13061);
nand U16875 (N_16875,N_14329,N_13591);
and U16876 (N_16876,N_13869,N_14330);
xnor U16877 (N_16877,N_11256,N_12164);
nand U16878 (N_16878,N_10915,N_14243);
or U16879 (N_16879,N_12818,N_13564);
and U16880 (N_16880,N_11131,N_13777);
or U16881 (N_16881,N_12591,N_12811);
xor U16882 (N_16882,N_12971,N_12015);
and U16883 (N_16883,N_11871,N_12644);
nor U16884 (N_16884,N_13429,N_11089);
or U16885 (N_16885,N_12787,N_13954);
xor U16886 (N_16886,N_14112,N_13008);
nand U16887 (N_16887,N_12580,N_10306);
nand U16888 (N_16888,N_12050,N_10475);
xor U16889 (N_16889,N_10602,N_10633);
nand U16890 (N_16890,N_12493,N_11804);
or U16891 (N_16891,N_14031,N_12760);
and U16892 (N_16892,N_14304,N_10298);
xnor U16893 (N_16893,N_12016,N_12608);
nor U16894 (N_16894,N_14427,N_10051);
xnor U16895 (N_16895,N_14434,N_14727);
and U16896 (N_16896,N_10758,N_12055);
and U16897 (N_16897,N_13776,N_14077);
and U16898 (N_16898,N_10309,N_13820);
and U16899 (N_16899,N_14998,N_14179);
xnor U16900 (N_16900,N_12709,N_11948);
or U16901 (N_16901,N_10060,N_11268);
or U16902 (N_16902,N_14913,N_13924);
nor U16903 (N_16903,N_14421,N_10368);
or U16904 (N_16904,N_11480,N_10318);
and U16905 (N_16905,N_13034,N_12341);
xor U16906 (N_16906,N_14576,N_13259);
and U16907 (N_16907,N_13884,N_11781);
or U16908 (N_16908,N_11242,N_11769);
nand U16909 (N_16909,N_14554,N_13309);
and U16910 (N_16910,N_12697,N_12682);
xnor U16911 (N_16911,N_12306,N_11890);
or U16912 (N_16912,N_12520,N_10643);
or U16913 (N_16913,N_11441,N_12043);
xor U16914 (N_16914,N_13242,N_10743);
or U16915 (N_16915,N_10402,N_12469);
and U16916 (N_16916,N_14126,N_11523);
nand U16917 (N_16917,N_11391,N_12085);
or U16918 (N_16918,N_13114,N_13463);
and U16919 (N_16919,N_14574,N_10240);
xnor U16920 (N_16920,N_14270,N_13294);
and U16921 (N_16921,N_14499,N_10929);
xor U16922 (N_16922,N_14939,N_14876);
or U16923 (N_16923,N_13391,N_12223);
or U16924 (N_16924,N_13849,N_14092);
xor U16925 (N_16925,N_13704,N_12702);
xor U16926 (N_16926,N_14361,N_13107);
nor U16927 (N_16927,N_13021,N_10140);
xnor U16928 (N_16928,N_10029,N_10644);
and U16929 (N_16929,N_10419,N_14026);
and U16930 (N_16930,N_11357,N_14257);
xor U16931 (N_16931,N_13505,N_11390);
nand U16932 (N_16932,N_13165,N_13712);
nand U16933 (N_16933,N_14291,N_13563);
nand U16934 (N_16934,N_11121,N_12205);
nand U16935 (N_16935,N_13437,N_13653);
and U16936 (N_16936,N_13089,N_14108);
or U16937 (N_16937,N_11318,N_14868);
nor U16938 (N_16938,N_14651,N_14564);
and U16939 (N_16939,N_12473,N_13651);
xor U16940 (N_16940,N_12285,N_12846);
or U16941 (N_16941,N_13551,N_14470);
nand U16942 (N_16942,N_13885,N_10597);
and U16943 (N_16943,N_12476,N_10322);
nor U16944 (N_16944,N_11271,N_10221);
xor U16945 (N_16945,N_11520,N_10607);
xor U16946 (N_16946,N_14018,N_11106);
or U16947 (N_16947,N_12895,N_14461);
and U16948 (N_16948,N_11457,N_11013);
nand U16949 (N_16949,N_10923,N_13537);
and U16950 (N_16950,N_11958,N_14256);
or U16951 (N_16951,N_13379,N_14962);
and U16952 (N_16952,N_12705,N_13638);
or U16953 (N_16953,N_11492,N_10209);
or U16954 (N_16954,N_10350,N_14334);
or U16955 (N_16955,N_14553,N_14294);
nand U16956 (N_16956,N_13540,N_12549);
nor U16957 (N_16957,N_13387,N_12571);
nor U16958 (N_16958,N_14140,N_11669);
nor U16959 (N_16959,N_13135,N_12598);
nand U16960 (N_16960,N_14844,N_10076);
xor U16961 (N_16961,N_14807,N_14767);
and U16962 (N_16962,N_14772,N_14675);
xnor U16963 (N_16963,N_10865,N_11570);
or U16964 (N_16964,N_10796,N_10834);
and U16965 (N_16965,N_10465,N_11356);
nand U16966 (N_16966,N_14788,N_12095);
xor U16967 (N_16967,N_10661,N_12742);
nor U16968 (N_16968,N_10015,N_11456);
and U16969 (N_16969,N_10830,N_11377);
xor U16970 (N_16970,N_14760,N_13546);
nor U16971 (N_16971,N_14165,N_11602);
xor U16972 (N_16972,N_11991,N_11585);
and U16973 (N_16973,N_14646,N_13647);
nor U16974 (N_16974,N_14594,N_14931);
and U16975 (N_16975,N_11791,N_11157);
xnor U16976 (N_16976,N_13485,N_12186);
nor U16977 (N_16977,N_14673,N_13600);
nor U16978 (N_16978,N_13261,N_12798);
nand U16979 (N_16979,N_11688,N_11276);
or U16980 (N_16980,N_13691,N_11971);
xor U16981 (N_16981,N_13654,N_10222);
or U16982 (N_16982,N_12867,N_11952);
and U16983 (N_16983,N_13875,N_10237);
or U16984 (N_16984,N_12854,N_10323);
xor U16985 (N_16985,N_12802,N_13404);
nor U16986 (N_16986,N_11996,N_13129);
xor U16987 (N_16987,N_13714,N_12502);
nand U16988 (N_16988,N_14202,N_10825);
or U16989 (N_16989,N_11111,N_12410);
nor U16990 (N_16990,N_10009,N_11660);
xnor U16991 (N_16991,N_13681,N_12458);
nand U16992 (N_16992,N_11533,N_11696);
nand U16993 (N_16993,N_12466,N_11592);
and U16994 (N_16994,N_14613,N_12304);
xor U16995 (N_16995,N_10391,N_13137);
or U16996 (N_16996,N_12949,N_10533);
and U16997 (N_16997,N_10386,N_13897);
nand U16998 (N_16998,N_11983,N_11858);
or U16999 (N_16999,N_12166,N_11928);
xor U17000 (N_17000,N_11026,N_10763);
nor U17001 (N_17001,N_12386,N_12062);
and U17002 (N_17002,N_12021,N_13801);
or U17003 (N_17003,N_12832,N_12180);
nand U17004 (N_17004,N_13645,N_12833);
or U17005 (N_17005,N_13161,N_11826);
xor U17006 (N_17006,N_11430,N_10981);
and U17007 (N_17007,N_14558,N_12668);
or U17008 (N_17008,N_12857,N_14234);
nand U17009 (N_17009,N_11886,N_12692);
and U17010 (N_17010,N_13043,N_10721);
nand U17011 (N_17011,N_12703,N_12468);
nor U17012 (N_17012,N_13857,N_13291);
and U17013 (N_17013,N_14580,N_14313);
nand U17014 (N_17014,N_13788,N_14484);
xnor U17015 (N_17015,N_11528,N_11607);
nand U17016 (N_17016,N_11161,N_12896);
xnor U17017 (N_17017,N_14820,N_11955);
nor U17018 (N_17018,N_11818,N_11603);
nor U17019 (N_17019,N_14136,N_14487);
xnor U17020 (N_17020,N_11935,N_12548);
xor U17021 (N_17021,N_11964,N_14855);
xnor U17022 (N_17022,N_12124,N_11762);
and U17023 (N_17023,N_14648,N_13217);
xor U17024 (N_17024,N_10385,N_13098);
nor U17025 (N_17025,N_14319,N_12427);
or U17026 (N_17026,N_12527,N_10749);
nor U17027 (N_17027,N_13104,N_14130);
nand U17028 (N_17028,N_13235,N_14002);
nand U17029 (N_17029,N_12848,N_12809);
and U17030 (N_17030,N_12961,N_11957);
nand U17031 (N_17031,N_10717,N_10001);
xnor U17032 (N_17032,N_10826,N_11240);
or U17033 (N_17033,N_10941,N_13208);
nand U17034 (N_17034,N_10978,N_10579);
xor U17035 (N_17035,N_14522,N_10044);
or U17036 (N_17036,N_13304,N_13435);
xor U17037 (N_17037,N_14248,N_11482);
or U17038 (N_17038,N_13773,N_11962);
xor U17039 (N_17039,N_11977,N_14671);
and U17040 (N_17040,N_11622,N_13358);
nand U17041 (N_17041,N_12189,N_12686);
nor U17042 (N_17042,N_10159,N_12475);
or U17043 (N_17043,N_13024,N_13728);
nor U17044 (N_17044,N_14196,N_11949);
or U17045 (N_17045,N_12739,N_11690);
xor U17046 (N_17046,N_12261,N_10809);
and U17047 (N_17047,N_11608,N_12791);
or U17048 (N_17048,N_14712,N_12744);
or U17049 (N_17049,N_10070,N_12779);
nand U17050 (N_17050,N_12039,N_10788);
or U17051 (N_17051,N_12417,N_13690);
nand U17052 (N_17052,N_12407,N_13076);
nand U17053 (N_17053,N_12743,N_11375);
xor U17054 (N_17054,N_14346,N_12574);
nand U17055 (N_17055,N_14260,N_14676);
nor U17056 (N_17056,N_14263,N_12788);
or U17057 (N_17057,N_10381,N_14360);
nand U17058 (N_17058,N_12710,N_10399);
nand U17059 (N_17059,N_11047,N_13195);
xnor U17060 (N_17060,N_13143,N_11076);
or U17061 (N_17061,N_14966,N_12945);
and U17062 (N_17062,N_13230,N_14793);
or U17063 (N_17063,N_13186,N_12204);
and U17064 (N_17064,N_12245,N_14000);
and U17065 (N_17065,N_10258,N_12649);
or U17066 (N_17066,N_13890,N_14176);
nor U17067 (N_17067,N_10178,N_12725);
xnor U17068 (N_17068,N_10423,N_12127);
xor U17069 (N_17069,N_11389,N_12504);
nand U17070 (N_17070,N_13048,N_14759);
xnor U17071 (N_17071,N_13721,N_12908);
xnor U17072 (N_17072,N_14930,N_11081);
nor U17073 (N_17073,N_11423,N_12312);
or U17074 (N_17074,N_13648,N_13926);
xor U17075 (N_17075,N_12316,N_11867);
nor U17076 (N_17076,N_13514,N_13030);
nand U17077 (N_17077,N_13779,N_10503);
and U17078 (N_17078,N_13081,N_10400);
nand U17079 (N_17079,N_11298,N_12862);
nor U17080 (N_17080,N_14333,N_10023);
nand U17081 (N_17081,N_11594,N_12830);
and U17082 (N_17082,N_12242,N_14064);
xor U17083 (N_17083,N_11908,N_11095);
and U17084 (N_17084,N_10135,N_11115);
and U17085 (N_17085,N_13778,N_12977);
nor U17086 (N_17086,N_10279,N_12719);
nand U17087 (N_17087,N_14865,N_12839);
nor U17088 (N_17088,N_12162,N_14289);
nand U17089 (N_17089,N_11238,N_10411);
nand U17090 (N_17090,N_12920,N_12639);
xnor U17091 (N_17091,N_13675,N_10453);
xnor U17092 (N_17092,N_14173,N_10534);
or U17093 (N_17093,N_11813,N_12425);
nor U17094 (N_17094,N_13498,N_14583);
or U17095 (N_17095,N_10663,N_11604);
or U17096 (N_17096,N_11750,N_12340);
nand U17097 (N_17097,N_12184,N_13623);
and U17098 (N_17098,N_13073,N_14152);
or U17099 (N_17099,N_11508,N_13670);
and U17100 (N_17100,N_12084,N_12196);
xor U17101 (N_17101,N_12122,N_11203);
xnor U17102 (N_17102,N_13833,N_14321);
or U17103 (N_17103,N_10152,N_11369);
xnor U17104 (N_17104,N_13944,N_14541);
and U17105 (N_17105,N_10272,N_13570);
and U17106 (N_17106,N_11163,N_11024);
and U17107 (N_17107,N_11005,N_11284);
and U17108 (N_17108,N_14225,N_14718);
or U17109 (N_17109,N_11973,N_10728);
or U17110 (N_17110,N_13122,N_11940);
or U17111 (N_17111,N_13940,N_13180);
or U17112 (N_17112,N_13448,N_10886);
nor U17113 (N_17113,N_11833,N_13385);
and U17114 (N_17114,N_13269,N_12228);
and U17115 (N_17115,N_12540,N_14358);
nor U17116 (N_17116,N_12755,N_13062);
and U17117 (N_17117,N_14937,N_11524);
xor U17118 (N_17118,N_14191,N_13863);
xor U17119 (N_17119,N_11579,N_11260);
and U17120 (N_17120,N_11336,N_13731);
or U17121 (N_17121,N_12056,N_10780);
or U17122 (N_17122,N_13458,N_11561);
or U17123 (N_17123,N_14616,N_11209);
nor U17124 (N_17124,N_12515,N_12346);
xor U17125 (N_17125,N_13555,N_12347);
nor U17126 (N_17126,N_10062,N_14422);
xnor U17127 (N_17127,N_12519,N_10069);
xor U17128 (N_17128,N_10086,N_11848);
nand U17129 (N_17129,N_14908,N_10527);
or U17130 (N_17130,N_10428,N_14479);
and U17131 (N_17131,N_11947,N_10677);
xor U17132 (N_17132,N_11264,N_14101);
xnor U17133 (N_17133,N_10157,N_13747);
nor U17134 (N_17134,N_13146,N_12380);
nand U17135 (N_17135,N_14030,N_11798);
nor U17136 (N_17136,N_10596,N_11668);
nor U17137 (N_17137,N_13321,N_11150);
nand U17138 (N_17138,N_12344,N_10708);
or U17139 (N_17139,N_11969,N_14545);
nand U17140 (N_17140,N_12349,N_10653);
xor U17141 (N_17141,N_13190,N_14481);
and U17142 (N_17142,N_10610,N_13688);
or U17143 (N_17143,N_11790,N_11295);
and U17144 (N_17144,N_14208,N_14860);
xnor U17145 (N_17145,N_11012,N_14062);
nand U17146 (N_17146,N_13562,N_11590);
nand U17147 (N_17147,N_14217,N_13257);
nand U17148 (N_17148,N_11146,N_12943);
xor U17149 (N_17149,N_12510,N_10967);
xor U17150 (N_17150,N_12662,N_11181);
and U17151 (N_17151,N_13070,N_13132);
nor U17152 (N_17152,N_12191,N_13693);
xnor U17153 (N_17153,N_12096,N_12128);
nand U17154 (N_17154,N_10478,N_10132);
nor U17155 (N_17155,N_10547,N_13518);
or U17156 (N_17156,N_14872,N_13466);
nand U17157 (N_17157,N_13400,N_14571);
xor U17158 (N_17158,N_14449,N_13784);
or U17159 (N_17159,N_10134,N_10504);
xnor U17160 (N_17160,N_14193,N_10851);
nor U17161 (N_17161,N_10329,N_14984);
and U17162 (N_17162,N_14394,N_13253);
and U17163 (N_17163,N_14953,N_13841);
and U17164 (N_17164,N_11173,N_13071);
nand U17165 (N_17165,N_13812,N_12489);
and U17166 (N_17166,N_11568,N_12607);
xnor U17167 (N_17167,N_10064,N_10071);
nand U17168 (N_17168,N_14997,N_14811);
nor U17169 (N_17169,N_13899,N_14033);
xor U17170 (N_17170,N_13014,N_13594);
and U17171 (N_17171,N_10936,N_11119);
nor U17172 (N_17172,N_13317,N_12665);
nor U17173 (N_17173,N_14710,N_13133);
and U17174 (N_17174,N_13372,N_14080);
or U17175 (N_17175,N_10444,N_11709);
and U17176 (N_17176,N_12771,N_13355);
nand U17177 (N_17177,N_14825,N_10467);
nand U17178 (N_17178,N_11736,N_14430);
xor U17179 (N_17179,N_14809,N_12898);
nor U17180 (N_17180,N_13529,N_14106);
xnor U17181 (N_17181,N_11006,N_10197);
xor U17182 (N_17182,N_13978,N_14254);
and U17183 (N_17183,N_12816,N_13711);
or U17184 (N_17184,N_10201,N_10546);
xnor U17185 (N_17185,N_14895,N_14709);
or U17186 (N_17186,N_13911,N_12342);
or U17187 (N_17187,N_12912,N_12603);
and U17188 (N_17188,N_10433,N_14465);
and U17189 (N_17189,N_13482,N_11694);
nor U17190 (N_17190,N_14529,N_14603);
or U17191 (N_17191,N_14875,N_11601);
xor U17192 (N_17192,N_12877,N_13218);
or U17193 (N_17193,N_10105,N_14752);
nand U17194 (N_17194,N_10470,N_14215);
and U17195 (N_17195,N_10061,N_10631);
and U17196 (N_17196,N_12865,N_10783);
nor U17197 (N_17197,N_14151,N_11098);
nor U17198 (N_17198,N_13501,N_14608);
and U17199 (N_17199,N_13677,N_10709);
or U17200 (N_17200,N_12335,N_10392);
or U17201 (N_17201,N_12613,N_12445);
or U17202 (N_17202,N_10155,N_14204);
xor U17203 (N_17203,N_13508,N_14296);
or U17204 (N_17204,N_13376,N_11639);
nand U17205 (N_17205,N_13605,N_10376);
nand U17206 (N_17206,N_14376,N_10127);
nor U17207 (N_17207,N_13334,N_11573);
nor U17208 (N_17208,N_14645,N_13985);
and U17209 (N_17209,N_10019,N_12408);
nor U17210 (N_17210,N_12594,N_10452);
nor U17211 (N_17211,N_11783,N_12331);
and U17212 (N_17212,N_14295,N_14107);
xnor U17213 (N_17213,N_14941,N_11819);
nor U17214 (N_17214,N_10768,N_13694);
and U17215 (N_17215,N_11689,N_14078);
and U17216 (N_17216,N_11124,N_13736);
and U17217 (N_17217,N_10821,N_10787);
xnor U17218 (N_17218,N_10761,N_12517);
xor U17219 (N_17219,N_14581,N_11252);
xor U17220 (N_17220,N_11854,N_10404);
xor U17221 (N_17221,N_13948,N_13973);
nand U17222 (N_17222,N_14735,N_12754);
nor U17223 (N_17223,N_14110,N_14169);
nand U17224 (N_17224,N_14326,N_13067);
nand U17225 (N_17225,N_12616,N_14359);
xnor U17226 (N_17226,N_11043,N_11581);
nor U17227 (N_17227,N_12264,N_12664);
or U17228 (N_17228,N_13486,N_12911);
and U17229 (N_17229,N_12770,N_10621);
nor U17230 (N_17230,N_11632,N_13395);
or U17231 (N_17231,N_10976,N_12762);
and U17232 (N_17232,N_12741,N_10089);
nand U17233 (N_17233,N_12653,N_11657);
nor U17234 (N_17234,N_13984,N_11953);
nor U17235 (N_17235,N_14262,N_11891);
and U17236 (N_17236,N_14079,N_12143);
xnor U17237 (N_17237,N_13075,N_14373);
xnor U17238 (N_17238,N_14011,N_10182);
nand U17239 (N_17239,N_14211,N_11330);
nor U17240 (N_17240,N_12428,N_14370);
or U17241 (N_17241,N_11894,N_10310);
and U17242 (N_17242,N_12670,N_13734);
xnor U17243 (N_17243,N_11127,N_14715);
xor U17244 (N_17244,N_12398,N_12976);
or U17245 (N_17245,N_14383,N_12656);
nor U17246 (N_17246,N_12348,N_11421);
nor U17247 (N_17247,N_13260,N_14091);
xor U17248 (N_17248,N_11231,N_14749);
nor U17249 (N_17249,N_14366,N_14940);
and U17250 (N_17250,N_11650,N_13078);
nor U17251 (N_17251,N_10296,N_12781);
nor U17252 (N_17252,N_12701,N_12400);
xor U17253 (N_17253,N_13534,N_13979);
or U17254 (N_17254,N_10905,N_14549);
or U17255 (N_17255,N_11873,N_10039);
nor U17256 (N_17256,N_10567,N_11510);
or U17257 (N_17257,N_10854,N_11158);
or U17258 (N_17258,N_14857,N_14124);
or U17259 (N_17259,N_14013,N_12900);
or U17260 (N_17260,N_12814,N_13789);
nor U17261 (N_17261,N_10084,N_12266);
and U17262 (N_17262,N_13467,N_10940);
nor U17263 (N_17263,N_13903,N_14625);
or U17264 (N_17264,N_10210,N_11397);
nor U17265 (N_17265,N_13955,N_10282);
or U17266 (N_17266,N_13388,N_13967);
xor U17267 (N_17267,N_12637,N_12586);
or U17268 (N_17268,N_12729,N_10698);
and U17269 (N_17269,N_14301,N_11045);
or U17270 (N_17270,N_13419,N_14670);
nand U17271 (N_17271,N_10888,N_14431);
or U17272 (N_17272,N_10388,N_11728);
nand U17273 (N_17273,N_11673,N_14926);
and U17274 (N_17274,N_11286,N_10993);
nor U17275 (N_17275,N_14385,N_14413);
or U17276 (N_17276,N_13554,N_11178);
and U17277 (N_17277,N_10514,N_13597);
xor U17278 (N_17278,N_11501,N_11934);
nor U17279 (N_17279,N_10145,N_14139);
xnor U17280 (N_17280,N_14779,N_11584);
nor U17281 (N_17281,N_13274,N_11541);
nor U17282 (N_17282,N_14052,N_11731);
xor U17283 (N_17283,N_14528,N_10984);
xor U17284 (N_17284,N_14828,N_14841);
nand U17285 (N_17285,N_12654,N_11447);
or U17286 (N_17286,N_10586,N_11509);
or U17287 (N_17287,N_10700,N_14999);
nand U17288 (N_17288,N_14232,N_12858);
and U17289 (N_17289,N_10891,N_10692);
and U17290 (N_17290,N_14699,N_12144);
xnor U17291 (N_17291,N_11052,N_14042);
or U17292 (N_17292,N_10770,N_13042);
nand U17293 (N_17293,N_10035,N_14588);
xnor U17294 (N_17294,N_11572,N_11007);
xnor U17295 (N_17295,N_10389,N_13511);
and U17296 (N_17296,N_13840,N_12140);
xor U17297 (N_17297,N_12903,N_11927);
nor U17298 (N_17298,N_11678,N_11063);
nor U17299 (N_17299,N_11042,N_10900);
and U17300 (N_17300,N_13326,N_11616);
nor U17301 (N_17301,N_12737,N_10862);
and U17302 (N_17302,N_12246,N_12385);
xor U17303 (N_17303,N_11705,N_13124);
and U17304 (N_17304,N_11988,N_13213);
or U17305 (N_17305,N_12984,N_11134);
nor U17306 (N_17306,N_11254,N_12923);
and U17307 (N_17307,N_10885,N_11112);
or U17308 (N_17308,N_11418,N_11320);
nor U17309 (N_17309,N_12777,N_10383);
and U17310 (N_17310,N_13090,N_12007);
nand U17311 (N_17311,N_12627,N_14523);
xor U17312 (N_17312,N_13914,N_10495);
nor U17313 (N_17313,N_14893,N_14622);
and U17314 (N_17314,N_10083,N_13548);
nor U17315 (N_17315,N_14039,N_14310);
or U17316 (N_17316,N_13120,N_14305);
nor U17317 (N_17317,N_13753,N_11469);
nand U17318 (N_17318,N_10634,N_10799);
nor U17319 (N_17319,N_14095,N_14061);
or U17320 (N_17320,N_11156,N_14463);
or U17321 (N_17321,N_13349,N_13687);
and U17322 (N_17322,N_11087,N_10757);
and U17323 (N_17323,N_11643,N_11939);
nand U17324 (N_17324,N_10252,N_14910);
or U17325 (N_17325,N_13187,N_12790);
xnor U17326 (N_17326,N_12452,N_11555);
nand U17327 (N_17327,N_11170,N_13800);
nor U17328 (N_17328,N_10379,N_13054);
nand U17329 (N_17329,N_12556,N_12980);
nand U17330 (N_17330,N_13697,N_11497);
nand U17331 (N_17331,N_13733,N_11453);
nor U17332 (N_17332,N_12073,N_11772);
or U17333 (N_17333,N_11693,N_14563);
or U17334 (N_17334,N_10482,N_10732);
nand U17335 (N_17335,N_12590,N_14199);
and U17336 (N_17336,N_11919,N_10337);
nor U17337 (N_17337,N_14424,N_10752);
or U17338 (N_17338,N_11767,N_13295);
or U17339 (N_17339,N_12040,N_11097);
xnor U17340 (N_17340,N_10706,N_11117);
and U17341 (N_17341,N_12946,N_10190);
nor U17342 (N_17342,N_14055,N_14219);
xor U17343 (N_17343,N_13946,N_11424);
nand U17344 (N_17344,N_12808,N_11378);
nand U17345 (N_17345,N_11475,N_12505);
nand U17346 (N_17346,N_14964,N_14916);
and U17347 (N_17347,N_10150,N_14762);
and U17348 (N_17348,N_11133,N_14830);
or U17349 (N_17349,N_11717,N_11597);
or U17350 (N_17350,N_11251,N_11704);
nor U17351 (N_17351,N_12234,N_10570);
or U17352 (N_17352,N_14221,N_13247);
or U17353 (N_17353,N_12957,N_14081);
nor U17354 (N_17354,N_11716,N_10494);
and U17355 (N_17355,N_10458,N_12136);
nand U17356 (N_17356,N_12573,N_11985);
xor U17357 (N_17357,N_11598,N_11785);
and U17358 (N_17358,N_14748,N_13826);
or U17359 (N_17359,N_12621,N_10794);
or U17360 (N_17360,N_13686,N_11887);
xnor U17361 (N_17361,N_14317,N_12111);
or U17362 (N_17362,N_14045,N_10842);
nor U17363 (N_17363,N_10156,N_13937);
and U17364 (N_17364,N_12260,N_11925);
nor U17365 (N_17365,N_12646,N_10056);
or U17366 (N_17366,N_12036,N_14929);
nor U17367 (N_17367,N_10651,N_11832);
or U17368 (N_17368,N_14278,N_12680);
and U17369 (N_17369,N_13855,N_10193);
xor U17370 (N_17370,N_10835,N_13191);
nand U17371 (N_17371,N_11332,N_14684);
nand U17372 (N_17372,N_12856,N_11549);
nand U17373 (N_17373,N_11053,N_11325);
nor U17374 (N_17374,N_10006,N_11984);
nor U17375 (N_17375,N_10255,N_11413);
xor U17376 (N_17376,N_12002,N_12330);
nand U17377 (N_17377,N_12630,N_10793);
and U17378 (N_17378,N_12369,N_14455);
and U17379 (N_17379,N_13276,N_14766);
xor U17380 (N_17380,N_11628,N_13629);
nand U17381 (N_17381,N_10573,N_14792);
nor U17382 (N_17382,N_10655,N_14344);
nor U17383 (N_17383,N_13639,N_11149);
nand U17384 (N_17384,N_14734,N_12894);
nor U17385 (N_17385,N_12843,N_12187);
and U17386 (N_17386,N_10207,N_12577);
nor U17387 (N_17387,N_12029,N_14157);
nor U17388 (N_17388,N_11419,N_12213);
nand U17389 (N_17389,N_11137,N_11893);
and U17390 (N_17390,N_13888,N_14503);
nand U17391 (N_17391,N_12792,N_13740);
and U17392 (N_17392,N_12108,N_13719);
nor U17393 (N_17393,N_14386,N_13798);
nand U17394 (N_17394,N_14742,N_12267);
or U17395 (N_17395,N_11576,N_13307);
xnor U17396 (N_17396,N_14186,N_14785);
and U17397 (N_17397,N_10099,N_11279);
xnor U17398 (N_17398,N_14864,N_12107);
xor U17399 (N_17399,N_11857,N_13339);
xor U17400 (N_17400,N_14005,N_10431);
and U17401 (N_17401,N_10493,N_12819);
or U17402 (N_17402,N_14981,N_10593);
xor U17403 (N_17403,N_12387,N_10669);
nand U17404 (N_17404,N_14685,N_12635);
xor U17405 (N_17405,N_11351,N_11402);
or U17406 (N_17406,N_14633,N_10394);
nor U17407 (N_17407,N_14513,N_10371);
xnor U17408 (N_17408,N_10234,N_14306);
and U17409 (N_17409,N_13296,N_14209);
nor U17410 (N_17410,N_14029,N_12465);
and U17411 (N_17411,N_11721,N_10317);
nand U17412 (N_17412,N_13118,N_13936);
or U17413 (N_17413,N_14565,N_14745);
nor U17414 (N_17414,N_12888,N_14814);
nand U17415 (N_17415,N_11422,N_14473);
or U17416 (N_17416,N_13988,N_12778);
and U17417 (N_17417,N_10184,N_14273);
nor U17418 (N_17418,N_14450,N_12009);
and U17419 (N_17419,N_13072,N_13053);
nor U17420 (N_17420,N_11180,N_10114);
and U17421 (N_17421,N_10776,N_11631);
or U17422 (N_17422,N_12528,N_11574);
nor U17423 (N_17423,N_13965,N_11636);
nor U17424 (N_17424,N_13414,N_13416);
nor U17425 (N_17425,N_12069,N_14288);
or U17426 (N_17426,N_12749,N_12258);
xor U17427 (N_17427,N_13036,N_13692);
nor U17428 (N_17428,N_11872,N_13982);
xnor U17429 (N_17429,N_12623,N_13708);
xor U17430 (N_17430,N_12509,N_10358);
nor U17431 (N_17431,N_11329,N_10471);
or U17432 (N_17432,N_14322,N_13096);
nand U17433 (N_17433,N_13838,N_11799);
nand U17434 (N_17434,N_12268,N_10192);
and U17435 (N_17435,N_14892,N_10289);
xor U17436 (N_17436,N_12844,N_11417);
or U17437 (N_17437,N_13625,N_11338);
and U17438 (N_17438,N_10874,N_12072);
and U17439 (N_17439,N_10049,N_14947);
nor U17440 (N_17440,N_10353,N_13493);
and U17441 (N_17441,N_10027,N_12883);
nor U17442 (N_17442,N_12170,N_10492);
xor U17443 (N_17443,N_13608,N_14183);
nor U17444 (N_17444,N_13791,N_11760);
nor U17445 (N_17445,N_12063,N_12720);
or U17446 (N_17446,N_14362,N_11428);
nand U17447 (N_17447,N_14543,N_12995);
nor U17448 (N_17448,N_14815,N_10005);
nand U17449 (N_17449,N_10113,N_12581);
nand U17450 (N_17450,N_10119,N_13614);
or U17451 (N_17451,N_13343,N_11381);
nor U17452 (N_17452,N_12780,N_14324);
nor U17453 (N_17453,N_12503,N_11125);
nor U17454 (N_17454,N_11474,N_11874);
nand U17455 (N_17455,N_11068,N_13209);
nand U17456 (N_17456,N_11741,N_10765);
or U17457 (N_17457,N_13406,N_10986);
xor U17458 (N_17458,N_10457,N_11583);
nand U17459 (N_17459,N_10829,N_12257);
nand U17460 (N_17460,N_10332,N_12969);
and U17461 (N_17461,N_13086,N_11747);
nand U17462 (N_17462,N_13666,N_11412);
nand U17463 (N_17463,N_12383,N_11801);
nor U17464 (N_17464,N_13284,N_12117);
nor U17465 (N_17465,N_13521,N_13808);
nand U17466 (N_17466,N_10137,N_11645);
nor U17467 (N_17467,N_11905,N_10521);
xnor U17468 (N_17468,N_11316,N_11779);
nor U17469 (N_17469,N_12291,N_13160);
xnor U17470 (N_17470,N_12157,N_13558);
nand U17471 (N_17471,N_11074,N_12679);
nand U17472 (N_17472,N_13665,N_12337);
nand U17473 (N_17473,N_13896,N_10922);
nor U17474 (N_17474,N_11359,N_11224);
xnor U17475 (N_17475,N_11420,N_13011);
or U17476 (N_17476,N_12273,N_10741);
nor U17477 (N_17477,N_11307,N_12177);
and U17478 (N_17478,N_13643,N_13610);
or U17479 (N_17479,N_10290,N_10552);
xor U17480 (N_17480,N_14642,N_13116);
or U17481 (N_17481,N_14922,N_11266);
or U17482 (N_17482,N_12048,N_14954);
or U17483 (N_17483,N_12031,N_10254);
or U17484 (N_17484,N_14621,N_13929);
and U17485 (N_17485,N_14923,N_12588);
and U17486 (N_17486,N_10268,N_11100);
xor U17487 (N_17487,N_10998,N_12093);
nor U17488 (N_17488,N_11435,N_13216);
nor U17489 (N_17489,N_11771,N_14626);
and U17490 (N_17490,N_10445,N_14720);
nor U17491 (N_17491,N_14599,N_13371);
or U17492 (N_17492,N_14488,N_10730);
xnor U17493 (N_17493,N_14530,N_10483);
and U17494 (N_17494,N_10030,N_13578);
xnor U17495 (N_17495,N_12756,N_14589);
and U17496 (N_17496,N_13041,N_12432);
xor U17497 (N_17497,N_14804,N_12173);
nand U17498 (N_17498,N_14355,N_14595);
or U17499 (N_17499,N_13156,N_14991);
nor U17500 (N_17500,N_12334,N_14278);
nand U17501 (N_17501,N_11271,N_11911);
nand U17502 (N_17502,N_10294,N_14025);
nor U17503 (N_17503,N_13992,N_10316);
xnor U17504 (N_17504,N_13052,N_12262);
nand U17505 (N_17505,N_11312,N_12086);
xnor U17506 (N_17506,N_14610,N_14267);
nand U17507 (N_17507,N_14813,N_12842);
or U17508 (N_17508,N_13046,N_13845);
nand U17509 (N_17509,N_11679,N_13532);
xnor U17510 (N_17510,N_13377,N_10225);
and U17511 (N_17511,N_10763,N_12241);
xnor U17512 (N_17512,N_12074,N_10740);
xor U17513 (N_17513,N_11786,N_13057);
xor U17514 (N_17514,N_10399,N_12417);
or U17515 (N_17515,N_12151,N_12822);
and U17516 (N_17516,N_12038,N_12878);
xor U17517 (N_17517,N_10724,N_11368);
nor U17518 (N_17518,N_13554,N_14711);
nor U17519 (N_17519,N_10807,N_13438);
xor U17520 (N_17520,N_14759,N_13816);
nand U17521 (N_17521,N_14100,N_14022);
nand U17522 (N_17522,N_11697,N_10716);
nor U17523 (N_17523,N_11916,N_12870);
nand U17524 (N_17524,N_12975,N_10355);
xnor U17525 (N_17525,N_11453,N_12265);
xnor U17526 (N_17526,N_13471,N_11734);
xor U17527 (N_17527,N_14985,N_11418);
or U17528 (N_17528,N_13890,N_14704);
or U17529 (N_17529,N_14694,N_14610);
xnor U17530 (N_17530,N_13994,N_11707);
or U17531 (N_17531,N_10812,N_10966);
nor U17532 (N_17532,N_13120,N_14622);
nor U17533 (N_17533,N_11220,N_10950);
and U17534 (N_17534,N_11785,N_10113);
xor U17535 (N_17535,N_10024,N_13737);
xnor U17536 (N_17536,N_13049,N_10530);
or U17537 (N_17537,N_14288,N_13835);
nand U17538 (N_17538,N_11851,N_13633);
nor U17539 (N_17539,N_14071,N_13256);
nand U17540 (N_17540,N_11863,N_14011);
or U17541 (N_17541,N_10123,N_13946);
nand U17542 (N_17542,N_13170,N_14135);
nor U17543 (N_17543,N_11022,N_12579);
xnor U17544 (N_17544,N_10208,N_13763);
and U17545 (N_17545,N_11700,N_11932);
or U17546 (N_17546,N_13380,N_13034);
or U17547 (N_17547,N_14494,N_13991);
nand U17548 (N_17548,N_13753,N_12135);
xor U17549 (N_17549,N_10976,N_12911);
and U17550 (N_17550,N_12604,N_14103);
and U17551 (N_17551,N_12616,N_10573);
or U17552 (N_17552,N_14460,N_14373);
nand U17553 (N_17553,N_13786,N_14046);
or U17554 (N_17554,N_10422,N_10804);
nor U17555 (N_17555,N_10654,N_13180);
xnor U17556 (N_17556,N_10327,N_11661);
or U17557 (N_17557,N_11597,N_10271);
nor U17558 (N_17558,N_11723,N_14673);
nand U17559 (N_17559,N_12144,N_13430);
or U17560 (N_17560,N_10762,N_10385);
xnor U17561 (N_17561,N_11087,N_12288);
or U17562 (N_17562,N_11690,N_13632);
nand U17563 (N_17563,N_14820,N_14959);
or U17564 (N_17564,N_10315,N_13149);
and U17565 (N_17565,N_10452,N_10826);
and U17566 (N_17566,N_13769,N_11551);
and U17567 (N_17567,N_12628,N_12392);
xor U17568 (N_17568,N_13037,N_11473);
and U17569 (N_17569,N_13375,N_11157);
and U17570 (N_17570,N_14971,N_11523);
nand U17571 (N_17571,N_13004,N_12126);
or U17572 (N_17572,N_13605,N_11977);
nand U17573 (N_17573,N_10391,N_11608);
xor U17574 (N_17574,N_12659,N_14015);
nor U17575 (N_17575,N_11482,N_14161);
or U17576 (N_17576,N_13224,N_13160);
xor U17577 (N_17577,N_10898,N_12861);
nor U17578 (N_17578,N_12846,N_12747);
nor U17579 (N_17579,N_13993,N_10431);
xor U17580 (N_17580,N_12210,N_12931);
nand U17581 (N_17581,N_12277,N_11239);
and U17582 (N_17582,N_12890,N_12939);
or U17583 (N_17583,N_10553,N_10857);
or U17584 (N_17584,N_12065,N_14550);
nand U17585 (N_17585,N_14590,N_11324);
xor U17586 (N_17586,N_14478,N_13715);
nor U17587 (N_17587,N_11831,N_13972);
nor U17588 (N_17588,N_12827,N_12214);
nand U17589 (N_17589,N_13451,N_14888);
nor U17590 (N_17590,N_11168,N_12794);
and U17591 (N_17591,N_10221,N_13452);
nand U17592 (N_17592,N_11065,N_11630);
nand U17593 (N_17593,N_12921,N_10163);
nand U17594 (N_17594,N_10784,N_14090);
xnor U17595 (N_17595,N_10503,N_10170);
nor U17596 (N_17596,N_11980,N_12796);
nand U17597 (N_17597,N_10720,N_12218);
and U17598 (N_17598,N_11205,N_13621);
nand U17599 (N_17599,N_14291,N_10794);
nand U17600 (N_17600,N_14430,N_13320);
xor U17601 (N_17601,N_10106,N_10181);
xor U17602 (N_17602,N_11711,N_11236);
nand U17603 (N_17603,N_10714,N_13884);
and U17604 (N_17604,N_12319,N_10032);
nand U17605 (N_17605,N_13497,N_12261);
nand U17606 (N_17606,N_13235,N_14494);
xor U17607 (N_17607,N_11784,N_14321);
or U17608 (N_17608,N_14412,N_11611);
and U17609 (N_17609,N_12869,N_12279);
nor U17610 (N_17610,N_11985,N_13685);
or U17611 (N_17611,N_14760,N_11326);
nand U17612 (N_17612,N_13177,N_14145);
or U17613 (N_17613,N_12902,N_13553);
or U17614 (N_17614,N_10572,N_10043);
and U17615 (N_17615,N_11981,N_14889);
and U17616 (N_17616,N_13774,N_11161);
and U17617 (N_17617,N_12344,N_14528);
and U17618 (N_17618,N_10960,N_12353);
nand U17619 (N_17619,N_11736,N_10314);
nor U17620 (N_17620,N_11482,N_11158);
nand U17621 (N_17621,N_11620,N_14907);
and U17622 (N_17622,N_14427,N_12353);
xor U17623 (N_17623,N_12208,N_14432);
or U17624 (N_17624,N_11883,N_13142);
xor U17625 (N_17625,N_13661,N_11209);
nor U17626 (N_17626,N_14585,N_13883);
nor U17627 (N_17627,N_13702,N_11379);
xor U17628 (N_17628,N_14812,N_10846);
or U17629 (N_17629,N_14039,N_10859);
nor U17630 (N_17630,N_11575,N_13664);
nand U17631 (N_17631,N_10450,N_14044);
xor U17632 (N_17632,N_14805,N_13582);
xor U17633 (N_17633,N_11334,N_11385);
or U17634 (N_17634,N_13913,N_11135);
or U17635 (N_17635,N_10162,N_12856);
and U17636 (N_17636,N_10206,N_12567);
xor U17637 (N_17637,N_11637,N_11949);
nand U17638 (N_17638,N_13296,N_13784);
nor U17639 (N_17639,N_14765,N_12650);
and U17640 (N_17640,N_12505,N_12838);
and U17641 (N_17641,N_12415,N_10163);
xnor U17642 (N_17642,N_11469,N_12903);
nand U17643 (N_17643,N_13422,N_13025);
nor U17644 (N_17644,N_14536,N_14839);
and U17645 (N_17645,N_10226,N_14576);
or U17646 (N_17646,N_14035,N_12185);
xnor U17647 (N_17647,N_10164,N_12608);
nand U17648 (N_17648,N_12671,N_13237);
nand U17649 (N_17649,N_10811,N_13375);
xor U17650 (N_17650,N_13524,N_10082);
nor U17651 (N_17651,N_14138,N_11834);
xnor U17652 (N_17652,N_14558,N_14524);
and U17653 (N_17653,N_11897,N_12463);
or U17654 (N_17654,N_10483,N_14164);
and U17655 (N_17655,N_14049,N_10473);
nor U17656 (N_17656,N_11491,N_11231);
nand U17657 (N_17657,N_10324,N_13368);
nand U17658 (N_17658,N_10967,N_11293);
nand U17659 (N_17659,N_13423,N_13941);
xnor U17660 (N_17660,N_14914,N_14401);
and U17661 (N_17661,N_12299,N_14747);
or U17662 (N_17662,N_11928,N_10508);
xor U17663 (N_17663,N_12404,N_12005);
and U17664 (N_17664,N_10791,N_12714);
or U17665 (N_17665,N_11789,N_12975);
xnor U17666 (N_17666,N_12780,N_10244);
or U17667 (N_17667,N_10732,N_10178);
nor U17668 (N_17668,N_13944,N_11312);
or U17669 (N_17669,N_10589,N_11328);
nor U17670 (N_17670,N_13131,N_12288);
or U17671 (N_17671,N_14897,N_14532);
xnor U17672 (N_17672,N_13819,N_13465);
xor U17673 (N_17673,N_11051,N_13506);
xor U17674 (N_17674,N_10762,N_13947);
or U17675 (N_17675,N_14888,N_10482);
and U17676 (N_17676,N_14506,N_12153);
and U17677 (N_17677,N_11502,N_12425);
or U17678 (N_17678,N_10581,N_10636);
or U17679 (N_17679,N_10718,N_12829);
nand U17680 (N_17680,N_14326,N_12002);
nor U17681 (N_17681,N_13866,N_14305);
or U17682 (N_17682,N_14696,N_13395);
or U17683 (N_17683,N_10779,N_10922);
and U17684 (N_17684,N_13692,N_14307);
nor U17685 (N_17685,N_13771,N_12166);
or U17686 (N_17686,N_13882,N_14388);
xor U17687 (N_17687,N_10076,N_10385);
xnor U17688 (N_17688,N_13543,N_14207);
or U17689 (N_17689,N_12261,N_11013);
nor U17690 (N_17690,N_11113,N_12183);
and U17691 (N_17691,N_12082,N_13406);
nand U17692 (N_17692,N_13947,N_11764);
nor U17693 (N_17693,N_11634,N_12251);
nand U17694 (N_17694,N_13573,N_11276);
nand U17695 (N_17695,N_13327,N_12744);
nor U17696 (N_17696,N_13449,N_13799);
or U17697 (N_17697,N_10473,N_10615);
xnor U17698 (N_17698,N_14961,N_13173);
nor U17699 (N_17699,N_11590,N_12468);
xor U17700 (N_17700,N_14173,N_12165);
or U17701 (N_17701,N_12245,N_14140);
xor U17702 (N_17702,N_11873,N_14905);
or U17703 (N_17703,N_10892,N_12742);
xor U17704 (N_17704,N_10884,N_11225);
and U17705 (N_17705,N_11937,N_11488);
and U17706 (N_17706,N_10075,N_12380);
or U17707 (N_17707,N_12527,N_11599);
nor U17708 (N_17708,N_14321,N_14698);
or U17709 (N_17709,N_12819,N_14770);
xor U17710 (N_17710,N_11204,N_11874);
xnor U17711 (N_17711,N_12531,N_10791);
or U17712 (N_17712,N_10935,N_13908);
and U17713 (N_17713,N_10798,N_14205);
nand U17714 (N_17714,N_14480,N_12620);
xnor U17715 (N_17715,N_11426,N_12709);
and U17716 (N_17716,N_14437,N_11375);
or U17717 (N_17717,N_10275,N_12748);
xor U17718 (N_17718,N_14147,N_14072);
xor U17719 (N_17719,N_10081,N_13600);
nand U17720 (N_17720,N_13232,N_14621);
xnor U17721 (N_17721,N_14532,N_12283);
and U17722 (N_17722,N_12091,N_11219);
xnor U17723 (N_17723,N_14918,N_11564);
and U17724 (N_17724,N_10863,N_12659);
nand U17725 (N_17725,N_14609,N_10007);
and U17726 (N_17726,N_14057,N_10379);
and U17727 (N_17727,N_10205,N_13227);
nor U17728 (N_17728,N_10428,N_12415);
xor U17729 (N_17729,N_11028,N_14002);
nor U17730 (N_17730,N_14267,N_13628);
nor U17731 (N_17731,N_12575,N_13419);
xor U17732 (N_17732,N_14825,N_13994);
or U17733 (N_17733,N_13555,N_12881);
and U17734 (N_17734,N_12559,N_10632);
nand U17735 (N_17735,N_12807,N_11689);
xor U17736 (N_17736,N_12773,N_11919);
nor U17737 (N_17737,N_14544,N_13205);
or U17738 (N_17738,N_13929,N_12717);
or U17739 (N_17739,N_14537,N_13229);
and U17740 (N_17740,N_10888,N_14652);
nor U17741 (N_17741,N_11784,N_13698);
or U17742 (N_17742,N_12813,N_14431);
nand U17743 (N_17743,N_12171,N_14318);
nor U17744 (N_17744,N_14345,N_14654);
and U17745 (N_17745,N_14547,N_12999);
xor U17746 (N_17746,N_11193,N_14992);
nand U17747 (N_17747,N_12892,N_14006);
or U17748 (N_17748,N_13590,N_11007);
or U17749 (N_17749,N_14653,N_14333);
and U17750 (N_17750,N_10598,N_11596);
nand U17751 (N_17751,N_10691,N_11060);
xor U17752 (N_17752,N_10569,N_13941);
xnor U17753 (N_17753,N_12559,N_10818);
xnor U17754 (N_17754,N_11317,N_13596);
nor U17755 (N_17755,N_12686,N_10047);
and U17756 (N_17756,N_10407,N_12250);
xor U17757 (N_17757,N_12127,N_11836);
nand U17758 (N_17758,N_10916,N_10454);
or U17759 (N_17759,N_13891,N_13342);
nand U17760 (N_17760,N_10356,N_13771);
and U17761 (N_17761,N_14974,N_11850);
nor U17762 (N_17762,N_10235,N_13134);
xnor U17763 (N_17763,N_14284,N_14609);
xnor U17764 (N_17764,N_14041,N_11215);
nor U17765 (N_17765,N_14818,N_13492);
xnor U17766 (N_17766,N_12746,N_11686);
or U17767 (N_17767,N_10805,N_11903);
nand U17768 (N_17768,N_12924,N_10755);
or U17769 (N_17769,N_14084,N_10037);
nor U17770 (N_17770,N_14717,N_14101);
and U17771 (N_17771,N_11274,N_10103);
xor U17772 (N_17772,N_11881,N_11310);
or U17773 (N_17773,N_12339,N_13471);
nand U17774 (N_17774,N_14630,N_10883);
nor U17775 (N_17775,N_13356,N_11750);
and U17776 (N_17776,N_12315,N_14111);
xor U17777 (N_17777,N_13500,N_12831);
nand U17778 (N_17778,N_10776,N_10282);
nor U17779 (N_17779,N_12595,N_13506);
nand U17780 (N_17780,N_12737,N_14705);
or U17781 (N_17781,N_13987,N_13719);
or U17782 (N_17782,N_10539,N_12972);
nand U17783 (N_17783,N_11442,N_11360);
xnor U17784 (N_17784,N_12499,N_12902);
or U17785 (N_17785,N_12707,N_11272);
xnor U17786 (N_17786,N_14308,N_11891);
nor U17787 (N_17787,N_11722,N_11298);
or U17788 (N_17788,N_13235,N_11896);
or U17789 (N_17789,N_10708,N_12776);
nand U17790 (N_17790,N_11261,N_10981);
or U17791 (N_17791,N_10937,N_14112);
or U17792 (N_17792,N_13931,N_12389);
nand U17793 (N_17793,N_11660,N_14577);
xor U17794 (N_17794,N_13382,N_14245);
nor U17795 (N_17795,N_11372,N_14250);
nor U17796 (N_17796,N_13911,N_10646);
and U17797 (N_17797,N_14306,N_12964);
nand U17798 (N_17798,N_14634,N_11895);
or U17799 (N_17799,N_10517,N_12727);
and U17800 (N_17800,N_14262,N_14028);
xor U17801 (N_17801,N_10470,N_13870);
and U17802 (N_17802,N_12572,N_13995);
and U17803 (N_17803,N_14437,N_13106);
and U17804 (N_17804,N_14529,N_13957);
or U17805 (N_17805,N_10603,N_11364);
and U17806 (N_17806,N_10386,N_12830);
xor U17807 (N_17807,N_10149,N_10838);
nand U17808 (N_17808,N_11090,N_11208);
nand U17809 (N_17809,N_14755,N_12880);
or U17810 (N_17810,N_11941,N_11352);
and U17811 (N_17811,N_10804,N_14345);
xnor U17812 (N_17812,N_12534,N_14104);
xnor U17813 (N_17813,N_12325,N_14009);
or U17814 (N_17814,N_12874,N_10038);
nand U17815 (N_17815,N_12523,N_13278);
xnor U17816 (N_17816,N_10379,N_14252);
and U17817 (N_17817,N_13688,N_10936);
or U17818 (N_17818,N_10938,N_13135);
and U17819 (N_17819,N_13477,N_13751);
or U17820 (N_17820,N_12180,N_10523);
xnor U17821 (N_17821,N_13161,N_12935);
or U17822 (N_17822,N_11724,N_13656);
nor U17823 (N_17823,N_13454,N_14010);
nand U17824 (N_17824,N_13416,N_11684);
nand U17825 (N_17825,N_11748,N_12578);
or U17826 (N_17826,N_13939,N_11026);
or U17827 (N_17827,N_14993,N_13938);
nor U17828 (N_17828,N_12765,N_11922);
nor U17829 (N_17829,N_12019,N_11306);
nor U17830 (N_17830,N_13471,N_14295);
nand U17831 (N_17831,N_10416,N_11241);
and U17832 (N_17832,N_11087,N_14271);
or U17833 (N_17833,N_11151,N_14742);
nand U17834 (N_17834,N_13996,N_10205);
and U17835 (N_17835,N_10187,N_11309);
xor U17836 (N_17836,N_14595,N_10974);
or U17837 (N_17837,N_13545,N_12030);
xor U17838 (N_17838,N_12396,N_11159);
nor U17839 (N_17839,N_10348,N_10316);
nand U17840 (N_17840,N_12894,N_10779);
nand U17841 (N_17841,N_10245,N_10797);
nor U17842 (N_17842,N_14738,N_11424);
nor U17843 (N_17843,N_11919,N_12421);
nand U17844 (N_17844,N_14112,N_10433);
and U17845 (N_17845,N_11802,N_12630);
and U17846 (N_17846,N_11462,N_13871);
and U17847 (N_17847,N_14327,N_10777);
or U17848 (N_17848,N_10123,N_12089);
and U17849 (N_17849,N_14248,N_11740);
xor U17850 (N_17850,N_11901,N_10303);
nor U17851 (N_17851,N_11551,N_11975);
xor U17852 (N_17852,N_10087,N_11511);
nor U17853 (N_17853,N_11751,N_12902);
nor U17854 (N_17854,N_13285,N_13936);
and U17855 (N_17855,N_14948,N_12074);
and U17856 (N_17856,N_10650,N_12798);
xor U17857 (N_17857,N_10483,N_13568);
xnor U17858 (N_17858,N_13108,N_12580);
nand U17859 (N_17859,N_12125,N_12283);
nor U17860 (N_17860,N_10564,N_12188);
or U17861 (N_17861,N_12149,N_13347);
or U17862 (N_17862,N_11785,N_14939);
nor U17863 (N_17863,N_13209,N_14958);
nor U17864 (N_17864,N_11076,N_12913);
xnor U17865 (N_17865,N_10869,N_14103);
xnor U17866 (N_17866,N_10350,N_13628);
nor U17867 (N_17867,N_10260,N_11564);
and U17868 (N_17868,N_14512,N_13055);
or U17869 (N_17869,N_13450,N_11635);
nor U17870 (N_17870,N_12552,N_10706);
nand U17871 (N_17871,N_12571,N_14292);
and U17872 (N_17872,N_12033,N_13242);
and U17873 (N_17873,N_13966,N_12685);
and U17874 (N_17874,N_13809,N_12287);
nor U17875 (N_17875,N_11017,N_13943);
nor U17876 (N_17876,N_14037,N_10969);
and U17877 (N_17877,N_12275,N_11223);
xnor U17878 (N_17878,N_13402,N_13688);
xnor U17879 (N_17879,N_12072,N_12724);
nor U17880 (N_17880,N_14511,N_14324);
and U17881 (N_17881,N_13867,N_11570);
xnor U17882 (N_17882,N_12999,N_12518);
nor U17883 (N_17883,N_13224,N_11042);
nand U17884 (N_17884,N_11401,N_14727);
or U17885 (N_17885,N_11184,N_12466);
or U17886 (N_17886,N_10748,N_11098);
and U17887 (N_17887,N_10028,N_12119);
nand U17888 (N_17888,N_14187,N_10287);
nand U17889 (N_17889,N_10193,N_11481);
xor U17890 (N_17890,N_12133,N_11734);
or U17891 (N_17891,N_12902,N_12528);
xnor U17892 (N_17892,N_12079,N_14009);
and U17893 (N_17893,N_13765,N_12287);
xor U17894 (N_17894,N_10760,N_11819);
or U17895 (N_17895,N_14210,N_13586);
nor U17896 (N_17896,N_13198,N_12514);
and U17897 (N_17897,N_13307,N_13902);
and U17898 (N_17898,N_14913,N_10049);
nor U17899 (N_17899,N_11663,N_12962);
or U17900 (N_17900,N_13787,N_12831);
nand U17901 (N_17901,N_14593,N_13614);
nor U17902 (N_17902,N_10850,N_11885);
nand U17903 (N_17903,N_13836,N_12842);
or U17904 (N_17904,N_12087,N_11907);
or U17905 (N_17905,N_10037,N_10637);
xor U17906 (N_17906,N_11069,N_11640);
xor U17907 (N_17907,N_11099,N_13892);
nor U17908 (N_17908,N_10663,N_13173);
nand U17909 (N_17909,N_12901,N_10585);
and U17910 (N_17910,N_13683,N_11550);
nor U17911 (N_17911,N_10603,N_10830);
nor U17912 (N_17912,N_10953,N_10591);
and U17913 (N_17913,N_10232,N_13307);
nand U17914 (N_17914,N_13346,N_12486);
nand U17915 (N_17915,N_13012,N_12050);
and U17916 (N_17916,N_12655,N_12707);
nand U17917 (N_17917,N_10449,N_11685);
and U17918 (N_17918,N_10054,N_11310);
and U17919 (N_17919,N_10658,N_14691);
and U17920 (N_17920,N_11714,N_11970);
nor U17921 (N_17921,N_11766,N_14615);
or U17922 (N_17922,N_12879,N_10563);
nor U17923 (N_17923,N_11167,N_13216);
xor U17924 (N_17924,N_14123,N_10056);
and U17925 (N_17925,N_10033,N_14448);
nand U17926 (N_17926,N_11570,N_11693);
and U17927 (N_17927,N_10408,N_10648);
xnor U17928 (N_17928,N_11567,N_10527);
or U17929 (N_17929,N_12664,N_13340);
nand U17930 (N_17930,N_12831,N_10250);
xnor U17931 (N_17931,N_11938,N_13252);
nand U17932 (N_17932,N_14425,N_13469);
nor U17933 (N_17933,N_13228,N_13808);
xnor U17934 (N_17934,N_11639,N_11534);
nand U17935 (N_17935,N_10923,N_13272);
xor U17936 (N_17936,N_10286,N_11549);
and U17937 (N_17937,N_12594,N_10403);
nand U17938 (N_17938,N_13640,N_14232);
or U17939 (N_17939,N_12383,N_12458);
nand U17940 (N_17940,N_13367,N_12557);
nand U17941 (N_17941,N_12217,N_10483);
or U17942 (N_17942,N_10939,N_13157);
or U17943 (N_17943,N_10234,N_14247);
or U17944 (N_17944,N_13787,N_12497);
xnor U17945 (N_17945,N_10090,N_11213);
or U17946 (N_17946,N_12967,N_14458);
xnor U17947 (N_17947,N_14539,N_10257);
nand U17948 (N_17948,N_14198,N_12512);
nand U17949 (N_17949,N_12124,N_14795);
or U17950 (N_17950,N_11796,N_11406);
nor U17951 (N_17951,N_13909,N_12097);
or U17952 (N_17952,N_14403,N_12869);
nor U17953 (N_17953,N_14727,N_11030);
nor U17954 (N_17954,N_10461,N_13306);
nand U17955 (N_17955,N_13184,N_13908);
or U17956 (N_17956,N_13386,N_12268);
and U17957 (N_17957,N_10801,N_12876);
and U17958 (N_17958,N_10959,N_10050);
nand U17959 (N_17959,N_13484,N_12378);
xnor U17960 (N_17960,N_14238,N_10095);
xnor U17961 (N_17961,N_10422,N_14308);
and U17962 (N_17962,N_12597,N_14757);
and U17963 (N_17963,N_10295,N_13292);
nor U17964 (N_17964,N_11449,N_13515);
or U17965 (N_17965,N_13900,N_14012);
nand U17966 (N_17966,N_11381,N_14246);
nor U17967 (N_17967,N_11390,N_13028);
and U17968 (N_17968,N_11154,N_12088);
or U17969 (N_17969,N_11886,N_12768);
and U17970 (N_17970,N_12752,N_14330);
and U17971 (N_17971,N_13435,N_14535);
nand U17972 (N_17972,N_10996,N_13595);
xor U17973 (N_17973,N_14182,N_14256);
nand U17974 (N_17974,N_10262,N_11110);
nor U17975 (N_17975,N_14302,N_13460);
nand U17976 (N_17976,N_11164,N_13473);
or U17977 (N_17977,N_12428,N_10803);
nand U17978 (N_17978,N_12569,N_12836);
and U17979 (N_17979,N_13672,N_14033);
nand U17980 (N_17980,N_10040,N_12083);
nand U17981 (N_17981,N_14107,N_13752);
or U17982 (N_17982,N_10776,N_14081);
nand U17983 (N_17983,N_14121,N_13542);
xor U17984 (N_17984,N_11465,N_13111);
nand U17985 (N_17985,N_14964,N_11944);
nor U17986 (N_17986,N_14548,N_10697);
and U17987 (N_17987,N_12264,N_10724);
nor U17988 (N_17988,N_11867,N_10544);
or U17989 (N_17989,N_14986,N_10339);
xor U17990 (N_17990,N_11762,N_10676);
and U17991 (N_17991,N_10905,N_13644);
and U17992 (N_17992,N_11320,N_14065);
xor U17993 (N_17993,N_10013,N_12583);
or U17994 (N_17994,N_11796,N_11849);
nand U17995 (N_17995,N_14926,N_14211);
nand U17996 (N_17996,N_11640,N_11501);
or U17997 (N_17997,N_14521,N_11206);
and U17998 (N_17998,N_11935,N_14342);
xor U17999 (N_17999,N_13888,N_12010);
xor U18000 (N_18000,N_10142,N_10175);
xor U18001 (N_18001,N_11055,N_12525);
xor U18002 (N_18002,N_10053,N_11121);
and U18003 (N_18003,N_10905,N_11587);
nand U18004 (N_18004,N_10727,N_12771);
nand U18005 (N_18005,N_12049,N_14846);
and U18006 (N_18006,N_14120,N_11031);
nand U18007 (N_18007,N_13366,N_11177);
xor U18008 (N_18008,N_14971,N_12343);
xor U18009 (N_18009,N_14865,N_14716);
xnor U18010 (N_18010,N_13721,N_12837);
or U18011 (N_18011,N_11200,N_12380);
nand U18012 (N_18012,N_12582,N_13231);
and U18013 (N_18013,N_14712,N_11110);
or U18014 (N_18014,N_11007,N_14866);
xor U18015 (N_18015,N_14439,N_11173);
nor U18016 (N_18016,N_11022,N_13283);
or U18017 (N_18017,N_13734,N_11627);
nand U18018 (N_18018,N_12926,N_11136);
xor U18019 (N_18019,N_10243,N_12283);
nor U18020 (N_18020,N_11785,N_10997);
or U18021 (N_18021,N_11007,N_13654);
nand U18022 (N_18022,N_12481,N_12170);
or U18023 (N_18023,N_13929,N_12594);
nand U18024 (N_18024,N_13442,N_12854);
or U18025 (N_18025,N_14364,N_12812);
nor U18026 (N_18026,N_14698,N_12824);
and U18027 (N_18027,N_10924,N_10424);
or U18028 (N_18028,N_12634,N_14882);
xnor U18029 (N_18029,N_13459,N_12043);
or U18030 (N_18030,N_11414,N_10874);
or U18031 (N_18031,N_11541,N_10077);
or U18032 (N_18032,N_11062,N_13885);
xnor U18033 (N_18033,N_11333,N_13358);
nor U18034 (N_18034,N_11051,N_13044);
nand U18035 (N_18035,N_12894,N_12754);
nand U18036 (N_18036,N_12707,N_10216);
or U18037 (N_18037,N_11479,N_13604);
or U18038 (N_18038,N_11926,N_11645);
nand U18039 (N_18039,N_10791,N_12738);
or U18040 (N_18040,N_10736,N_14492);
nor U18041 (N_18041,N_14490,N_13006);
or U18042 (N_18042,N_12330,N_13680);
and U18043 (N_18043,N_12792,N_14182);
nand U18044 (N_18044,N_11765,N_11426);
nor U18045 (N_18045,N_11675,N_14250);
nor U18046 (N_18046,N_10106,N_13492);
xor U18047 (N_18047,N_11651,N_10340);
nand U18048 (N_18048,N_10760,N_11537);
nor U18049 (N_18049,N_12410,N_11046);
or U18050 (N_18050,N_12302,N_13090);
nor U18051 (N_18051,N_13991,N_13424);
or U18052 (N_18052,N_13961,N_11268);
nor U18053 (N_18053,N_14382,N_14334);
xor U18054 (N_18054,N_11202,N_13054);
xnor U18055 (N_18055,N_13890,N_12292);
and U18056 (N_18056,N_12503,N_10018);
xnor U18057 (N_18057,N_14354,N_13051);
nor U18058 (N_18058,N_12863,N_11670);
nor U18059 (N_18059,N_11096,N_13474);
or U18060 (N_18060,N_10770,N_12291);
and U18061 (N_18061,N_10463,N_10107);
nand U18062 (N_18062,N_10938,N_13393);
nor U18063 (N_18063,N_10756,N_13968);
and U18064 (N_18064,N_11569,N_14164);
or U18065 (N_18065,N_14595,N_14949);
and U18066 (N_18066,N_14681,N_13361);
nand U18067 (N_18067,N_10061,N_14278);
or U18068 (N_18068,N_13492,N_14012);
or U18069 (N_18069,N_12847,N_14883);
or U18070 (N_18070,N_13413,N_13357);
nor U18071 (N_18071,N_12604,N_10923);
and U18072 (N_18072,N_11349,N_10516);
nor U18073 (N_18073,N_10719,N_11349);
nor U18074 (N_18074,N_13249,N_13085);
nor U18075 (N_18075,N_10939,N_12080);
and U18076 (N_18076,N_14762,N_11148);
xnor U18077 (N_18077,N_11305,N_12118);
and U18078 (N_18078,N_14719,N_12257);
nand U18079 (N_18079,N_12435,N_11472);
xnor U18080 (N_18080,N_14170,N_14115);
nor U18081 (N_18081,N_14904,N_14689);
or U18082 (N_18082,N_10444,N_10952);
xnor U18083 (N_18083,N_12684,N_13899);
nand U18084 (N_18084,N_14123,N_13335);
xnor U18085 (N_18085,N_12293,N_13922);
xor U18086 (N_18086,N_13341,N_14883);
or U18087 (N_18087,N_11694,N_10875);
xnor U18088 (N_18088,N_12300,N_12040);
nand U18089 (N_18089,N_14195,N_13171);
or U18090 (N_18090,N_12514,N_10539);
xor U18091 (N_18091,N_12639,N_13706);
nand U18092 (N_18092,N_14530,N_13263);
xor U18093 (N_18093,N_13958,N_10329);
nor U18094 (N_18094,N_11674,N_13592);
or U18095 (N_18095,N_12070,N_12505);
nand U18096 (N_18096,N_13752,N_11788);
or U18097 (N_18097,N_11414,N_10123);
or U18098 (N_18098,N_12747,N_13601);
or U18099 (N_18099,N_14769,N_13371);
nand U18100 (N_18100,N_11064,N_13120);
and U18101 (N_18101,N_10567,N_14866);
nand U18102 (N_18102,N_13734,N_12097);
nor U18103 (N_18103,N_14641,N_13946);
nand U18104 (N_18104,N_13069,N_13007);
and U18105 (N_18105,N_14805,N_14499);
nand U18106 (N_18106,N_11089,N_10112);
nand U18107 (N_18107,N_13216,N_13355);
nor U18108 (N_18108,N_12001,N_13803);
nor U18109 (N_18109,N_10531,N_12881);
or U18110 (N_18110,N_12684,N_13229);
nand U18111 (N_18111,N_14625,N_14671);
or U18112 (N_18112,N_14247,N_13457);
or U18113 (N_18113,N_12251,N_11408);
or U18114 (N_18114,N_14108,N_10489);
or U18115 (N_18115,N_12167,N_14660);
or U18116 (N_18116,N_13455,N_11069);
or U18117 (N_18117,N_12419,N_13085);
or U18118 (N_18118,N_11353,N_13319);
or U18119 (N_18119,N_11701,N_14086);
or U18120 (N_18120,N_13439,N_14138);
or U18121 (N_18121,N_12943,N_12976);
and U18122 (N_18122,N_12736,N_13889);
xor U18123 (N_18123,N_14032,N_13800);
xor U18124 (N_18124,N_11694,N_14147);
nand U18125 (N_18125,N_10152,N_14865);
or U18126 (N_18126,N_14036,N_13634);
xor U18127 (N_18127,N_10431,N_12920);
xor U18128 (N_18128,N_11201,N_12011);
nor U18129 (N_18129,N_11033,N_10230);
xor U18130 (N_18130,N_13788,N_10253);
nor U18131 (N_18131,N_12911,N_11991);
nor U18132 (N_18132,N_12273,N_13253);
nand U18133 (N_18133,N_11207,N_11141);
and U18134 (N_18134,N_11734,N_10361);
or U18135 (N_18135,N_12471,N_10098);
or U18136 (N_18136,N_13708,N_14071);
or U18137 (N_18137,N_11212,N_10992);
nand U18138 (N_18138,N_13941,N_12471);
nor U18139 (N_18139,N_13073,N_14190);
and U18140 (N_18140,N_10414,N_10870);
or U18141 (N_18141,N_12758,N_12840);
or U18142 (N_18142,N_14077,N_12000);
nand U18143 (N_18143,N_10581,N_12974);
nor U18144 (N_18144,N_14424,N_11866);
or U18145 (N_18145,N_10076,N_13119);
and U18146 (N_18146,N_14946,N_13907);
nand U18147 (N_18147,N_11420,N_14713);
nor U18148 (N_18148,N_13612,N_13340);
xnor U18149 (N_18149,N_14907,N_10513);
nor U18150 (N_18150,N_10328,N_14497);
xnor U18151 (N_18151,N_13417,N_11996);
nand U18152 (N_18152,N_11341,N_11109);
and U18153 (N_18153,N_12744,N_10868);
nor U18154 (N_18154,N_11452,N_14863);
or U18155 (N_18155,N_14086,N_10865);
or U18156 (N_18156,N_12411,N_12910);
or U18157 (N_18157,N_14149,N_11163);
nand U18158 (N_18158,N_11824,N_13680);
nor U18159 (N_18159,N_13344,N_11364);
nand U18160 (N_18160,N_11146,N_12811);
xor U18161 (N_18161,N_13877,N_11024);
xor U18162 (N_18162,N_14852,N_12006);
or U18163 (N_18163,N_11449,N_11884);
xor U18164 (N_18164,N_11762,N_14524);
nand U18165 (N_18165,N_11266,N_10645);
and U18166 (N_18166,N_12854,N_14447);
xnor U18167 (N_18167,N_11421,N_14807);
nor U18168 (N_18168,N_12794,N_10264);
nand U18169 (N_18169,N_13947,N_10503);
nand U18170 (N_18170,N_13833,N_14345);
xnor U18171 (N_18171,N_11179,N_14426);
nand U18172 (N_18172,N_13367,N_14040);
xor U18173 (N_18173,N_13178,N_11568);
nand U18174 (N_18174,N_12315,N_13231);
nand U18175 (N_18175,N_13760,N_10887);
nand U18176 (N_18176,N_11242,N_14221);
or U18177 (N_18177,N_10905,N_12469);
nor U18178 (N_18178,N_14988,N_13154);
xor U18179 (N_18179,N_14837,N_11615);
nor U18180 (N_18180,N_12319,N_11355);
nor U18181 (N_18181,N_13257,N_12949);
xnor U18182 (N_18182,N_13017,N_12565);
xnor U18183 (N_18183,N_11622,N_13280);
nand U18184 (N_18184,N_11446,N_12890);
and U18185 (N_18185,N_11091,N_11575);
and U18186 (N_18186,N_10449,N_12454);
nand U18187 (N_18187,N_10086,N_11823);
or U18188 (N_18188,N_14023,N_11737);
or U18189 (N_18189,N_11535,N_13070);
nand U18190 (N_18190,N_13858,N_13479);
nand U18191 (N_18191,N_10992,N_14945);
or U18192 (N_18192,N_11188,N_10583);
nor U18193 (N_18193,N_12950,N_12601);
nor U18194 (N_18194,N_10297,N_12436);
and U18195 (N_18195,N_11572,N_13065);
or U18196 (N_18196,N_12907,N_11429);
and U18197 (N_18197,N_14384,N_10183);
nor U18198 (N_18198,N_11173,N_11911);
nor U18199 (N_18199,N_10821,N_14144);
xor U18200 (N_18200,N_12719,N_13633);
and U18201 (N_18201,N_13524,N_11874);
nor U18202 (N_18202,N_14106,N_14581);
nand U18203 (N_18203,N_10785,N_13486);
nor U18204 (N_18204,N_11388,N_13013);
nor U18205 (N_18205,N_10874,N_11332);
nand U18206 (N_18206,N_10635,N_13901);
nor U18207 (N_18207,N_13586,N_11321);
nor U18208 (N_18208,N_12483,N_11205);
nand U18209 (N_18209,N_11524,N_10490);
nor U18210 (N_18210,N_10765,N_10299);
xor U18211 (N_18211,N_12098,N_12748);
nor U18212 (N_18212,N_13027,N_10274);
nand U18213 (N_18213,N_13351,N_13012);
nor U18214 (N_18214,N_10741,N_11543);
or U18215 (N_18215,N_14552,N_14809);
xor U18216 (N_18216,N_10671,N_12756);
or U18217 (N_18217,N_13315,N_12430);
or U18218 (N_18218,N_11265,N_11930);
xnor U18219 (N_18219,N_10828,N_13102);
xor U18220 (N_18220,N_10098,N_13398);
nand U18221 (N_18221,N_11706,N_12591);
nor U18222 (N_18222,N_11050,N_13066);
nand U18223 (N_18223,N_10633,N_13342);
nand U18224 (N_18224,N_12859,N_14580);
and U18225 (N_18225,N_13441,N_12527);
nand U18226 (N_18226,N_12936,N_13385);
xnor U18227 (N_18227,N_12214,N_11690);
or U18228 (N_18228,N_14657,N_13419);
nor U18229 (N_18229,N_10776,N_10639);
or U18230 (N_18230,N_13996,N_13546);
nand U18231 (N_18231,N_12638,N_11549);
nand U18232 (N_18232,N_11790,N_13318);
nor U18233 (N_18233,N_12519,N_10524);
nand U18234 (N_18234,N_11083,N_14462);
or U18235 (N_18235,N_14199,N_12892);
and U18236 (N_18236,N_13803,N_12554);
or U18237 (N_18237,N_10569,N_14869);
nand U18238 (N_18238,N_12542,N_11036);
or U18239 (N_18239,N_14596,N_11802);
xor U18240 (N_18240,N_14071,N_10348);
xnor U18241 (N_18241,N_10224,N_10005);
nand U18242 (N_18242,N_12821,N_14139);
nor U18243 (N_18243,N_13671,N_11668);
xnor U18244 (N_18244,N_14795,N_14494);
or U18245 (N_18245,N_12638,N_11957);
nand U18246 (N_18246,N_14896,N_11442);
and U18247 (N_18247,N_12217,N_13518);
nand U18248 (N_18248,N_12797,N_10551);
xnor U18249 (N_18249,N_11444,N_10512);
xor U18250 (N_18250,N_10619,N_11144);
nand U18251 (N_18251,N_10438,N_13672);
or U18252 (N_18252,N_13167,N_11593);
and U18253 (N_18253,N_11362,N_11251);
or U18254 (N_18254,N_13150,N_13358);
xor U18255 (N_18255,N_10075,N_10723);
or U18256 (N_18256,N_14275,N_10964);
and U18257 (N_18257,N_14945,N_13107);
nor U18258 (N_18258,N_13835,N_10262);
and U18259 (N_18259,N_12147,N_14397);
nand U18260 (N_18260,N_14007,N_11437);
or U18261 (N_18261,N_13834,N_13399);
or U18262 (N_18262,N_14360,N_14502);
nand U18263 (N_18263,N_13413,N_13728);
and U18264 (N_18264,N_14201,N_12707);
and U18265 (N_18265,N_12135,N_14445);
xnor U18266 (N_18266,N_14064,N_11563);
nor U18267 (N_18267,N_10080,N_14921);
nor U18268 (N_18268,N_14632,N_14368);
xnor U18269 (N_18269,N_11932,N_11519);
or U18270 (N_18270,N_14268,N_11499);
xor U18271 (N_18271,N_12133,N_10522);
and U18272 (N_18272,N_14486,N_11635);
nand U18273 (N_18273,N_13783,N_14964);
xor U18274 (N_18274,N_14866,N_10124);
nand U18275 (N_18275,N_10440,N_10388);
or U18276 (N_18276,N_12219,N_11315);
or U18277 (N_18277,N_14243,N_10808);
xnor U18278 (N_18278,N_14145,N_11466);
nor U18279 (N_18279,N_10174,N_12473);
nor U18280 (N_18280,N_12498,N_11502);
xnor U18281 (N_18281,N_14737,N_14617);
nor U18282 (N_18282,N_12365,N_14951);
and U18283 (N_18283,N_13993,N_11255);
or U18284 (N_18284,N_11324,N_11441);
and U18285 (N_18285,N_12850,N_14861);
nor U18286 (N_18286,N_11209,N_12271);
and U18287 (N_18287,N_14207,N_11541);
and U18288 (N_18288,N_12295,N_13605);
and U18289 (N_18289,N_11670,N_12478);
nor U18290 (N_18290,N_14900,N_12477);
nand U18291 (N_18291,N_13970,N_14990);
xnor U18292 (N_18292,N_14293,N_12042);
nor U18293 (N_18293,N_10283,N_11583);
nand U18294 (N_18294,N_11588,N_12595);
xnor U18295 (N_18295,N_10807,N_11372);
or U18296 (N_18296,N_14766,N_13733);
or U18297 (N_18297,N_13641,N_14272);
xor U18298 (N_18298,N_11720,N_13803);
nand U18299 (N_18299,N_13041,N_11569);
or U18300 (N_18300,N_13822,N_14463);
and U18301 (N_18301,N_12301,N_14189);
xor U18302 (N_18302,N_12680,N_13051);
and U18303 (N_18303,N_10396,N_13393);
xnor U18304 (N_18304,N_12937,N_13663);
or U18305 (N_18305,N_12583,N_13959);
xor U18306 (N_18306,N_11911,N_11734);
or U18307 (N_18307,N_14644,N_13970);
nor U18308 (N_18308,N_11826,N_13878);
or U18309 (N_18309,N_13782,N_14914);
and U18310 (N_18310,N_11239,N_10760);
and U18311 (N_18311,N_10788,N_14110);
and U18312 (N_18312,N_10670,N_10922);
or U18313 (N_18313,N_13470,N_13922);
and U18314 (N_18314,N_13101,N_11859);
nor U18315 (N_18315,N_13051,N_13604);
nor U18316 (N_18316,N_12555,N_12940);
and U18317 (N_18317,N_14888,N_10427);
nand U18318 (N_18318,N_11837,N_13649);
nand U18319 (N_18319,N_10794,N_13226);
nor U18320 (N_18320,N_11043,N_10851);
and U18321 (N_18321,N_11663,N_11270);
nand U18322 (N_18322,N_14112,N_12009);
xor U18323 (N_18323,N_11829,N_14795);
nand U18324 (N_18324,N_10280,N_11658);
nand U18325 (N_18325,N_11371,N_14775);
or U18326 (N_18326,N_14264,N_11266);
nor U18327 (N_18327,N_10369,N_12651);
or U18328 (N_18328,N_11561,N_10659);
nor U18329 (N_18329,N_14980,N_13051);
nand U18330 (N_18330,N_13890,N_14351);
xnor U18331 (N_18331,N_13049,N_12938);
xor U18332 (N_18332,N_11760,N_11284);
or U18333 (N_18333,N_12156,N_14921);
nand U18334 (N_18334,N_13278,N_14015);
and U18335 (N_18335,N_12302,N_13547);
xor U18336 (N_18336,N_14576,N_11251);
nand U18337 (N_18337,N_11628,N_13293);
and U18338 (N_18338,N_12463,N_13088);
and U18339 (N_18339,N_10045,N_11740);
and U18340 (N_18340,N_11349,N_10372);
xnor U18341 (N_18341,N_11353,N_13932);
nor U18342 (N_18342,N_11872,N_10531);
nor U18343 (N_18343,N_14200,N_14859);
nor U18344 (N_18344,N_12452,N_12983);
nor U18345 (N_18345,N_10511,N_10070);
nand U18346 (N_18346,N_14976,N_12663);
or U18347 (N_18347,N_13090,N_10889);
and U18348 (N_18348,N_14342,N_13312);
or U18349 (N_18349,N_10886,N_12586);
nor U18350 (N_18350,N_14364,N_13835);
and U18351 (N_18351,N_14053,N_14593);
xnor U18352 (N_18352,N_14902,N_14171);
nor U18353 (N_18353,N_14209,N_10193);
xor U18354 (N_18354,N_10371,N_12357);
nand U18355 (N_18355,N_14710,N_14346);
xor U18356 (N_18356,N_14718,N_12607);
and U18357 (N_18357,N_13623,N_12150);
nor U18358 (N_18358,N_13002,N_14684);
nand U18359 (N_18359,N_14201,N_12958);
or U18360 (N_18360,N_13763,N_11179);
nor U18361 (N_18361,N_10186,N_11859);
and U18362 (N_18362,N_10092,N_14983);
nor U18363 (N_18363,N_10056,N_13921);
nand U18364 (N_18364,N_12080,N_10819);
or U18365 (N_18365,N_12958,N_10289);
nand U18366 (N_18366,N_14411,N_13316);
xor U18367 (N_18367,N_10447,N_14273);
xor U18368 (N_18368,N_14274,N_13044);
or U18369 (N_18369,N_10575,N_14639);
xor U18370 (N_18370,N_10842,N_12492);
nand U18371 (N_18371,N_10789,N_11450);
xnor U18372 (N_18372,N_12826,N_13436);
and U18373 (N_18373,N_14717,N_13718);
and U18374 (N_18374,N_14888,N_14042);
nor U18375 (N_18375,N_14256,N_10008);
and U18376 (N_18376,N_11963,N_12179);
or U18377 (N_18377,N_12135,N_10528);
nand U18378 (N_18378,N_13578,N_14647);
nor U18379 (N_18379,N_10886,N_12326);
or U18380 (N_18380,N_12740,N_10770);
nor U18381 (N_18381,N_12803,N_10871);
and U18382 (N_18382,N_11759,N_14621);
xnor U18383 (N_18383,N_13286,N_10726);
xnor U18384 (N_18384,N_11678,N_14449);
nand U18385 (N_18385,N_13826,N_14982);
nor U18386 (N_18386,N_14655,N_14837);
and U18387 (N_18387,N_12273,N_10991);
or U18388 (N_18388,N_10181,N_11161);
nand U18389 (N_18389,N_12742,N_12143);
nand U18390 (N_18390,N_14788,N_14992);
or U18391 (N_18391,N_10771,N_10952);
xor U18392 (N_18392,N_13481,N_11694);
or U18393 (N_18393,N_14625,N_14183);
nand U18394 (N_18394,N_12132,N_12379);
and U18395 (N_18395,N_12117,N_11059);
or U18396 (N_18396,N_11235,N_13200);
and U18397 (N_18397,N_13183,N_14435);
xnor U18398 (N_18398,N_13125,N_10347);
xor U18399 (N_18399,N_14803,N_11858);
or U18400 (N_18400,N_13409,N_11842);
and U18401 (N_18401,N_11784,N_11636);
nor U18402 (N_18402,N_14940,N_10698);
nor U18403 (N_18403,N_14291,N_13349);
and U18404 (N_18404,N_11861,N_11475);
xnor U18405 (N_18405,N_10104,N_11208);
nor U18406 (N_18406,N_12993,N_14244);
nand U18407 (N_18407,N_12292,N_14454);
nand U18408 (N_18408,N_13187,N_11648);
xnor U18409 (N_18409,N_11744,N_10955);
or U18410 (N_18410,N_10122,N_13350);
or U18411 (N_18411,N_10328,N_11753);
or U18412 (N_18412,N_14891,N_14067);
or U18413 (N_18413,N_13469,N_13327);
or U18414 (N_18414,N_11336,N_11380);
nor U18415 (N_18415,N_10067,N_10945);
nand U18416 (N_18416,N_10347,N_11981);
or U18417 (N_18417,N_14159,N_10920);
xor U18418 (N_18418,N_10253,N_13655);
nand U18419 (N_18419,N_14691,N_13837);
nand U18420 (N_18420,N_13807,N_10508);
xnor U18421 (N_18421,N_12030,N_13238);
nand U18422 (N_18422,N_13259,N_13660);
xnor U18423 (N_18423,N_13618,N_13865);
or U18424 (N_18424,N_10296,N_12056);
and U18425 (N_18425,N_14912,N_11581);
and U18426 (N_18426,N_12198,N_14775);
and U18427 (N_18427,N_14108,N_11760);
nand U18428 (N_18428,N_10824,N_10306);
nor U18429 (N_18429,N_11017,N_11453);
or U18430 (N_18430,N_12420,N_12227);
xnor U18431 (N_18431,N_11190,N_10680);
xor U18432 (N_18432,N_13056,N_10557);
nor U18433 (N_18433,N_13308,N_11387);
nor U18434 (N_18434,N_14195,N_10039);
xor U18435 (N_18435,N_14923,N_12038);
or U18436 (N_18436,N_10718,N_14542);
nand U18437 (N_18437,N_11616,N_13270);
nor U18438 (N_18438,N_11801,N_13817);
and U18439 (N_18439,N_11193,N_11767);
nand U18440 (N_18440,N_13022,N_13578);
or U18441 (N_18441,N_10912,N_13175);
nand U18442 (N_18442,N_12329,N_13534);
nand U18443 (N_18443,N_11453,N_14680);
and U18444 (N_18444,N_10587,N_10270);
nand U18445 (N_18445,N_11510,N_12954);
or U18446 (N_18446,N_11764,N_12322);
and U18447 (N_18447,N_14555,N_10068);
nand U18448 (N_18448,N_10470,N_11250);
nand U18449 (N_18449,N_11206,N_10406);
and U18450 (N_18450,N_13736,N_12811);
or U18451 (N_18451,N_14575,N_11839);
nand U18452 (N_18452,N_14925,N_10518);
nand U18453 (N_18453,N_10383,N_12659);
or U18454 (N_18454,N_12586,N_11668);
or U18455 (N_18455,N_13580,N_14130);
xor U18456 (N_18456,N_11609,N_11153);
or U18457 (N_18457,N_13404,N_12218);
and U18458 (N_18458,N_11323,N_14062);
and U18459 (N_18459,N_10566,N_11926);
xor U18460 (N_18460,N_14668,N_12458);
nor U18461 (N_18461,N_13415,N_12275);
and U18462 (N_18462,N_10035,N_12850);
and U18463 (N_18463,N_12631,N_11722);
and U18464 (N_18464,N_14154,N_12652);
and U18465 (N_18465,N_11966,N_10982);
or U18466 (N_18466,N_10182,N_10175);
nand U18467 (N_18467,N_13548,N_12285);
and U18468 (N_18468,N_10855,N_14630);
or U18469 (N_18469,N_10187,N_14103);
or U18470 (N_18470,N_12404,N_10003);
nor U18471 (N_18471,N_12176,N_10114);
xnor U18472 (N_18472,N_13572,N_10409);
nor U18473 (N_18473,N_12997,N_10694);
nand U18474 (N_18474,N_13884,N_12024);
nor U18475 (N_18475,N_12914,N_10852);
xor U18476 (N_18476,N_13729,N_13609);
nor U18477 (N_18477,N_11684,N_12250);
nor U18478 (N_18478,N_14762,N_13370);
and U18479 (N_18479,N_10102,N_13234);
and U18480 (N_18480,N_12622,N_14839);
nand U18481 (N_18481,N_10706,N_14756);
nor U18482 (N_18482,N_10190,N_12055);
or U18483 (N_18483,N_13076,N_14594);
nand U18484 (N_18484,N_12011,N_12512);
xnor U18485 (N_18485,N_12720,N_10465);
or U18486 (N_18486,N_14758,N_11842);
or U18487 (N_18487,N_12466,N_10989);
nor U18488 (N_18488,N_11988,N_14009);
nor U18489 (N_18489,N_12309,N_13419);
nor U18490 (N_18490,N_12397,N_10690);
or U18491 (N_18491,N_12062,N_10684);
or U18492 (N_18492,N_11801,N_11211);
nor U18493 (N_18493,N_12404,N_10475);
nor U18494 (N_18494,N_10845,N_10112);
nor U18495 (N_18495,N_12616,N_10747);
nand U18496 (N_18496,N_13530,N_12861);
or U18497 (N_18497,N_10525,N_11928);
and U18498 (N_18498,N_14175,N_12140);
or U18499 (N_18499,N_10590,N_13413);
nor U18500 (N_18500,N_10015,N_11333);
and U18501 (N_18501,N_12113,N_14224);
or U18502 (N_18502,N_10164,N_11156);
nand U18503 (N_18503,N_10635,N_11830);
xor U18504 (N_18504,N_12465,N_13995);
nor U18505 (N_18505,N_12704,N_14276);
and U18506 (N_18506,N_12180,N_14254);
nand U18507 (N_18507,N_13624,N_13009);
nor U18508 (N_18508,N_14650,N_10521);
or U18509 (N_18509,N_13095,N_11044);
nor U18510 (N_18510,N_14992,N_13728);
or U18511 (N_18511,N_13980,N_14840);
nor U18512 (N_18512,N_10567,N_13153);
and U18513 (N_18513,N_11708,N_10850);
nand U18514 (N_18514,N_11313,N_13202);
or U18515 (N_18515,N_10703,N_14669);
or U18516 (N_18516,N_11001,N_12012);
and U18517 (N_18517,N_10691,N_10664);
xor U18518 (N_18518,N_10089,N_14354);
and U18519 (N_18519,N_13066,N_11495);
nand U18520 (N_18520,N_11795,N_10410);
xor U18521 (N_18521,N_10985,N_12895);
or U18522 (N_18522,N_11712,N_10461);
nand U18523 (N_18523,N_12102,N_14330);
or U18524 (N_18524,N_11634,N_12791);
nand U18525 (N_18525,N_10045,N_11545);
or U18526 (N_18526,N_11781,N_13825);
xnor U18527 (N_18527,N_14457,N_10887);
and U18528 (N_18528,N_11144,N_10136);
and U18529 (N_18529,N_13030,N_14660);
or U18530 (N_18530,N_14795,N_13208);
nor U18531 (N_18531,N_10876,N_10386);
nor U18532 (N_18532,N_14340,N_13441);
nor U18533 (N_18533,N_13144,N_12099);
nand U18534 (N_18534,N_13551,N_14763);
or U18535 (N_18535,N_14277,N_14722);
nand U18536 (N_18536,N_14282,N_12658);
nand U18537 (N_18537,N_13112,N_10947);
xor U18538 (N_18538,N_10552,N_13289);
and U18539 (N_18539,N_14921,N_12577);
nor U18540 (N_18540,N_11722,N_11883);
nand U18541 (N_18541,N_11610,N_10292);
or U18542 (N_18542,N_14761,N_11177);
or U18543 (N_18543,N_11624,N_10914);
nand U18544 (N_18544,N_11082,N_12989);
nand U18545 (N_18545,N_13067,N_11972);
xnor U18546 (N_18546,N_14833,N_14798);
nand U18547 (N_18547,N_14148,N_14449);
xor U18548 (N_18548,N_14068,N_11562);
nor U18549 (N_18549,N_13880,N_10869);
xnor U18550 (N_18550,N_10015,N_12539);
xnor U18551 (N_18551,N_13650,N_11954);
and U18552 (N_18552,N_13916,N_13849);
and U18553 (N_18553,N_14828,N_10413);
xor U18554 (N_18554,N_10300,N_10367);
and U18555 (N_18555,N_12262,N_11409);
nor U18556 (N_18556,N_13469,N_12766);
nand U18557 (N_18557,N_10220,N_12816);
xnor U18558 (N_18558,N_11418,N_13357);
nor U18559 (N_18559,N_13229,N_10064);
xnor U18560 (N_18560,N_11767,N_13484);
nand U18561 (N_18561,N_13253,N_13080);
nand U18562 (N_18562,N_14009,N_13571);
nor U18563 (N_18563,N_11767,N_14936);
xnor U18564 (N_18564,N_14919,N_10358);
xor U18565 (N_18565,N_13623,N_12029);
xnor U18566 (N_18566,N_10870,N_13097);
nor U18567 (N_18567,N_14787,N_11331);
xnor U18568 (N_18568,N_11792,N_10564);
xor U18569 (N_18569,N_12783,N_10042);
or U18570 (N_18570,N_14018,N_13401);
xor U18571 (N_18571,N_14526,N_11970);
xor U18572 (N_18572,N_14636,N_11127);
xor U18573 (N_18573,N_13645,N_12501);
or U18574 (N_18574,N_14473,N_10982);
or U18575 (N_18575,N_12882,N_14819);
or U18576 (N_18576,N_11554,N_11016);
and U18577 (N_18577,N_12993,N_14317);
xor U18578 (N_18578,N_12870,N_13472);
or U18579 (N_18579,N_13515,N_11460);
or U18580 (N_18580,N_14925,N_12274);
or U18581 (N_18581,N_14928,N_12803);
or U18582 (N_18582,N_10945,N_13425);
nor U18583 (N_18583,N_14093,N_10424);
or U18584 (N_18584,N_13152,N_10393);
xnor U18585 (N_18585,N_12353,N_12730);
or U18586 (N_18586,N_12209,N_11965);
nand U18587 (N_18587,N_13705,N_10725);
or U18588 (N_18588,N_12889,N_12051);
nor U18589 (N_18589,N_13196,N_12399);
nand U18590 (N_18590,N_14433,N_14197);
and U18591 (N_18591,N_11449,N_13796);
nor U18592 (N_18592,N_13083,N_11769);
nor U18593 (N_18593,N_11124,N_14219);
and U18594 (N_18594,N_11273,N_11311);
or U18595 (N_18595,N_10929,N_13888);
nor U18596 (N_18596,N_14105,N_14184);
nand U18597 (N_18597,N_10801,N_10233);
xnor U18598 (N_18598,N_12731,N_14828);
and U18599 (N_18599,N_12442,N_14433);
nand U18600 (N_18600,N_10806,N_13754);
xor U18601 (N_18601,N_10331,N_13594);
nor U18602 (N_18602,N_10019,N_11528);
nand U18603 (N_18603,N_14710,N_12488);
or U18604 (N_18604,N_14824,N_14746);
and U18605 (N_18605,N_11461,N_10602);
or U18606 (N_18606,N_13480,N_11521);
or U18607 (N_18607,N_12701,N_10042);
xnor U18608 (N_18608,N_12145,N_11782);
or U18609 (N_18609,N_13106,N_14152);
nand U18610 (N_18610,N_12306,N_10862);
and U18611 (N_18611,N_11590,N_11033);
nor U18612 (N_18612,N_14486,N_12796);
nand U18613 (N_18613,N_11689,N_10979);
and U18614 (N_18614,N_13261,N_12992);
and U18615 (N_18615,N_10924,N_10741);
or U18616 (N_18616,N_14469,N_10248);
nor U18617 (N_18617,N_11205,N_13926);
xnor U18618 (N_18618,N_14569,N_10995);
nand U18619 (N_18619,N_13744,N_10290);
nand U18620 (N_18620,N_10708,N_10344);
or U18621 (N_18621,N_13684,N_12923);
nor U18622 (N_18622,N_13736,N_14523);
and U18623 (N_18623,N_11885,N_13296);
nand U18624 (N_18624,N_10349,N_12207);
and U18625 (N_18625,N_10735,N_11315);
or U18626 (N_18626,N_13463,N_13148);
nor U18627 (N_18627,N_11975,N_11991);
nor U18628 (N_18628,N_12771,N_13208);
nand U18629 (N_18629,N_14625,N_11709);
nor U18630 (N_18630,N_13341,N_14300);
and U18631 (N_18631,N_14897,N_13664);
and U18632 (N_18632,N_11034,N_12145);
and U18633 (N_18633,N_14195,N_14036);
nor U18634 (N_18634,N_10550,N_14123);
or U18635 (N_18635,N_11037,N_10531);
nand U18636 (N_18636,N_13371,N_13353);
or U18637 (N_18637,N_14183,N_12976);
nor U18638 (N_18638,N_14552,N_13430);
or U18639 (N_18639,N_10906,N_10282);
or U18640 (N_18640,N_13164,N_14865);
nor U18641 (N_18641,N_11120,N_10769);
nand U18642 (N_18642,N_13456,N_10295);
and U18643 (N_18643,N_12501,N_11292);
nor U18644 (N_18644,N_10578,N_12069);
nor U18645 (N_18645,N_10355,N_14713);
nand U18646 (N_18646,N_11534,N_10625);
and U18647 (N_18647,N_12718,N_10318);
and U18648 (N_18648,N_12290,N_12527);
xor U18649 (N_18649,N_14558,N_12214);
or U18650 (N_18650,N_11204,N_14174);
or U18651 (N_18651,N_11127,N_12518);
nor U18652 (N_18652,N_13271,N_13432);
nor U18653 (N_18653,N_11451,N_11475);
and U18654 (N_18654,N_13000,N_13342);
or U18655 (N_18655,N_13515,N_13537);
or U18656 (N_18656,N_12250,N_13682);
nand U18657 (N_18657,N_13578,N_12762);
nand U18658 (N_18658,N_11897,N_12160);
or U18659 (N_18659,N_11442,N_10351);
xnor U18660 (N_18660,N_10137,N_11438);
and U18661 (N_18661,N_13813,N_10615);
and U18662 (N_18662,N_14938,N_11988);
xor U18663 (N_18663,N_13902,N_11861);
or U18664 (N_18664,N_13200,N_10589);
or U18665 (N_18665,N_11169,N_14770);
and U18666 (N_18666,N_14564,N_11386);
or U18667 (N_18667,N_14057,N_12828);
or U18668 (N_18668,N_14983,N_10454);
and U18669 (N_18669,N_14001,N_14422);
nand U18670 (N_18670,N_12987,N_10751);
and U18671 (N_18671,N_11482,N_13112);
xnor U18672 (N_18672,N_10265,N_13817);
nor U18673 (N_18673,N_12404,N_11828);
nand U18674 (N_18674,N_13683,N_12706);
nand U18675 (N_18675,N_10061,N_10342);
and U18676 (N_18676,N_10355,N_14807);
and U18677 (N_18677,N_14397,N_12939);
and U18678 (N_18678,N_14693,N_11788);
nand U18679 (N_18679,N_12745,N_13395);
xnor U18680 (N_18680,N_12218,N_10189);
nor U18681 (N_18681,N_12944,N_13491);
or U18682 (N_18682,N_14659,N_14912);
xnor U18683 (N_18683,N_14271,N_13544);
nand U18684 (N_18684,N_13871,N_12496);
nor U18685 (N_18685,N_14977,N_13202);
and U18686 (N_18686,N_13067,N_10244);
xor U18687 (N_18687,N_13603,N_14003);
and U18688 (N_18688,N_11109,N_14541);
nor U18689 (N_18689,N_14113,N_11343);
and U18690 (N_18690,N_11510,N_12729);
nor U18691 (N_18691,N_12984,N_11015);
or U18692 (N_18692,N_11563,N_10628);
nor U18693 (N_18693,N_10930,N_10443);
xnor U18694 (N_18694,N_11046,N_13957);
xnor U18695 (N_18695,N_11031,N_11029);
nand U18696 (N_18696,N_10518,N_13323);
or U18697 (N_18697,N_13283,N_11965);
nor U18698 (N_18698,N_12054,N_12301);
xor U18699 (N_18699,N_12974,N_11481);
or U18700 (N_18700,N_11378,N_14461);
or U18701 (N_18701,N_14906,N_13640);
xnor U18702 (N_18702,N_14263,N_13153);
nor U18703 (N_18703,N_11262,N_13576);
nor U18704 (N_18704,N_11380,N_13892);
nand U18705 (N_18705,N_14108,N_10281);
xnor U18706 (N_18706,N_11943,N_14298);
xor U18707 (N_18707,N_12243,N_11812);
or U18708 (N_18708,N_12254,N_11389);
or U18709 (N_18709,N_13499,N_11813);
and U18710 (N_18710,N_10927,N_14279);
nor U18711 (N_18711,N_14384,N_10776);
and U18712 (N_18712,N_14400,N_11825);
xnor U18713 (N_18713,N_14424,N_12764);
xnor U18714 (N_18714,N_13823,N_14555);
xnor U18715 (N_18715,N_10321,N_11260);
nor U18716 (N_18716,N_11562,N_13402);
nor U18717 (N_18717,N_14899,N_14796);
nand U18718 (N_18718,N_12676,N_13542);
xnor U18719 (N_18719,N_10631,N_11828);
or U18720 (N_18720,N_13608,N_12852);
and U18721 (N_18721,N_10283,N_10080);
or U18722 (N_18722,N_10982,N_11619);
and U18723 (N_18723,N_11882,N_12304);
nor U18724 (N_18724,N_10930,N_11189);
and U18725 (N_18725,N_13905,N_14188);
nor U18726 (N_18726,N_13822,N_12588);
xor U18727 (N_18727,N_12437,N_10346);
xnor U18728 (N_18728,N_12401,N_11591);
nand U18729 (N_18729,N_14113,N_11739);
and U18730 (N_18730,N_14616,N_14631);
and U18731 (N_18731,N_11228,N_13275);
xnor U18732 (N_18732,N_14121,N_11579);
xnor U18733 (N_18733,N_11085,N_12815);
nor U18734 (N_18734,N_11153,N_12194);
and U18735 (N_18735,N_11818,N_11455);
nand U18736 (N_18736,N_12233,N_13248);
or U18737 (N_18737,N_10687,N_13636);
or U18738 (N_18738,N_13368,N_12369);
and U18739 (N_18739,N_10183,N_11460);
xnor U18740 (N_18740,N_11999,N_13850);
xnor U18741 (N_18741,N_11557,N_11126);
and U18742 (N_18742,N_10225,N_14797);
xor U18743 (N_18743,N_14602,N_13824);
or U18744 (N_18744,N_10578,N_12257);
xor U18745 (N_18745,N_10929,N_14733);
nor U18746 (N_18746,N_14051,N_14495);
nor U18747 (N_18747,N_12091,N_11677);
xor U18748 (N_18748,N_13134,N_13730);
nor U18749 (N_18749,N_13649,N_14999);
or U18750 (N_18750,N_10804,N_14672);
xnor U18751 (N_18751,N_11820,N_14714);
and U18752 (N_18752,N_14443,N_12648);
xnor U18753 (N_18753,N_11014,N_12474);
nor U18754 (N_18754,N_13542,N_14275);
nand U18755 (N_18755,N_12221,N_13436);
and U18756 (N_18756,N_14875,N_13351);
nand U18757 (N_18757,N_12398,N_14216);
nor U18758 (N_18758,N_13171,N_13651);
and U18759 (N_18759,N_13174,N_14453);
or U18760 (N_18760,N_10461,N_13643);
nor U18761 (N_18761,N_11568,N_12290);
nor U18762 (N_18762,N_11738,N_11084);
xor U18763 (N_18763,N_13845,N_13409);
and U18764 (N_18764,N_10242,N_12150);
or U18765 (N_18765,N_12702,N_12846);
xnor U18766 (N_18766,N_13337,N_14928);
and U18767 (N_18767,N_11766,N_13479);
nor U18768 (N_18768,N_11134,N_11204);
and U18769 (N_18769,N_10726,N_11480);
or U18770 (N_18770,N_13379,N_10050);
nand U18771 (N_18771,N_13436,N_13328);
xnor U18772 (N_18772,N_12002,N_12229);
and U18773 (N_18773,N_12604,N_10593);
nand U18774 (N_18774,N_14032,N_14214);
nor U18775 (N_18775,N_14495,N_11084);
or U18776 (N_18776,N_12024,N_11941);
nor U18777 (N_18777,N_11120,N_10571);
or U18778 (N_18778,N_12475,N_12921);
or U18779 (N_18779,N_11094,N_10203);
and U18780 (N_18780,N_10703,N_13587);
xor U18781 (N_18781,N_13197,N_13608);
nor U18782 (N_18782,N_12464,N_10159);
nand U18783 (N_18783,N_12533,N_12171);
nand U18784 (N_18784,N_14711,N_14394);
nor U18785 (N_18785,N_12268,N_14252);
and U18786 (N_18786,N_10663,N_14785);
nand U18787 (N_18787,N_14738,N_14158);
xor U18788 (N_18788,N_13602,N_14224);
nand U18789 (N_18789,N_11561,N_10372);
and U18790 (N_18790,N_12225,N_14431);
or U18791 (N_18791,N_12575,N_13590);
nand U18792 (N_18792,N_13556,N_10204);
nand U18793 (N_18793,N_11850,N_10319);
and U18794 (N_18794,N_10033,N_14319);
xnor U18795 (N_18795,N_11565,N_12920);
xor U18796 (N_18796,N_12981,N_11696);
xnor U18797 (N_18797,N_13674,N_10418);
or U18798 (N_18798,N_10849,N_11441);
nand U18799 (N_18799,N_13795,N_11783);
or U18800 (N_18800,N_13572,N_13671);
or U18801 (N_18801,N_14898,N_14729);
nor U18802 (N_18802,N_11842,N_11698);
and U18803 (N_18803,N_13900,N_11351);
nand U18804 (N_18804,N_13728,N_11849);
nor U18805 (N_18805,N_10785,N_14397);
nor U18806 (N_18806,N_11499,N_14236);
nand U18807 (N_18807,N_10808,N_14006);
nor U18808 (N_18808,N_10943,N_14357);
nand U18809 (N_18809,N_11161,N_10058);
and U18810 (N_18810,N_14421,N_13709);
and U18811 (N_18811,N_11831,N_13331);
xnor U18812 (N_18812,N_12853,N_14217);
xnor U18813 (N_18813,N_13090,N_13187);
xor U18814 (N_18814,N_14011,N_14780);
xor U18815 (N_18815,N_13846,N_11731);
nand U18816 (N_18816,N_12877,N_11320);
nor U18817 (N_18817,N_14871,N_12109);
and U18818 (N_18818,N_10780,N_12537);
xor U18819 (N_18819,N_11379,N_14323);
nor U18820 (N_18820,N_14772,N_12992);
or U18821 (N_18821,N_13467,N_11126);
xor U18822 (N_18822,N_10852,N_12413);
nor U18823 (N_18823,N_13657,N_12603);
xor U18824 (N_18824,N_14059,N_13974);
nand U18825 (N_18825,N_14653,N_14513);
and U18826 (N_18826,N_11814,N_12749);
nor U18827 (N_18827,N_14679,N_13537);
or U18828 (N_18828,N_14570,N_14858);
and U18829 (N_18829,N_12116,N_13668);
xor U18830 (N_18830,N_12404,N_12659);
xor U18831 (N_18831,N_14505,N_12500);
xnor U18832 (N_18832,N_10212,N_12359);
or U18833 (N_18833,N_11742,N_13808);
and U18834 (N_18834,N_12081,N_12065);
or U18835 (N_18835,N_14257,N_13085);
or U18836 (N_18836,N_14495,N_11581);
nor U18837 (N_18837,N_11361,N_11493);
and U18838 (N_18838,N_11971,N_11653);
or U18839 (N_18839,N_12221,N_11017);
or U18840 (N_18840,N_14814,N_14999);
nor U18841 (N_18841,N_10986,N_14147);
and U18842 (N_18842,N_13793,N_14007);
or U18843 (N_18843,N_10922,N_14919);
or U18844 (N_18844,N_11755,N_11186);
xnor U18845 (N_18845,N_13678,N_13031);
and U18846 (N_18846,N_13509,N_14848);
and U18847 (N_18847,N_11992,N_10547);
and U18848 (N_18848,N_14375,N_11347);
and U18849 (N_18849,N_13887,N_14118);
and U18850 (N_18850,N_14236,N_10213);
or U18851 (N_18851,N_12481,N_14057);
nor U18852 (N_18852,N_14266,N_12153);
xnor U18853 (N_18853,N_10924,N_12235);
nor U18854 (N_18854,N_11743,N_14721);
nand U18855 (N_18855,N_12270,N_12666);
xor U18856 (N_18856,N_10033,N_14773);
nand U18857 (N_18857,N_14513,N_12083);
xor U18858 (N_18858,N_12052,N_10836);
or U18859 (N_18859,N_13834,N_12765);
nand U18860 (N_18860,N_11792,N_14510);
or U18861 (N_18861,N_12735,N_12266);
nor U18862 (N_18862,N_12362,N_11513);
or U18863 (N_18863,N_11457,N_14726);
nor U18864 (N_18864,N_13958,N_13102);
and U18865 (N_18865,N_10846,N_10163);
and U18866 (N_18866,N_12645,N_13918);
nor U18867 (N_18867,N_12199,N_10576);
and U18868 (N_18868,N_10970,N_12255);
nor U18869 (N_18869,N_14360,N_12110);
or U18870 (N_18870,N_12300,N_11935);
nor U18871 (N_18871,N_11463,N_14354);
nand U18872 (N_18872,N_12548,N_13723);
xor U18873 (N_18873,N_13323,N_10307);
nor U18874 (N_18874,N_11397,N_11851);
or U18875 (N_18875,N_11244,N_12510);
nor U18876 (N_18876,N_10225,N_10245);
xnor U18877 (N_18877,N_14229,N_12271);
nand U18878 (N_18878,N_13910,N_10457);
nor U18879 (N_18879,N_10277,N_11763);
and U18880 (N_18880,N_12844,N_14876);
nor U18881 (N_18881,N_11661,N_14055);
xor U18882 (N_18882,N_10216,N_10040);
nand U18883 (N_18883,N_13791,N_14589);
and U18884 (N_18884,N_11376,N_12645);
and U18885 (N_18885,N_13520,N_14906);
nand U18886 (N_18886,N_11899,N_13384);
or U18887 (N_18887,N_14534,N_12950);
or U18888 (N_18888,N_14350,N_14228);
or U18889 (N_18889,N_14016,N_13620);
xnor U18890 (N_18890,N_13757,N_14318);
nor U18891 (N_18891,N_13750,N_12666);
and U18892 (N_18892,N_11812,N_11282);
nand U18893 (N_18893,N_13225,N_12799);
nand U18894 (N_18894,N_12222,N_14564);
nor U18895 (N_18895,N_12166,N_10554);
xor U18896 (N_18896,N_13210,N_11359);
and U18897 (N_18897,N_11191,N_14427);
nand U18898 (N_18898,N_14637,N_11622);
nor U18899 (N_18899,N_12958,N_12086);
xnor U18900 (N_18900,N_11081,N_11516);
nor U18901 (N_18901,N_13673,N_10898);
and U18902 (N_18902,N_13920,N_12371);
and U18903 (N_18903,N_14563,N_14739);
nor U18904 (N_18904,N_11820,N_10833);
nor U18905 (N_18905,N_11739,N_11744);
nand U18906 (N_18906,N_11112,N_13180);
and U18907 (N_18907,N_13881,N_13400);
xor U18908 (N_18908,N_14270,N_12584);
nor U18909 (N_18909,N_14597,N_12615);
nor U18910 (N_18910,N_14759,N_12770);
nor U18911 (N_18911,N_12217,N_13409);
and U18912 (N_18912,N_11767,N_11366);
nor U18913 (N_18913,N_14829,N_14718);
and U18914 (N_18914,N_11433,N_11287);
and U18915 (N_18915,N_13325,N_11195);
nor U18916 (N_18916,N_13072,N_14216);
and U18917 (N_18917,N_11640,N_12173);
or U18918 (N_18918,N_13130,N_11867);
nor U18919 (N_18919,N_13157,N_13034);
xor U18920 (N_18920,N_12663,N_13053);
and U18921 (N_18921,N_10122,N_13468);
xor U18922 (N_18922,N_12926,N_10118);
or U18923 (N_18923,N_14467,N_14082);
nand U18924 (N_18924,N_10689,N_14827);
nor U18925 (N_18925,N_11197,N_14621);
and U18926 (N_18926,N_12906,N_14561);
or U18927 (N_18927,N_10875,N_11200);
xnor U18928 (N_18928,N_13254,N_10936);
nor U18929 (N_18929,N_10890,N_10480);
and U18930 (N_18930,N_14181,N_11221);
nor U18931 (N_18931,N_10439,N_11502);
xor U18932 (N_18932,N_10302,N_13028);
nand U18933 (N_18933,N_13200,N_13746);
or U18934 (N_18934,N_11273,N_14834);
and U18935 (N_18935,N_12381,N_11757);
and U18936 (N_18936,N_13992,N_12399);
xor U18937 (N_18937,N_10382,N_14910);
xor U18938 (N_18938,N_14020,N_12778);
xor U18939 (N_18939,N_12416,N_14278);
nor U18940 (N_18940,N_14268,N_13539);
or U18941 (N_18941,N_13873,N_11425);
and U18942 (N_18942,N_12662,N_11120);
or U18943 (N_18943,N_13643,N_14516);
xor U18944 (N_18944,N_12573,N_13714);
nor U18945 (N_18945,N_14327,N_10198);
nor U18946 (N_18946,N_13005,N_10659);
nand U18947 (N_18947,N_11039,N_13477);
nand U18948 (N_18948,N_10321,N_14602);
and U18949 (N_18949,N_10102,N_14343);
xnor U18950 (N_18950,N_14831,N_14843);
xnor U18951 (N_18951,N_14459,N_11854);
nor U18952 (N_18952,N_13103,N_12021);
nand U18953 (N_18953,N_14215,N_13333);
and U18954 (N_18954,N_10349,N_10915);
nand U18955 (N_18955,N_10185,N_10943);
and U18956 (N_18956,N_13499,N_10640);
xnor U18957 (N_18957,N_10954,N_10390);
xnor U18958 (N_18958,N_12187,N_11322);
nand U18959 (N_18959,N_12387,N_14649);
nor U18960 (N_18960,N_14851,N_11593);
and U18961 (N_18961,N_10212,N_11538);
xor U18962 (N_18962,N_14085,N_14430);
nand U18963 (N_18963,N_12705,N_10118);
xor U18964 (N_18964,N_13205,N_10709);
xor U18965 (N_18965,N_12555,N_13413);
nor U18966 (N_18966,N_14127,N_12772);
xnor U18967 (N_18967,N_13427,N_11570);
nand U18968 (N_18968,N_11689,N_12906);
and U18969 (N_18969,N_11474,N_12461);
nor U18970 (N_18970,N_12841,N_14145);
or U18971 (N_18971,N_11972,N_14930);
nand U18972 (N_18972,N_11427,N_12169);
nand U18973 (N_18973,N_14533,N_14765);
and U18974 (N_18974,N_12438,N_12763);
nand U18975 (N_18975,N_13452,N_11988);
nand U18976 (N_18976,N_12690,N_12773);
and U18977 (N_18977,N_11861,N_13818);
nor U18978 (N_18978,N_10822,N_11896);
nor U18979 (N_18979,N_11786,N_10925);
nand U18980 (N_18980,N_11172,N_12128);
or U18981 (N_18981,N_11611,N_13294);
and U18982 (N_18982,N_11444,N_11871);
and U18983 (N_18983,N_11213,N_11162);
or U18984 (N_18984,N_12565,N_11471);
nor U18985 (N_18985,N_14170,N_13794);
nand U18986 (N_18986,N_10122,N_10001);
and U18987 (N_18987,N_11323,N_11070);
or U18988 (N_18988,N_13489,N_10724);
xor U18989 (N_18989,N_12939,N_11842);
nor U18990 (N_18990,N_11669,N_12990);
nand U18991 (N_18991,N_11568,N_14842);
xor U18992 (N_18992,N_14018,N_14812);
nor U18993 (N_18993,N_14383,N_11976);
and U18994 (N_18994,N_10062,N_11093);
xor U18995 (N_18995,N_14455,N_11060);
nor U18996 (N_18996,N_12142,N_10833);
or U18997 (N_18997,N_10134,N_14221);
or U18998 (N_18998,N_10879,N_11851);
and U18999 (N_18999,N_11284,N_13963);
or U19000 (N_19000,N_13545,N_14445);
or U19001 (N_19001,N_11250,N_13818);
xnor U19002 (N_19002,N_11783,N_11162);
and U19003 (N_19003,N_11127,N_11948);
nand U19004 (N_19004,N_12715,N_10210);
nor U19005 (N_19005,N_14210,N_11646);
xnor U19006 (N_19006,N_12773,N_12302);
and U19007 (N_19007,N_10203,N_11766);
xor U19008 (N_19008,N_13159,N_11292);
xor U19009 (N_19009,N_10141,N_14446);
nor U19010 (N_19010,N_12245,N_14229);
or U19011 (N_19011,N_13107,N_11715);
nor U19012 (N_19012,N_11186,N_12077);
nand U19013 (N_19013,N_11731,N_13542);
or U19014 (N_19014,N_12861,N_11285);
xnor U19015 (N_19015,N_10127,N_11315);
nor U19016 (N_19016,N_14222,N_12287);
and U19017 (N_19017,N_11552,N_12206);
nand U19018 (N_19018,N_11962,N_13274);
xor U19019 (N_19019,N_12839,N_11378);
nand U19020 (N_19020,N_12998,N_12264);
xnor U19021 (N_19021,N_14343,N_14574);
xnor U19022 (N_19022,N_11773,N_14709);
or U19023 (N_19023,N_12306,N_13650);
nand U19024 (N_19024,N_12653,N_10273);
and U19025 (N_19025,N_12635,N_11532);
nand U19026 (N_19026,N_11237,N_10516);
nand U19027 (N_19027,N_14140,N_11318);
or U19028 (N_19028,N_10690,N_13597);
nand U19029 (N_19029,N_14592,N_14730);
nand U19030 (N_19030,N_14913,N_14916);
nand U19031 (N_19031,N_11976,N_13384);
and U19032 (N_19032,N_14241,N_11821);
and U19033 (N_19033,N_12637,N_14482);
xnor U19034 (N_19034,N_14192,N_13704);
or U19035 (N_19035,N_14451,N_10349);
nand U19036 (N_19036,N_11043,N_12638);
xnor U19037 (N_19037,N_10511,N_12312);
and U19038 (N_19038,N_12527,N_14410);
nand U19039 (N_19039,N_13051,N_11521);
and U19040 (N_19040,N_12760,N_12041);
nand U19041 (N_19041,N_14355,N_10289);
nand U19042 (N_19042,N_10872,N_10980);
nor U19043 (N_19043,N_13714,N_10384);
nor U19044 (N_19044,N_11673,N_14139);
or U19045 (N_19045,N_14029,N_10285);
or U19046 (N_19046,N_14539,N_14946);
or U19047 (N_19047,N_11074,N_14348);
xnor U19048 (N_19048,N_12369,N_12812);
and U19049 (N_19049,N_13328,N_11118);
nor U19050 (N_19050,N_11644,N_12595);
xnor U19051 (N_19051,N_12352,N_10500);
nand U19052 (N_19052,N_12754,N_10614);
or U19053 (N_19053,N_13095,N_13527);
and U19054 (N_19054,N_10838,N_13902);
nor U19055 (N_19055,N_11404,N_14562);
and U19056 (N_19056,N_13375,N_10163);
or U19057 (N_19057,N_10862,N_13174);
and U19058 (N_19058,N_10590,N_10365);
nor U19059 (N_19059,N_13642,N_13609);
or U19060 (N_19060,N_13417,N_13978);
nor U19061 (N_19061,N_12008,N_13450);
or U19062 (N_19062,N_10654,N_14113);
or U19063 (N_19063,N_12062,N_14648);
or U19064 (N_19064,N_11726,N_13415);
and U19065 (N_19065,N_13333,N_12462);
xor U19066 (N_19066,N_12735,N_13004);
xor U19067 (N_19067,N_14456,N_14283);
and U19068 (N_19068,N_14850,N_14401);
nor U19069 (N_19069,N_10539,N_11310);
and U19070 (N_19070,N_12025,N_10482);
nor U19071 (N_19071,N_14317,N_12482);
nor U19072 (N_19072,N_12024,N_11250);
nand U19073 (N_19073,N_11343,N_13808);
nor U19074 (N_19074,N_13765,N_13301);
or U19075 (N_19075,N_10736,N_12816);
xor U19076 (N_19076,N_10452,N_13902);
xor U19077 (N_19077,N_13920,N_10873);
xnor U19078 (N_19078,N_14131,N_12633);
nor U19079 (N_19079,N_12537,N_10068);
xnor U19080 (N_19080,N_10212,N_11322);
nand U19081 (N_19081,N_13169,N_12803);
or U19082 (N_19082,N_12411,N_12754);
or U19083 (N_19083,N_12940,N_14910);
nand U19084 (N_19084,N_13816,N_11188);
or U19085 (N_19085,N_12472,N_11186);
xnor U19086 (N_19086,N_11801,N_12258);
nor U19087 (N_19087,N_12290,N_11703);
and U19088 (N_19088,N_13651,N_12798);
and U19089 (N_19089,N_12545,N_14352);
and U19090 (N_19090,N_12260,N_10094);
xor U19091 (N_19091,N_14722,N_12437);
and U19092 (N_19092,N_13077,N_14265);
nand U19093 (N_19093,N_12391,N_11756);
xnor U19094 (N_19094,N_12834,N_14327);
or U19095 (N_19095,N_10334,N_14163);
nor U19096 (N_19096,N_14773,N_10320);
nand U19097 (N_19097,N_13284,N_14213);
nor U19098 (N_19098,N_14045,N_11416);
xor U19099 (N_19099,N_12365,N_13109);
and U19100 (N_19100,N_12144,N_13892);
and U19101 (N_19101,N_12820,N_14643);
xor U19102 (N_19102,N_13080,N_13125);
xnor U19103 (N_19103,N_11906,N_13070);
and U19104 (N_19104,N_11711,N_11945);
or U19105 (N_19105,N_12543,N_14346);
xnor U19106 (N_19106,N_14732,N_14044);
or U19107 (N_19107,N_11359,N_13670);
xnor U19108 (N_19108,N_10939,N_13858);
xnor U19109 (N_19109,N_11340,N_10063);
xnor U19110 (N_19110,N_10932,N_13291);
and U19111 (N_19111,N_14036,N_10216);
and U19112 (N_19112,N_12093,N_12776);
and U19113 (N_19113,N_11413,N_10715);
nor U19114 (N_19114,N_12048,N_10051);
or U19115 (N_19115,N_10553,N_11020);
nor U19116 (N_19116,N_13654,N_13175);
nand U19117 (N_19117,N_14910,N_12845);
and U19118 (N_19118,N_13214,N_12103);
xor U19119 (N_19119,N_14175,N_14649);
or U19120 (N_19120,N_14155,N_14087);
nand U19121 (N_19121,N_14044,N_11024);
nor U19122 (N_19122,N_13906,N_11761);
nor U19123 (N_19123,N_10422,N_11775);
nor U19124 (N_19124,N_12937,N_13615);
nor U19125 (N_19125,N_14002,N_14833);
or U19126 (N_19126,N_13878,N_12936);
and U19127 (N_19127,N_11489,N_13898);
xnor U19128 (N_19128,N_10619,N_11447);
xnor U19129 (N_19129,N_11418,N_11552);
nand U19130 (N_19130,N_12054,N_12190);
xor U19131 (N_19131,N_12732,N_11877);
nand U19132 (N_19132,N_12475,N_11785);
or U19133 (N_19133,N_12743,N_11653);
nor U19134 (N_19134,N_10822,N_10026);
and U19135 (N_19135,N_14682,N_13339);
or U19136 (N_19136,N_14797,N_10576);
or U19137 (N_19137,N_11147,N_13632);
nor U19138 (N_19138,N_14425,N_13809);
nand U19139 (N_19139,N_10542,N_13694);
or U19140 (N_19140,N_12417,N_10554);
xor U19141 (N_19141,N_10927,N_13062);
or U19142 (N_19142,N_11973,N_12743);
and U19143 (N_19143,N_12335,N_14016);
nand U19144 (N_19144,N_11516,N_12989);
and U19145 (N_19145,N_11267,N_13398);
nor U19146 (N_19146,N_12963,N_12592);
nor U19147 (N_19147,N_10865,N_11790);
or U19148 (N_19148,N_13083,N_13992);
or U19149 (N_19149,N_10512,N_10976);
xnor U19150 (N_19150,N_14115,N_13384);
and U19151 (N_19151,N_14213,N_11317);
or U19152 (N_19152,N_11094,N_14506);
nor U19153 (N_19153,N_14575,N_14063);
and U19154 (N_19154,N_12867,N_11804);
xor U19155 (N_19155,N_11108,N_11987);
nor U19156 (N_19156,N_14442,N_12888);
and U19157 (N_19157,N_12206,N_11819);
and U19158 (N_19158,N_13246,N_12229);
nand U19159 (N_19159,N_10616,N_12264);
or U19160 (N_19160,N_13970,N_12505);
nor U19161 (N_19161,N_14234,N_13803);
nor U19162 (N_19162,N_11132,N_10943);
xnor U19163 (N_19163,N_13685,N_11698);
nand U19164 (N_19164,N_12243,N_12298);
and U19165 (N_19165,N_14422,N_11669);
xor U19166 (N_19166,N_11142,N_11800);
nor U19167 (N_19167,N_12698,N_12661);
nand U19168 (N_19168,N_12707,N_12380);
or U19169 (N_19169,N_14438,N_12648);
or U19170 (N_19170,N_10263,N_11041);
nand U19171 (N_19171,N_10837,N_12300);
and U19172 (N_19172,N_12702,N_14723);
nand U19173 (N_19173,N_10353,N_11169);
nor U19174 (N_19174,N_14822,N_12225);
or U19175 (N_19175,N_14489,N_10325);
nand U19176 (N_19176,N_13067,N_11261);
xor U19177 (N_19177,N_11227,N_13547);
nand U19178 (N_19178,N_14648,N_11465);
xor U19179 (N_19179,N_14867,N_13323);
nand U19180 (N_19180,N_10894,N_13188);
xnor U19181 (N_19181,N_14638,N_13460);
xor U19182 (N_19182,N_11554,N_12383);
nand U19183 (N_19183,N_10695,N_11202);
nand U19184 (N_19184,N_12021,N_12824);
or U19185 (N_19185,N_11867,N_10022);
nor U19186 (N_19186,N_13237,N_10862);
and U19187 (N_19187,N_14343,N_11479);
or U19188 (N_19188,N_13277,N_12603);
or U19189 (N_19189,N_11705,N_12816);
and U19190 (N_19190,N_12744,N_11886);
or U19191 (N_19191,N_10059,N_14390);
or U19192 (N_19192,N_10764,N_10005);
nor U19193 (N_19193,N_14027,N_13484);
xnor U19194 (N_19194,N_13406,N_10992);
nor U19195 (N_19195,N_14330,N_14864);
nor U19196 (N_19196,N_12710,N_11332);
xor U19197 (N_19197,N_11110,N_13260);
and U19198 (N_19198,N_14844,N_12648);
xnor U19199 (N_19199,N_12597,N_11137);
nand U19200 (N_19200,N_10597,N_12125);
nand U19201 (N_19201,N_11958,N_10698);
or U19202 (N_19202,N_11615,N_13628);
or U19203 (N_19203,N_13192,N_13456);
or U19204 (N_19204,N_12270,N_13308);
nand U19205 (N_19205,N_13842,N_12041);
nand U19206 (N_19206,N_10732,N_13248);
nor U19207 (N_19207,N_12760,N_12238);
and U19208 (N_19208,N_11597,N_12783);
xor U19209 (N_19209,N_14226,N_11177);
xor U19210 (N_19210,N_14444,N_11666);
or U19211 (N_19211,N_10721,N_14259);
or U19212 (N_19212,N_10891,N_11137);
and U19213 (N_19213,N_11897,N_12444);
and U19214 (N_19214,N_11819,N_13590);
nand U19215 (N_19215,N_11513,N_12587);
nand U19216 (N_19216,N_10019,N_11827);
nor U19217 (N_19217,N_13513,N_12466);
nand U19218 (N_19218,N_14195,N_14518);
nor U19219 (N_19219,N_10614,N_10005);
or U19220 (N_19220,N_12293,N_11614);
nand U19221 (N_19221,N_14154,N_11527);
or U19222 (N_19222,N_14588,N_10608);
or U19223 (N_19223,N_10333,N_12795);
nor U19224 (N_19224,N_14250,N_11944);
nor U19225 (N_19225,N_13011,N_13206);
nand U19226 (N_19226,N_10271,N_13899);
and U19227 (N_19227,N_14401,N_10744);
or U19228 (N_19228,N_11783,N_10660);
and U19229 (N_19229,N_11702,N_10395);
nor U19230 (N_19230,N_10495,N_13757);
nor U19231 (N_19231,N_13224,N_10210);
and U19232 (N_19232,N_14764,N_13314);
nand U19233 (N_19233,N_10187,N_12916);
nand U19234 (N_19234,N_14955,N_10200);
and U19235 (N_19235,N_13914,N_10478);
xnor U19236 (N_19236,N_11574,N_11655);
and U19237 (N_19237,N_13196,N_11862);
nand U19238 (N_19238,N_13618,N_13398);
nand U19239 (N_19239,N_14797,N_13804);
xor U19240 (N_19240,N_10184,N_13393);
nor U19241 (N_19241,N_11610,N_13579);
nor U19242 (N_19242,N_14906,N_10580);
nor U19243 (N_19243,N_10142,N_12235);
and U19244 (N_19244,N_13968,N_10880);
or U19245 (N_19245,N_13994,N_12891);
nor U19246 (N_19246,N_14679,N_10460);
nor U19247 (N_19247,N_12399,N_13599);
or U19248 (N_19248,N_10688,N_13516);
nor U19249 (N_19249,N_12393,N_11075);
nand U19250 (N_19250,N_12324,N_14487);
or U19251 (N_19251,N_12160,N_12609);
and U19252 (N_19252,N_11742,N_12822);
xnor U19253 (N_19253,N_11053,N_11151);
or U19254 (N_19254,N_12720,N_10733);
xor U19255 (N_19255,N_13474,N_10863);
and U19256 (N_19256,N_11908,N_12218);
or U19257 (N_19257,N_13456,N_14401);
and U19258 (N_19258,N_14953,N_10790);
and U19259 (N_19259,N_14956,N_10043);
nand U19260 (N_19260,N_14697,N_12424);
or U19261 (N_19261,N_12803,N_13988);
nor U19262 (N_19262,N_14849,N_10896);
xnor U19263 (N_19263,N_13689,N_10746);
and U19264 (N_19264,N_10524,N_11307);
xor U19265 (N_19265,N_14168,N_10709);
or U19266 (N_19266,N_12721,N_14410);
xnor U19267 (N_19267,N_13803,N_13904);
nand U19268 (N_19268,N_14824,N_10888);
xnor U19269 (N_19269,N_12896,N_12361);
nor U19270 (N_19270,N_13700,N_11764);
xor U19271 (N_19271,N_11011,N_11494);
xnor U19272 (N_19272,N_12999,N_10240);
and U19273 (N_19273,N_14037,N_11734);
or U19274 (N_19274,N_10520,N_10296);
nand U19275 (N_19275,N_13441,N_13817);
and U19276 (N_19276,N_14002,N_11743);
nor U19277 (N_19277,N_12637,N_13315);
nand U19278 (N_19278,N_13203,N_13182);
xnor U19279 (N_19279,N_13338,N_14551);
or U19280 (N_19280,N_14022,N_12683);
and U19281 (N_19281,N_10589,N_12068);
nor U19282 (N_19282,N_13926,N_10235);
nor U19283 (N_19283,N_12876,N_13121);
and U19284 (N_19284,N_11563,N_11566);
or U19285 (N_19285,N_12005,N_14971);
xor U19286 (N_19286,N_13814,N_14325);
nand U19287 (N_19287,N_14475,N_12350);
or U19288 (N_19288,N_14425,N_11298);
and U19289 (N_19289,N_12394,N_13785);
or U19290 (N_19290,N_11629,N_10971);
and U19291 (N_19291,N_12127,N_14467);
nor U19292 (N_19292,N_12567,N_10783);
nand U19293 (N_19293,N_12945,N_13490);
xor U19294 (N_19294,N_10054,N_10181);
and U19295 (N_19295,N_13648,N_14524);
or U19296 (N_19296,N_14474,N_13906);
nand U19297 (N_19297,N_13851,N_11027);
xnor U19298 (N_19298,N_12608,N_13324);
or U19299 (N_19299,N_14939,N_14528);
xor U19300 (N_19300,N_13238,N_11218);
nand U19301 (N_19301,N_14037,N_12991);
nand U19302 (N_19302,N_10660,N_14471);
nand U19303 (N_19303,N_14302,N_14885);
and U19304 (N_19304,N_14613,N_11972);
and U19305 (N_19305,N_10875,N_13130);
and U19306 (N_19306,N_11374,N_12683);
nor U19307 (N_19307,N_14643,N_12949);
nor U19308 (N_19308,N_13513,N_12066);
nand U19309 (N_19309,N_14169,N_14660);
and U19310 (N_19310,N_14125,N_13856);
xnor U19311 (N_19311,N_14704,N_11623);
or U19312 (N_19312,N_11486,N_14473);
or U19313 (N_19313,N_10616,N_14790);
and U19314 (N_19314,N_12645,N_12565);
nand U19315 (N_19315,N_13512,N_11243);
nand U19316 (N_19316,N_12459,N_13476);
or U19317 (N_19317,N_14488,N_12894);
nor U19318 (N_19318,N_10735,N_14920);
xnor U19319 (N_19319,N_13936,N_13149);
nor U19320 (N_19320,N_13425,N_14038);
xor U19321 (N_19321,N_13191,N_11317);
or U19322 (N_19322,N_14530,N_11157);
nor U19323 (N_19323,N_13011,N_14078);
xnor U19324 (N_19324,N_13692,N_11543);
nand U19325 (N_19325,N_11716,N_12328);
or U19326 (N_19326,N_13393,N_12942);
nand U19327 (N_19327,N_13133,N_10283);
nor U19328 (N_19328,N_13959,N_13000);
or U19329 (N_19329,N_10818,N_13528);
nand U19330 (N_19330,N_13562,N_11934);
nand U19331 (N_19331,N_13715,N_14987);
and U19332 (N_19332,N_11964,N_14575);
and U19333 (N_19333,N_12686,N_10671);
nor U19334 (N_19334,N_12713,N_13424);
nand U19335 (N_19335,N_10707,N_11473);
or U19336 (N_19336,N_13357,N_10116);
or U19337 (N_19337,N_13876,N_14012);
xnor U19338 (N_19338,N_10086,N_12266);
and U19339 (N_19339,N_11309,N_10204);
nand U19340 (N_19340,N_11974,N_12694);
and U19341 (N_19341,N_10035,N_13893);
nor U19342 (N_19342,N_12736,N_14799);
nand U19343 (N_19343,N_13699,N_13049);
nand U19344 (N_19344,N_11805,N_13817);
nand U19345 (N_19345,N_13693,N_10748);
xor U19346 (N_19346,N_12104,N_13505);
or U19347 (N_19347,N_10696,N_13391);
xor U19348 (N_19348,N_12133,N_12638);
and U19349 (N_19349,N_12511,N_11069);
nor U19350 (N_19350,N_11346,N_10407);
or U19351 (N_19351,N_10003,N_13824);
nand U19352 (N_19352,N_14204,N_10354);
nor U19353 (N_19353,N_14931,N_11307);
and U19354 (N_19354,N_10138,N_14152);
nand U19355 (N_19355,N_13696,N_12962);
nand U19356 (N_19356,N_10669,N_12570);
xor U19357 (N_19357,N_13653,N_14159);
and U19358 (N_19358,N_14848,N_14223);
nand U19359 (N_19359,N_13326,N_13889);
xnor U19360 (N_19360,N_13761,N_14499);
nor U19361 (N_19361,N_12221,N_13944);
xor U19362 (N_19362,N_13302,N_14847);
nand U19363 (N_19363,N_12164,N_13998);
or U19364 (N_19364,N_10394,N_13147);
or U19365 (N_19365,N_14688,N_12749);
xnor U19366 (N_19366,N_12555,N_11543);
nor U19367 (N_19367,N_12474,N_12028);
xor U19368 (N_19368,N_14371,N_12529);
xor U19369 (N_19369,N_10121,N_10050);
or U19370 (N_19370,N_12328,N_13057);
nor U19371 (N_19371,N_11244,N_14760);
nor U19372 (N_19372,N_10621,N_11028);
or U19373 (N_19373,N_14648,N_10855);
or U19374 (N_19374,N_11378,N_10105);
xor U19375 (N_19375,N_12717,N_13039);
or U19376 (N_19376,N_11505,N_13394);
xnor U19377 (N_19377,N_11878,N_12992);
and U19378 (N_19378,N_11034,N_13291);
or U19379 (N_19379,N_12087,N_13115);
xor U19380 (N_19380,N_14412,N_12945);
and U19381 (N_19381,N_11045,N_11101);
nand U19382 (N_19382,N_13545,N_12158);
xor U19383 (N_19383,N_13085,N_10765);
or U19384 (N_19384,N_11444,N_14475);
nand U19385 (N_19385,N_12126,N_12276);
nand U19386 (N_19386,N_13058,N_14634);
nand U19387 (N_19387,N_13615,N_13286);
xor U19388 (N_19388,N_14613,N_14201);
nand U19389 (N_19389,N_14199,N_14477);
or U19390 (N_19390,N_13994,N_13712);
nor U19391 (N_19391,N_14824,N_11124);
nand U19392 (N_19392,N_11216,N_12716);
and U19393 (N_19393,N_14095,N_13406);
xnor U19394 (N_19394,N_14484,N_11330);
or U19395 (N_19395,N_14715,N_13145);
or U19396 (N_19396,N_11460,N_12887);
nor U19397 (N_19397,N_10201,N_12322);
or U19398 (N_19398,N_13874,N_10945);
xnor U19399 (N_19399,N_10079,N_13424);
and U19400 (N_19400,N_13690,N_11626);
xnor U19401 (N_19401,N_10614,N_14710);
or U19402 (N_19402,N_13861,N_14820);
or U19403 (N_19403,N_12095,N_10034);
nor U19404 (N_19404,N_10395,N_12437);
xnor U19405 (N_19405,N_14433,N_11893);
and U19406 (N_19406,N_11811,N_10204);
and U19407 (N_19407,N_10062,N_10855);
and U19408 (N_19408,N_10729,N_14080);
xor U19409 (N_19409,N_11107,N_11320);
or U19410 (N_19410,N_14589,N_10844);
or U19411 (N_19411,N_10171,N_10229);
xnor U19412 (N_19412,N_14509,N_13108);
nand U19413 (N_19413,N_11082,N_13886);
nand U19414 (N_19414,N_10720,N_11661);
nand U19415 (N_19415,N_12117,N_12723);
and U19416 (N_19416,N_12757,N_11177);
nor U19417 (N_19417,N_14179,N_14912);
and U19418 (N_19418,N_12376,N_11383);
nor U19419 (N_19419,N_14971,N_10098);
nor U19420 (N_19420,N_10004,N_10863);
nor U19421 (N_19421,N_13159,N_14797);
and U19422 (N_19422,N_11366,N_11641);
or U19423 (N_19423,N_11653,N_11224);
and U19424 (N_19424,N_11760,N_12655);
nand U19425 (N_19425,N_14137,N_14660);
xor U19426 (N_19426,N_12092,N_12406);
and U19427 (N_19427,N_12887,N_13693);
or U19428 (N_19428,N_13102,N_13159);
or U19429 (N_19429,N_10503,N_14405);
nand U19430 (N_19430,N_11431,N_13263);
nor U19431 (N_19431,N_12930,N_14619);
or U19432 (N_19432,N_14583,N_12427);
xnor U19433 (N_19433,N_14104,N_11192);
or U19434 (N_19434,N_12755,N_11176);
nand U19435 (N_19435,N_12081,N_10980);
nor U19436 (N_19436,N_10408,N_10096);
xor U19437 (N_19437,N_12164,N_11244);
nand U19438 (N_19438,N_13199,N_13406);
nand U19439 (N_19439,N_14231,N_11639);
and U19440 (N_19440,N_14630,N_13025);
and U19441 (N_19441,N_12238,N_14195);
and U19442 (N_19442,N_10714,N_11053);
or U19443 (N_19443,N_10667,N_12356);
xnor U19444 (N_19444,N_12877,N_14456);
nor U19445 (N_19445,N_12451,N_10687);
xnor U19446 (N_19446,N_14877,N_12205);
nand U19447 (N_19447,N_11596,N_12374);
nor U19448 (N_19448,N_11746,N_14621);
or U19449 (N_19449,N_12660,N_12312);
xnor U19450 (N_19450,N_11679,N_12270);
nor U19451 (N_19451,N_14716,N_12178);
nor U19452 (N_19452,N_11398,N_12051);
nor U19453 (N_19453,N_11286,N_11646);
xor U19454 (N_19454,N_14139,N_12848);
and U19455 (N_19455,N_11143,N_13101);
xnor U19456 (N_19456,N_12432,N_10644);
xor U19457 (N_19457,N_10103,N_12485);
or U19458 (N_19458,N_14668,N_10663);
or U19459 (N_19459,N_14913,N_14421);
or U19460 (N_19460,N_11984,N_11417);
nor U19461 (N_19461,N_10152,N_10789);
nor U19462 (N_19462,N_10546,N_10400);
nand U19463 (N_19463,N_10166,N_11810);
and U19464 (N_19464,N_13682,N_12380);
or U19465 (N_19465,N_10482,N_11624);
or U19466 (N_19466,N_12895,N_13062);
and U19467 (N_19467,N_11013,N_13492);
or U19468 (N_19468,N_10937,N_13574);
nand U19469 (N_19469,N_14986,N_11115);
xor U19470 (N_19470,N_12287,N_14413);
xnor U19471 (N_19471,N_11326,N_12402);
nor U19472 (N_19472,N_13441,N_12480);
xor U19473 (N_19473,N_10806,N_13646);
nand U19474 (N_19474,N_10824,N_11821);
or U19475 (N_19475,N_11960,N_13902);
nor U19476 (N_19476,N_12326,N_13391);
or U19477 (N_19477,N_11481,N_12404);
nor U19478 (N_19478,N_12869,N_10640);
xor U19479 (N_19479,N_14843,N_10502);
and U19480 (N_19480,N_11892,N_11669);
nand U19481 (N_19481,N_13705,N_13669);
nor U19482 (N_19482,N_13960,N_13780);
or U19483 (N_19483,N_12200,N_11858);
nand U19484 (N_19484,N_11971,N_10604);
nand U19485 (N_19485,N_13424,N_14137);
xor U19486 (N_19486,N_11568,N_14215);
xnor U19487 (N_19487,N_11507,N_14146);
and U19488 (N_19488,N_13959,N_13666);
nand U19489 (N_19489,N_13802,N_12560);
nor U19490 (N_19490,N_11975,N_11150);
and U19491 (N_19491,N_11475,N_12900);
and U19492 (N_19492,N_11941,N_14488);
nand U19493 (N_19493,N_13171,N_14074);
nor U19494 (N_19494,N_10795,N_10748);
nor U19495 (N_19495,N_10929,N_14595);
nand U19496 (N_19496,N_13529,N_14970);
nand U19497 (N_19497,N_10035,N_11058);
nor U19498 (N_19498,N_13251,N_14112);
and U19499 (N_19499,N_13472,N_10259);
xor U19500 (N_19500,N_12446,N_12506);
xnor U19501 (N_19501,N_13625,N_14470);
nor U19502 (N_19502,N_12392,N_14516);
xnor U19503 (N_19503,N_10035,N_13353);
and U19504 (N_19504,N_12448,N_10174);
and U19505 (N_19505,N_12078,N_11368);
or U19506 (N_19506,N_14716,N_13251);
nand U19507 (N_19507,N_14451,N_14947);
nand U19508 (N_19508,N_13024,N_11593);
and U19509 (N_19509,N_14512,N_14499);
and U19510 (N_19510,N_10532,N_12227);
nor U19511 (N_19511,N_11211,N_12092);
and U19512 (N_19512,N_10729,N_14243);
nand U19513 (N_19513,N_14452,N_10325);
nand U19514 (N_19514,N_13127,N_10481);
and U19515 (N_19515,N_14791,N_13830);
or U19516 (N_19516,N_12728,N_14124);
and U19517 (N_19517,N_12216,N_13448);
nand U19518 (N_19518,N_13198,N_12973);
xnor U19519 (N_19519,N_10324,N_11747);
nor U19520 (N_19520,N_10498,N_14611);
nand U19521 (N_19521,N_13140,N_14598);
nand U19522 (N_19522,N_10321,N_12732);
nor U19523 (N_19523,N_12159,N_12544);
or U19524 (N_19524,N_13867,N_10190);
nor U19525 (N_19525,N_11320,N_11195);
or U19526 (N_19526,N_14898,N_11588);
xor U19527 (N_19527,N_14959,N_10430);
nand U19528 (N_19528,N_10055,N_11050);
and U19529 (N_19529,N_14809,N_12089);
nor U19530 (N_19530,N_13831,N_11623);
and U19531 (N_19531,N_11801,N_10069);
and U19532 (N_19532,N_13133,N_11024);
nor U19533 (N_19533,N_14209,N_12142);
and U19534 (N_19534,N_12853,N_11290);
nand U19535 (N_19535,N_14131,N_10089);
or U19536 (N_19536,N_13592,N_12179);
xnor U19537 (N_19537,N_10732,N_14543);
or U19538 (N_19538,N_10872,N_11978);
or U19539 (N_19539,N_11459,N_13717);
or U19540 (N_19540,N_10853,N_11491);
and U19541 (N_19541,N_11694,N_12389);
nand U19542 (N_19542,N_13225,N_14544);
nor U19543 (N_19543,N_11427,N_13680);
and U19544 (N_19544,N_12832,N_14352);
and U19545 (N_19545,N_12355,N_10750);
xnor U19546 (N_19546,N_12503,N_10269);
nand U19547 (N_19547,N_12143,N_11798);
or U19548 (N_19548,N_14825,N_12054);
and U19549 (N_19549,N_13581,N_13912);
nor U19550 (N_19550,N_14141,N_10761);
and U19551 (N_19551,N_11267,N_14602);
or U19552 (N_19552,N_11229,N_12042);
nor U19553 (N_19553,N_14133,N_14661);
nand U19554 (N_19554,N_14050,N_10250);
and U19555 (N_19555,N_14695,N_13281);
and U19556 (N_19556,N_12985,N_11334);
nand U19557 (N_19557,N_12161,N_10958);
or U19558 (N_19558,N_14873,N_11500);
nand U19559 (N_19559,N_14938,N_10458);
nand U19560 (N_19560,N_11024,N_11534);
nor U19561 (N_19561,N_11129,N_14821);
xor U19562 (N_19562,N_12858,N_13723);
xnor U19563 (N_19563,N_10185,N_14531);
or U19564 (N_19564,N_10732,N_11926);
nand U19565 (N_19565,N_11567,N_11673);
nand U19566 (N_19566,N_10839,N_13199);
nor U19567 (N_19567,N_10549,N_10428);
xor U19568 (N_19568,N_11953,N_11227);
nor U19569 (N_19569,N_10085,N_14390);
xnor U19570 (N_19570,N_11461,N_11384);
xor U19571 (N_19571,N_14400,N_11766);
xor U19572 (N_19572,N_11817,N_13715);
and U19573 (N_19573,N_14057,N_10548);
and U19574 (N_19574,N_14986,N_12540);
xnor U19575 (N_19575,N_11102,N_11062);
nor U19576 (N_19576,N_12520,N_14234);
nor U19577 (N_19577,N_11411,N_12560);
nor U19578 (N_19578,N_12743,N_12713);
nor U19579 (N_19579,N_12164,N_12390);
or U19580 (N_19580,N_12470,N_11463);
nand U19581 (N_19581,N_14188,N_10344);
nor U19582 (N_19582,N_11005,N_11944);
and U19583 (N_19583,N_12612,N_11465);
and U19584 (N_19584,N_13363,N_10430);
or U19585 (N_19585,N_14556,N_10114);
and U19586 (N_19586,N_12966,N_10024);
xnor U19587 (N_19587,N_12037,N_12435);
or U19588 (N_19588,N_13034,N_13636);
nand U19589 (N_19589,N_11098,N_12652);
xnor U19590 (N_19590,N_14044,N_13173);
or U19591 (N_19591,N_11775,N_11842);
or U19592 (N_19592,N_11089,N_10496);
xnor U19593 (N_19593,N_11689,N_14449);
nand U19594 (N_19594,N_14964,N_14233);
and U19595 (N_19595,N_11773,N_10823);
xor U19596 (N_19596,N_13370,N_10736);
nor U19597 (N_19597,N_11939,N_12112);
or U19598 (N_19598,N_12834,N_10690);
nor U19599 (N_19599,N_11367,N_13080);
or U19600 (N_19600,N_13200,N_12578);
or U19601 (N_19601,N_10756,N_13612);
or U19602 (N_19602,N_14760,N_14568);
or U19603 (N_19603,N_12172,N_10757);
nor U19604 (N_19604,N_11164,N_13566);
nor U19605 (N_19605,N_14660,N_14202);
nand U19606 (N_19606,N_12639,N_12417);
xnor U19607 (N_19607,N_13335,N_10257);
and U19608 (N_19608,N_10832,N_14318);
nor U19609 (N_19609,N_11600,N_12695);
nor U19610 (N_19610,N_12747,N_10757);
and U19611 (N_19611,N_13201,N_11909);
xor U19612 (N_19612,N_11809,N_14276);
nor U19613 (N_19613,N_14951,N_13122);
xnor U19614 (N_19614,N_11280,N_13209);
and U19615 (N_19615,N_14942,N_14927);
or U19616 (N_19616,N_12206,N_10499);
or U19617 (N_19617,N_11499,N_12779);
nor U19618 (N_19618,N_12908,N_14274);
xnor U19619 (N_19619,N_12377,N_12062);
or U19620 (N_19620,N_11784,N_10017);
nand U19621 (N_19621,N_10934,N_14321);
nand U19622 (N_19622,N_12207,N_11828);
nor U19623 (N_19623,N_14887,N_14120);
xor U19624 (N_19624,N_13335,N_14758);
and U19625 (N_19625,N_13980,N_11543);
or U19626 (N_19626,N_12603,N_12040);
nand U19627 (N_19627,N_14093,N_11980);
xor U19628 (N_19628,N_12086,N_10556);
and U19629 (N_19629,N_10364,N_14474);
and U19630 (N_19630,N_13741,N_12836);
and U19631 (N_19631,N_10475,N_12001);
or U19632 (N_19632,N_11290,N_10278);
xnor U19633 (N_19633,N_11280,N_13288);
or U19634 (N_19634,N_11018,N_14695);
nor U19635 (N_19635,N_12011,N_12827);
nor U19636 (N_19636,N_13926,N_14422);
nand U19637 (N_19637,N_10976,N_10294);
nand U19638 (N_19638,N_13818,N_12660);
nor U19639 (N_19639,N_12384,N_10785);
or U19640 (N_19640,N_13266,N_13386);
xor U19641 (N_19641,N_14290,N_14195);
nor U19642 (N_19642,N_14386,N_13688);
and U19643 (N_19643,N_10971,N_10964);
nor U19644 (N_19644,N_13422,N_10872);
nor U19645 (N_19645,N_13165,N_11041);
nand U19646 (N_19646,N_11395,N_10726);
nand U19647 (N_19647,N_12627,N_12372);
nand U19648 (N_19648,N_13073,N_11956);
xnor U19649 (N_19649,N_10065,N_13958);
and U19650 (N_19650,N_10481,N_10535);
nand U19651 (N_19651,N_14400,N_10299);
nand U19652 (N_19652,N_12851,N_10499);
nand U19653 (N_19653,N_13459,N_11656);
nand U19654 (N_19654,N_10670,N_11231);
nand U19655 (N_19655,N_10076,N_13017);
xnor U19656 (N_19656,N_13057,N_14127);
or U19657 (N_19657,N_13355,N_13832);
xnor U19658 (N_19658,N_12805,N_13244);
xor U19659 (N_19659,N_11396,N_10376);
or U19660 (N_19660,N_10246,N_12689);
nor U19661 (N_19661,N_10147,N_14074);
and U19662 (N_19662,N_13058,N_10530);
or U19663 (N_19663,N_13410,N_13467);
nor U19664 (N_19664,N_13144,N_12943);
and U19665 (N_19665,N_12917,N_14994);
or U19666 (N_19666,N_10513,N_12926);
xnor U19667 (N_19667,N_13265,N_13678);
or U19668 (N_19668,N_14418,N_13091);
and U19669 (N_19669,N_11420,N_12991);
nor U19670 (N_19670,N_14844,N_12294);
xor U19671 (N_19671,N_12420,N_10419);
or U19672 (N_19672,N_11321,N_13783);
nor U19673 (N_19673,N_12681,N_12832);
or U19674 (N_19674,N_13723,N_14405);
nor U19675 (N_19675,N_10875,N_14711);
nand U19676 (N_19676,N_13283,N_11078);
nand U19677 (N_19677,N_14253,N_10390);
and U19678 (N_19678,N_14845,N_13418);
or U19679 (N_19679,N_12980,N_12866);
nand U19680 (N_19680,N_10173,N_11686);
nor U19681 (N_19681,N_10816,N_11286);
nand U19682 (N_19682,N_12822,N_14903);
xnor U19683 (N_19683,N_14246,N_11137);
and U19684 (N_19684,N_14348,N_11175);
nand U19685 (N_19685,N_11029,N_13477);
nor U19686 (N_19686,N_12934,N_11312);
xor U19687 (N_19687,N_14470,N_12495);
nand U19688 (N_19688,N_10330,N_11707);
xnor U19689 (N_19689,N_14618,N_13083);
xnor U19690 (N_19690,N_11474,N_10730);
xor U19691 (N_19691,N_11281,N_13982);
and U19692 (N_19692,N_12253,N_11366);
or U19693 (N_19693,N_13223,N_14681);
and U19694 (N_19694,N_10739,N_14629);
and U19695 (N_19695,N_11488,N_10148);
nand U19696 (N_19696,N_11263,N_10856);
nand U19697 (N_19697,N_10745,N_11901);
nor U19698 (N_19698,N_11337,N_13169);
nor U19699 (N_19699,N_10127,N_14064);
and U19700 (N_19700,N_10797,N_14106);
nand U19701 (N_19701,N_12747,N_13360);
or U19702 (N_19702,N_13339,N_11492);
nand U19703 (N_19703,N_13878,N_10813);
and U19704 (N_19704,N_11243,N_10111);
and U19705 (N_19705,N_14360,N_14328);
nand U19706 (N_19706,N_12458,N_14433);
and U19707 (N_19707,N_11366,N_10394);
or U19708 (N_19708,N_14117,N_14481);
nor U19709 (N_19709,N_10679,N_10979);
nor U19710 (N_19710,N_14216,N_14020);
and U19711 (N_19711,N_14642,N_13931);
nor U19712 (N_19712,N_12757,N_13128);
nand U19713 (N_19713,N_10426,N_10918);
or U19714 (N_19714,N_11746,N_11883);
nor U19715 (N_19715,N_12195,N_14799);
or U19716 (N_19716,N_11677,N_12603);
nor U19717 (N_19717,N_10985,N_11570);
xnor U19718 (N_19718,N_10145,N_13766);
xnor U19719 (N_19719,N_10456,N_12419);
nand U19720 (N_19720,N_13974,N_12667);
or U19721 (N_19721,N_11918,N_10686);
nor U19722 (N_19722,N_10339,N_11527);
xor U19723 (N_19723,N_10493,N_13041);
and U19724 (N_19724,N_10592,N_11408);
or U19725 (N_19725,N_13087,N_11058);
or U19726 (N_19726,N_10226,N_11793);
or U19727 (N_19727,N_10692,N_13450);
nor U19728 (N_19728,N_12187,N_14290);
and U19729 (N_19729,N_10672,N_12529);
or U19730 (N_19730,N_11063,N_11028);
or U19731 (N_19731,N_12917,N_12832);
or U19732 (N_19732,N_14651,N_10796);
and U19733 (N_19733,N_13791,N_12920);
or U19734 (N_19734,N_13787,N_13585);
or U19735 (N_19735,N_14688,N_10021);
nand U19736 (N_19736,N_10781,N_13821);
xnor U19737 (N_19737,N_13644,N_14653);
nand U19738 (N_19738,N_12160,N_12161);
or U19739 (N_19739,N_10751,N_13439);
nor U19740 (N_19740,N_10766,N_14285);
or U19741 (N_19741,N_13446,N_11137);
and U19742 (N_19742,N_10528,N_14509);
nand U19743 (N_19743,N_10682,N_14044);
xor U19744 (N_19744,N_14889,N_10560);
or U19745 (N_19745,N_12973,N_13227);
and U19746 (N_19746,N_12648,N_14476);
or U19747 (N_19747,N_14640,N_14312);
and U19748 (N_19748,N_10979,N_11984);
xnor U19749 (N_19749,N_13294,N_10937);
nor U19750 (N_19750,N_14509,N_14898);
nor U19751 (N_19751,N_10267,N_12424);
nand U19752 (N_19752,N_11224,N_13047);
xnor U19753 (N_19753,N_13307,N_13039);
nor U19754 (N_19754,N_11611,N_11944);
and U19755 (N_19755,N_11753,N_10021);
and U19756 (N_19756,N_12710,N_10582);
nor U19757 (N_19757,N_12210,N_12068);
and U19758 (N_19758,N_11875,N_12348);
xor U19759 (N_19759,N_12386,N_13348);
xnor U19760 (N_19760,N_13875,N_14690);
or U19761 (N_19761,N_11243,N_14888);
and U19762 (N_19762,N_10421,N_11580);
or U19763 (N_19763,N_10071,N_13515);
or U19764 (N_19764,N_12696,N_13496);
nor U19765 (N_19765,N_11279,N_12975);
or U19766 (N_19766,N_12975,N_10943);
nand U19767 (N_19767,N_13815,N_14196);
and U19768 (N_19768,N_10076,N_12103);
nor U19769 (N_19769,N_14079,N_11831);
nor U19770 (N_19770,N_12469,N_10037);
nor U19771 (N_19771,N_13707,N_11704);
xnor U19772 (N_19772,N_12734,N_14416);
xor U19773 (N_19773,N_10159,N_13663);
nand U19774 (N_19774,N_10896,N_10387);
xnor U19775 (N_19775,N_14569,N_14241);
or U19776 (N_19776,N_12812,N_10114);
nor U19777 (N_19777,N_12110,N_14844);
xnor U19778 (N_19778,N_11213,N_10846);
or U19779 (N_19779,N_12671,N_11590);
or U19780 (N_19780,N_10245,N_10049);
and U19781 (N_19781,N_13967,N_13831);
xnor U19782 (N_19782,N_10888,N_13148);
nand U19783 (N_19783,N_10657,N_12992);
or U19784 (N_19784,N_12070,N_14659);
xor U19785 (N_19785,N_11052,N_11814);
nor U19786 (N_19786,N_13131,N_10942);
nor U19787 (N_19787,N_12246,N_14737);
or U19788 (N_19788,N_14508,N_14665);
nor U19789 (N_19789,N_14313,N_11350);
nor U19790 (N_19790,N_13269,N_14437);
and U19791 (N_19791,N_11870,N_11254);
nand U19792 (N_19792,N_12080,N_14506);
xor U19793 (N_19793,N_10569,N_14779);
or U19794 (N_19794,N_13551,N_11365);
nor U19795 (N_19795,N_10259,N_12557);
xnor U19796 (N_19796,N_10827,N_12674);
or U19797 (N_19797,N_14865,N_13016);
nor U19798 (N_19798,N_14566,N_11906);
and U19799 (N_19799,N_11433,N_10500);
nand U19800 (N_19800,N_13201,N_11304);
nand U19801 (N_19801,N_11208,N_10171);
nor U19802 (N_19802,N_13612,N_13192);
or U19803 (N_19803,N_10066,N_13161);
xnor U19804 (N_19804,N_12274,N_10691);
and U19805 (N_19805,N_11957,N_11187);
nor U19806 (N_19806,N_14653,N_10675);
nor U19807 (N_19807,N_13929,N_10575);
xor U19808 (N_19808,N_13956,N_13937);
or U19809 (N_19809,N_14380,N_12323);
nand U19810 (N_19810,N_13901,N_13343);
or U19811 (N_19811,N_12692,N_11845);
or U19812 (N_19812,N_10642,N_13399);
nand U19813 (N_19813,N_12084,N_12351);
or U19814 (N_19814,N_10145,N_14479);
xor U19815 (N_19815,N_10270,N_10718);
nand U19816 (N_19816,N_13005,N_11225);
nand U19817 (N_19817,N_12276,N_13829);
nor U19818 (N_19818,N_12205,N_14569);
nand U19819 (N_19819,N_12263,N_11590);
xor U19820 (N_19820,N_12132,N_14638);
nor U19821 (N_19821,N_13696,N_12246);
xnor U19822 (N_19822,N_11105,N_11736);
and U19823 (N_19823,N_13270,N_10469);
nor U19824 (N_19824,N_11992,N_10673);
nor U19825 (N_19825,N_12240,N_14807);
or U19826 (N_19826,N_10587,N_13460);
xor U19827 (N_19827,N_10222,N_13023);
nor U19828 (N_19828,N_13416,N_11509);
and U19829 (N_19829,N_13831,N_13738);
xor U19830 (N_19830,N_14632,N_12921);
nand U19831 (N_19831,N_14315,N_10400);
or U19832 (N_19832,N_13491,N_12982);
and U19833 (N_19833,N_14857,N_13273);
nand U19834 (N_19834,N_12207,N_13676);
nand U19835 (N_19835,N_14377,N_11063);
and U19836 (N_19836,N_12791,N_13083);
and U19837 (N_19837,N_10051,N_12523);
nor U19838 (N_19838,N_13178,N_14066);
nor U19839 (N_19839,N_14726,N_11000);
xor U19840 (N_19840,N_13379,N_11375);
nor U19841 (N_19841,N_13590,N_14412);
xor U19842 (N_19842,N_11462,N_10388);
nor U19843 (N_19843,N_12278,N_14721);
and U19844 (N_19844,N_10490,N_13474);
nand U19845 (N_19845,N_13084,N_12771);
or U19846 (N_19846,N_13726,N_11656);
nand U19847 (N_19847,N_10352,N_11189);
or U19848 (N_19848,N_14583,N_11231);
nor U19849 (N_19849,N_10716,N_14692);
or U19850 (N_19850,N_12929,N_10550);
nand U19851 (N_19851,N_14826,N_11336);
or U19852 (N_19852,N_13643,N_14075);
nand U19853 (N_19853,N_13536,N_13932);
and U19854 (N_19854,N_11004,N_10925);
xnor U19855 (N_19855,N_10995,N_14760);
or U19856 (N_19856,N_10915,N_14844);
nor U19857 (N_19857,N_12066,N_11532);
or U19858 (N_19858,N_11417,N_13219);
and U19859 (N_19859,N_12653,N_11484);
and U19860 (N_19860,N_14108,N_14215);
xor U19861 (N_19861,N_12275,N_10822);
nor U19862 (N_19862,N_13952,N_11933);
and U19863 (N_19863,N_11324,N_11846);
xor U19864 (N_19864,N_14931,N_13637);
xor U19865 (N_19865,N_10509,N_10957);
and U19866 (N_19866,N_13606,N_14846);
xor U19867 (N_19867,N_13368,N_11994);
nand U19868 (N_19868,N_14972,N_13002);
and U19869 (N_19869,N_10760,N_13729);
nor U19870 (N_19870,N_12437,N_13803);
nor U19871 (N_19871,N_10920,N_13984);
xor U19872 (N_19872,N_12934,N_14393);
or U19873 (N_19873,N_14750,N_14906);
xor U19874 (N_19874,N_14207,N_10082);
and U19875 (N_19875,N_11059,N_14282);
or U19876 (N_19876,N_11693,N_14505);
and U19877 (N_19877,N_13752,N_10956);
or U19878 (N_19878,N_12093,N_11121);
xor U19879 (N_19879,N_11225,N_12589);
or U19880 (N_19880,N_10246,N_10104);
nand U19881 (N_19881,N_10800,N_10400);
and U19882 (N_19882,N_10336,N_10410);
xor U19883 (N_19883,N_11364,N_13310);
and U19884 (N_19884,N_10011,N_12609);
nor U19885 (N_19885,N_13303,N_10836);
and U19886 (N_19886,N_14828,N_12728);
or U19887 (N_19887,N_14077,N_14738);
nand U19888 (N_19888,N_11279,N_12184);
or U19889 (N_19889,N_14774,N_14824);
nand U19890 (N_19890,N_14091,N_10121);
and U19891 (N_19891,N_10718,N_14062);
or U19892 (N_19892,N_10403,N_14696);
nor U19893 (N_19893,N_10323,N_12247);
and U19894 (N_19894,N_12192,N_11097);
xnor U19895 (N_19895,N_11267,N_10699);
and U19896 (N_19896,N_12170,N_13131);
and U19897 (N_19897,N_13412,N_11106);
or U19898 (N_19898,N_10979,N_10772);
and U19899 (N_19899,N_11512,N_13398);
and U19900 (N_19900,N_11693,N_14634);
nor U19901 (N_19901,N_11508,N_10799);
xor U19902 (N_19902,N_12367,N_14264);
nand U19903 (N_19903,N_13913,N_10195);
nand U19904 (N_19904,N_14901,N_14297);
nand U19905 (N_19905,N_10640,N_12304);
and U19906 (N_19906,N_14998,N_11718);
xnor U19907 (N_19907,N_11129,N_11469);
nand U19908 (N_19908,N_10234,N_13608);
or U19909 (N_19909,N_11456,N_11726);
or U19910 (N_19910,N_11966,N_13841);
nor U19911 (N_19911,N_14129,N_13576);
xor U19912 (N_19912,N_14760,N_13918);
nand U19913 (N_19913,N_14914,N_11691);
nand U19914 (N_19914,N_11797,N_14087);
or U19915 (N_19915,N_14580,N_10596);
nor U19916 (N_19916,N_13066,N_10188);
or U19917 (N_19917,N_10818,N_13556);
nor U19918 (N_19918,N_12761,N_10543);
nand U19919 (N_19919,N_13339,N_10623);
xor U19920 (N_19920,N_14538,N_14400);
and U19921 (N_19921,N_12489,N_14655);
and U19922 (N_19922,N_11118,N_10190);
nor U19923 (N_19923,N_12871,N_12632);
and U19924 (N_19924,N_10949,N_13004);
and U19925 (N_19925,N_12747,N_10221);
nor U19926 (N_19926,N_11299,N_12219);
or U19927 (N_19927,N_14124,N_13329);
or U19928 (N_19928,N_10861,N_11544);
and U19929 (N_19929,N_11058,N_10756);
and U19930 (N_19930,N_11519,N_13654);
xnor U19931 (N_19931,N_13047,N_10752);
nor U19932 (N_19932,N_12730,N_12629);
nor U19933 (N_19933,N_12425,N_14769);
xnor U19934 (N_19934,N_13858,N_12880);
and U19935 (N_19935,N_12569,N_13096);
nor U19936 (N_19936,N_11025,N_10816);
nand U19937 (N_19937,N_13357,N_12204);
nand U19938 (N_19938,N_14657,N_10419);
and U19939 (N_19939,N_11497,N_12708);
nor U19940 (N_19940,N_12622,N_13323);
nand U19941 (N_19941,N_14448,N_14993);
nand U19942 (N_19942,N_14686,N_12593);
xnor U19943 (N_19943,N_14237,N_14656);
and U19944 (N_19944,N_10249,N_11720);
nor U19945 (N_19945,N_12603,N_10716);
and U19946 (N_19946,N_11785,N_12994);
or U19947 (N_19947,N_13012,N_12026);
or U19948 (N_19948,N_13034,N_13082);
nand U19949 (N_19949,N_12354,N_13063);
or U19950 (N_19950,N_12507,N_10757);
and U19951 (N_19951,N_12207,N_14507);
or U19952 (N_19952,N_11837,N_13287);
xor U19953 (N_19953,N_10705,N_12186);
and U19954 (N_19954,N_13752,N_13717);
nand U19955 (N_19955,N_11492,N_13043);
and U19956 (N_19956,N_14358,N_12944);
nor U19957 (N_19957,N_14925,N_14904);
or U19958 (N_19958,N_14617,N_12063);
xor U19959 (N_19959,N_13592,N_13718);
nor U19960 (N_19960,N_14255,N_10475);
or U19961 (N_19961,N_14145,N_11240);
xnor U19962 (N_19962,N_14784,N_10719);
nor U19963 (N_19963,N_14554,N_14740);
nand U19964 (N_19964,N_14330,N_14257);
and U19965 (N_19965,N_11541,N_10044);
xor U19966 (N_19966,N_13071,N_13982);
xnor U19967 (N_19967,N_11287,N_11591);
or U19968 (N_19968,N_12938,N_14958);
or U19969 (N_19969,N_10906,N_12937);
nand U19970 (N_19970,N_14594,N_13452);
nor U19971 (N_19971,N_10327,N_14119);
xnor U19972 (N_19972,N_10589,N_12816);
nor U19973 (N_19973,N_14519,N_13305);
and U19974 (N_19974,N_10474,N_12033);
or U19975 (N_19975,N_12550,N_11863);
nor U19976 (N_19976,N_12458,N_12771);
nand U19977 (N_19977,N_14799,N_13455);
xnor U19978 (N_19978,N_14086,N_12444);
nor U19979 (N_19979,N_13747,N_11706);
and U19980 (N_19980,N_10072,N_11429);
xor U19981 (N_19981,N_10615,N_12387);
or U19982 (N_19982,N_12075,N_14530);
nand U19983 (N_19983,N_14090,N_11183);
nand U19984 (N_19984,N_10881,N_14959);
nand U19985 (N_19985,N_11390,N_14589);
nor U19986 (N_19986,N_13048,N_13437);
nand U19987 (N_19987,N_10636,N_12431);
or U19988 (N_19988,N_10262,N_12025);
nor U19989 (N_19989,N_12440,N_14252);
xnor U19990 (N_19990,N_13791,N_10465);
or U19991 (N_19991,N_11726,N_13815);
or U19992 (N_19992,N_14167,N_10498);
nand U19993 (N_19993,N_13371,N_13813);
and U19994 (N_19994,N_10381,N_14371);
xor U19995 (N_19995,N_11398,N_14424);
nand U19996 (N_19996,N_11221,N_11517);
or U19997 (N_19997,N_10218,N_14587);
and U19998 (N_19998,N_10988,N_13616);
nor U19999 (N_19999,N_12752,N_14826);
and U20000 (N_20000,N_17857,N_18777);
xor U20001 (N_20001,N_17038,N_15480);
and U20002 (N_20002,N_19225,N_18369);
nand U20003 (N_20003,N_19244,N_18375);
xnor U20004 (N_20004,N_18938,N_15910);
and U20005 (N_20005,N_15628,N_16950);
nand U20006 (N_20006,N_15732,N_17212);
xnor U20007 (N_20007,N_17607,N_18531);
and U20008 (N_20008,N_15265,N_18289);
xor U20009 (N_20009,N_15777,N_18579);
xor U20010 (N_20010,N_19195,N_19300);
xnor U20011 (N_20011,N_15414,N_19174);
xnor U20012 (N_20012,N_17064,N_16337);
nand U20013 (N_20013,N_17577,N_15392);
and U20014 (N_20014,N_15338,N_17154);
nand U20015 (N_20015,N_19950,N_19559);
and U20016 (N_20016,N_18167,N_19947);
xor U20017 (N_20017,N_15035,N_17364);
nand U20018 (N_20018,N_17337,N_19290);
and U20019 (N_20019,N_16104,N_19065);
or U20020 (N_20020,N_15409,N_17391);
or U20021 (N_20021,N_16647,N_18552);
nor U20022 (N_20022,N_17077,N_18488);
or U20023 (N_20023,N_18765,N_16288);
or U20024 (N_20024,N_15303,N_16149);
nand U20025 (N_20025,N_15433,N_15679);
or U20026 (N_20026,N_18239,N_17168);
nand U20027 (N_20027,N_19203,N_16001);
nand U20028 (N_20028,N_16776,N_19068);
nand U20029 (N_20029,N_19025,N_19308);
nand U20030 (N_20030,N_19094,N_15030);
xnor U20031 (N_20031,N_18386,N_17535);
nand U20032 (N_20032,N_18557,N_17494);
and U20033 (N_20033,N_16694,N_15872);
or U20034 (N_20034,N_19901,N_17061);
nand U20035 (N_20035,N_15370,N_17914);
and U20036 (N_20036,N_18370,N_15168);
xnor U20037 (N_20037,N_15192,N_15682);
and U20038 (N_20038,N_19824,N_15499);
xnor U20039 (N_20039,N_17604,N_18277);
nor U20040 (N_20040,N_18588,N_18930);
nand U20041 (N_20041,N_16918,N_17449);
and U20042 (N_20042,N_19304,N_17120);
nor U20043 (N_20043,N_19525,N_18798);
nand U20044 (N_20044,N_19513,N_16510);
or U20045 (N_20045,N_19965,N_15927);
or U20046 (N_20046,N_15888,N_16002);
nand U20047 (N_20047,N_19579,N_17576);
nand U20048 (N_20048,N_15521,N_18584);
nand U20049 (N_20049,N_19788,N_19792);
nand U20050 (N_20050,N_16812,N_15333);
nor U20051 (N_20051,N_19782,N_17016);
nand U20052 (N_20052,N_15875,N_19204);
and U20053 (N_20053,N_17111,N_19015);
or U20054 (N_20054,N_16489,N_18011);
nor U20055 (N_20055,N_17868,N_19795);
nand U20056 (N_20056,N_19623,N_17605);
nor U20057 (N_20057,N_15269,N_18231);
nand U20058 (N_20058,N_15427,N_15725);
or U20059 (N_20059,N_15759,N_19903);
or U20060 (N_20060,N_19866,N_19004);
nor U20061 (N_20061,N_17144,N_16701);
and U20062 (N_20062,N_18511,N_19982);
nor U20063 (N_20063,N_15250,N_17558);
nand U20064 (N_20064,N_16749,N_17821);
nand U20065 (N_20065,N_15787,N_19742);
nand U20066 (N_20066,N_15490,N_18091);
nor U20067 (N_20067,N_19109,N_17982);
and U20068 (N_20068,N_15771,N_18600);
xor U20069 (N_20069,N_15190,N_17525);
and U20070 (N_20070,N_16517,N_16369);
nand U20071 (N_20071,N_15273,N_18536);
nor U20072 (N_20072,N_16471,N_17112);
xnor U20073 (N_20073,N_16128,N_15425);
xnor U20074 (N_20074,N_16263,N_15102);
nand U20075 (N_20075,N_19231,N_19744);
nor U20076 (N_20076,N_15707,N_19191);
xor U20077 (N_20077,N_18684,N_19755);
and U20078 (N_20078,N_17999,N_15712);
and U20079 (N_20079,N_17370,N_17871);
nand U20080 (N_20080,N_17615,N_19937);
xnor U20081 (N_20081,N_19233,N_16589);
and U20082 (N_20082,N_17553,N_17170);
and U20083 (N_20083,N_15600,N_16525);
nor U20084 (N_20084,N_16081,N_15123);
xor U20085 (N_20085,N_18691,N_15554);
and U20086 (N_20086,N_18810,N_16506);
nor U20087 (N_20087,N_18731,N_15428);
xnor U20088 (N_20088,N_15642,N_16898);
xor U20089 (N_20089,N_17331,N_18363);
nor U20090 (N_20090,N_16815,N_16590);
and U20091 (N_20091,N_15640,N_19749);
xnor U20092 (N_20092,N_19692,N_17712);
and U20093 (N_20093,N_16367,N_16714);
nand U20094 (N_20094,N_16177,N_17555);
and U20095 (N_20095,N_18248,N_16200);
or U20096 (N_20096,N_16915,N_17841);
nand U20097 (N_20097,N_19269,N_15698);
nor U20098 (N_20098,N_16285,N_17932);
or U20099 (N_20099,N_17595,N_15589);
nand U20100 (N_20100,N_15797,N_17973);
xnor U20101 (N_20101,N_18967,N_19898);
nand U20102 (N_20102,N_15505,N_18583);
xnor U20103 (N_20103,N_18595,N_18829);
xor U20104 (N_20104,N_17183,N_16453);
and U20105 (N_20105,N_19962,N_18893);
or U20106 (N_20106,N_16171,N_16700);
nor U20107 (N_20107,N_17197,N_19565);
or U20108 (N_20108,N_15268,N_15743);
xor U20109 (N_20109,N_18636,N_19650);
xnor U20110 (N_20110,N_15384,N_18179);
or U20111 (N_20111,N_16225,N_16341);
nand U20112 (N_20112,N_16187,N_18449);
xor U20113 (N_20113,N_15789,N_18433);
nor U20114 (N_20114,N_18549,N_17368);
nor U20115 (N_20115,N_19176,N_16325);
nor U20116 (N_20116,N_18198,N_17946);
xnor U20117 (N_20117,N_15005,N_19315);
nand U20118 (N_20118,N_19006,N_15949);
and U20119 (N_20119,N_17019,N_16595);
or U20120 (N_20120,N_18696,N_17078);
nand U20121 (N_20121,N_19138,N_16791);
xor U20122 (N_20122,N_19709,N_16680);
nand U20123 (N_20123,N_17560,N_16227);
nor U20124 (N_20124,N_16264,N_18577);
and U20125 (N_20125,N_19802,N_15072);
and U20126 (N_20126,N_15101,N_16523);
or U20127 (N_20127,N_16644,N_18215);
xor U20128 (N_20128,N_15568,N_17412);
xor U20129 (N_20129,N_19633,N_17386);
or U20130 (N_20130,N_17313,N_18516);
nand U20131 (N_20131,N_18352,N_16443);
xor U20132 (N_20132,N_15987,N_19083);
nand U20133 (N_20133,N_17282,N_18382);
nand U20134 (N_20134,N_19930,N_18233);
or U20135 (N_20135,N_17659,N_16097);
nor U20136 (N_20136,N_16555,N_19121);
and U20137 (N_20137,N_15919,N_19759);
xor U20138 (N_20138,N_18790,N_15671);
nor U20139 (N_20139,N_19710,N_16474);
xor U20140 (N_20140,N_19575,N_17749);
or U20141 (N_20141,N_17708,N_17457);
nand U20142 (N_20142,N_18517,N_16927);
xnor U20143 (N_20143,N_18946,N_18146);
and U20144 (N_20144,N_18243,N_17741);
or U20145 (N_20145,N_15112,N_17783);
and U20146 (N_20146,N_17900,N_15256);
or U20147 (N_20147,N_17715,N_16848);
or U20148 (N_20148,N_17498,N_15780);
nand U20149 (N_20149,N_15355,N_18408);
nor U20150 (N_20150,N_17452,N_17430);
or U20151 (N_20151,N_15196,N_19028);
or U20152 (N_20152,N_16014,N_16465);
nand U20153 (N_20153,N_15178,N_19154);
nor U20154 (N_20154,N_18926,N_19378);
nand U20155 (N_20155,N_19098,N_19684);
nand U20156 (N_20156,N_18418,N_19757);
nor U20157 (N_20157,N_17125,N_18532);
nand U20158 (N_20158,N_18415,N_18148);
nand U20159 (N_20159,N_16683,N_18786);
nand U20160 (N_20160,N_19527,N_18237);
or U20161 (N_20161,N_19890,N_15952);
or U20162 (N_20162,N_18384,N_17159);
and U20163 (N_20163,N_17311,N_19563);
nor U20164 (N_20164,N_17419,N_15633);
nand U20165 (N_20165,N_18041,N_19752);
and U20166 (N_20166,N_15177,N_19354);
or U20167 (N_20167,N_16747,N_19221);
and U20168 (N_20168,N_17163,N_18441);
nand U20169 (N_20169,N_16179,N_16188);
nor U20170 (N_20170,N_16573,N_16382);
and U20171 (N_20171,N_16737,N_18285);
and U20172 (N_20172,N_19251,N_16221);
and U20173 (N_20173,N_18365,N_18149);
nand U20174 (N_20174,N_18085,N_15217);
nand U20175 (N_20175,N_18013,N_16193);
nor U20176 (N_20176,N_15948,N_16882);
nand U20177 (N_20177,N_19564,N_18722);
nor U20178 (N_20178,N_19413,N_19417);
xnor U20179 (N_20179,N_18524,N_15233);
nor U20180 (N_20180,N_17438,N_19035);
or U20181 (N_20181,N_17556,N_18079);
and U20182 (N_20182,N_18301,N_17347);
xor U20183 (N_20183,N_18891,N_16141);
and U20184 (N_20184,N_17819,N_16302);
or U20185 (N_20185,N_19566,N_17845);
nand U20186 (N_20186,N_16342,N_19783);
nand U20187 (N_20187,N_18554,N_15654);
nor U20188 (N_20188,N_15489,N_18349);
or U20189 (N_20189,N_18681,N_17149);
nor U20190 (N_20190,N_15661,N_15764);
and U20191 (N_20191,N_19870,N_17538);
nand U20192 (N_20192,N_15594,N_18279);
nand U20193 (N_20193,N_17917,N_19119);
nand U20194 (N_20194,N_19241,N_16062);
nand U20195 (N_20195,N_19701,N_18097);
nor U20196 (N_20196,N_16396,N_19080);
nand U20197 (N_20197,N_18473,N_15717);
or U20198 (N_20198,N_19326,N_15260);
nand U20199 (N_20199,N_15807,N_16486);
xnor U20200 (N_20200,N_16088,N_18499);
or U20201 (N_20201,N_17596,N_18269);
nand U20202 (N_20202,N_15213,N_17619);
nor U20203 (N_20203,N_19586,N_19546);
xor U20204 (N_20204,N_17587,N_17543);
nand U20205 (N_20205,N_18306,N_18051);
and U20206 (N_20206,N_16482,N_17451);
and U20207 (N_20207,N_17667,N_15039);
or U20208 (N_20208,N_15198,N_18420);
and U20209 (N_20209,N_18741,N_18840);
or U20210 (N_20210,N_17432,N_19092);
nand U20211 (N_20211,N_18435,N_16360);
nand U20212 (N_20212,N_15110,N_18181);
and U20213 (N_20213,N_17084,N_19143);
or U20214 (N_20214,N_19186,N_16874);
nor U20215 (N_20215,N_19472,N_16261);
nand U20216 (N_20216,N_17924,N_17469);
nor U20217 (N_20217,N_17006,N_15267);
or U20218 (N_20218,N_15093,N_19307);
nand U20219 (N_20219,N_17931,N_17955);
or U20220 (N_20220,N_15348,N_16638);
nor U20221 (N_20221,N_17592,N_15465);
nor U20222 (N_20222,N_15484,N_18980);
and U20223 (N_20223,N_15538,N_17192);
nand U20224 (N_20224,N_16295,N_17651);
xnor U20225 (N_20225,N_18800,N_15106);
or U20226 (N_20226,N_19569,N_15630);
nand U20227 (N_20227,N_15530,N_17358);
nor U20228 (N_20228,N_15091,N_17756);
nand U20229 (N_20229,N_17897,N_15843);
nand U20230 (N_20230,N_16111,N_19626);
or U20231 (N_20231,N_19531,N_19368);
or U20232 (N_20232,N_17961,N_19522);
xnor U20233 (N_20233,N_17540,N_17864);
nor U20234 (N_20234,N_19858,N_16702);
or U20235 (N_20235,N_19777,N_15165);
nor U20236 (N_20236,N_19851,N_19311);
and U20237 (N_20237,N_18389,N_17929);
and U20238 (N_20238,N_17586,N_19722);
nand U20239 (N_20239,N_16715,N_18987);
nand U20240 (N_20240,N_16593,N_19706);
nor U20241 (N_20241,N_16576,N_19585);
or U20242 (N_20242,N_17122,N_16755);
nor U20243 (N_20243,N_15517,N_17272);
nand U20244 (N_20244,N_15728,N_15398);
and U20245 (N_20245,N_16330,N_18200);
and U20246 (N_20246,N_16828,N_19699);
nor U20247 (N_20247,N_15914,N_18721);
and U20248 (N_20248,N_16730,N_17017);
nand U20249 (N_20249,N_19625,N_18468);
nand U20250 (N_20250,N_15090,N_16024);
nor U20251 (N_20251,N_16960,N_15758);
xor U20252 (N_20252,N_16331,N_17926);
nor U20253 (N_20253,N_17348,N_18502);
and U20254 (N_20254,N_16826,N_18672);
xnor U20255 (N_20255,N_16228,N_16375);
nand U20256 (N_20256,N_16671,N_16266);
xnor U20257 (N_20257,N_15040,N_16237);
xor U20258 (N_20258,N_17504,N_16243);
xor U20259 (N_20259,N_17557,N_18015);
nor U20260 (N_20260,N_17970,N_18388);
or U20261 (N_20261,N_16952,N_19117);
nor U20262 (N_20262,N_16378,N_17859);
nand U20263 (N_20263,N_19881,N_18560);
xor U20264 (N_20264,N_16026,N_17207);
nand U20265 (N_20265,N_16911,N_18916);
nor U20266 (N_20266,N_19369,N_17645);
nor U20267 (N_20267,N_19578,N_17026);
or U20268 (N_20268,N_15850,N_19276);
xnor U20269 (N_20269,N_18142,N_17940);
nand U20270 (N_20270,N_16183,N_19761);
nor U20271 (N_20271,N_19988,N_19935);
nand U20272 (N_20272,N_19164,N_17184);
nand U20273 (N_20273,N_15244,N_18644);
nand U20274 (N_20274,N_18400,N_16254);
nor U20275 (N_20275,N_19443,N_15786);
or U20276 (N_20276,N_18050,N_19172);
or U20277 (N_20277,N_18302,N_17883);
nand U20278 (N_20278,N_18609,N_16257);
xnor U20279 (N_20279,N_15898,N_16125);
and U20280 (N_20280,N_16716,N_17918);
nand U20281 (N_20281,N_18804,N_18642);
or U20282 (N_20282,N_16793,N_17690);
or U20283 (N_20283,N_19708,N_15611);
nand U20284 (N_20284,N_19153,N_16640);
or U20285 (N_20285,N_15070,N_19665);
and U20286 (N_20286,N_16387,N_16122);
xnor U20287 (N_20287,N_15374,N_17182);
xor U20288 (N_20288,N_17660,N_19856);
nor U20289 (N_20289,N_19689,N_19053);
and U20290 (N_20290,N_18197,N_18346);
and U20291 (N_20291,N_15316,N_18839);
and U20292 (N_20292,N_19345,N_15009);
and U20293 (N_20293,N_17385,N_18378);
xor U20294 (N_20294,N_18640,N_17123);
and U20295 (N_20295,N_18212,N_15904);
or U20296 (N_20296,N_15537,N_18304);
and U20297 (N_20297,N_15666,N_18712);
and U20298 (N_20298,N_18876,N_18907);
nor U20299 (N_20299,N_17088,N_17700);
xor U20300 (N_20300,N_19885,N_19646);
or U20301 (N_20301,N_18870,N_18170);
nand U20302 (N_20302,N_18300,N_18906);
xor U20303 (N_20303,N_16194,N_16980);
nor U20304 (N_20304,N_19057,N_16604);
and U20305 (N_20305,N_19132,N_18358);
nor U20306 (N_20306,N_17133,N_17099);
or U20307 (N_20307,N_18463,N_18929);
nor U20308 (N_20308,N_15432,N_16448);
or U20309 (N_20309,N_15004,N_16211);
or U20310 (N_20310,N_16923,N_16881);
or U20311 (N_20311,N_17481,N_17794);
nand U20312 (N_20312,N_16279,N_19246);
and U20313 (N_20313,N_18944,N_18796);
and U20314 (N_20314,N_17701,N_17761);
and U20315 (N_20315,N_16912,N_15491);
nor U20316 (N_20316,N_18496,N_18716);
and U20317 (N_20317,N_17601,N_15601);
or U20318 (N_20318,N_19543,N_19632);
and U20319 (N_20319,N_15175,N_19591);
nor U20320 (N_20320,N_15917,N_19404);
nor U20321 (N_20321,N_16854,N_19674);
xor U20322 (N_20322,N_16428,N_16891);
nand U20323 (N_20323,N_17698,N_18625);
xor U20324 (N_20324,N_19334,N_18785);
nor U20325 (N_20325,N_15638,N_17721);
nor U20326 (N_20326,N_18002,N_17625);
or U20327 (N_20327,N_16823,N_19495);
or U20328 (N_20328,N_15125,N_15691);
nor U20329 (N_20329,N_17409,N_16229);
xnor U20330 (N_20330,N_17008,N_16032);
or U20331 (N_20331,N_19341,N_15367);
nand U20332 (N_20332,N_17421,N_19484);
and U20333 (N_20333,N_16042,N_16837);
nor U20334 (N_20334,N_16588,N_19726);
nand U20335 (N_20335,N_17166,N_16144);
or U20336 (N_20336,N_17140,N_18127);
or U20337 (N_20337,N_19298,N_17442);
and U20338 (N_20338,N_15603,N_15580);
and U20339 (N_20339,N_19616,N_19147);
nand U20340 (N_20340,N_17983,N_15403);
nand U20341 (N_20341,N_15581,N_15080);
or U20342 (N_20342,N_17366,N_17589);
and U20343 (N_20343,N_19451,N_19691);
nor U20344 (N_20344,N_15120,N_16729);
nand U20345 (N_20345,N_15647,N_15117);
and U20346 (N_20346,N_19075,N_17908);
nand U20347 (N_20347,N_15905,N_16920);
or U20348 (N_20348,N_16087,N_17969);
nor U20349 (N_20349,N_19806,N_18303);
nor U20350 (N_20350,N_17742,N_16623);
or U20351 (N_20351,N_15306,N_19405);
nand U20352 (N_20352,N_19801,N_19485);
and U20353 (N_20353,N_18479,N_17005);
nand U20354 (N_20354,N_17851,N_15939);
nand U20355 (N_20355,N_15363,N_19009);
and U20356 (N_20356,N_16078,N_15736);
and U20357 (N_20357,N_16620,N_17893);
nor U20358 (N_20358,N_16413,N_19707);
or U20359 (N_20359,N_18529,N_17580);
xor U20360 (N_20360,N_17217,N_19395);
or U20361 (N_20361,N_17633,N_15584);
and U20362 (N_20362,N_15225,N_18882);
xor U20363 (N_20363,N_18066,N_15562);
or U20364 (N_20364,N_17433,N_16584);
or U20365 (N_20365,N_17478,N_18868);
nand U20366 (N_20366,N_19313,N_18989);
nand U20367 (N_20367,N_19322,N_18006);
and U20368 (N_20368,N_15902,N_19996);
nor U20369 (N_20369,N_18328,N_15776);
and U20370 (N_20370,N_18635,N_15082);
nor U20371 (N_20371,N_18090,N_16528);
or U20372 (N_20372,N_15279,N_16132);
and U20373 (N_20373,N_15632,N_18646);
and U20374 (N_20374,N_18802,N_19100);
nor U20375 (N_20375,N_16675,N_15286);
xor U20376 (N_20376,N_15551,N_18522);
nand U20377 (N_20377,N_17549,N_18617);
xor U20378 (N_20378,N_19540,N_19581);
and U20379 (N_20379,N_16344,N_15720);
or U20380 (N_20380,N_18847,N_15596);
xnor U20381 (N_20381,N_18183,N_19779);
nand U20382 (N_20382,N_18586,N_16697);
or U20383 (N_20383,N_18470,N_15578);
nor U20384 (N_20384,N_15909,N_15969);
nand U20385 (N_20385,N_16648,N_17569);
xnor U20386 (N_20386,N_16880,N_19904);
nor U20387 (N_20387,N_18224,N_18497);
xor U20388 (N_20388,N_16505,N_15417);
or U20389 (N_20389,N_15767,N_16735);
xor U20390 (N_20390,N_19274,N_19651);
xnor U20391 (N_20391,N_17669,N_16296);
nand U20392 (N_20392,N_16585,N_17734);
nand U20393 (N_20393,N_17617,N_17920);
nor U20394 (N_20394,N_15752,N_19515);
xnor U20395 (N_20395,N_19349,N_18422);
and U20396 (N_20396,N_17722,N_19401);
nand U20397 (N_20397,N_15135,N_17025);
nor U20398 (N_20398,N_16318,N_15038);
xor U20399 (N_20399,N_18659,N_16391);
xnor U20400 (N_20400,N_15295,N_17208);
or U20401 (N_20401,N_19964,N_16819);
nor U20402 (N_20402,N_16779,N_15907);
or U20403 (N_20403,N_15227,N_16343);
or U20404 (N_20404,N_18707,N_15372);
nand U20405 (N_20405,N_16821,N_17551);
nor U20406 (N_20406,N_19677,N_17263);
or U20407 (N_20407,N_19848,N_18728);
nor U20408 (N_20408,N_19643,N_17839);
nand U20409 (N_20409,N_18357,N_15547);
nor U20410 (N_20410,N_19201,N_17583);
nand U20411 (N_20411,N_15754,N_18272);
nand U20412 (N_20412,N_18461,N_17675);
xnor U20413 (N_20413,N_15404,N_16870);
xor U20414 (N_20414,N_19849,N_15219);
nor U20415 (N_20415,N_19679,N_19729);
and U20416 (N_20416,N_17502,N_17731);
xnor U20417 (N_20417,N_16722,N_18106);
xor U20418 (N_20418,N_19590,N_17817);
nand U20419 (N_20419,N_16797,N_15446);
and U20420 (N_20420,N_17823,N_17995);
and U20421 (N_20421,N_15958,N_15692);
or U20422 (N_20422,N_15027,N_19460);
or U20423 (N_20423,N_16594,N_15294);
and U20424 (N_20424,N_15650,N_15173);
nand U20425 (N_20425,N_16196,N_19774);
nand U20426 (N_20426,N_18897,N_15516);
xor U20427 (N_20427,N_15186,N_16503);
or U20428 (N_20428,N_17243,N_16332);
nor U20429 (N_20429,N_17349,N_16514);
or U20430 (N_20430,N_19573,N_16490);
nand U20431 (N_20431,N_16885,N_17379);
and U20432 (N_20432,N_17608,N_17226);
nand U20433 (N_20433,N_17162,N_17703);
and U20434 (N_20434,N_15335,N_17332);
or U20435 (N_20435,N_15284,N_19867);
xnor U20436 (N_20436,N_15890,N_17648);
or U20437 (N_20437,N_15270,N_16925);
xnor U20438 (N_20438,N_16669,N_15634);
nand U20439 (N_20439,N_15445,N_17739);
nand U20440 (N_20440,N_19514,N_17966);
and U20441 (N_20441,N_18665,N_18585);
and U20442 (N_20442,N_19713,N_18207);
nand U20443 (N_20443,N_16452,N_15688);
nor U20444 (N_20444,N_15867,N_15968);
nor U20445 (N_20445,N_18874,N_16255);
nand U20446 (N_20446,N_15183,N_18682);
nand U20447 (N_20447,N_18219,N_18782);
and U20448 (N_20448,N_15886,N_17777);
nand U20449 (N_20449,N_16287,N_17980);
nand U20450 (N_20450,N_16904,N_16770);
xor U20451 (N_20451,N_17262,N_16617);
nand U20452 (N_20452,N_19029,N_19198);
and U20453 (N_20453,N_17004,N_18784);
nand U20454 (N_20454,N_18787,N_15320);
and U20455 (N_20455,N_19022,N_19456);
and U20456 (N_20456,N_17156,N_17414);
xor U20457 (N_20457,N_19287,N_17867);
or U20458 (N_20458,N_15723,N_17958);
nor U20459 (N_20459,N_17629,N_16077);
nand U20460 (N_20460,N_16075,N_19812);
and U20461 (N_20461,N_16061,N_19628);
or U20462 (N_20462,N_18995,N_18683);
and U20463 (N_20463,N_18689,N_15437);
and U20464 (N_20464,N_15689,N_16892);
or U20465 (N_20465,N_17674,N_18706);
or U20466 (N_20466,N_18092,N_16049);
nand U20467 (N_20467,N_16532,N_19089);
and U20468 (N_20468,N_15853,N_15142);
nor U20469 (N_20469,N_18291,N_15223);
nand U20470 (N_20470,N_16074,N_18112);
nand U20471 (N_20471,N_19469,N_15696);
and U20472 (N_20472,N_16928,N_17664);
nor U20473 (N_20473,N_15032,N_17820);
nor U20474 (N_20474,N_17631,N_19220);
nor U20475 (N_20475,N_15096,N_16426);
and U20476 (N_20476,N_15871,N_16571);
and U20477 (N_20477,N_16771,N_17101);
nand U20478 (N_20478,N_19283,N_19592);
xor U20479 (N_20479,N_17776,N_15181);
xnor U20480 (N_20480,N_18169,N_16878);
nor U20481 (N_20481,N_16563,N_19086);
nor U20482 (N_20482,N_17406,N_18189);
and U20483 (N_20483,N_16516,N_19482);
xor U20484 (N_20484,N_16629,N_19832);
xor U20485 (N_20485,N_19256,N_19427);
or U20486 (N_20486,N_19464,N_18992);
and U20487 (N_20487,N_15327,N_17107);
or U20488 (N_20488,N_15699,N_15237);
or U20489 (N_20489,N_17216,N_17933);
or U20490 (N_20490,N_16395,N_18052);
or U20491 (N_20491,N_15702,N_17344);
nor U20492 (N_20492,N_18740,N_15734);
nor U20493 (N_20493,N_18620,N_18493);
and U20494 (N_20494,N_17997,N_16513);
nand U20495 (N_20495,N_16053,N_17275);
or U20496 (N_20496,N_18699,N_19855);
xnor U20497 (N_20497,N_17146,N_18736);
xnor U20498 (N_20498,N_15228,N_16829);
nor U20499 (N_20499,N_15148,N_19811);
or U20500 (N_20500,N_18571,N_19175);
nand U20501 (N_20501,N_19069,N_16143);
nand U20502 (N_20502,N_19768,N_15662);
and U20503 (N_20503,N_18593,N_15412);
nor U20504 (N_20504,N_16873,N_16795);
nor U20505 (N_20505,N_16526,N_19805);
and U20506 (N_20506,N_15990,N_19810);
and U20507 (N_20507,N_15812,N_19853);
and U20508 (N_20508,N_18982,N_18668);
or U20509 (N_20509,N_15556,N_18923);
nand U20510 (N_20510,N_16639,N_18454);
and U20511 (N_20511,N_18564,N_19895);
nand U20512 (N_20512,N_19775,N_17719);
and U20513 (N_20513,N_18203,N_17288);
or U20514 (N_20514,N_16041,N_15976);
and U20515 (N_20515,N_19305,N_16723);
or U20516 (N_20516,N_17373,N_18514);
or U20517 (N_20517,N_15230,N_16043);
nor U20518 (N_20518,N_17733,N_19001);
xnor U20519 (N_20519,N_15152,N_19258);
nand U20520 (N_20520,N_18698,N_15208);
nor U20521 (N_20521,N_17322,N_15806);
nor U20522 (N_20522,N_18236,N_19668);
nor U20523 (N_20523,N_15302,N_19847);
or U20524 (N_20524,N_15724,N_19126);
xnor U20525 (N_20525,N_15681,N_15486);
or U20526 (N_20526,N_17100,N_17899);
and U20527 (N_20527,N_15627,N_17662);
nor U20528 (N_20528,N_19297,N_18794);
nand U20529 (N_20529,N_17098,N_19398);
nor U20530 (N_20530,N_18037,N_17812);
nor U20531 (N_20531,N_15560,N_15705);
and U20532 (N_20532,N_17874,N_16006);
and U20533 (N_20533,N_18402,N_19925);
xor U20534 (N_20534,N_15733,N_16762);
or U20535 (N_20535,N_16662,N_17178);
or U20536 (N_20536,N_19008,N_19224);
nor U20537 (N_20537,N_19502,N_16300);
nor U20538 (N_20538,N_16174,N_16007);
nor U20539 (N_20539,N_15121,N_17167);
and U20540 (N_20540,N_19010,N_17071);
xor U20541 (N_20541,N_17251,N_19868);
or U20542 (N_20542,N_17080,N_16052);
nor U20543 (N_20543,N_16400,N_18438);
or U20544 (N_20544,N_16371,N_15378);
xnor U20545 (N_20545,N_15388,N_17422);
nor U20546 (N_20546,N_19597,N_16252);
nor U20547 (N_20547,N_15829,N_17239);
and U20548 (N_20548,N_19636,N_17278);
nor U20549 (N_20549,N_19149,N_15804);
xor U20550 (N_20550,N_15245,N_15677);
and U20551 (N_20551,N_17896,N_19447);
nand U20552 (N_20552,N_15848,N_18242);
and U20553 (N_20553,N_16023,N_19205);
xor U20554 (N_20554,N_19393,N_17530);
nor U20555 (N_20555,N_19917,N_18833);
nand U20556 (N_20556,N_17027,N_16462);
or U20557 (N_20557,N_15906,N_19661);
nand U20558 (N_20558,N_19066,N_16769);
and U20559 (N_20559,N_18184,N_17427);
nand U20560 (N_20560,N_16767,N_15587);
and U20561 (N_20561,N_19350,N_16092);
nor U20562 (N_20562,N_15229,N_16470);
and U20563 (N_20563,N_15645,N_18019);
and U20564 (N_20564,N_16085,N_15021);
nor U20565 (N_20565,N_15672,N_19196);
and U20566 (N_20566,N_17890,N_19905);
or U20567 (N_20567,N_19237,N_17470);
and U20568 (N_20568,N_18812,N_17060);
nand U20569 (N_20569,N_19356,N_19183);
nor U20570 (N_20570,N_19902,N_17497);
nand U20571 (N_20571,N_19444,N_17547);
xor U20572 (N_20572,N_19470,N_18459);
nor U20573 (N_20573,N_15305,N_15343);
nor U20574 (N_20574,N_15071,N_15053);
nor U20575 (N_20575,N_19946,N_19989);
nor U20576 (N_20576,N_16760,N_17467);
or U20577 (N_20577,N_17032,N_15998);
nor U20578 (N_20578,N_16238,N_15003);
nor U20579 (N_20579,N_15299,N_15609);
nor U20580 (N_20580,N_19542,N_19963);
or U20581 (N_20581,N_19091,N_15795);
nor U20582 (N_20582,N_15095,N_18774);
nand U20583 (N_20583,N_19278,N_18674);
nor U20584 (N_20584,N_19202,N_15167);
nor U20585 (N_20585,N_18972,N_18191);
nor U20586 (N_20586,N_18316,N_17335);
and U20587 (N_20587,N_16399,N_18270);
and U20588 (N_20588,N_17124,N_17516);
nand U20589 (N_20589,N_16549,N_19532);
nor U20590 (N_20590,N_19861,N_16139);
xnor U20591 (N_20591,N_16977,N_19766);
or U20592 (N_20592,N_17475,N_17934);
xor U20593 (N_20593,N_15394,N_16724);
and U20594 (N_20594,N_16564,N_15644);
nor U20595 (N_20595,N_15985,N_18743);
nand U20596 (N_20596,N_16556,N_17378);
nor U20597 (N_20597,N_19418,N_17264);
or U20598 (N_20598,N_19177,N_19099);
nor U20599 (N_20599,N_17987,N_19449);
or U20600 (N_20600,N_15089,N_18824);
or U20601 (N_20601,N_19271,N_17713);
nor U20602 (N_20602,N_16844,N_15471);
nor U20603 (N_20603,N_15441,N_18652);
nor U20604 (N_20604,N_15264,N_18278);
xnor U20605 (N_20605,N_16384,N_15391);
nand U20606 (N_20606,N_18596,N_16996);
nor U20607 (N_20607,N_16872,N_15304);
nand U20608 (N_20608,N_16319,N_15463);
nand U20609 (N_20609,N_16083,N_17056);
nor U20610 (N_20610,N_17772,N_17334);
nand U20611 (N_20611,N_15766,N_17753);
nor U20612 (N_20612,N_19785,N_19975);
xor U20613 (N_20613,N_17822,N_15874);
nand U20614 (N_20614,N_16630,N_19376);
nand U20615 (N_20615,N_15986,N_17585);
nor U20616 (N_20616,N_16094,N_18150);
and U20617 (N_20617,N_18979,N_15711);
nor U20618 (N_20618,N_16560,N_16045);
and U20619 (N_20619,N_18581,N_15818);
or U20620 (N_20620,N_19997,N_16364);
nand U20621 (N_20621,N_15133,N_17573);
xnor U20622 (N_20622,N_17431,N_17345);
xnor U20623 (N_20623,N_17301,N_16794);
xor U20624 (N_20624,N_19512,N_18007);
xor U20625 (N_20625,N_16637,N_16333);
and U20626 (N_20626,N_17831,N_16982);
nand U20627 (N_20627,N_16070,N_19266);
nand U20628 (N_20628,N_18759,N_17299);
xnor U20629 (N_20629,N_19402,N_19430);
nor U20630 (N_20630,N_15790,N_16863);
xnor U20631 (N_20631,N_16558,N_17750);
or U20632 (N_20632,N_19941,N_15314);
or U20633 (N_20633,N_17042,N_16412);
or U20634 (N_20634,N_19926,N_15138);
or U20635 (N_20635,N_15092,N_18160);
or U20636 (N_20636,N_18024,N_19945);
nor U20637 (N_20637,N_16419,N_15535);
or U20638 (N_20638,N_18263,N_16297);
or U20639 (N_20639,N_18808,N_17186);
or U20640 (N_20640,N_16226,N_18241);
and U20641 (N_20641,N_19245,N_15659);
or U20642 (N_20642,N_16710,N_16191);
or U20643 (N_20643,N_15452,N_19052);
nand U20644 (N_20644,N_19455,N_18448);
or U20645 (N_20645,N_17179,N_15389);
nor U20646 (N_20646,N_18877,N_19296);
nor U20647 (N_20647,N_17757,N_17280);
or U20648 (N_20648,N_18362,N_15532);
and U20649 (N_20649,N_16929,N_16274);
and U20650 (N_20650,N_18818,N_19445);
xnor U20651 (N_20651,N_17109,N_17474);
and U20652 (N_20652,N_15149,N_17744);
and U20653 (N_20653,N_16789,N_15994);
or U20654 (N_20654,N_16845,N_15860);
or U20655 (N_20655,N_18273,N_16491);
or U20656 (N_20656,N_15438,N_18779);
or U20657 (N_20657,N_17465,N_17425);
nand U20658 (N_20658,N_15066,N_17643);
and U20659 (N_20659,N_18902,N_18262);
or U20660 (N_20660,N_16046,N_19051);
nor U20661 (N_20661,N_16401,N_19259);
and U20662 (N_20662,N_16322,N_17351);
nor U20663 (N_20663,N_18455,N_16890);
nor U20664 (N_20664,N_18044,N_15664);
nand U20665 (N_20665,N_18309,N_19005);
xnor U20666 (N_20666,N_18708,N_16015);
nor U20667 (N_20667,N_16627,N_17150);
or U20668 (N_20668,N_19310,N_18159);
and U20669 (N_20669,N_19108,N_18151);
xor U20670 (N_20670,N_19864,N_17325);
nor U20671 (N_20671,N_18144,N_17290);
xor U20672 (N_20672,N_18857,N_18942);
and U20673 (N_20673,N_19776,N_17130);
nor U20674 (N_20674,N_17229,N_16734);
or U20675 (N_20675,N_15319,N_15016);
nor U20676 (N_20676,N_17837,N_18440);
nor U20677 (N_20677,N_18098,N_15118);
nand U20678 (N_20678,N_16922,N_15513);
xor U20679 (N_20679,N_19388,N_19574);
xnor U20680 (N_20680,N_19223,N_17047);
xnor U20681 (N_20681,N_15155,N_18315);
nor U20682 (N_20682,N_18582,N_18017);
nand U20683 (N_20683,N_18922,N_17287);
nor U20684 (N_20684,N_17909,N_18719);
nor U20685 (N_20685,N_19182,N_18361);
and U20686 (N_20686,N_18673,N_19658);
nand U20687 (N_20687,N_19714,N_15376);
or U20688 (N_20688,N_16250,N_18837);
nor U20689 (N_20689,N_17488,N_18483);
nand U20690 (N_20690,N_18457,N_18558);
nor U20691 (N_20691,N_15188,N_15478);
nand U20692 (N_20692,N_18484,N_17956);
nand U20693 (N_20693,N_18758,N_15328);
xnor U20694 (N_20694,N_17443,N_17256);
or U20695 (N_20695,N_16393,N_16059);
or U20696 (N_20696,N_19107,N_17670);
or U20697 (N_20697,N_18310,N_18261);
xnor U20698 (N_20698,N_19538,N_18020);
nor U20699 (N_20699,N_17730,N_15243);
nor U20700 (N_20700,N_17418,N_15126);
nand U20701 (N_20701,N_19375,N_18095);
and U20702 (N_20702,N_17702,N_19837);
and U20703 (N_20703,N_19551,N_17834);
nor U20704 (N_20704,N_16899,N_18783);
and U20705 (N_20705,N_15278,N_15653);
nor U20706 (N_20706,N_17528,N_17141);
or U20707 (N_20707,N_18210,N_19718);
nand U20708 (N_20708,N_19739,N_17339);
nand U20709 (N_20709,N_18534,N_16135);
nor U20710 (N_20710,N_15467,N_17018);
and U20711 (N_20711,N_17402,N_16543);
nor U20712 (N_20712,N_19060,N_18955);
nor U20713 (N_20713,N_16358,N_18761);
nand U20714 (N_20714,N_18566,N_19031);
nand U20715 (N_20715,N_17070,N_16622);
xor U20716 (N_20716,N_15310,N_15393);
or U20717 (N_20717,N_19167,N_18725);
or U20718 (N_20718,N_18383,N_16231);
nand U20719 (N_20719,N_19784,N_15342);
or U20720 (N_20720,N_18825,N_17395);
and U20721 (N_20721,N_18676,N_18768);
nand U20722 (N_20722,N_18062,N_17872);
or U20723 (N_20723,N_15882,N_17472);
xor U20724 (N_20724,N_18744,N_17135);
nor U20725 (N_20725,N_18578,N_19353);
nor U20726 (N_20726,N_18605,N_15041);
nor U20727 (N_20727,N_16473,N_16197);
xor U20728 (N_20728,N_15730,N_18040);
nand U20729 (N_20729,N_17487,N_19084);
and U20730 (N_20730,N_15259,N_19827);
nand U20731 (N_20731,N_19758,N_16608);
nor U20732 (N_20732,N_19803,N_19748);
and U20733 (N_20733,N_16145,N_16783);
nand U20734 (N_20734,N_19419,N_17416);
and U20735 (N_20735,N_16368,N_15934);
and U20736 (N_20736,N_18234,N_18196);
nand U20737 (N_20737,N_18747,N_16668);
nand U20738 (N_20738,N_15756,N_18228);
xor U20739 (N_20739,N_16600,N_18900);
nand U20740 (N_20740,N_15201,N_16066);
and U20741 (N_20741,N_18750,N_15447);
xor U20742 (N_20742,N_15346,N_18351);
nand U20743 (N_20743,N_18249,N_17889);
nand U20744 (N_20744,N_17976,N_15064);
or U20745 (N_20745,N_17618,N_18940);
nor U20746 (N_20746,N_16997,N_17858);
nor U20747 (N_20747,N_15891,N_16843);
nand U20748 (N_20748,N_19994,N_18244);
nor U20749 (N_20749,N_18947,N_17672);
and U20750 (N_20750,N_17410,N_17314);
or U20751 (N_20751,N_16834,N_17572);
xnor U20752 (N_20752,N_15205,N_19613);
nor U20753 (N_20753,N_19745,N_17471);
nor U20754 (N_20754,N_19943,N_17767);
nand U20755 (N_20755,N_16282,N_18456);
or U20756 (N_20756,N_17978,N_18070);
nand U20757 (N_20757,N_16324,N_16430);
nand U20758 (N_20758,N_19365,N_17447);
or U20759 (N_20759,N_16067,N_16582);
nand U20760 (N_20760,N_18976,N_16449);
nor U20761 (N_20761,N_15179,N_16501);
and U20762 (N_20762,N_16981,N_19063);
or U20763 (N_20763,N_19016,N_18108);
xor U20764 (N_20764,N_18500,N_17537);
nand U20765 (N_20765,N_16787,N_19772);
nor U20766 (N_20766,N_19712,N_19312);
xor U20767 (N_20767,N_16209,N_17594);
xnor U20768 (N_20768,N_19972,N_19200);
xor U20769 (N_20769,N_17392,N_16386);
or U20770 (N_20770,N_17145,N_17881);
nand U20771 (N_20771,N_19580,N_18592);
or U20772 (N_20772,N_15830,N_16704);
nor U20773 (N_20773,N_15169,N_18405);
nand U20774 (N_20774,N_19897,N_18012);
nor U20775 (N_20775,N_19385,N_19918);
xor U20776 (N_20776,N_16105,N_15176);
xnor U20777 (N_20777,N_15504,N_18873);
and U20778 (N_20778,N_16699,N_19642);
nor U20779 (N_20779,N_18852,N_18849);
nor U20780 (N_20780,N_19406,N_18655);
nand U20781 (N_20781,N_19736,N_16803);
nor U20782 (N_20782,N_18647,N_19372);
and U20783 (N_20783,N_19415,N_15762);
or U20784 (N_20784,N_16612,N_18222);
nor U20785 (N_20785,N_17876,N_15718);
nor U20786 (N_20786,N_18274,N_16973);
nand U20787 (N_20787,N_16677,N_19507);
xor U20788 (N_20788,N_17746,N_16314);
nor U20789 (N_20789,N_19044,N_17114);
xor U20790 (N_20790,N_17638,N_18447);
nor U20791 (N_20791,N_18956,N_19934);
or U20792 (N_20792,N_18133,N_15344);
xnor U20793 (N_20793,N_15920,N_17554);
nor U20794 (N_20794,N_18205,N_19833);
and U20795 (N_20795,N_19886,N_15159);
or U20796 (N_20796,N_17210,N_16178);
and U20797 (N_20797,N_17875,N_16365);
and U20798 (N_20798,N_16292,N_17259);
and U20799 (N_20799,N_15512,N_19351);
and U20800 (N_20800,N_16385,N_17965);
nor U20801 (N_20801,N_16862,N_17289);
and U20802 (N_20802,N_16799,N_16207);
nand U20803 (N_20803,N_18726,N_18426);
nand U20804 (N_20804,N_16148,N_15954);
xor U20805 (N_20805,N_16804,N_15262);
nor U20806 (N_20806,N_16645,N_16435);
nand U20807 (N_20807,N_19433,N_18147);
nand U20808 (N_20808,N_16467,N_15922);
nor U20809 (N_20809,N_15395,N_19206);
nor U20810 (N_20810,N_19670,N_16220);
and U20811 (N_20811,N_17223,N_18476);
xnor U20812 (N_20812,N_17759,N_18446);
nor U20813 (N_20813,N_17816,N_17201);
nor U20814 (N_20814,N_18981,N_17341);
nor U20815 (N_20815,N_15147,N_17132);
and U20816 (N_20816,N_17190,N_19872);
and U20817 (N_20817,N_17261,N_18757);
and U20818 (N_20818,N_16359,N_16987);
or U20819 (N_20819,N_18844,N_16404);
and U20820 (N_20820,N_19358,N_15060);
nand U20821 (N_20821,N_19762,N_19991);
nor U20822 (N_20822,N_15143,N_16667);
and U20823 (N_20823,N_15880,N_18086);
xor U20824 (N_20824,N_17584,N_16970);
nor U20825 (N_20825,N_17486,N_17950);
nor U20826 (N_20826,N_18700,N_19249);
nor U20827 (N_20827,N_15023,N_17495);
and U20828 (N_20828,N_18084,N_17877);
and U20829 (N_20829,N_15402,N_16832);
nand U20830 (N_20830,N_15199,N_15635);
xor U20831 (N_20831,N_17599,N_15729);
xor U20832 (N_20832,N_18053,N_15362);
nor U20833 (N_20833,N_15862,N_17514);
nor U20834 (N_20834,N_15020,N_17652);
and U20835 (N_20835,N_16583,N_18917);
and U20836 (N_20836,N_19227,N_19056);
and U20837 (N_20837,N_19103,N_16504);
xor U20838 (N_20838,N_16961,N_19329);
and U20839 (N_20839,N_17879,N_19948);
nor U20840 (N_20840,N_19352,N_15983);
or U20841 (N_20841,N_19698,N_15894);
nor U20842 (N_20842,N_16746,N_19047);
xnor U20843 (N_20843,N_17840,N_16478);
nor U20844 (N_20844,N_15300,N_19032);
nor U20845 (N_20845,N_18390,N_18997);
and U20846 (N_20846,N_16485,N_17075);
xnor U20847 (N_20847,N_19055,N_17523);
xor U20848 (N_20848,N_15180,N_16561);
and U20849 (N_20849,N_19026,N_19281);
nor U20850 (N_20850,N_18528,N_19199);
nor U20851 (N_20851,N_15876,N_16836);
nand U20852 (N_20852,N_17195,N_15022);
nand U20853 (N_20853,N_16858,N_17244);
xnor U20854 (N_20854,N_18094,N_18687);
and U20855 (N_20855,N_15553,N_18697);
nand U20856 (N_20856,N_17501,N_19448);
or U20857 (N_20857,N_19318,N_16036);
and U20858 (N_20858,N_19828,N_15145);
or U20859 (N_20859,N_17974,N_16293);
nor U20860 (N_20860,N_15622,N_16184);
xnor U20861 (N_20861,N_18226,N_17854);
or U20862 (N_20862,N_16777,N_17155);
or U20863 (N_20863,N_16192,N_17763);
and U20864 (N_20864,N_18021,N_19809);
or U20865 (N_20865,N_18161,N_17220);
nand U20866 (N_20866,N_17628,N_18255);
xor U20867 (N_20867,N_16720,N_16058);
nand U20868 (N_20868,N_19074,N_16711);
nor U20869 (N_20869,N_16869,N_15926);
xor U20870 (N_20870,N_15313,N_19571);
xor U20871 (N_20871,N_17116,N_19548);
nor U20872 (N_20872,N_16312,N_18004);
nand U20873 (N_20873,N_17458,N_17398);
xnor U20874 (N_20874,N_19959,N_15828);
and U20875 (N_20875,N_17013,N_19553);
and U20876 (N_20876,N_16664,N_16230);
nand U20877 (N_20877,N_18886,N_16972);
nand U20878 (N_20878,N_15775,N_17892);
and U20879 (N_20879,N_17009,N_16566);
nor U20880 (N_20880,N_18677,N_18353);
or U20881 (N_20881,N_15113,N_19914);
nor U20882 (N_20882,N_19682,N_16806);
and U20883 (N_20883,N_17515,N_16056);
xor U20884 (N_20884,N_18045,N_15330);
xnor U20885 (N_20885,N_18965,N_16456);
or U20886 (N_20886,N_15407,N_19263);
or U20887 (N_20887,N_18526,N_15132);
nor U20888 (N_20888,N_19382,N_18396);
nand U20889 (N_20889,N_18265,N_16992);
xnor U20890 (N_20890,N_17306,N_19131);
and U20891 (N_20891,N_16744,N_17981);
and U20892 (N_20892,N_18332,N_17784);
nor U20893 (N_20893,N_15351,N_18933);
nand U20894 (N_20894,N_15819,N_15784);
xor U20895 (N_20895,N_17901,N_18909);
or U20896 (N_20896,N_17119,N_15945);
xnor U20897 (N_20897,N_16515,N_19877);
xor U20898 (N_20898,N_19309,N_15119);
and U20899 (N_20899,N_17745,N_15592);
or U20900 (N_20900,N_18486,N_17824);
nor U20901 (N_20901,N_16773,N_16130);
xnor U20902 (N_20902,N_15406,N_19473);
xnor U20903 (N_20903,N_17143,N_19961);
nor U20904 (N_20904,N_18114,N_15293);
nor U20905 (N_20905,N_16190,N_16020);
xor U20906 (N_20906,N_19267,N_18401);
or U20907 (N_20907,N_15913,N_19038);
nor U20908 (N_20908,N_17010,N_18324);
xnor U20909 (N_20909,N_17975,N_17117);
or U20910 (N_20910,N_18788,N_15814);
nor U20911 (N_20911,N_15864,N_19361);
xor U20912 (N_20912,N_16956,N_18797);
nand U20913 (N_20913,N_17793,N_18046);
or U20914 (N_20914,N_17118,N_17603);
xor U20915 (N_20915,N_15488,N_18993);
nand U20916 (N_20916,N_17836,N_18478);
nand U20917 (N_20917,N_15656,N_18911);
or U20918 (N_20918,N_18292,N_15195);
nor U20919 (N_20919,N_18685,N_15024);
nand U20920 (N_20920,N_17346,N_17531);
or U20921 (N_20921,N_17319,N_15740);
xnor U20922 (N_20922,N_15354,N_17561);
or U20923 (N_20923,N_16377,N_18730);
or U20924 (N_20924,N_18589,N_19887);
xor U20925 (N_20925,N_16199,N_18887);
xor U20926 (N_20926,N_15283,N_19261);
xor U20927 (N_20927,N_16672,N_15938);
xnor U20928 (N_20928,N_18845,N_16065);
xnor U20929 (N_20929,N_17428,N_17021);
nor U20930 (N_20930,N_17552,N_19171);
and U20931 (N_20931,N_19452,N_17829);
and U20932 (N_20932,N_19831,N_17067);
and U20933 (N_20933,N_16866,N_15487);
nor U20934 (N_20934,N_17085,N_15385);
nor U20935 (N_20935,N_16271,N_15193);
nand U20936 (N_20936,N_15895,N_15339);
and U20937 (N_20937,N_15059,N_16095);
xor U20938 (N_20938,N_18284,N_16841);
and U20939 (N_20939,N_15868,N_17455);
nand U20940 (N_20940,N_17397,N_18680);
xnor U20941 (N_20941,N_16138,N_19319);
and U20942 (N_20942,N_17590,N_17298);
and U20943 (N_20943,N_19663,N_15235);
xor U20944 (N_20944,N_16276,N_18080);
or U20945 (N_20945,N_15825,N_16937);
or U20946 (N_20946,N_18314,N_18022);
or U20947 (N_20947,N_17737,N_15708);
xor U20948 (N_20948,N_17720,N_15823);
nor U20949 (N_20949,N_18259,N_16650);
or U20950 (N_20950,N_19192,N_17866);
or U20951 (N_20951,N_19627,N_19984);
or U20952 (N_20952,N_19794,N_19468);
xor U20953 (N_20953,N_16444,N_16352);
and U20954 (N_20954,N_15252,N_17040);
nor U20955 (N_20955,N_16437,N_19093);
nor U20956 (N_20956,N_16926,N_17434);
nor U20957 (N_20957,N_17002,N_15741);
nor U20958 (N_20958,N_17813,N_15111);
nor U20959 (N_20959,N_16752,N_16055);
and U20960 (N_20960,N_15869,N_17110);
nand U20961 (N_20961,N_18690,N_19478);
nor U20962 (N_20962,N_15216,N_15054);
nand U20963 (N_20963,N_18492,N_16093);
nor U20964 (N_20964,N_17305,N_17022);
or U20965 (N_20965,N_18125,N_16450);
xnor U20966 (N_20966,N_15572,N_17891);
xnor U20967 (N_20967,N_16850,N_19859);
nor U20968 (N_20968,N_19500,N_15494);
and U20969 (N_20969,N_15911,N_18059);
xor U20970 (N_20970,N_17635,N_15835);
nand U20971 (N_20971,N_19510,N_15482);
nor U20972 (N_20972,N_16551,N_19477);
nand U20973 (N_20973,N_19288,N_17566);
nand U20974 (N_20974,N_15131,N_15697);
or U20975 (N_20975,N_19952,N_16446);
and U20976 (N_20976,N_18201,N_17225);
and U20977 (N_20977,N_17945,N_15029);
xor U20978 (N_20978,N_15585,N_17482);
and U20979 (N_20979,N_17581,N_16653);
and U20980 (N_20980,N_15197,N_18559);
and U20981 (N_20981,N_18501,N_15241);
nand U20982 (N_20982,N_18988,N_18126);
nor U20983 (N_20983,N_15309,N_18381);
or U20984 (N_20984,N_16247,N_19325);
nor U20985 (N_20985,N_18429,N_19070);
and U20986 (N_20986,N_19741,N_19230);
xnor U20987 (N_20987,N_15065,N_15277);
nor U20988 (N_20988,N_18953,N_19840);
xor U20989 (N_20989,N_17988,N_18294);
or U20990 (N_20990,N_19265,N_15714);
nor U20991 (N_20991,N_17907,N_18927);
xnor U20992 (N_20992,N_18391,N_18703);
or U20993 (N_20993,N_17496,N_15846);
xnor U20994 (N_20994,N_17972,N_18111);
or U20995 (N_20995,N_18264,N_16975);
nor U20996 (N_20996,N_15454,N_16380);
and U20997 (N_20997,N_18614,N_17127);
nor U20998 (N_20998,N_16481,N_15161);
nand U20999 (N_20999,N_19683,N_16660);
and U21000 (N_21000,N_18561,N_19607);
xor U21001 (N_21001,N_15222,N_16965);
and U21002 (N_21002,N_19549,N_18238);
nand U21003 (N_21003,N_16461,N_19425);
or U21004 (N_21004,N_16575,N_15364);
or U21005 (N_21005,N_18372,N_16546);
nor U21006 (N_21006,N_15308,N_18898);
nand U21007 (N_21007,N_18490,N_16554);
and U21008 (N_21008,N_19157,N_18137);
and U21009 (N_21009,N_19913,N_16294);
xor U21010 (N_21010,N_19320,N_18889);
xor U21011 (N_21011,N_17194,N_16643);
and U21012 (N_21012,N_17415,N_19475);
nand U21013 (N_21013,N_15422,N_18936);
xnor U21014 (N_21014,N_15361,N_15575);
nor U21015 (N_21015,N_16313,N_16244);
and U21016 (N_21016,N_16060,N_15386);
and U21017 (N_21017,N_18064,N_18778);
or U21018 (N_21018,N_15129,N_17074);
nor U21019 (N_21019,N_15280,N_16047);
nand U21020 (N_21020,N_18057,N_16652);
nand U21021 (N_21021,N_19400,N_16597);
and U21022 (N_21022,N_18968,N_19818);
nand U21023 (N_21023,N_15105,N_15415);
or U21024 (N_21024,N_15651,N_18465);
nand U21025 (N_21025,N_15573,N_18299);
and U21026 (N_21026,N_17699,N_18669);
and U21027 (N_21027,N_18853,N_16012);
and U21028 (N_21028,N_15988,N_19421);
nand U21029 (N_21029,N_16438,N_19161);
or U21030 (N_21030,N_16106,N_18280);
nor U21031 (N_21031,N_19252,N_15542);
nor U21032 (N_21032,N_18425,N_15301);
and U21033 (N_21033,N_19014,N_16157);
nor U21034 (N_21034,N_16270,N_18442);
xnor U21035 (N_21035,N_19434,N_17575);
nand U21036 (N_21036,N_16818,N_16816);
and U21037 (N_21037,N_15242,N_17048);
nand U21038 (N_21038,N_17727,N_15947);
and U21039 (N_21039,N_16414,N_16820);
nor U21040 (N_21040,N_18996,N_15514);
nor U21041 (N_21041,N_15586,N_15076);
nor U21042 (N_21042,N_15646,N_18208);
and U21043 (N_21043,N_17885,N_19407);
or U21044 (N_21044,N_15873,N_16236);
nor U21045 (N_21045,N_16176,N_15365);
and U21046 (N_21046,N_19145,N_17686);
or U21047 (N_21047,N_15769,N_19560);
nand U21048 (N_21048,N_19096,N_16784);
and U21049 (N_21049,N_19438,N_19110);
nor U21050 (N_21050,N_18510,N_15033);
and U21051 (N_21051,N_18434,N_18307);
nor U21052 (N_21052,N_19414,N_16219);
xnor U21053 (N_21053,N_18471,N_18240);
xnor U21054 (N_21054,N_16283,N_16126);
xor U21055 (N_21055,N_19931,N_19279);
nor U21056 (N_21056,N_16805,N_18168);
and U21057 (N_21057,N_16121,N_19286);
nand U21058 (N_21058,N_18028,N_17138);
and U21059 (N_21059,N_18958,N_16917);
and U21060 (N_21060,N_19291,N_17882);
and U21061 (N_21061,N_16788,N_16924);
xor U21062 (N_21062,N_19253,N_15527);
xnor U21063 (N_21063,N_18724,N_19584);
nor U21064 (N_21064,N_18099,N_17338);
nand U21065 (N_21065,N_18791,N_16936);
nand U21066 (N_21066,N_16864,N_19874);
xnor U21067 (N_21067,N_15549,N_19232);
nor U21068 (N_21068,N_19150,N_19629);
xnor U21069 (N_21069,N_17807,N_16488);
nand U21070 (N_21070,N_19076,N_18268);
nand U21071 (N_21071,N_16852,N_16649);
nand U21072 (N_21072,N_15291,N_15765);
and U21073 (N_21073,N_17265,N_17260);
or U21074 (N_21074,N_19033,N_18991);
or U21075 (N_21075,N_16406,N_19067);
nand U21076 (N_21076,N_18154,N_16091);
nor U21077 (N_21077,N_17198,N_17562);
nand U21078 (N_21078,N_16550,N_17296);
xor U21079 (N_21079,N_17214,N_19474);
xor U21080 (N_21080,N_17241,N_15483);
xnor U21081 (N_21081,N_19921,N_17303);
nor U21082 (N_21082,N_18960,N_18275);
and U21083 (N_21083,N_16402,N_17637);
and U21084 (N_21084,N_18866,N_17718);
and U21085 (N_21085,N_19883,N_16214);
nand U21086 (N_21086,N_16774,N_15368);
xor U21087 (N_21087,N_18974,N_15435);
nor U21088 (N_21088,N_19112,N_15704);
and U21089 (N_21089,N_15017,N_16398);
nand U21090 (N_21090,N_19390,N_17001);
nand U21091 (N_21091,N_15536,N_15773);
xnor U21092 (N_21092,N_18821,N_17691);
xor U21093 (N_21093,N_19292,N_18631);
xnor U21094 (N_21094,N_16817,N_15008);
or U21095 (N_21095,N_17464,N_15358);
xnor U21096 (N_21096,N_17446,N_19118);
nand U21097 (N_21097,N_15084,N_19550);
and U21098 (N_21098,N_18427,N_18838);
and U21099 (N_21099,N_18867,N_17527);
or U21100 (N_21100,N_16458,N_18036);
nand U21101 (N_21101,N_17234,N_18515);
nand U21102 (N_21102,N_19547,N_18545);
xnor U21103 (N_21103,N_16477,N_15824);
nand U21104 (N_21104,N_17723,N_18512);
nor U21105 (N_21105,N_15613,N_15163);
and U21106 (N_21106,N_17726,N_16883);
and U21107 (N_21107,N_15085,N_17043);
nand U21108 (N_21108,N_17014,N_19134);
xnor U21109 (N_21109,N_19799,N_19704);
and U21110 (N_21110,N_16173,N_16240);
nor U21111 (N_21111,N_18335,N_16495);
xnor U21112 (N_21112,N_19410,N_16394);
xor U21113 (N_21113,N_17316,N_16530);
or U21114 (N_21114,N_15263,N_17732);
and U21115 (N_21115,N_18213,N_19019);
and U21116 (N_21116,N_19081,N_16625);
xnor U21117 (N_21117,N_16146,N_17328);
nand U21118 (N_21118,N_17171,N_19179);
and U21119 (N_21119,N_19327,N_19703);
xor U21120 (N_21120,N_15971,N_15918);
xnor U21121 (N_21121,N_15234,N_15116);
nor U21122 (N_21122,N_16309,N_19211);
or U21123 (N_21123,N_15670,N_17189);
nand U21124 (N_21124,N_17493,N_19798);
and U21125 (N_21125,N_16242,N_19040);
nand U21126 (N_21126,N_16253,N_16748);
nor U21127 (N_21127,N_15506,N_17697);
nor U21128 (N_21128,N_15042,N_19995);
or U21129 (N_21129,N_18952,N_16842);
and U21130 (N_21130,N_18141,N_15803);
xnor U21131 (N_21131,N_16761,N_16539);
xnor U21132 (N_21132,N_18027,N_19125);
nand U21133 (N_21133,N_17271,N_16658);
nand U21134 (N_21134,N_17717,N_18961);
nor U21135 (N_21135,N_19912,N_18860);
nor U21136 (N_21136,N_18450,N_16089);
nand U21137 (N_21137,N_17097,N_15345);
nor U21138 (N_21138,N_15251,N_19583);
nand U21139 (N_21139,N_15476,N_15204);
nand U21140 (N_21140,N_18166,N_15620);
and U21141 (N_21141,N_15298,N_15893);
or U21142 (N_21142,N_16591,N_19711);
or U21143 (N_21143,N_19371,N_15510);
nand U21144 (N_21144,N_19197,N_17588);
or U21145 (N_21145,N_19624,N_18751);
or U21146 (N_21146,N_16512,N_18749);
xnor U21147 (N_21147,N_18252,N_15856);
xor U21148 (N_21148,N_17160,N_19980);
nand U21149 (N_21149,N_19234,N_15598);
and U21150 (N_21150,N_17460,N_17405);
nand U21151 (N_21151,N_17743,N_19841);
nand U21152 (N_21152,N_18340,N_18042);
and U21153 (N_21153,N_18619,N_18766);
nor U21154 (N_21154,N_19135,N_15974);
xnor U21155 (N_21155,N_15063,N_19556);
or U21156 (N_21156,N_17147,N_15212);
xor U21157 (N_21157,N_17209,N_19133);
or U21158 (N_21158,N_16657,N_16522);
and U21159 (N_21159,N_19970,N_15055);
xnor U21160 (N_21160,N_16631,N_18039);
and U21161 (N_21161,N_17513,N_16889);
nand U21162 (N_21162,N_15282,N_19653);
xnor U21163 (N_21163,N_15944,N_15977);
or U21164 (N_21164,N_16463,N_19807);
and U21165 (N_21165,N_15884,N_16733);
and U21166 (N_21166,N_18970,N_19238);
or U21167 (N_21167,N_15610,N_16133);
nor U21168 (N_21168,N_16742,N_19882);
or U21169 (N_21169,N_17281,N_15629);
or U21170 (N_21170,N_15207,N_18523);
nor U21171 (N_21171,N_17318,N_17565);
and U21172 (N_21172,N_18816,N_18667);
nand U21173 (N_21173,N_18404,N_16547);
and U21174 (N_21174,N_15617,N_16957);
nor U21175 (N_21175,N_17408,N_17626);
xor U21176 (N_21176,N_19724,N_16935);
xor U21177 (N_21177,N_16198,N_19634);
xnor U21178 (N_21178,N_19020,N_19728);
xor U21179 (N_21179,N_19387,N_15798);
or U21180 (N_21180,N_18305,N_15086);
nor U21181 (N_21181,N_16479,N_15056);
or U21182 (N_21182,N_16897,N_15957);
xor U21183 (N_21183,N_16086,N_16536);
nor U21184 (N_21184,N_19339,N_19097);
and U21185 (N_21185,N_19391,N_16635);
xnor U21186 (N_21186,N_15324,N_17237);
or U21187 (N_21187,N_19330,N_15411);
and U21188 (N_21188,N_17353,N_17424);
and U21189 (N_21189,N_16217,N_19878);
and U21190 (N_21190,N_15323,N_16117);
and U21191 (N_21191,N_16988,N_15182);
xnor U21192 (N_21192,N_17862,N_17036);
nor U21193 (N_21193,N_15185,N_19717);
nor U21194 (N_21194,N_16186,N_16853);
and U21195 (N_21195,N_19411,N_15191);
nand U21196 (N_21196,N_19496,N_15546);
nand U21197 (N_21197,N_19212,N_16717);
or U21198 (N_21198,N_19716,N_17947);
nor U21199 (N_21199,N_15805,N_15341);
nand U21200 (N_21200,N_18336,N_15464);
or U21201 (N_21201,N_17187,N_18814);
and U21202 (N_21202,N_19957,N_19808);
and U21203 (N_21203,N_18005,N_17203);
and U21204 (N_21204,N_19127,N_19731);
or U21205 (N_21205,N_17454,N_19896);
xor U21206 (N_21206,N_15940,N_16415);
and U21207 (N_21207,N_18190,N_15716);
and U21208 (N_21208,N_16079,N_18320);
and U21209 (N_21209,N_18354,N_17838);
nor U21210 (N_21210,N_18083,N_16310);
nand U21211 (N_21211,N_17245,N_19852);
xor U21212 (N_21212,N_15087,N_15285);
xnor U21213 (N_21213,N_17312,N_17710);
and U21214 (N_21214,N_19397,N_15569);
nor U21215 (N_21215,N_19082,N_17128);
xor U21216 (N_21216,N_17326,N_16118);
and U21217 (N_21217,N_18089,N_18764);
and U21218 (N_21218,N_18348,N_18610);
and U21219 (N_21219,N_15051,N_17444);
and U21220 (N_21220,N_19743,N_17102);
and U21221 (N_21221,N_17399,N_17705);
and U21222 (N_21222,N_17191,N_17058);
or U21223 (N_21223,N_17687,N_18225);
xor U21224 (N_21224,N_15124,N_17967);
or U21225 (N_21225,N_18174,N_17752);
and U21226 (N_21226,N_18548,N_15544);
nand U21227 (N_21227,N_17413,N_19137);
xnor U21228 (N_21228,N_19412,N_19384);
or U21229 (N_21229,N_15436,N_18695);
or U21230 (N_21230,N_19544,N_19804);
or U21231 (N_21231,N_15533,N_15266);
nor U21232 (N_21232,N_18482,N_16335);
and U21233 (N_21233,N_17529,N_17049);
xor U21234 (N_21234,N_18670,N_17957);
nor U21235 (N_21235,N_15676,N_16725);
or U21236 (N_21236,N_18347,N_17853);
xor U21237 (N_21237,N_15602,N_19645);
and U21238 (N_21238,N_15817,N_19462);
xor U21239 (N_21239,N_19045,N_17835);
xor U21240 (N_21240,N_18163,N_18678);
nor U21241 (N_21241,N_16436,N_19239);
xor U21242 (N_21242,N_15667,N_19953);
and U21243 (N_21243,N_17548,N_19641);
nor U21244 (N_21244,N_17676,N_17367);
nor U21245 (N_21245,N_17696,N_17407);
or U21246 (N_21246,N_16578,N_19236);
xor U21247 (N_21247,N_18507,N_19523);
nand U21248 (N_21248,N_18880,N_18811);
or U21249 (N_21249,N_17436,N_17065);
or U21250 (N_21250,N_18407,N_19424);
or U21251 (N_21251,N_16933,N_17053);
nand U21252 (N_21252,N_17329,N_15451);
nand U21253 (N_21253,N_16976,N_16614);
xor U21254 (N_21254,N_18494,N_16165);
or U21255 (N_21255,N_18910,N_15290);
xnor U21256 (N_21256,N_19077,N_15493);
nor U21257 (N_21257,N_16765,N_18630);
nand U21258 (N_21258,N_18504,N_17321);
or U21259 (N_21259,N_17254,N_16822);
nand U21260 (N_21260,N_18319,N_17663);
nor U21261 (N_21261,N_18805,N_19243);
and U21262 (N_21262,N_18949,N_17359);
nor U21263 (N_21263,N_17964,N_15831);
and U21264 (N_21264,N_17843,N_18637);
nor U21265 (N_21265,N_16351,N_19723);
nand U21266 (N_21266,N_18738,N_18487);
or U21267 (N_21267,N_15079,N_19218);
or U21268 (N_21268,N_17740,N_18366);
or U21269 (N_21269,N_19409,N_17771);
xor U21270 (N_21270,N_16031,N_19987);
or U21271 (N_21271,N_18869,N_15749);
or U21272 (N_21272,N_15660,N_19545);
nand U21273 (N_21273,N_15474,N_18820);
and U21274 (N_21274,N_16705,N_18058);
nor U21275 (N_21275,N_18903,N_16008);
nand U21276 (N_21276,N_15458,N_16407);
or U21277 (N_21277,N_17848,N_17196);
nand U21278 (N_21278,N_18608,N_17052);
nand U21279 (N_21279,N_17015,N_18337);
xor U21280 (N_21280,N_17805,N_18394);
or U21281 (N_21281,N_19676,N_15637);
and U21282 (N_21282,N_18928,N_17941);
xor U21283 (N_21283,N_19681,N_16609);
xor U21284 (N_21284,N_19595,N_17653);
and U21285 (N_21285,N_16905,N_15418);
xnor U21286 (N_21286,N_19152,N_19979);
and U21287 (N_21287,N_18851,N_18879);
and U21288 (N_21288,N_18563,N_16388);
nand U21289 (N_21289,N_15122,N_15865);
nor U21290 (N_21290,N_19790,N_17033);
nand U21291 (N_21291,N_19875,N_18373);
or U21292 (N_21292,N_15081,N_18436);
xnor U21293 (N_21293,N_17185,N_15861);
nor U21294 (N_21294,N_18591,N_15900);
and U21295 (N_21295,N_15915,N_18071);
xor U21296 (N_21296,N_16289,N_19486);
or U21297 (N_21297,N_16944,N_19465);
or U21298 (N_21298,N_16738,N_18530);
and U21299 (N_21299,N_15755,N_16796);
nor U21300 (N_21300,N_19842,N_15810);
nand U21301 (N_21301,N_15496,N_16039);
xor U21302 (N_21302,N_19649,N_17545);
xnor U21303 (N_21303,N_16159,N_15993);
nor U21304 (N_21304,N_19535,N_17435);
and U21305 (N_21305,N_18437,N_18131);
and U21306 (N_21306,N_18128,N_18192);
nor U21307 (N_21307,N_17927,N_18713);
nand U21308 (N_21308,N_19013,N_17894);
or U21309 (N_21309,N_16120,N_17979);
and U21310 (N_21310,N_16586,N_18343);
nand U21311 (N_21311,N_16524,N_15073);
xnor U21312 (N_21312,N_17613,N_19193);
nand U21313 (N_21313,N_17921,N_19120);
or U21314 (N_21314,N_19884,N_18067);
nor U21315 (N_21315,N_18663,N_15416);
and U21316 (N_21316,N_18948,N_19919);
xor U21317 (N_21317,N_16224,N_18905);
xnor U21318 (N_21318,N_16017,N_17089);
xor U21319 (N_21319,N_16492,N_17169);
nand U21320 (N_21320,N_18061,N_19606);
or U21321 (N_21321,N_18195,N_19366);
or U21322 (N_21322,N_17086,N_16304);
xor U21323 (N_21323,N_16827,N_16718);
xnor U21324 (N_21324,N_15738,N_15094);
or U21325 (N_21325,N_16562,N_19721);
or U21326 (N_21326,N_17020,N_17273);
nand U21327 (N_21327,N_18379,N_19567);
and U21328 (N_21328,N_15468,N_19042);
nor U21329 (N_21329,N_18312,N_19719);
nor U21330 (N_21330,N_18789,N_17977);
nor U21331 (N_21331,N_18629,N_18410);
and U21332 (N_21332,N_19769,N_19392);
xnor U21333 (N_21333,N_17087,N_19602);
nand U21334 (N_21334,N_17108,N_18653);
nand U21335 (N_21335,N_16830,N_17463);
or U21336 (N_21336,N_19208,N_18999);
and U21337 (N_21337,N_16665,N_17439);
nor U21338 (N_21338,N_18387,N_17096);
nand U21339 (N_21339,N_17804,N_18694);
and U21340 (N_21340,N_15377,N_18611);
nor U21341 (N_21341,N_16301,N_17971);
and U21342 (N_21342,N_16496,N_17591);
xor U21343 (N_21343,N_17636,N_15844);
nor U21344 (N_21344,N_16497,N_18313);
or U21345 (N_21345,N_16064,N_16519);
nand U21346 (N_21346,N_19294,N_19317);
nand U21347 (N_21347,N_15608,N_19986);
xor U21348 (N_21348,N_15540,N_15567);
nor U21349 (N_21349,N_18287,N_19054);
nor U21350 (N_21350,N_16372,N_16751);
or U21351 (N_21351,N_16455,N_16778);
nand U21352 (N_21352,N_19617,N_16206);
nand U21353 (N_21353,N_19738,N_19458);
nor U21354 (N_21354,N_16603,N_17459);
nand U21355 (N_21355,N_19920,N_16025);
or U21356 (N_21356,N_15034,N_19285);
and U21357 (N_21357,N_16849,N_16559);
nand U21358 (N_21358,N_19604,N_15928);
or U21359 (N_21359,N_17729,N_16508);
and U21360 (N_21360,N_15822,N_16598);
and U21361 (N_21361,N_19420,N_18597);
nand U21362 (N_21362,N_16707,N_18704);
nor U21363 (N_21363,N_15220,N_19386);
nor U21364 (N_21364,N_15816,N_18129);
or U21365 (N_21365,N_16258,N_15231);
nor U21366 (N_21366,N_15737,N_16107);
nand U21367 (N_21367,N_18010,N_19506);
and U21368 (N_21368,N_15942,N_17559);
and U21369 (N_21369,N_18286,N_17880);
and U21370 (N_21370,N_16170,N_15329);
or U21371 (N_21371,N_16142,N_17094);
xnor U21372 (N_21372,N_18247,N_19949);
nand U21373 (N_21373,N_17308,N_17246);
nor U21374 (N_21374,N_19911,N_17911);
nand U21375 (N_21375,N_15811,N_16901);
and U21376 (N_21376,N_16241,N_18220);
nand U21377 (N_21377,N_16676,N_17873);
nor U21378 (N_21378,N_18964,N_18919);
or U21379 (N_21379,N_18297,N_17055);
nand U21380 (N_21380,N_17847,N_15967);
xor U21381 (N_21381,N_18920,N_16535);
nor U21382 (N_21382,N_18145,N_19215);
nand U21383 (N_21383,N_18439,N_18109);
xnor U21384 (N_21384,N_15157,N_17059);
xnor U21385 (N_21385,N_17510,N_17294);
or U21386 (N_21386,N_18525,N_17779);
xor U21387 (N_21387,N_17270,N_19610);
nand U21388 (N_21388,N_19695,N_15526);
nor U21389 (N_21389,N_19754,N_19188);
or U21390 (N_21390,N_16447,N_15352);
nand U21391 (N_21391,N_17320,N_15453);
and U21392 (N_21392,N_18171,N_18078);
or U21393 (N_21393,N_17621,N_17602);
or U21394 (N_21394,N_18858,N_17327);
or U21395 (N_21395,N_18533,N_15706);
or U21396 (N_21396,N_16114,N_19439);
nand U21397 (N_21397,N_18834,N_15791);
or U21398 (N_21398,N_17054,N_16057);
nor U21399 (N_21399,N_16687,N_17340);
xor U21400 (N_21400,N_16115,N_16172);
nor U21401 (N_21401,N_18729,N_19380);
and U21402 (N_21402,N_15955,N_17310);
xnor U21403 (N_21403,N_15400,N_17760);
nor U21404 (N_21404,N_18251,N_19932);
nand U21405 (N_21405,N_18718,N_19760);
nand U21406 (N_21406,N_16896,N_16906);
nor U21407 (N_21407,N_16839,N_17655);
xor U21408 (N_21408,N_17656,N_15744);
or U21409 (N_21409,N_16914,N_15037);
and U21410 (N_21410,N_17177,N_18325);
nand U21411 (N_21411,N_17948,N_15966);
nor U21412 (N_21412,N_15470,N_18049);
xnor U21413 (N_21413,N_16740,N_18477);
and U21414 (N_21414,N_15356,N_17826);
or U21415 (N_21415,N_17499,N_15690);
nor U21416 (N_21416,N_19751,N_19454);
xnor U21417 (N_21417,N_18892,N_16048);
nor U21418 (N_21418,N_19036,N_16267);
and U21419 (N_21419,N_18555,N_15943);
nor U21420 (N_21420,N_17860,N_18520);
nor U21421 (N_21421,N_15077,N_15826);
xor U21422 (N_21422,N_15639,N_16758);
nor U21423 (N_21423,N_19598,N_19173);
and U21424 (N_21424,N_16953,N_17795);
nand U21425 (N_21425,N_16895,N_18671);
or U21426 (N_21426,N_18861,N_18048);
and U21427 (N_21427,N_17830,N_18986);
nand U21428 (N_21428,N_16698,N_17380);
xnor U21429 (N_21429,N_19770,N_17028);
or U21430 (N_21430,N_15648,N_18350);
nor U21431 (N_21431,N_18445,N_19379);
or U21432 (N_21432,N_17420,N_16781);
nand U21433 (N_21433,N_18648,N_16745);
and U21434 (N_21434,N_18660,N_19457);
or U21435 (N_21435,N_16893,N_19156);
and U21436 (N_21436,N_17942,N_16876);
and U21437 (N_21437,N_15657,N_15457);
nor U21438 (N_21438,N_19170,N_16968);
and U21439 (N_21439,N_15715,N_16131);
nor U21440 (N_21440,N_17445,N_17692);
and U21441 (N_21441,N_18809,N_15621);
nor U21442 (N_21442,N_18650,N_19503);
xor U21443 (N_21443,N_18377,N_15783);
and U21444 (N_21444,N_15215,N_15420);
nand U21445 (N_21445,N_16621,N_15989);
nor U21446 (N_21446,N_15695,N_15624);
xnor U21447 (N_21447,N_17292,N_19476);
xnor U21448 (N_21448,N_15336,N_19346);
nor U21449 (N_21449,N_19720,N_15978);
nor U21450 (N_21450,N_15781,N_17199);
nor U21451 (N_21451,N_18443,N_17222);
nand U21452 (N_21452,N_18826,N_15735);
and U21453 (N_21453,N_19436,N_19303);
nor U21454 (N_21454,N_16284,N_15597);
nor U21455 (N_21455,N_16286,N_16938);
nand U21456 (N_21456,N_16249,N_16423);
nor U21457 (N_21457,N_17828,N_17134);
nor U21458 (N_21458,N_16641,N_15574);
xnor U21459 (N_21459,N_19034,N_19422);
and U21460 (N_21460,N_17372,N_18431);
nor U21461 (N_21461,N_19873,N_19771);
xnor U21462 (N_21462,N_18344,N_16782);
and U21463 (N_21463,N_15150,N_16370);
xor U21464 (N_21464,N_18835,N_19488);
nor U21465 (N_21465,N_19446,N_15636);
xnor U21466 (N_21466,N_16248,N_17382);
or U21467 (N_21467,N_15164,N_18081);
nand U21468 (N_21468,N_18639,N_18717);
or U21469 (N_21469,N_16421,N_19072);
or U21470 (N_21470,N_16756,N_16666);
xnor U21471 (N_21471,N_19018,N_19219);
nor U21472 (N_21472,N_18481,N_19530);
nand U21473 (N_21473,N_15469,N_15799);
nand U21474 (N_21474,N_16831,N_19588);
nor U21475 (N_21475,N_17193,N_16811);
and U21476 (N_21476,N_18063,N_18187);
and U21477 (N_21477,N_18194,N_18884);
nand U21478 (N_21478,N_18943,N_17627);
and U21479 (N_21479,N_17360,N_15534);
xor U21480 (N_21480,N_17083,N_18983);
nor U21481 (N_21481,N_15500,N_16084);
and U21482 (N_21482,N_18994,N_18657);
and U21483 (N_21483,N_16416,N_17844);
or U21484 (N_21484,N_16531,N_16969);
nor U21485 (N_21485,N_18293,N_19825);
or U21486 (N_21486,N_18093,N_18822);
xnor U21487 (N_21487,N_15423,N_17105);
xor U21488 (N_21488,N_17333,N_16754);
nor U21489 (N_21489,N_15218,N_16080);
nor U21490 (N_21490,N_15014,N_18267);
or U21491 (N_21491,N_19373,N_18209);
and U21492 (N_21492,N_18074,N_15524);
and U21493 (N_21493,N_19342,N_15134);
xnor U21494 (N_21494,N_16538,N_16712);
or U21495 (N_21495,N_18836,N_18662);
nor U21496 (N_21496,N_16422,N_19942);
or U21497 (N_21497,N_18755,N_18356);
xor U21498 (N_21498,N_16581,N_15318);
nor U21499 (N_21499,N_15078,N_15839);
or U21500 (N_21500,N_19678,N_16440);
nor U21501 (N_21501,N_17343,N_18742);
nand U21502 (N_21502,N_15903,N_17236);
and U21503 (N_21503,N_17279,N_18918);
nand U21504 (N_21504,N_19102,N_17748);
nand U21505 (N_21505,N_17782,N_19940);
nand U21506 (N_21506,N_18538,N_18380);
nor U21507 (N_21507,N_19687,N_15649);
or U21508 (N_21508,N_18551,N_15680);
or U21509 (N_21509,N_16802,N_16541);
nand U21510 (N_21510,N_17242,N_17814);
nand U21511 (N_21511,N_15595,N_17401);
nand U21512 (N_21512,N_19539,N_18828);
nor U21513 (N_21513,N_15061,N_19331);
nor U21514 (N_21514,N_18739,N_18116);
or U21515 (N_21515,N_17129,N_19666);
and U21516 (N_21516,N_17511,N_15272);
xnor U21517 (N_21517,N_17818,N_19640);
and U21518 (N_21518,N_19106,N_18120);
xnor U21519 (N_21519,N_17791,N_15921);
and U21520 (N_21520,N_17666,N_18135);
and U21521 (N_21521,N_19435,N_19637);
nor U21522 (N_21522,N_18218,N_18568);
xor U21523 (N_21523,N_16721,N_17773);
nor U21524 (N_21524,N_15745,N_16825);
nor U21525 (N_21525,N_17072,N_15961);
xor U21526 (N_21526,N_15887,N_16619);
nor U21527 (N_21527,N_15214,N_17073);
xnor U21528 (N_21528,N_15100,N_19951);
and U21529 (N_21529,N_19101,N_16277);
nand U21530 (N_21530,N_19324,N_15258);
and U21531 (N_21531,N_15761,N_16381);
nand U21532 (N_21532,N_18088,N_19377);
xor U21533 (N_21533,N_19740,N_19340);
nor U21534 (N_21534,N_19593,N_16994);
nand U21535 (N_21535,N_17161,N_19459);
nor U21536 (N_21536,N_16010,N_19248);
xnor U21537 (N_21537,N_15951,N_18178);
or U21538 (N_21538,N_18518,N_16150);
nor U21539 (N_21539,N_15583,N_17505);
nand U21540 (N_21540,N_15036,N_16182);
xor U21541 (N_21541,N_15130,N_16634);
nor U21542 (N_21542,N_17247,N_18087);
and U21543 (N_21543,N_19216,N_16951);
xnor U21544 (N_21544,N_19483,N_15068);
nand U21545 (N_21545,N_18573,N_19993);
or U21546 (N_21546,N_18355,N_18732);
and U21547 (N_21547,N_15931,N_16262);
and U21548 (N_21548,N_17902,N_17126);
nor U21549 (N_21549,N_15331,N_15815);
and U21550 (N_21550,N_18031,N_15366);
xnor U21551 (N_21551,N_15430,N_18430);
and U21552 (N_21552,N_18474,N_18626);
nand U21553 (N_21553,N_15933,N_16859);
nand U21554 (N_21554,N_19983,N_16124);
and U21555 (N_21555,N_19295,N_18924);
nor U21556 (N_21556,N_16181,N_19370);
xor U21557 (N_21557,N_15827,N_18266);
nor U21558 (N_21558,N_19059,N_17568);
nand U21559 (N_21559,N_15693,N_19000);
nand U21560 (N_21560,N_19166,N_17800);
nand U21561 (N_21561,N_19461,N_15410);
xor U21562 (N_21562,N_17915,N_19027);
or U21563 (N_21563,N_16022,N_16308);
nand U21564 (N_21564,N_17375,N_17598);
or U21565 (N_21565,N_15337,N_19922);
or U21566 (N_21566,N_16540,N_19836);
nand U21567 (N_21567,N_15984,N_18621);
or U21568 (N_21568,N_18256,N_16353);
nor U21569 (N_21569,N_17448,N_15257);
nor U21570 (N_21570,N_16411,N_17387);
xor U21571 (N_21571,N_19854,N_17762);
and U21572 (N_21572,N_19374,N_18754);
nor U21573 (N_21573,N_19521,N_19440);
xnor U21574 (N_21574,N_16599,N_19146);
and U21575 (N_21575,N_15694,N_16786);
nand U21576 (N_21576,N_19638,N_19958);
nor U21577 (N_21577,N_16766,N_15007);
nand U21578 (N_21578,N_17483,N_16983);
nand U21579 (N_21579,N_15380,N_17563);
or U21580 (N_21580,N_17437,N_19289);
nor U21581 (N_21581,N_15722,N_16940);
nand U21582 (N_21582,N_18752,N_19675);
and U21583 (N_21583,N_19050,N_15515);
xnor U21584 (N_21584,N_17491,N_18118);
nor U21585 (N_21585,N_18984,N_18688);
nor U21586 (N_21586,N_15528,N_17224);
xnor U21587 (N_21587,N_15896,N_15739);
nor U21588 (N_21588,N_16345,N_16299);
xnor U21589 (N_21589,N_18542,N_18134);
nand U21590 (N_21590,N_15253,N_19529);
nand U21591 (N_21591,N_18803,N_18998);
xor U21592 (N_21592,N_19631,N_17213);
nand U21593 (N_21593,N_17684,N_19235);
and U21594 (N_21594,N_18572,N_17564);
or U21595 (N_21595,N_19429,N_15144);
nor U21596 (N_21596,N_17986,N_18643);
or U21597 (N_21597,N_19648,N_17526);
nor U21598 (N_21598,N_16347,N_18132);
and U21599 (N_21599,N_16846,N_17173);
nand U21600 (N_21600,N_16272,N_19518);
or U21601 (N_21601,N_15721,N_15908);
or U21602 (N_21602,N_16127,N_19936);
or U21603 (N_21603,N_19764,N_19787);
xor U21604 (N_21604,N_17668,N_18932);
nand U21605 (N_21605,N_18130,N_15460);
nor U21606 (N_21606,N_17695,N_17825);
xor U21607 (N_21607,N_16233,N_15511);
or U21608 (N_21608,N_18409,N_18899);
and U21609 (N_21609,N_15485,N_17115);
nand U21610 (N_21610,N_15999,N_18735);
xnor U21611 (N_21611,N_16633,N_17994);
xor U21612 (N_21612,N_18341,N_18175);
nor U21613 (N_21613,N_15652,N_19857);
nand U21614 (N_21614,N_19647,N_16234);
nor U21615 (N_21615,N_16861,N_15570);
or U21616 (N_21616,N_17610,N_19428);
nor U21617 (N_21617,N_16273,N_15387);
nand U21618 (N_21618,N_17716,N_15591);
nor U21619 (N_21619,N_15187,N_19894);
and U21620 (N_21620,N_18318,N_18495);
nor U21621 (N_21621,N_19062,N_18069);
xor U21622 (N_21622,N_19876,N_15442);
and U21623 (N_21623,N_17895,N_17888);
nor U21624 (N_21624,N_15047,N_16038);
xor U21625 (N_21625,N_18934,N_17365);
xnor U21626 (N_21626,N_17884,N_16354);
nand U21627 (N_21627,N_17506,N_16357);
xor U21628 (N_21628,N_18153,N_16908);
and U21629 (N_21629,N_18056,N_16507);
xor U21630 (N_21630,N_16161,N_19589);
nor U21631 (N_21631,N_17574,N_19214);
nor U21632 (N_21632,N_18199,N_19021);
xor U21633 (N_21633,N_19184,N_16418);
xnor U21634 (N_21634,N_19733,N_19403);
xnor U21635 (N_21635,N_15833,N_17300);
or U21636 (N_21636,N_17253,N_18915);
or U21637 (N_21637,N_15019,N_16679);
nand U21638 (N_21638,N_17172,N_18931);
nand U21639 (N_21639,N_15221,N_18623);
or U21640 (N_21640,N_15325,N_18638);
nor U21641 (N_21641,N_15851,N_19113);
nor U21642 (N_21642,N_19815,N_15800);
or U21643 (N_21643,N_15726,N_16618);
nor U21644 (N_21644,N_15495,N_15669);
nor U21645 (N_21645,N_17751,N_16439);
xnor U21646 (N_21646,N_18977,N_17685);
nor U21647 (N_21647,N_16569,N_17904);
and U21648 (N_21648,N_16103,N_15970);
xor U21649 (N_21649,N_18544,N_19148);
nor U21650 (N_21650,N_17188,N_17898);
and U21651 (N_21651,N_17624,N_16596);
and U21652 (N_21652,N_16743,N_17959);
and U21653 (N_21653,N_15834,N_18859);
xor U21654 (N_21654,N_18003,N_18330);
nand U21655 (N_21655,N_15953,N_16974);
nor U21656 (N_21656,N_19966,N_17400);
and U21657 (N_21657,N_18864,N_19981);
nor U21658 (N_21658,N_17788,N_19463);
nor U21659 (N_21659,N_16628,N_19789);
xnor U21660 (N_21660,N_17811,N_16306);
nor U21661 (N_21661,N_17991,N_16693);
and U21662 (N_21662,N_15026,N_19399);
xnor U21663 (N_21663,N_16984,N_17774);
and U21664 (N_21664,N_19247,N_16934);
nand U21665 (N_21665,N_19688,N_17268);
or U21666 (N_21666,N_16856,N_18574);
xnor U21667 (N_21667,N_17091,N_15424);
nand U21668 (N_21668,N_19690,N_15979);
nor U21669 (N_21669,N_16003,N_16013);
nor U21670 (N_21670,N_15808,N_18509);
xnor U21671 (N_21671,N_17377,N_15889);
or U21672 (N_21672,N_16119,N_18556);
and U21673 (N_21673,N_17850,N_15997);
xor U21674 (N_21674,N_18806,N_19275);
and U21675 (N_21675,N_19814,N_18101);
or U21676 (N_21676,N_15275,N_19336);
or U21677 (N_21677,N_15396,N_15238);
or U21678 (N_21678,N_19909,N_19554);
nor U21679 (N_21679,N_17801,N_19505);
and U21680 (N_21680,N_15172,N_18295);
xor U21681 (N_21681,N_18508,N_17833);
and U21682 (N_21682,N_18506,N_19111);
or U21683 (N_21683,N_16813,N_17910);
or U21684 (N_21684,N_16189,N_16116);
or U21685 (N_21685,N_18323,N_19222);
and U21686 (N_21686,N_18374,N_15162);
xnor U21687 (N_21687,N_19321,N_16040);
or U21688 (N_21688,N_17524,N_19049);
nor U21689 (N_21689,N_18985,N_18908);
and U21690 (N_21690,N_16451,N_15127);
or U21691 (N_21691,N_17063,N_15271);
and U21692 (N_21692,N_15809,N_18232);
and U21693 (N_21693,N_15590,N_18748);
or U21694 (N_21694,N_19599,N_17521);
nand U21695 (N_21695,N_18594,N_16037);
and U21696 (N_21696,N_15002,N_17057);
xnor U21697 (N_21697,N_18872,N_17755);
and U21698 (N_21698,N_16580,N_16417);
or U21699 (N_21699,N_19071,N_19046);
nand U21700 (N_21700,N_17462,N_15930);
xor U21701 (N_21701,N_16011,N_15748);
xor U21702 (N_21702,N_15062,N_17735);
xnor U21703 (N_21703,N_18206,N_15461);
or U21704 (N_21704,N_16136,N_18246);
nand U21705 (N_21705,N_17985,N_18854);
xnor U21706 (N_21706,N_18883,N_16068);
nor U21707 (N_21707,N_16916,N_19316);
nor U21708 (N_21708,N_17796,N_17693);
and U21709 (N_21709,N_18376,N_19572);
xor U21710 (N_21710,N_18102,N_17388);
nand U21711 (N_21711,N_16741,N_16167);
nand U21712 (N_21712,N_19207,N_17283);
nor U21713 (N_21713,N_19432,N_19869);
or U21714 (N_21714,N_17870,N_16082);
nor U21715 (N_21715,N_17792,N_15742);
nand U21716 (N_21716,N_18715,N_17381);
nor U21717 (N_21717,N_16775,N_18155);
xor U21718 (N_21718,N_15932,N_17677);
and U21719 (N_21719,N_16703,N_16494);
xor U21720 (N_21720,N_16268,N_15747);
or U21721 (N_21721,N_18417,N_19190);
or U21722 (N_21722,N_15497,N_18317);
nand U21723 (N_21723,N_18217,N_18885);
nor U21724 (N_21724,N_17369,N_16005);
or U21725 (N_21725,N_15794,N_18223);
xnor U21726 (N_21726,N_17709,N_17579);
nor U21727 (N_21727,N_18480,N_17103);
xnor U21728 (N_21728,N_18815,N_16567);
nor U21729 (N_21729,N_19846,N_17775);
nor U21730 (N_21730,N_18819,N_16884);
and U21731 (N_21731,N_18807,N_19491);
or U21732 (N_21732,N_15419,N_18308);
nand U21733 (N_21733,N_17938,N_17567);
xnor U21734 (N_21734,N_19956,N_19694);
nand U21735 (N_21735,N_17520,N_19088);
nor U21736 (N_21736,N_16278,N_16780);
or U21737 (N_21737,N_18709,N_16123);
nand U21738 (N_21738,N_16348,N_16109);
nor U21739 (N_21739,N_16019,N_18801);
nand U21740 (N_21740,N_17724,N_15801);
nand U21741 (N_21741,N_16303,N_16673);
nand U21742 (N_21742,N_19715,N_19978);
nor U21743 (N_21743,N_15641,N_16445);
and U21744 (N_21744,N_18491,N_16545);
nor U21745 (N_21745,N_15552,N_15841);
nor U21746 (N_21746,N_15254,N_15782);
nor U21747 (N_21747,N_15296,N_17468);
or U21748 (N_21748,N_18122,N_16500);
nor U21749 (N_21749,N_15057,N_17799);
nor U21750 (N_21750,N_19816,N_17081);
xor U21751 (N_21751,N_18878,N_16110);
nor U21752 (N_21752,N_15686,N_19002);
xor U21753 (N_21753,N_19078,N_16995);
nor U21754 (N_21754,N_19023,N_17376);
and U21755 (N_21755,N_17484,N_17277);
nand U21756 (N_21756,N_15792,N_17736);
nor U21757 (N_21757,N_16246,N_19394);
nand U21758 (N_21758,N_19562,N_17050);
or U21759 (N_21759,N_19660,N_15274);
nor U21760 (N_21760,N_15980,N_19899);
and U21761 (N_21761,N_15973,N_19747);
and U21762 (N_21762,N_18627,N_16910);
and U21763 (N_21763,N_15678,N_16410);
or U21764 (N_21764,N_18769,N_16468);
or U21765 (N_21765,N_16099,N_17276);
xnor U21766 (N_21766,N_18360,N_19582);
or U21767 (N_21767,N_16328,N_16919);
xor U21768 (N_21768,N_17682,N_17661);
nor U21769 (N_21769,N_16480,N_15288);
xnor U21770 (N_21770,N_18406,N_18937);
nor U21771 (N_21771,N_16433,N_17512);
or U21772 (N_21772,N_16708,N_15793);
and U21773 (N_21773,N_19555,N_15710);
and U21774 (N_21774,N_19501,N_16979);
and U21775 (N_21775,N_18973,N_19314);
nand U21776 (N_21776,N_16801,N_18760);
nor U21777 (N_21777,N_15001,N_17536);
xor U21778 (N_21778,N_15901,N_19826);
and U21779 (N_21779,N_15000,N_18547);
nor U21780 (N_21780,N_17508,N_16327);
and U21781 (N_21781,N_18414,N_17998);
xor U21782 (N_21782,N_16315,N_15709);
and U21783 (N_21783,N_18580,N_17045);
and U21784 (N_21784,N_18009,N_16454);
nor U21785 (N_21785,N_19697,N_17550);
nand U21786 (N_21786,N_18781,N_17477);
nor U21787 (N_21787,N_18421,N_17647);
nor U21788 (N_21788,N_17228,N_15836);
and U21789 (N_21789,N_16565,N_17142);
or U21790 (N_21790,N_16054,N_19168);
nor U21791 (N_21791,N_18282,N_16682);
or U21792 (N_21792,N_15472,N_17051);
xor U21793 (N_21793,N_18072,N_15845);
nand U21794 (N_21794,N_17342,N_18527);
nand U21795 (N_21795,N_16601,N_16959);
nand U21796 (N_21796,N_17630,N_15307);
nand U21797 (N_21797,N_18321,N_18622);
nor U21798 (N_21798,N_15475,N_18871);
and U21799 (N_21799,N_15643,N_17000);
xor U21800 (N_21800,N_18227,N_19123);
and U21801 (N_21801,N_16855,N_16613);
nor U21802 (N_21802,N_17039,N_17728);
nand U21803 (N_21803,N_19187,N_15727);
and U21804 (N_21804,N_15760,N_16986);
nand U21805 (N_21805,N_16877,N_16259);
xnor U21806 (N_21806,N_19608,N_16939);
and U21807 (N_21807,N_18615,N_17250);
and U21808 (N_21808,N_17518,N_16548);
nand U21809 (N_21809,N_18115,N_18392);
and U21810 (N_21810,N_19888,N_17024);
xnor U21811 (N_21811,N_16692,N_17389);
and U21812 (N_21812,N_19159,N_16719);
xnor U21813 (N_21813,N_17649,N_19702);
nor U21814 (N_21814,N_18001,N_18519);
nor U21815 (N_21815,N_15383,N_19693);
xor U21816 (N_21816,N_18954,N_15359);
nor U21817 (N_21817,N_16408,N_19416);
or U21818 (N_21818,N_17996,N_18978);
nor U21819 (N_21819,N_17939,N_18055);
xor U21820 (N_21820,N_17542,N_19910);
and U21821 (N_21821,N_16732,N_18060);
nand U21822 (N_21822,N_16160,N_15075);
nand U21823 (N_21823,N_16689,N_18881);
and U21824 (N_21824,N_17747,N_18565);
or U21825 (N_21825,N_18913,N_16655);
or U21826 (N_21826,N_15381,N_17164);
nand U21827 (N_21827,N_16642,N_15675);
nor U21828 (N_21828,N_16321,N_17258);
nand U21829 (N_21829,N_18711,N_18339);
and U21830 (N_21830,N_16076,N_16670);
and U21831 (N_21831,N_15991,N_15564);
and U21832 (N_21832,N_19667,N_19242);
nor U21833 (N_21833,N_17480,N_15612);
nand U21834 (N_21834,N_15964,N_16871);
or U21835 (N_21835,N_17928,N_18601);
and U21836 (N_21836,N_16656,N_18419);
nor U21837 (N_21837,N_17200,N_18156);
xor U21838 (N_21838,N_18462,N_16930);
nand U21839 (N_21839,N_19915,N_16824);
nand U21840 (N_21840,N_15599,N_16941);
or U21841 (N_21841,N_18413,N_19635);
nor U21842 (N_21842,N_17165,N_17842);
nor U21843 (N_21843,N_16810,N_15099);
or U21844 (N_21844,N_17992,N_19618);
nand U21845 (N_21845,N_16155,N_15674);
nand U21846 (N_21846,N_19621,N_15184);
xnor U21847 (N_21847,N_19124,N_15326);
or U21848 (N_21848,N_15778,N_17221);
or U21849 (N_21849,N_18345,N_15440);
nand U21850 (N_21850,N_16487,N_18065);
nand U21851 (N_21851,N_16185,N_19990);
xor U21852 (N_21852,N_16484,N_17106);
nor U21853 (N_21853,N_18334,N_17363);
or U21854 (N_21854,N_19871,N_19526);
nor U21855 (N_21855,N_19865,N_19095);
nand U21856 (N_21856,N_19924,N_17711);
or U21857 (N_21857,N_16223,N_18966);
nand U21858 (N_21858,N_17362,N_18543);
and U21859 (N_21859,N_15509,N_18342);
nor U21860 (N_21860,N_15631,N_19644);
or U21861 (N_21861,N_15240,N_19144);
and U21862 (N_21862,N_16009,N_16695);
xnor U21863 (N_21863,N_16553,N_16156);
and U21864 (N_21864,N_17252,N_18634);
nand U21865 (N_21865,N_18152,N_15995);
nor U21866 (N_21866,N_18831,N_18896);
xor U21867 (N_21867,N_19254,N_18576);
or U21868 (N_21868,N_19007,N_19822);
or U21869 (N_21869,N_17151,N_18073);
xor U21870 (N_21870,N_18123,N_18734);
nor U21871 (N_21871,N_18962,N_16275);
or U21872 (N_21872,N_16814,N_18395);
xnor U21873 (N_21873,N_16432,N_15555);
xor U21874 (N_21874,N_15371,N_19323);
nor U21875 (N_21875,N_19778,N_16690);
nor U21876 (N_21876,N_16731,N_19796);
or U21877 (N_21877,N_17355,N_17654);
and U21878 (N_21878,N_17582,N_16269);
nor U21879 (N_21879,N_18632,N_18775);
nand U21880 (N_21880,N_18505,N_17204);
nor U21881 (N_21881,N_16835,N_18368);
or U21882 (N_21882,N_19976,N_18204);
or U21883 (N_21883,N_15200,N_19821);
or U21884 (N_21884,N_19730,N_16420);
or U21885 (N_21885,N_19359,N_16990);
xor U21886 (N_21886,N_17937,N_17534);
or U21887 (N_21887,N_16098,N_17658);
nor U21888 (N_21888,N_17681,N_16798);
xnor U21889 (N_21889,N_18651,N_19048);
xnor U21890 (N_21890,N_18034,N_15975);
nand U21891 (N_21891,N_18035,N_19213);
nor U21892 (N_21892,N_16425,N_16659);
xor U21893 (N_21893,N_16654,N_16971);
nand U21894 (N_21894,N_15982,N_15571);
nand U21895 (N_21895,N_18921,N_16998);
or U21896 (N_21896,N_18843,N_19534);
and U21897 (N_21897,N_16175,N_17205);
nand U21898 (N_21898,N_19891,N_17953);
or U21899 (N_21899,N_19680,N_18258);
nor U21900 (N_21900,N_15996,N_19226);
or U21901 (N_21901,N_15849,N_17678);
and U21902 (N_21902,N_16542,N_19160);
nand U21903 (N_21903,N_18398,N_16999);
or U21904 (N_21904,N_15334,N_16320);
nor U21905 (N_21905,N_18100,N_15481);
or U21906 (N_21906,N_19024,N_15746);
nand U21907 (N_21907,N_16018,N_17612);
nor U21908 (N_21908,N_19823,N_17394);
or U21909 (N_21909,N_15340,N_18113);
nor U21910 (N_21910,N_15785,N_15541);
xor U21911 (N_21911,N_18271,N_18550);
nor U21912 (N_21912,N_15897,N_15615);
nand U21913 (N_21913,N_17827,N_16570);
nor U21914 (N_21914,N_17989,N_16424);
nand U21915 (N_21915,N_19367,N_18641);
nor U21916 (N_21916,N_19907,N_16379);
xor U21917 (N_21917,N_15972,N_15232);
nor U21918 (N_21918,N_18793,N_18411);
nor U21919 (N_21919,N_18770,N_16029);
and U21920 (N_21920,N_17810,N_16210);
and U21921 (N_21921,N_15840,N_17485);
xor U21922 (N_21922,N_18971,N_18173);
xor U21923 (N_21923,N_16947,N_18562);
or U21924 (N_21924,N_17541,N_17330);
nand U21925 (N_21925,N_15397,N_16035);
nand U21926 (N_21926,N_17758,N_19860);
nor U21927 (N_21927,N_17657,N_18180);
and U21928 (N_21928,N_15719,N_19282);
nor U21929 (N_21929,N_15559,N_16840);
nor U21930 (N_21930,N_16907,N_15456);
or U21931 (N_21931,N_16533,N_17865);
nand U21932 (N_21932,N_16305,N_18823);
xnor U21933 (N_21933,N_15507,N_15619);
nand U21934 (N_21934,N_17429,N_16800);
or U21935 (N_21935,N_18082,N_18096);
nor U21936 (N_21936,N_19085,N_17317);
nor U21937 (N_21937,N_17121,N_16431);
nor U21938 (N_21938,N_19793,N_19487);
xor U21939 (N_21939,N_19587,N_16978);
nor U21940 (N_21940,N_18862,N_15607);
or U21941 (N_21941,N_15466,N_19104);
and U21942 (N_21942,N_17802,N_16646);
and U21943 (N_21943,N_15519,N_15912);
or U21944 (N_21944,N_15317,N_17919);
or U21945 (N_21945,N_19892,N_18950);
xor U21946 (N_21946,N_16728,N_16100);
nand U21947 (N_21947,N_16706,N_17984);
or U21948 (N_21948,N_17679,N_18540);
and U21949 (N_21949,N_16281,N_18322);
xor U21950 (N_21950,N_19906,N_18485);
xnor U21951 (N_21951,N_16727,N_18539);
or U21952 (N_21952,N_17440,N_16028);
nor U21953 (N_21953,N_16568,N_19654);
nor U21954 (N_21954,N_19229,N_19845);
and U21955 (N_21955,N_15960,N_17490);
nor U21956 (N_21956,N_15523,N_17640);
or U21957 (N_21957,N_15543,N_15616);
or U21958 (N_21958,N_19960,N_15347);
nand U21959 (N_21959,N_16879,N_16493);
nor U21960 (N_21960,N_15855,N_16592);
and U21961 (N_21961,N_17037,N_18616);
xnor U21962 (N_21962,N_16833,N_17174);
and U21963 (N_21963,N_17798,N_19797);
and U21964 (N_21964,N_16785,N_18827);
xnor U21965 (N_21965,N_15010,N_19944);
and U21966 (N_21966,N_18329,N_17704);
or U21967 (N_21967,N_19656,N_16790);
nor U21968 (N_21968,N_18038,N_16757);
or U21969 (N_21969,N_19337,N_18458);
nor U21970 (N_21970,N_17936,N_15434);
and U21971 (N_21971,N_18590,N_19041);
xnor U21972 (N_21972,N_16684,N_18032);
nor U21973 (N_21973,N_15160,N_15899);
xnor U21974 (N_21974,N_15311,N_15606);
nand U21975 (N_21975,N_19732,N_16954);
and U21976 (N_21976,N_16663,N_19408);
nand U21977 (N_21977,N_19348,N_15074);
nor U21978 (N_21978,N_17396,N_19273);
nor U21979 (N_21979,N_19209,N_19939);
xnor U21980 (N_21980,N_18298,N_19037);
nor U21981 (N_21981,N_19992,N_19158);
or U21982 (N_21982,N_15838,N_17066);
and U21983 (N_21983,N_16222,N_16964);
or U21984 (N_21984,N_16709,N_19264);
and U21985 (N_21985,N_18856,N_18767);
nand U21986 (N_21986,N_19489,N_16004);
and U21987 (N_21987,N_15098,N_15408);
nor U21988 (N_21988,N_18830,N_15103);
nor U21989 (N_21989,N_15104,N_19985);
xor U21990 (N_21990,N_17815,N_16587);
and U21991 (N_21991,N_17456,N_15625);
nand U21992 (N_21992,N_17738,N_19423);
nand U21993 (N_21993,N_18733,N_19509);
and U21994 (N_21994,N_18990,N_15796);
and U21995 (N_21995,N_15429,N_16993);
xnor U21996 (N_21996,N_15031,N_16326);
nand U21997 (N_21997,N_18423,N_16027);
xnor U21998 (N_21998,N_18901,N_16215);
xnor U21999 (N_21999,N_17507,N_19927);
nand U22000 (N_22000,N_15753,N_18117);
nand U22001 (N_22001,N_16346,N_16809);
xor U22002 (N_22002,N_18043,N_16942);
nor U22003 (N_22003,N_18633,N_15015);
or U22004 (N_22004,N_15390,N_17215);
and U22005 (N_22005,N_19900,N_16967);
nand U22006 (N_22006,N_15924,N_15141);
xor U22007 (N_22007,N_15255,N_17768);
nand U22008 (N_22008,N_15401,N_15870);
nor U22009 (N_22009,N_15431,N_16051);
xor U22010 (N_22010,N_18397,N_16317);
nand U22011 (N_22011,N_19011,N_18780);
and U22012 (N_22012,N_16334,N_16985);
nor U22013 (N_22013,N_17092,N_17925);
and U22014 (N_22014,N_15462,N_18664);
and U22015 (N_22015,N_17390,N_17644);
nor U22016 (N_22016,N_18331,N_17393);
and U22017 (N_22017,N_18776,N_16260);
xnor U22018 (N_22018,N_16033,N_15751);
nor U22019 (N_22019,N_16071,N_19967);
or U22020 (N_22020,N_16886,N_17231);
nand U22021 (N_22021,N_16427,N_17570);
xnor U22022 (N_22022,N_15443,N_19479);
or U22023 (N_22023,N_15209,N_19938);
xnor U22024 (N_22024,N_18107,N_15139);
and U22025 (N_22025,N_19396,N_16527);
nand U22026 (N_22026,N_15012,N_16030);
nor U22027 (N_22027,N_17906,N_18466);
nor U22028 (N_22028,N_19605,N_16626);
nor U22029 (N_22029,N_17046,N_19471);
nand U22030 (N_22030,N_15045,N_19058);
xnor U22031 (N_22031,N_17293,N_18177);
nor U22032 (N_22032,N_17249,N_18176);
nand U22033 (N_22033,N_18211,N_15028);
xor U22034 (N_22034,N_16472,N_19834);
nor U22035 (N_22035,N_16611,N_17031);
and U22036 (N_22036,N_19493,N_19043);
or U22037 (N_22037,N_16218,N_19685);
xnor U22038 (N_22038,N_17374,N_19185);
and U22039 (N_22039,N_19850,N_17284);
nand U22040 (N_22040,N_16792,N_16162);
or U22041 (N_22041,N_16475,N_18018);
nand U22042 (N_22042,N_18537,N_17935);
nor U22043 (N_22043,N_16316,N_15859);
or U22044 (N_22044,N_15684,N_18221);
nand U22045 (N_22045,N_15750,N_16900);
nand U22046 (N_22046,N_19843,N_19519);
xnor U22047 (N_22047,N_17302,N_16574);
nand U22048 (N_22048,N_16113,N_17806);
xnor U22049 (N_22049,N_15473,N_17476);
nor U22050 (N_22050,N_17849,N_19612);
or U22051 (N_22051,N_19497,N_18110);
and U22052 (N_22052,N_17003,N_18753);
nand U22053 (N_22053,N_18855,N_18393);
and U22054 (N_22054,N_17180,N_15174);
nand U22055 (N_22055,N_18848,N_16887);
or U22056 (N_22056,N_19669,N_17766);
or U22057 (N_22057,N_16397,N_17855);
and U22058 (N_22058,N_19039,N_17371);
xor U22059 (N_22059,N_17257,N_16868);
nand U22060 (N_22060,N_18737,N_17616);
or U22061 (N_22061,N_16857,N_15522);
xor U22062 (N_22062,N_17269,N_19272);
xor U22063 (N_22063,N_18472,N_16529);
or U22064 (N_22064,N_15768,N_18656);
nand U22065 (N_22065,N_19355,N_15448);
or U22066 (N_22066,N_16340,N_18281);
nand U22067 (N_22067,N_18705,N_17754);
xnor U22068 (N_22068,N_18945,N_18498);
xnor U22069 (N_22069,N_15067,N_17218);
or U22070 (N_22070,N_17285,N_17034);
and U22071 (N_22071,N_19466,N_19601);
and U22072 (N_22072,N_15956,N_16063);
xor U22073 (N_22073,N_19630,N_19923);
and U22074 (N_22074,N_18541,N_17954);
or U22075 (N_22075,N_19178,N_19622);
nand U22076 (N_22076,N_17148,N_17361);
xnor U22077 (N_22077,N_17949,N_16875);
or U22078 (N_22078,N_15959,N_15052);
and U22079 (N_22079,N_15156,N_19293);
xor U22080 (N_22080,N_15115,N_16323);
nor U22081 (N_22081,N_15069,N_18745);
nand U22082 (N_22082,N_15261,N_19596);
xnor U22083 (N_22083,N_18165,N_19659);
or U22084 (N_22084,N_18075,N_15626);
nor U22085 (N_22085,N_16251,N_17960);
nand U22086 (N_22086,N_16137,N_18569);
xnor U22087 (N_22087,N_18957,N_18260);
and U22088 (N_22088,N_17778,N_16736);
nor U22089 (N_22089,N_15224,N_18453);
nor U22090 (N_22090,N_15892,N_16245);
nor U22091 (N_22091,N_18385,N_15878);
nor U22092 (N_22092,N_16949,N_17202);
or U22093 (N_22093,N_19725,N_18606);
nor U22094 (N_22094,N_17886,N_16154);
xor U22095 (N_22095,N_18912,N_19332);
nand U22096 (N_22096,N_18813,N_19030);
xnor U22097 (N_22097,N_15965,N_16147);
nor U22098 (N_22098,N_17725,N_19552);
xor U22099 (N_22099,N_17532,N_16374);
or U22100 (N_22100,N_18701,N_15153);
and U22101 (N_22101,N_17069,N_18773);
xnor U22102 (N_22102,N_19977,N_17943);
or U22103 (N_22103,N_15048,N_19756);
or U22104 (N_22104,N_17951,N_15866);
or U22105 (N_22105,N_16963,N_15382);
nor U22106 (N_22106,N_16636,N_15937);
nor U22107 (N_22107,N_18253,N_19973);
xor U22108 (N_22108,N_17153,N_17291);
and U22109 (N_22109,N_17764,N_16072);
xor U22110 (N_22110,N_15929,N_18842);
and U22111 (N_22111,N_16838,N_18424);
nor U22112 (N_22112,N_19844,N_16134);
nand U22113 (N_22113,N_16373,N_18521);
nor U22114 (N_22114,N_17688,N_17780);
xor U22115 (N_22115,N_19568,N_17503);
xnor U22116 (N_22116,N_18904,N_17113);
and U22117 (N_22117,N_17403,N_19615);
nand U22118 (N_22118,N_19347,N_16681);
nor U22119 (N_22119,N_16112,N_17356);
or U22120 (N_22120,N_15685,N_19763);
nor U22121 (N_22121,N_19791,N_18016);
nor U22122 (N_22122,N_19536,N_17809);
or U22123 (N_22123,N_18158,N_15108);
nand U22124 (N_22124,N_17641,N_18513);
xnor U22125 (N_22125,N_18661,N_18054);
xor U22126 (N_22126,N_15248,N_19999);
and U22127 (N_22127,N_15136,N_16685);
or U22128 (N_22128,N_18503,N_17274);
nor U22129 (N_22129,N_17181,N_15992);
nand U22130 (N_22130,N_16163,N_18720);
xor U22131 (N_22131,N_19169,N_17539);
xnor U22132 (N_22132,N_17206,N_18567);
and U22133 (N_22133,N_17611,N_19122);
nand U22134 (N_22134,N_15772,N_15502);
xnor U22135 (N_22135,N_17404,N_19210);
nor U22136 (N_22136,N_18604,N_15788);
nand U22137 (N_22137,N_18371,N_15877);
and U22138 (N_22138,N_16460,N_16888);
and U22139 (N_22139,N_19727,N_19270);
and U22140 (N_22140,N_17878,N_18939);
and U22141 (N_22141,N_16034,N_15879);
and U22142 (N_22142,N_15357,N_16552);
nor U22143 (N_22143,N_18157,N_18008);
and U22144 (N_22144,N_17639,N_17152);
or U22145 (N_22145,N_19163,N_15049);
and U22146 (N_22146,N_19450,N_16579);
and U22147 (N_22147,N_19657,N_17905);
nor U22148 (N_22148,N_19879,N_15821);
xnor U22149 (N_22149,N_19969,N_15044);
and U22150 (N_22150,N_16989,N_19974);
and U22151 (N_22151,N_19262,N_15857);
and U22152 (N_22152,N_19520,N_17384);
or U22153 (N_22153,N_15700,N_15941);
or U22154 (N_22154,N_19498,N_15276);
and U22155 (N_22155,N_18000,N_19363);
and U22156 (N_22156,N_16948,N_18587);
xor U22157 (N_22157,N_17797,N_19639);
nand U22158 (N_22158,N_16534,N_15107);
nor U22159 (N_22159,N_16469,N_19453);
and U22160 (N_22160,N_18795,N_18975);
nor U22161 (N_22161,N_19889,N_16772);
nor U22162 (N_22162,N_15421,N_19576);
and U22163 (N_22163,N_18403,N_17990);
nor U22164 (N_22164,N_16688,N_17007);
nor U22165 (N_22165,N_15369,N_18138);
xnor U22166 (N_22166,N_15088,N_16966);
nor U22167 (N_22167,N_18799,N_17786);
nand U22168 (N_22168,N_17597,N_17227);
and U22169 (N_22169,N_19140,N_18628);
nand U22170 (N_22170,N_19773,N_18792);
nor U22171 (N_22171,N_16108,N_16202);
or U22172 (N_22172,N_17441,N_19090);
nand U22173 (N_22173,N_19511,N_19333);
xnor U22174 (N_22174,N_19299,N_16903);
nand U22175 (N_22175,N_19968,N_18846);
xor U22176 (N_22176,N_18602,N_19328);
or U22177 (N_22177,N_16403,N_17023);
xnor U22178 (N_22178,N_18140,N_17131);
or U22179 (N_22179,N_16457,N_19105);
and U22180 (N_22180,N_17029,N_17176);
or U22181 (N_22181,N_15557,N_17600);
or U22182 (N_22182,N_15852,N_17076);
or U22183 (N_22183,N_15236,N_18895);
or U22184 (N_22184,N_18452,N_17944);
nor U22185 (N_22185,N_16356,N_18290);
xor U22186 (N_22186,N_18763,N_17450);
xnor U22187 (N_22187,N_15550,N_19357);
xor U22188 (N_22188,N_19614,N_15837);
xor U22189 (N_22189,N_16307,N_17952);
nor U22190 (N_22190,N_18475,N_16502);
xnor U22191 (N_22191,N_18288,N_17079);
xor U22192 (N_22192,N_17913,N_15379);
and U22193 (N_22193,N_16544,N_15614);
nor U22194 (N_22194,N_15058,N_16298);
xor U22195 (N_22195,N_16537,N_16511);
or U22196 (N_22196,N_19753,N_17903);
and U22197 (N_22197,N_19557,N_16615);
and U22198 (N_22198,N_15563,N_16696);
xnor U22199 (N_22199,N_18963,N_15508);
or U22200 (N_22200,N_16847,N_19381);
and U22201 (N_22201,N_17706,N_16336);
or U22202 (N_22202,N_16280,N_16713);
nor U22203 (N_22203,N_18023,N_18692);
nor U22204 (N_22204,N_17646,N_15577);
nor U22205 (N_22205,N_15292,N_16256);
xnor U22206 (N_22206,N_18464,N_15950);
xor U22207 (N_22207,N_16764,N_16674);
nor U22208 (N_22208,N_17267,N_16521);
or U22209 (N_22209,N_17671,N_18143);
or U22210 (N_22210,N_15025,N_17489);
nand U22211 (N_22211,N_17593,N_15492);
or U22212 (N_22212,N_19442,N_15687);
and U22213 (N_22213,N_18658,N_17707);
and U22214 (N_22214,N_17158,N_15146);
or U22215 (N_22215,N_18951,N_17683);
xor U22216 (N_22216,N_19115,N_19528);
xor U22217 (N_22217,N_17694,N_17968);
or U22218 (N_22218,N_15663,N_15854);
nor U22219 (N_22219,N_16158,N_15703);
nor U22220 (N_22220,N_18399,N_17622);
xnor U22221 (N_22221,N_15779,N_15083);
nand U22222 (N_22222,N_17963,N_17785);
or U22223 (N_22223,N_17922,N_18326);
xor U22224 (N_22224,N_15459,N_18276);
nor U22225 (N_22225,N_16678,N_15665);
or U22226 (N_22226,N_17680,N_18451);
and U22227 (N_22227,N_19155,N_17770);
or U22228 (N_22228,N_17856,N_15151);
xnor U22229 (N_22229,N_15439,N_18033);
or U22230 (N_22230,N_18612,N_19561);
and U22231 (N_22231,N_15618,N_19819);
xnor U22232 (N_22232,N_19151,N_16102);
or U22233 (N_22233,N_16152,N_15673);
and U22234 (N_22234,N_15604,N_19362);
xnor U22235 (N_22235,N_18599,N_18444);
nand U22236 (N_22236,N_19194,N_19343);
nand U22237 (N_22237,N_15802,N_18762);
or U22238 (N_22238,N_19129,N_17012);
xor U22239 (N_22239,N_15858,N_19737);
and U22240 (N_22240,N_18467,N_15501);
nor U22241 (N_22241,N_15962,N_19577);
nand U22242 (N_22242,N_17248,N_19603);
nor U22243 (N_22243,N_18185,N_18727);
and U22244 (N_22244,N_17417,N_19228);
nor U22245 (N_22245,N_16476,N_19389);
nor U22246 (N_22246,N_16069,N_16483);
nand U22247 (N_22247,N_15593,N_15561);
nor U22248 (N_22248,N_19955,N_18068);
or U22249 (N_22249,N_15373,N_18214);
and U22250 (N_22250,N_16203,N_16943);
or U22251 (N_22251,N_15246,N_18603);
and U22252 (N_22252,N_16759,N_15588);
xnor U22253 (N_22253,N_15226,N_18890);
nand U22254 (N_22254,N_19426,N_16768);
or U22255 (N_22255,N_17336,N_18469);
xor U22256 (N_22256,N_16610,N_18364);
and U22257 (N_22257,N_17350,N_17923);
or U22258 (N_22258,N_17887,N_19746);
nand U22259 (N_22259,N_17863,N_18675);
or U22260 (N_22260,N_15576,N_18841);
and U22261 (N_22261,N_18959,N_17044);
xor U22262 (N_22262,N_18257,N_16894);
or U22263 (N_22263,N_15166,N_19954);
xor U22264 (N_22264,N_17765,N_15281);
or U22265 (N_22265,N_19813,N_17175);
and U22266 (N_22266,N_18164,N_19257);
nor U22267 (N_22267,N_15206,N_19284);
or U22268 (N_22268,N_19338,N_16073);
nand U22269 (N_22269,N_18935,N_17832);
and U22270 (N_22270,N_19750,N_19268);
xor U22271 (N_22271,N_17137,N_17255);
and U22272 (N_22272,N_18077,N_16867);
nand U22273 (N_22273,N_15658,N_15529);
nand U22274 (N_22274,N_15321,N_16239);
nand U22275 (N_22275,N_16651,N_19467);
nand U22276 (N_22276,N_16932,N_15565);
nand U22277 (N_22277,N_16366,N_17035);
and U22278 (N_22278,N_18489,N_15202);
xor U22279 (N_22279,N_15763,N_18105);
and U22280 (N_22280,N_19181,N_15287);
and U22281 (N_22281,N_19664,N_16632);
nor U22282 (N_22282,N_19508,N_16235);
and U22283 (N_22283,N_17473,N_16361);
or U22284 (N_22284,N_15413,N_15479);
xor U22285 (N_22285,N_15353,N_17665);
and U22286 (N_22286,N_17062,N_16180);
or U22287 (N_22287,N_19655,N_16750);
xor U22288 (N_22288,N_15525,N_17962);
nand U22289 (N_22289,N_18172,N_16958);
nor U22290 (N_22290,N_16763,N_19835);
and U22291 (N_22291,N_18250,N_15114);
and U22292 (N_22292,N_15455,N_17352);
nand U22293 (N_22293,N_15847,N_16459);
and U22294 (N_22294,N_17519,N_17411);
or U22295 (N_22295,N_18546,N_19908);
and U22296 (N_22296,N_16753,N_16509);
or U22297 (N_22297,N_19302,N_15189);
nand U22298 (N_22298,N_15043,N_16466);
xnor U22299 (N_22299,N_17219,N_17324);
nor U22300 (N_22300,N_18710,N_17571);
nand U22301 (N_22301,N_19064,N_19880);
nor U22302 (N_22302,N_19499,N_18575);
nor U22303 (N_22303,N_18162,N_16955);
nor U22304 (N_22304,N_15194,N_16169);
or U22305 (N_22305,N_17673,N_18235);
xor U22306 (N_22306,N_16265,N_16499);
nand U22307 (N_22307,N_19306,N_19517);
nand U22308 (N_22308,N_15539,N_18772);
xor U22309 (N_22309,N_15668,N_15963);
or U22310 (N_22310,N_19558,N_19734);
nand U22311 (N_22311,N_16921,N_19087);
and U22312 (N_22312,N_18613,N_19765);
and U22313 (N_22313,N_16349,N_17323);
nor U22314 (N_22314,N_18832,N_16168);
xnor U22315 (N_22315,N_17232,N_18311);
or U22316 (N_22316,N_19541,N_15128);
and U22317 (N_22317,N_17606,N_16945);
nor U22318 (N_22318,N_19611,N_19280);
nand U22319 (N_22319,N_16913,N_16000);
nor U22320 (N_22320,N_19652,N_19700);
and U22321 (N_22321,N_19820,N_16355);
or U22322 (N_22322,N_15426,N_16865);
and U22323 (N_22323,N_16044,N_19916);
or U22324 (N_22324,N_19431,N_17304);
or U22325 (N_22325,N_15109,N_16991);
or U22326 (N_22326,N_15558,N_19609);
nor U22327 (N_22327,N_16151,N_19524);
nand U22328 (N_22328,N_18229,N_15770);
nand U22329 (N_22329,N_16166,N_17789);
or U22330 (N_22330,N_15623,N_19335);
nor U22331 (N_22331,N_15605,N_16096);
and U22332 (N_22332,N_17634,N_18714);
xnor U22333 (N_22333,N_19839,N_19673);
nand U22334 (N_22334,N_16602,N_15249);
nor U22335 (N_22335,N_18025,N_15210);
nand U22336 (N_22336,N_17852,N_15399);
and U22337 (N_22337,N_15360,N_17614);
or U22338 (N_22338,N_18969,N_18283);
nor U22339 (N_22339,N_19142,N_19533);
nand U22340 (N_22340,N_17383,N_18925);
or U22341 (N_22341,N_18746,N_19480);
or U22342 (N_22342,N_15247,N_17578);
and U22343 (N_22343,N_15713,N_16691);
and U22344 (N_22344,N_18029,N_19364);
nand U22345 (N_22345,N_17500,N_18428);
and U22346 (N_22346,N_19672,N_18645);
nor U22347 (N_22347,N_16661,N_19017);
or U22348 (N_22348,N_18535,N_17461);
and U22349 (N_22349,N_19383,N_18327);
nor U22350 (N_22350,N_17295,N_16807);
xor U22351 (N_22351,N_18654,N_15916);
nand U22352 (N_22352,N_18894,N_19817);
and U22353 (N_22353,N_16624,N_18359);
or U22354 (N_22354,N_18863,N_18914);
xor U22355 (N_22355,N_18367,N_18245);
nand U22356 (N_22356,N_19441,N_16290);
xnor U22357 (N_22357,N_17544,N_19662);
xnor U22358 (N_22358,N_15774,N_18014);
nor U22359 (N_22359,N_16931,N_15518);
nand U22360 (N_22360,N_17787,N_17093);
or U22361 (N_22361,N_15655,N_15140);
xnor U22362 (N_22362,N_16946,N_17790);
nor U22363 (N_22363,N_16739,N_19862);
nand U22364 (N_22364,N_19003,N_16498);
xnor U22365 (N_22365,N_15349,N_15925);
or U22366 (N_22366,N_18182,N_16208);
xnor U22367 (N_22367,N_18618,N_18338);
and U22368 (N_22368,N_17912,N_16153);
nand U22369 (N_22369,N_19128,N_16860);
nand U22370 (N_22370,N_18570,N_18188);
nand U22371 (N_22371,N_16726,N_18124);
or U22372 (N_22372,N_19217,N_19116);
xor U22373 (N_22373,N_16409,N_17769);
and U22374 (N_22374,N_19301,N_17309);
nor U22375 (N_22375,N_16607,N_16383);
or U22376 (N_22376,N_15375,N_15477);
xor U22377 (N_22377,N_17266,N_18756);
nor U22378 (N_22378,N_15350,N_16050);
and U22379 (N_22379,N_18104,N_15405);
nor U22380 (N_22380,N_16232,N_16363);
and U22381 (N_22381,N_16572,N_17993);
xor U22382 (N_22382,N_17642,N_17233);
nand U22383 (N_22383,N_19504,N_19735);
xor U22384 (N_22384,N_16291,N_16213);
nand U22385 (N_22385,N_16518,N_17357);
or U22386 (N_22386,N_19516,N_16606);
xor U22387 (N_22387,N_19130,N_17238);
nand U22388 (N_22388,N_17453,N_16902);
and U22389 (N_22389,N_16140,N_19971);
and U22390 (N_22390,N_17623,N_19620);
or U22391 (N_22391,N_17423,N_15820);
and U22392 (N_22392,N_17479,N_15881);
nor U22393 (N_22393,N_15946,N_15923);
nor U22394 (N_22394,N_17139,N_17620);
or U22395 (N_22395,N_15545,N_18624);
and U22396 (N_22396,N_15498,N_15315);
nor U22397 (N_22397,N_15449,N_19786);
nor U22398 (N_22398,N_15137,N_18119);
xor U22399 (N_22399,N_15842,N_18202);
xor U22400 (N_22400,N_17082,N_16557);
nor U22401 (N_22401,N_17808,N_16362);
and U22402 (N_22402,N_17861,N_18103);
nand U22403 (N_22403,N_18193,N_19481);
nand U22404 (N_22404,N_18723,N_15548);
xnor U22405 (N_22405,N_19619,N_16201);
xor U22406 (N_22406,N_15297,N_16205);
nand U22407 (N_22407,N_19933,N_16350);
and U22408 (N_22408,N_19570,N_18598);
or U22409 (N_22409,N_17230,N_18649);
and U22410 (N_22410,N_15013,N_16389);
and U22411 (N_22411,N_15863,N_16021);
nor U22412 (N_22412,N_15832,N_17041);
nand U22413 (N_22413,N_16390,N_18432);
or U22414 (N_22414,N_16376,N_16605);
or U22415 (N_22415,N_18693,N_18030);
nor U22416 (N_22416,N_19494,N_17689);
nand U22417 (N_22417,N_15935,N_19830);
nor U22418 (N_22418,N_19180,N_16434);
and U22419 (N_22419,N_17509,N_19594);
nor U22420 (N_22420,N_19250,N_19800);
nor U22421 (N_22421,N_19136,N_15701);
and U22422 (N_22422,N_16616,N_19360);
xor U22423 (N_22423,N_15883,N_16339);
or U22424 (N_22424,N_17522,N_17609);
and U22425 (N_22425,N_19114,N_18865);
nor U22426 (N_22426,N_15050,N_17846);
nor U22427 (N_22427,N_17517,N_19705);
and U22428 (N_22428,N_16962,N_18333);
xor U22429 (N_22429,N_15006,N_19781);
and U22430 (N_22430,N_15531,N_17211);
or U22431 (N_22431,N_18686,N_18817);
xnor U22432 (N_22432,N_19863,N_16392);
xnor U22433 (N_22433,N_19162,N_17546);
or U22434 (N_22434,N_17030,N_15936);
and U22435 (N_22435,N_18121,N_18553);
or U22436 (N_22436,N_17803,N_15171);
and U22437 (N_22437,N_18607,N_16129);
or U22438 (N_22438,N_15289,N_17632);
or U22439 (N_22439,N_16442,N_17916);
nor U22440 (N_22440,N_19079,N_19490);
nand U22441 (N_22441,N_16204,N_15579);
xor U22442 (N_22442,N_17315,N_18850);
nand U22443 (N_22443,N_18047,N_15813);
or U22444 (N_22444,N_16195,N_15885);
or U22445 (N_22445,N_17240,N_15444);
xnor U22446 (N_22446,N_16520,N_17781);
and U22447 (N_22447,N_17235,N_15312);
nor U22448 (N_22448,N_16338,N_19928);
and U22449 (N_22449,N_15981,N_15011);
xor U22450 (N_22450,N_19255,N_19696);
xnor U22451 (N_22451,N_16405,N_18026);
nor U22452 (N_22452,N_18254,N_16212);
and U22453 (N_22453,N_16464,N_18296);
nand U22454 (N_22454,N_16016,N_16429);
nand U22455 (N_22455,N_15582,N_16808);
nand U22456 (N_22456,N_18679,N_15211);
xnor U22457 (N_22457,N_16686,N_16441);
or U22458 (N_22458,N_17492,N_17286);
and U22459 (N_22459,N_18941,N_17136);
or U22460 (N_22460,N_19344,N_17354);
xnor U22461 (N_22461,N_19165,N_15239);
xor U22462 (N_22462,N_16329,N_18460);
xnor U22463 (N_22463,N_15503,N_18416);
xor U22464 (N_22464,N_19537,N_19240);
nor U22465 (N_22465,N_19141,N_15158);
and U22466 (N_22466,N_19767,N_15170);
nor U22467 (N_22467,N_19061,N_17930);
xnor U22468 (N_22468,N_19012,N_19073);
nor U22469 (N_22469,N_15203,N_15731);
nand U22470 (N_22470,N_19838,N_17307);
nor U22471 (N_22471,N_18875,N_18216);
nor U22472 (N_22472,N_18412,N_16851);
or U22473 (N_22473,N_19277,N_17714);
xor U22474 (N_22474,N_16216,N_15322);
and U22475 (N_22475,N_17426,N_19829);
nor U22476 (N_22476,N_15520,N_17297);
and U22477 (N_22477,N_17011,N_18888);
nor U22478 (N_22478,N_15154,N_17466);
nor U22479 (N_22479,N_17650,N_18076);
xor U22480 (N_22480,N_19260,N_19671);
and U22481 (N_22481,N_19893,N_15097);
nand U22482 (N_22482,N_19437,N_17157);
xor U22483 (N_22483,N_19686,N_18186);
nand U22484 (N_22484,N_15332,N_17068);
and U22485 (N_22485,N_15566,N_15683);
and U22486 (N_22486,N_18230,N_16090);
xor U22487 (N_22487,N_16909,N_18666);
xnor U22488 (N_22488,N_19780,N_18771);
nor U22489 (N_22489,N_19139,N_19998);
nand U22490 (N_22490,N_18139,N_17533);
xnor U22491 (N_22491,N_17090,N_16311);
xor U22492 (N_22492,N_15757,N_19600);
or U22493 (N_22493,N_19189,N_16577);
nor U22494 (N_22494,N_17095,N_15450);
nand U22495 (N_22495,N_17869,N_19492);
xor U22496 (N_22496,N_15018,N_15046);
and U22497 (N_22497,N_17104,N_18702);
nor U22498 (N_22498,N_16101,N_16164);
xor U22499 (N_22499,N_19929,N_18136);
nor U22500 (N_22500,N_17247,N_17867);
nor U22501 (N_22501,N_18785,N_19752);
and U22502 (N_22502,N_18786,N_15038);
xnor U22503 (N_22503,N_15447,N_19106);
or U22504 (N_22504,N_15168,N_18977);
xor U22505 (N_22505,N_15155,N_18372);
xnor U22506 (N_22506,N_15614,N_19742);
or U22507 (N_22507,N_15175,N_15771);
xor U22508 (N_22508,N_15213,N_19352);
and U22509 (N_22509,N_18453,N_18418);
and U22510 (N_22510,N_15565,N_15761);
or U22511 (N_22511,N_18938,N_19906);
or U22512 (N_22512,N_16676,N_19220);
nand U22513 (N_22513,N_18791,N_15109);
xnor U22514 (N_22514,N_17564,N_15541);
nand U22515 (N_22515,N_15704,N_15850);
or U22516 (N_22516,N_19072,N_19677);
nor U22517 (N_22517,N_18404,N_16677);
nor U22518 (N_22518,N_19470,N_17204);
nor U22519 (N_22519,N_15676,N_19341);
nand U22520 (N_22520,N_15503,N_16086);
nor U22521 (N_22521,N_15501,N_16026);
nand U22522 (N_22522,N_16033,N_16245);
or U22523 (N_22523,N_17979,N_15454);
xor U22524 (N_22524,N_17386,N_16247);
xor U22525 (N_22525,N_19710,N_19161);
or U22526 (N_22526,N_17424,N_18452);
nor U22527 (N_22527,N_18281,N_19411);
and U22528 (N_22528,N_17003,N_19073);
xnor U22529 (N_22529,N_15385,N_15545);
or U22530 (N_22530,N_15916,N_16586);
or U22531 (N_22531,N_19818,N_18513);
nand U22532 (N_22532,N_18552,N_15650);
xnor U22533 (N_22533,N_18614,N_16981);
and U22534 (N_22534,N_16255,N_16146);
nor U22535 (N_22535,N_17905,N_16283);
nor U22536 (N_22536,N_16851,N_19191);
and U22537 (N_22537,N_17503,N_16583);
xnor U22538 (N_22538,N_19979,N_17560);
nor U22539 (N_22539,N_18322,N_17067);
or U22540 (N_22540,N_17716,N_16712);
xnor U22541 (N_22541,N_16906,N_18949);
nor U22542 (N_22542,N_19351,N_16118);
xnor U22543 (N_22543,N_18490,N_18957);
or U22544 (N_22544,N_15067,N_15546);
nor U22545 (N_22545,N_16937,N_17764);
nor U22546 (N_22546,N_17734,N_16640);
or U22547 (N_22547,N_15094,N_16674);
and U22548 (N_22548,N_18414,N_19068);
or U22549 (N_22549,N_17996,N_16680);
xnor U22550 (N_22550,N_16495,N_16078);
or U22551 (N_22551,N_18322,N_16032);
nor U22552 (N_22552,N_15418,N_16751);
or U22553 (N_22553,N_17800,N_17229);
xnor U22554 (N_22554,N_17837,N_16259);
nand U22555 (N_22555,N_19439,N_15357);
or U22556 (N_22556,N_18091,N_17483);
and U22557 (N_22557,N_17343,N_17852);
nand U22558 (N_22558,N_19150,N_15567);
nor U22559 (N_22559,N_15087,N_15575);
nor U22560 (N_22560,N_15404,N_18078);
nand U22561 (N_22561,N_18565,N_18341);
or U22562 (N_22562,N_18844,N_18529);
and U22563 (N_22563,N_18565,N_15989);
xnor U22564 (N_22564,N_18112,N_15238);
nand U22565 (N_22565,N_16909,N_16954);
nor U22566 (N_22566,N_17330,N_15407);
or U22567 (N_22567,N_15151,N_18210);
and U22568 (N_22568,N_19007,N_15991);
nor U22569 (N_22569,N_19811,N_16866);
nand U22570 (N_22570,N_15293,N_15927);
and U22571 (N_22571,N_17090,N_19291);
xor U22572 (N_22572,N_18509,N_15980);
nand U22573 (N_22573,N_19703,N_15635);
nor U22574 (N_22574,N_15734,N_15258);
xor U22575 (N_22575,N_18065,N_19170);
and U22576 (N_22576,N_15942,N_15648);
nand U22577 (N_22577,N_18560,N_16963);
nor U22578 (N_22578,N_17153,N_19715);
or U22579 (N_22579,N_18126,N_17225);
xnor U22580 (N_22580,N_19825,N_16913);
xor U22581 (N_22581,N_19228,N_16963);
nand U22582 (N_22582,N_15407,N_19550);
xor U22583 (N_22583,N_16641,N_18426);
or U22584 (N_22584,N_16309,N_18267);
and U22585 (N_22585,N_18757,N_16079);
nand U22586 (N_22586,N_18618,N_19774);
nor U22587 (N_22587,N_16551,N_15207);
nor U22588 (N_22588,N_18130,N_16556);
nand U22589 (N_22589,N_15713,N_18788);
nand U22590 (N_22590,N_15702,N_16483);
nor U22591 (N_22591,N_19437,N_19415);
nand U22592 (N_22592,N_16757,N_19274);
nand U22593 (N_22593,N_18885,N_18566);
nand U22594 (N_22594,N_18266,N_17152);
nand U22595 (N_22595,N_15815,N_19481);
nor U22596 (N_22596,N_18011,N_17346);
xor U22597 (N_22597,N_19624,N_15434);
nand U22598 (N_22598,N_16153,N_19181);
nand U22599 (N_22599,N_17244,N_16369);
nand U22600 (N_22600,N_16576,N_16492);
and U22601 (N_22601,N_18293,N_18559);
and U22602 (N_22602,N_15621,N_16736);
xnor U22603 (N_22603,N_15141,N_18070);
and U22604 (N_22604,N_19038,N_18534);
nand U22605 (N_22605,N_19388,N_17898);
and U22606 (N_22606,N_15526,N_17558);
or U22607 (N_22607,N_16915,N_16293);
nor U22608 (N_22608,N_17284,N_18319);
xnor U22609 (N_22609,N_15928,N_16422);
and U22610 (N_22610,N_19966,N_17852);
nor U22611 (N_22611,N_16005,N_16236);
nand U22612 (N_22612,N_15430,N_16427);
and U22613 (N_22613,N_18963,N_15769);
nor U22614 (N_22614,N_19419,N_16302);
nor U22615 (N_22615,N_16104,N_17101);
nor U22616 (N_22616,N_15408,N_15334);
and U22617 (N_22617,N_18188,N_18791);
xor U22618 (N_22618,N_15224,N_17035);
nor U22619 (N_22619,N_16547,N_17303);
and U22620 (N_22620,N_15499,N_16754);
nor U22621 (N_22621,N_16577,N_15158);
nor U22622 (N_22622,N_18564,N_17573);
xnor U22623 (N_22623,N_18536,N_18285);
nand U22624 (N_22624,N_19064,N_15739);
nor U22625 (N_22625,N_18852,N_18221);
xor U22626 (N_22626,N_16820,N_17789);
nor U22627 (N_22627,N_18458,N_18308);
and U22628 (N_22628,N_17125,N_18557);
and U22629 (N_22629,N_16193,N_19852);
or U22630 (N_22630,N_19580,N_19198);
and U22631 (N_22631,N_19115,N_17400);
nand U22632 (N_22632,N_16537,N_16395);
xnor U22633 (N_22633,N_17658,N_16345);
nand U22634 (N_22634,N_17128,N_15126);
nand U22635 (N_22635,N_18377,N_18718);
xnor U22636 (N_22636,N_16765,N_15318);
or U22637 (N_22637,N_17158,N_16862);
and U22638 (N_22638,N_16999,N_19785);
or U22639 (N_22639,N_16638,N_16705);
xnor U22640 (N_22640,N_18278,N_17093);
xnor U22641 (N_22641,N_15948,N_19183);
nor U22642 (N_22642,N_16637,N_19333);
or U22643 (N_22643,N_16643,N_19086);
or U22644 (N_22644,N_15751,N_17431);
and U22645 (N_22645,N_15855,N_15314);
nand U22646 (N_22646,N_19328,N_16326);
and U22647 (N_22647,N_16379,N_19153);
xor U22648 (N_22648,N_16575,N_19656);
or U22649 (N_22649,N_15181,N_18888);
xor U22650 (N_22650,N_16690,N_15865);
nand U22651 (N_22651,N_19841,N_15182);
or U22652 (N_22652,N_15129,N_19933);
xor U22653 (N_22653,N_17921,N_19808);
nand U22654 (N_22654,N_15746,N_17232);
or U22655 (N_22655,N_19471,N_15885);
and U22656 (N_22656,N_19301,N_16931);
nor U22657 (N_22657,N_18290,N_17589);
and U22658 (N_22658,N_19823,N_19222);
nor U22659 (N_22659,N_18386,N_16406);
xnor U22660 (N_22660,N_18572,N_16362);
nor U22661 (N_22661,N_17878,N_16833);
xor U22662 (N_22662,N_19030,N_16610);
and U22663 (N_22663,N_17816,N_15481);
and U22664 (N_22664,N_19095,N_16741);
and U22665 (N_22665,N_18227,N_16839);
nor U22666 (N_22666,N_15782,N_17363);
or U22667 (N_22667,N_18268,N_16440);
or U22668 (N_22668,N_15891,N_17397);
nand U22669 (N_22669,N_18910,N_18960);
nor U22670 (N_22670,N_15116,N_18458);
nand U22671 (N_22671,N_16686,N_19141);
or U22672 (N_22672,N_17723,N_17260);
nor U22673 (N_22673,N_17177,N_18204);
and U22674 (N_22674,N_18990,N_18565);
nor U22675 (N_22675,N_16954,N_17458);
and U22676 (N_22676,N_15356,N_17038);
and U22677 (N_22677,N_19468,N_17523);
or U22678 (N_22678,N_15672,N_15542);
nand U22679 (N_22679,N_19934,N_15371);
nor U22680 (N_22680,N_17113,N_16232);
nand U22681 (N_22681,N_18311,N_16083);
nor U22682 (N_22682,N_16159,N_17540);
nor U22683 (N_22683,N_16633,N_19219);
or U22684 (N_22684,N_17946,N_16353);
or U22685 (N_22685,N_15786,N_18918);
nor U22686 (N_22686,N_16728,N_15196);
xnor U22687 (N_22687,N_15127,N_19107);
xnor U22688 (N_22688,N_15323,N_19481);
and U22689 (N_22689,N_18789,N_16761);
nand U22690 (N_22690,N_15060,N_15627);
nor U22691 (N_22691,N_18131,N_15597);
nor U22692 (N_22692,N_15523,N_17924);
nand U22693 (N_22693,N_17426,N_18607);
nand U22694 (N_22694,N_19937,N_16386);
nor U22695 (N_22695,N_16906,N_17460);
xnor U22696 (N_22696,N_19002,N_17062);
nand U22697 (N_22697,N_18691,N_19934);
nand U22698 (N_22698,N_16085,N_15208);
nor U22699 (N_22699,N_16746,N_17364);
nand U22700 (N_22700,N_19692,N_16204);
nand U22701 (N_22701,N_18498,N_19841);
nor U22702 (N_22702,N_18582,N_19194);
or U22703 (N_22703,N_15089,N_16375);
and U22704 (N_22704,N_18658,N_17841);
nand U22705 (N_22705,N_17043,N_19080);
or U22706 (N_22706,N_16148,N_18226);
or U22707 (N_22707,N_17744,N_17568);
nor U22708 (N_22708,N_17627,N_17093);
nor U22709 (N_22709,N_17588,N_19760);
nor U22710 (N_22710,N_19273,N_19940);
xor U22711 (N_22711,N_16338,N_16681);
nand U22712 (N_22712,N_17454,N_15926);
xnor U22713 (N_22713,N_18155,N_15887);
or U22714 (N_22714,N_15106,N_19777);
nand U22715 (N_22715,N_17447,N_16553);
or U22716 (N_22716,N_15285,N_17398);
or U22717 (N_22717,N_17046,N_16428);
xor U22718 (N_22718,N_17292,N_17853);
and U22719 (N_22719,N_16615,N_16047);
nand U22720 (N_22720,N_17370,N_15088);
nor U22721 (N_22721,N_18175,N_18918);
xor U22722 (N_22722,N_19931,N_15708);
or U22723 (N_22723,N_17189,N_15054);
or U22724 (N_22724,N_17236,N_17092);
nand U22725 (N_22725,N_19147,N_18997);
nor U22726 (N_22726,N_18868,N_17413);
and U22727 (N_22727,N_19659,N_16507);
and U22728 (N_22728,N_19809,N_16420);
nand U22729 (N_22729,N_18412,N_15266);
nor U22730 (N_22730,N_15177,N_19492);
nor U22731 (N_22731,N_18730,N_18615);
and U22732 (N_22732,N_16688,N_15638);
xor U22733 (N_22733,N_16444,N_15226);
nor U22734 (N_22734,N_19007,N_16333);
or U22735 (N_22735,N_16791,N_16279);
or U22736 (N_22736,N_16069,N_15122);
and U22737 (N_22737,N_18416,N_16624);
xnor U22738 (N_22738,N_18968,N_16196);
nor U22739 (N_22739,N_18469,N_19753);
and U22740 (N_22740,N_16379,N_17137);
nor U22741 (N_22741,N_16727,N_15955);
xor U22742 (N_22742,N_17578,N_16503);
or U22743 (N_22743,N_19717,N_19297);
and U22744 (N_22744,N_19673,N_15808);
nor U22745 (N_22745,N_17856,N_19050);
nand U22746 (N_22746,N_18747,N_19017);
nand U22747 (N_22747,N_16344,N_16311);
nor U22748 (N_22748,N_15888,N_16639);
or U22749 (N_22749,N_18304,N_17785);
nand U22750 (N_22750,N_19968,N_19992);
xor U22751 (N_22751,N_19045,N_19738);
or U22752 (N_22752,N_18995,N_16949);
and U22753 (N_22753,N_17689,N_17692);
xor U22754 (N_22754,N_15580,N_19018);
xor U22755 (N_22755,N_19412,N_16000);
and U22756 (N_22756,N_15885,N_18556);
xor U22757 (N_22757,N_17025,N_15718);
and U22758 (N_22758,N_15911,N_19484);
and U22759 (N_22759,N_16765,N_17878);
nand U22760 (N_22760,N_17279,N_18856);
and U22761 (N_22761,N_15307,N_17212);
or U22762 (N_22762,N_19320,N_18848);
xor U22763 (N_22763,N_17696,N_19062);
and U22764 (N_22764,N_18115,N_19829);
and U22765 (N_22765,N_16347,N_15135);
nor U22766 (N_22766,N_15238,N_16967);
and U22767 (N_22767,N_19402,N_19327);
or U22768 (N_22768,N_16436,N_16471);
or U22769 (N_22769,N_15143,N_19912);
or U22770 (N_22770,N_16665,N_15623);
xor U22771 (N_22771,N_17284,N_17521);
or U22772 (N_22772,N_19371,N_17472);
or U22773 (N_22773,N_17098,N_16219);
or U22774 (N_22774,N_18820,N_15442);
or U22775 (N_22775,N_18890,N_18808);
xor U22776 (N_22776,N_15501,N_17877);
xnor U22777 (N_22777,N_16063,N_17711);
and U22778 (N_22778,N_17299,N_18357);
or U22779 (N_22779,N_17887,N_16266);
or U22780 (N_22780,N_18018,N_16229);
nand U22781 (N_22781,N_16538,N_16075);
nand U22782 (N_22782,N_18934,N_19139);
xnor U22783 (N_22783,N_15972,N_16177);
or U22784 (N_22784,N_15284,N_16456);
or U22785 (N_22785,N_16490,N_17206);
nand U22786 (N_22786,N_16969,N_19105);
nor U22787 (N_22787,N_15102,N_15764);
nand U22788 (N_22788,N_16650,N_19238);
xor U22789 (N_22789,N_17007,N_16225);
nor U22790 (N_22790,N_17090,N_19719);
or U22791 (N_22791,N_15109,N_19305);
nor U22792 (N_22792,N_15428,N_17895);
nand U22793 (N_22793,N_19492,N_15592);
nor U22794 (N_22794,N_17905,N_16254);
or U22795 (N_22795,N_18324,N_18430);
or U22796 (N_22796,N_19995,N_17762);
nand U22797 (N_22797,N_19524,N_19747);
nand U22798 (N_22798,N_18285,N_15985);
nor U22799 (N_22799,N_17282,N_17750);
and U22800 (N_22800,N_16462,N_15055);
xnor U22801 (N_22801,N_18915,N_15014);
nor U22802 (N_22802,N_19962,N_16733);
xnor U22803 (N_22803,N_19773,N_16470);
or U22804 (N_22804,N_15358,N_15006);
and U22805 (N_22805,N_18944,N_16082);
xor U22806 (N_22806,N_16418,N_15811);
nand U22807 (N_22807,N_17257,N_17746);
xnor U22808 (N_22808,N_19844,N_17444);
xnor U22809 (N_22809,N_15794,N_15020);
or U22810 (N_22810,N_19871,N_19287);
or U22811 (N_22811,N_16564,N_18079);
and U22812 (N_22812,N_18677,N_19948);
nand U22813 (N_22813,N_16588,N_18143);
and U22814 (N_22814,N_17199,N_17181);
nor U22815 (N_22815,N_19938,N_19642);
nor U22816 (N_22816,N_15280,N_17628);
nand U22817 (N_22817,N_17222,N_18732);
nand U22818 (N_22818,N_15415,N_18923);
nand U22819 (N_22819,N_16748,N_16307);
nand U22820 (N_22820,N_17308,N_17418);
nand U22821 (N_22821,N_15363,N_15909);
nand U22822 (N_22822,N_18912,N_19328);
and U22823 (N_22823,N_17953,N_16582);
xnor U22824 (N_22824,N_15932,N_15757);
nand U22825 (N_22825,N_15198,N_19710);
nand U22826 (N_22826,N_15203,N_17938);
xor U22827 (N_22827,N_18265,N_18908);
xnor U22828 (N_22828,N_19167,N_19333);
nand U22829 (N_22829,N_19588,N_18777);
nor U22830 (N_22830,N_17873,N_17962);
nand U22831 (N_22831,N_16371,N_17467);
nand U22832 (N_22832,N_16430,N_17742);
nand U22833 (N_22833,N_19278,N_15288);
or U22834 (N_22834,N_16546,N_15341);
xnor U22835 (N_22835,N_16380,N_19076);
nand U22836 (N_22836,N_16507,N_18563);
and U22837 (N_22837,N_18365,N_16521);
xor U22838 (N_22838,N_19865,N_16727);
and U22839 (N_22839,N_16058,N_18441);
xnor U22840 (N_22840,N_19656,N_18383);
xnor U22841 (N_22841,N_18019,N_16593);
and U22842 (N_22842,N_16538,N_19777);
or U22843 (N_22843,N_15073,N_16413);
or U22844 (N_22844,N_16952,N_19994);
or U22845 (N_22845,N_16897,N_19528);
nor U22846 (N_22846,N_16766,N_17961);
and U22847 (N_22847,N_15713,N_19005);
nor U22848 (N_22848,N_16728,N_16057);
or U22849 (N_22849,N_17164,N_19462);
xnor U22850 (N_22850,N_17164,N_15861);
nand U22851 (N_22851,N_18425,N_17998);
nand U22852 (N_22852,N_16436,N_16157);
or U22853 (N_22853,N_17329,N_19526);
nor U22854 (N_22854,N_16846,N_17923);
nor U22855 (N_22855,N_15644,N_18139);
nor U22856 (N_22856,N_17406,N_15910);
nand U22857 (N_22857,N_18601,N_18327);
nor U22858 (N_22858,N_16428,N_15182);
xor U22859 (N_22859,N_17527,N_19944);
nor U22860 (N_22860,N_16757,N_15416);
or U22861 (N_22861,N_19918,N_16352);
nor U22862 (N_22862,N_16093,N_19590);
nand U22863 (N_22863,N_16482,N_18336);
and U22864 (N_22864,N_16908,N_18968);
nor U22865 (N_22865,N_18912,N_17081);
nand U22866 (N_22866,N_19927,N_18578);
nor U22867 (N_22867,N_18452,N_19698);
xnor U22868 (N_22868,N_15779,N_15028);
or U22869 (N_22869,N_15217,N_17353);
or U22870 (N_22870,N_19915,N_15218);
nor U22871 (N_22871,N_17815,N_16566);
nor U22872 (N_22872,N_17700,N_18946);
and U22873 (N_22873,N_19305,N_15591);
or U22874 (N_22874,N_19360,N_17016);
xor U22875 (N_22875,N_16794,N_16130);
xnor U22876 (N_22876,N_16930,N_16474);
xor U22877 (N_22877,N_15419,N_17501);
or U22878 (N_22878,N_17645,N_17853);
xnor U22879 (N_22879,N_17722,N_17211);
nor U22880 (N_22880,N_16890,N_16364);
nand U22881 (N_22881,N_17736,N_15562);
xnor U22882 (N_22882,N_17418,N_16419);
or U22883 (N_22883,N_15301,N_18377);
nor U22884 (N_22884,N_19245,N_18651);
nor U22885 (N_22885,N_15435,N_18430);
and U22886 (N_22886,N_18656,N_17487);
and U22887 (N_22887,N_17607,N_18025);
xnor U22888 (N_22888,N_18636,N_19878);
xor U22889 (N_22889,N_17516,N_15811);
and U22890 (N_22890,N_17496,N_15590);
or U22891 (N_22891,N_16261,N_16724);
nor U22892 (N_22892,N_18371,N_17038);
and U22893 (N_22893,N_19773,N_19575);
nand U22894 (N_22894,N_15244,N_19103);
and U22895 (N_22895,N_19849,N_16483);
and U22896 (N_22896,N_16843,N_19739);
or U22897 (N_22897,N_15386,N_16945);
nor U22898 (N_22898,N_18846,N_19358);
xor U22899 (N_22899,N_19418,N_16776);
or U22900 (N_22900,N_19984,N_18938);
or U22901 (N_22901,N_19949,N_17733);
and U22902 (N_22902,N_17264,N_17463);
nand U22903 (N_22903,N_19197,N_19874);
or U22904 (N_22904,N_18994,N_16426);
nand U22905 (N_22905,N_16101,N_18456);
nor U22906 (N_22906,N_18005,N_18342);
nor U22907 (N_22907,N_19785,N_17010);
or U22908 (N_22908,N_19073,N_15488);
nand U22909 (N_22909,N_16305,N_15779);
or U22910 (N_22910,N_18885,N_19661);
and U22911 (N_22911,N_16358,N_15521);
nand U22912 (N_22912,N_15088,N_15850);
nor U22913 (N_22913,N_15275,N_17553);
or U22914 (N_22914,N_15175,N_17125);
and U22915 (N_22915,N_17067,N_15993);
nor U22916 (N_22916,N_16970,N_19683);
or U22917 (N_22917,N_17380,N_15524);
nor U22918 (N_22918,N_17943,N_19457);
xnor U22919 (N_22919,N_19264,N_19740);
or U22920 (N_22920,N_19245,N_15371);
or U22921 (N_22921,N_17883,N_17372);
or U22922 (N_22922,N_18807,N_18338);
nor U22923 (N_22923,N_19517,N_19701);
and U22924 (N_22924,N_18176,N_15968);
xnor U22925 (N_22925,N_19850,N_18238);
or U22926 (N_22926,N_15319,N_19877);
nor U22927 (N_22927,N_18534,N_19801);
nand U22928 (N_22928,N_15204,N_16891);
xnor U22929 (N_22929,N_17286,N_15250);
and U22930 (N_22930,N_17200,N_15616);
or U22931 (N_22931,N_16750,N_19118);
and U22932 (N_22932,N_15418,N_16416);
and U22933 (N_22933,N_18854,N_19163);
xor U22934 (N_22934,N_15083,N_16803);
xnor U22935 (N_22935,N_18987,N_18661);
or U22936 (N_22936,N_19081,N_15510);
nor U22937 (N_22937,N_17693,N_16889);
or U22938 (N_22938,N_17425,N_16815);
and U22939 (N_22939,N_17244,N_18925);
nand U22940 (N_22940,N_15856,N_18774);
and U22941 (N_22941,N_16509,N_18889);
nor U22942 (N_22942,N_15602,N_15812);
xnor U22943 (N_22943,N_17833,N_16587);
or U22944 (N_22944,N_18341,N_17358);
or U22945 (N_22945,N_18775,N_19678);
nand U22946 (N_22946,N_19959,N_15694);
xnor U22947 (N_22947,N_17753,N_19339);
nor U22948 (N_22948,N_18963,N_17786);
nand U22949 (N_22949,N_19740,N_16919);
nand U22950 (N_22950,N_16910,N_16060);
and U22951 (N_22951,N_19958,N_19212);
or U22952 (N_22952,N_19708,N_16496);
or U22953 (N_22953,N_17889,N_17402);
xor U22954 (N_22954,N_17692,N_17825);
or U22955 (N_22955,N_15278,N_18183);
and U22956 (N_22956,N_18577,N_17801);
and U22957 (N_22957,N_16588,N_18291);
and U22958 (N_22958,N_18585,N_17111);
nor U22959 (N_22959,N_15196,N_16805);
or U22960 (N_22960,N_19619,N_17322);
and U22961 (N_22961,N_17040,N_18172);
xnor U22962 (N_22962,N_15302,N_18238);
nor U22963 (N_22963,N_15773,N_16006);
xor U22964 (N_22964,N_17974,N_17056);
and U22965 (N_22965,N_17239,N_16246);
or U22966 (N_22966,N_18481,N_16083);
nor U22967 (N_22967,N_16605,N_17562);
nor U22968 (N_22968,N_15194,N_18284);
nor U22969 (N_22969,N_17773,N_16036);
and U22970 (N_22970,N_19990,N_16774);
xor U22971 (N_22971,N_19312,N_17462);
and U22972 (N_22972,N_18681,N_17925);
or U22973 (N_22973,N_19391,N_18019);
or U22974 (N_22974,N_15189,N_16149);
and U22975 (N_22975,N_17741,N_15598);
nor U22976 (N_22976,N_17332,N_18676);
xnor U22977 (N_22977,N_19500,N_19677);
and U22978 (N_22978,N_17239,N_15389);
nand U22979 (N_22979,N_19727,N_15420);
nand U22980 (N_22980,N_18398,N_15139);
nor U22981 (N_22981,N_15924,N_15163);
xnor U22982 (N_22982,N_15742,N_16821);
or U22983 (N_22983,N_18454,N_16848);
nand U22984 (N_22984,N_17588,N_15336);
nor U22985 (N_22985,N_19542,N_15433);
nor U22986 (N_22986,N_17749,N_19075);
xnor U22987 (N_22987,N_16278,N_18439);
nor U22988 (N_22988,N_18581,N_16597);
xnor U22989 (N_22989,N_15471,N_18287);
and U22990 (N_22990,N_18576,N_18648);
xnor U22991 (N_22991,N_17959,N_15674);
xnor U22992 (N_22992,N_16675,N_18106);
xor U22993 (N_22993,N_18811,N_19599);
and U22994 (N_22994,N_18478,N_18282);
xnor U22995 (N_22995,N_16276,N_15190);
xor U22996 (N_22996,N_16820,N_19933);
or U22997 (N_22997,N_18138,N_15279);
nand U22998 (N_22998,N_17425,N_18720);
nor U22999 (N_22999,N_17380,N_18329);
nor U23000 (N_23000,N_16590,N_18942);
nor U23001 (N_23001,N_15700,N_17676);
nor U23002 (N_23002,N_18792,N_17945);
and U23003 (N_23003,N_17861,N_19761);
and U23004 (N_23004,N_19557,N_18981);
nor U23005 (N_23005,N_16072,N_17128);
nand U23006 (N_23006,N_17718,N_18613);
nor U23007 (N_23007,N_18806,N_19270);
and U23008 (N_23008,N_19763,N_15688);
nand U23009 (N_23009,N_19538,N_19066);
xnor U23010 (N_23010,N_17706,N_19209);
and U23011 (N_23011,N_15585,N_17310);
or U23012 (N_23012,N_17494,N_19039);
and U23013 (N_23013,N_18488,N_19176);
nand U23014 (N_23014,N_19290,N_17366);
xor U23015 (N_23015,N_16369,N_19892);
xor U23016 (N_23016,N_15805,N_15224);
or U23017 (N_23017,N_15050,N_18363);
nand U23018 (N_23018,N_15081,N_16268);
or U23019 (N_23019,N_18987,N_17862);
and U23020 (N_23020,N_16849,N_15588);
or U23021 (N_23021,N_15303,N_15627);
or U23022 (N_23022,N_17668,N_16578);
and U23023 (N_23023,N_17913,N_17488);
nand U23024 (N_23024,N_18804,N_15539);
nand U23025 (N_23025,N_15087,N_16807);
nand U23026 (N_23026,N_19106,N_15045);
and U23027 (N_23027,N_16440,N_17507);
or U23028 (N_23028,N_17320,N_18074);
xnor U23029 (N_23029,N_17295,N_18433);
or U23030 (N_23030,N_15776,N_19939);
or U23031 (N_23031,N_16601,N_15428);
nand U23032 (N_23032,N_16218,N_16302);
xor U23033 (N_23033,N_18134,N_19882);
xnor U23034 (N_23034,N_17495,N_16180);
nand U23035 (N_23035,N_19790,N_19209);
or U23036 (N_23036,N_15556,N_17727);
and U23037 (N_23037,N_18454,N_15358);
or U23038 (N_23038,N_18955,N_18468);
xor U23039 (N_23039,N_19066,N_15975);
nor U23040 (N_23040,N_15512,N_15226);
nand U23041 (N_23041,N_15707,N_17820);
nand U23042 (N_23042,N_17479,N_18406);
nand U23043 (N_23043,N_19663,N_15708);
or U23044 (N_23044,N_16305,N_19215);
and U23045 (N_23045,N_19832,N_18958);
nand U23046 (N_23046,N_16470,N_16093);
xor U23047 (N_23047,N_19532,N_16453);
xnor U23048 (N_23048,N_18147,N_15834);
and U23049 (N_23049,N_19645,N_19560);
nand U23050 (N_23050,N_19247,N_15543);
xnor U23051 (N_23051,N_16485,N_15610);
and U23052 (N_23052,N_15663,N_15672);
or U23053 (N_23053,N_19205,N_15327);
or U23054 (N_23054,N_18722,N_18422);
or U23055 (N_23055,N_17174,N_16942);
and U23056 (N_23056,N_19049,N_16380);
nand U23057 (N_23057,N_17994,N_17631);
and U23058 (N_23058,N_19613,N_19369);
xnor U23059 (N_23059,N_19142,N_18201);
xnor U23060 (N_23060,N_15888,N_16797);
xor U23061 (N_23061,N_19469,N_18639);
and U23062 (N_23062,N_19269,N_18864);
and U23063 (N_23063,N_18936,N_17676);
and U23064 (N_23064,N_16133,N_18066);
and U23065 (N_23065,N_17201,N_18893);
and U23066 (N_23066,N_18626,N_16408);
or U23067 (N_23067,N_17755,N_17966);
xnor U23068 (N_23068,N_16279,N_17065);
xor U23069 (N_23069,N_18566,N_18583);
and U23070 (N_23070,N_18343,N_15639);
nor U23071 (N_23071,N_18047,N_19713);
nand U23072 (N_23072,N_16464,N_15888);
nand U23073 (N_23073,N_19717,N_17856);
nor U23074 (N_23074,N_17569,N_15735);
nand U23075 (N_23075,N_18415,N_18510);
or U23076 (N_23076,N_18808,N_18006);
nor U23077 (N_23077,N_17121,N_16594);
nand U23078 (N_23078,N_19374,N_16181);
or U23079 (N_23079,N_17435,N_16670);
or U23080 (N_23080,N_17579,N_18900);
xor U23081 (N_23081,N_19759,N_17922);
and U23082 (N_23082,N_15380,N_19939);
xnor U23083 (N_23083,N_15645,N_15621);
nand U23084 (N_23084,N_19900,N_16806);
nor U23085 (N_23085,N_19895,N_16611);
nand U23086 (N_23086,N_15170,N_17563);
and U23087 (N_23087,N_18848,N_15811);
xor U23088 (N_23088,N_15427,N_19215);
nand U23089 (N_23089,N_18100,N_15130);
xnor U23090 (N_23090,N_16878,N_15614);
or U23091 (N_23091,N_15092,N_16796);
or U23092 (N_23092,N_15013,N_16399);
nand U23093 (N_23093,N_15544,N_18380);
or U23094 (N_23094,N_19857,N_15946);
nand U23095 (N_23095,N_15939,N_15619);
or U23096 (N_23096,N_15952,N_15738);
or U23097 (N_23097,N_15597,N_19685);
nand U23098 (N_23098,N_17119,N_16307);
or U23099 (N_23099,N_16092,N_18340);
nor U23100 (N_23100,N_17004,N_17018);
and U23101 (N_23101,N_17750,N_16082);
nand U23102 (N_23102,N_16540,N_16068);
xor U23103 (N_23103,N_18755,N_16092);
xor U23104 (N_23104,N_16692,N_15427);
nand U23105 (N_23105,N_19923,N_16279);
nand U23106 (N_23106,N_18986,N_17603);
or U23107 (N_23107,N_18744,N_17234);
xor U23108 (N_23108,N_16520,N_17032);
or U23109 (N_23109,N_19909,N_17790);
and U23110 (N_23110,N_19089,N_19682);
nand U23111 (N_23111,N_19059,N_19029);
xnor U23112 (N_23112,N_15105,N_16458);
nor U23113 (N_23113,N_16709,N_18114);
nor U23114 (N_23114,N_15155,N_16498);
xnor U23115 (N_23115,N_16036,N_17770);
nand U23116 (N_23116,N_16778,N_19246);
or U23117 (N_23117,N_19978,N_16321);
nor U23118 (N_23118,N_15670,N_16264);
nand U23119 (N_23119,N_18219,N_17680);
nand U23120 (N_23120,N_16965,N_19503);
nand U23121 (N_23121,N_19053,N_19477);
nand U23122 (N_23122,N_17717,N_18500);
nand U23123 (N_23123,N_19118,N_18997);
or U23124 (N_23124,N_15731,N_15644);
xnor U23125 (N_23125,N_15505,N_18979);
or U23126 (N_23126,N_17764,N_16562);
xor U23127 (N_23127,N_15632,N_15901);
nand U23128 (N_23128,N_18742,N_19704);
and U23129 (N_23129,N_17091,N_18868);
nand U23130 (N_23130,N_18027,N_16286);
and U23131 (N_23131,N_17997,N_17371);
nor U23132 (N_23132,N_17992,N_17558);
or U23133 (N_23133,N_19599,N_19056);
nand U23134 (N_23134,N_16157,N_16831);
or U23135 (N_23135,N_19502,N_17974);
nor U23136 (N_23136,N_19826,N_16356);
nand U23137 (N_23137,N_18066,N_17852);
xor U23138 (N_23138,N_15929,N_16716);
xor U23139 (N_23139,N_18508,N_19914);
xnor U23140 (N_23140,N_19065,N_17280);
or U23141 (N_23141,N_16378,N_17087);
and U23142 (N_23142,N_15641,N_17561);
xnor U23143 (N_23143,N_18971,N_18335);
nor U23144 (N_23144,N_18340,N_18113);
nor U23145 (N_23145,N_17954,N_17808);
nor U23146 (N_23146,N_17340,N_18500);
nand U23147 (N_23147,N_18260,N_19784);
or U23148 (N_23148,N_18647,N_15677);
xor U23149 (N_23149,N_15778,N_19890);
or U23150 (N_23150,N_15533,N_15578);
xnor U23151 (N_23151,N_18131,N_18062);
or U23152 (N_23152,N_15289,N_17497);
or U23153 (N_23153,N_16536,N_18767);
xnor U23154 (N_23154,N_19142,N_15508);
nor U23155 (N_23155,N_19362,N_15804);
and U23156 (N_23156,N_17518,N_18446);
and U23157 (N_23157,N_19787,N_19966);
or U23158 (N_23158,N_19268,N_15714);
or U23159 (N_23159,N_18485,N_19980);
nor U23160 (N_23160,N_18191,N_15166);
or U23161 (N_23161,N_16137,N_17839);
nor U23162 (N_23162,N_16531,N_18697);
and U23163 (N_23163,N_17138,N_18927);
nand U23164 (N_23164,N_18997,N_17619);
xnor U23165 (N_23165,N_19312,N_17666);
nor U23166 (N_23166,N_15907,N_16825);
nor U23167 (N_23167,N_15949,N_16884);
and U23168 (N_23168,N_18566,N_16926);
nor U23169 (N_23169,N_19524,N_19485);
xor U23170 (N_23170,N_19752,N_16827);
nand U23171 (N_23171,N_16887,N_18340);
nand U23172 (N_23172,N_16754,N_18422);
nand U23173 (N_23173,N_17950,N_18529);
and U23174 (N_23174,N_17605,N_16780);
xor U23175 (N_23175,N_17102,N_19677);
nor U23176 (N_23176,N_15754,N_18444);
nor U23177 (N_23177,N_16094,N_15645);
or U23178 (N_23178,N_18277,N_19438);
nor U23179 (N_23179,N_19441,N_19579);
nand U23180 (N_23180,N_15947,N_18585);
or U23181 (N_23181,N_15243,N_17807);
or U23182 (N_23182,N_15490,N_19861);
nor U23183 (N_23183,N_15927,N_19416);
nor U23184 (N_23184,N_15901,N_17950);
xor U23185 (N_23185,N_17805,N_17540);
xor U23186 (N_23186,N_17081,N_17857);
and U23187 (N_23187,N_16869,N_17771);
xnor U23188 (N_23188,N_18784,N_18587);
nor U23189 (N_23189,N_17897,N_15243);
or U23190 (N_23190,N_17950,N_17716);
nor U23191 (N_23191,N_16454,N_16312);
nor U23192 (N_23192,N_17750,N_16250);
and U23193 (N_23193,N_15609,N_17179);
nor U23194 (N_23194,N_17508,N_18048);
nand U23195 (N_23195,N_19733,N_15501);
or U23196 (N_23196,N_19610,N_16485);
nand U23197 (N_23197,N_19027,N_15049);
or U23198 (N_23198,N_16741,N_18205);
nor U23199 (N_23199,N_15299,N_15228);
nor U23200 (N_23200,N_16089,N_18090);
nor U23201 (N_23201,N_17898,N_16873);
and U23202 (N_23202,N_17163,N_18453);
nand U23203 (N_23203,N_16272,N_18383);
nor U23204 (N_23204,N_19563,N_17736);
xnor U23205 (N_23205,N_18764,N_17477);
and U23206 (N_23206,N_16314,N_17279);
and U23207 (N_23207,N_18685,N_16972);
xor U23208 (N_23208,N_15701,N_16130);
nand U23209 (N_23209,N_19445,N_15215);
nor U23210 (N_23210,N_17482,N_19221);
nor U23211 (N_23211,N_16101,N_16479);
or U23212 (N_23212,N_16151,N_16693);
nand U23213 (N_23213,N_16838,N_16489);
and U23214 (N_23214,N_15374,N_17610);
and U23215 (N_23215,N_15627,N_16896);
xor U23216 (N_23216,N_15341,N_18840);
nor U23217 (N_23217,N_15480,N_17062);
xor U23218 (N_23218,N_16638,N_16681);
nand U23219 (N_23219,N_18738,N_19460);
and U23220 (N_23220,N_16559,N_16933);
or U23221 (N_23221,N_19469,N_16178);
and U23222 (N_23222,N_17097,N_15809);
nor U23223 (N_23223,N_15703,N_16824);
xnor U23224 (N_23224,N_18027,N_18445);
nor U23225 (N_23225,N_15445,N_15059);
or U23226 (N_23226,N_19057,N_18631);
and U23227 (N_23227,N_16866,N_15671);
xor U23228 (N_23228,N_15616,N_16735);
or U23229 (N_23229,N_15507,N_18133);
and U23230 (N_23230,N_18584,N_18963);
nand U23231 (N_23231,N_16681,N_16354);
nor U23232 (N_23232,N_18839,N_16998);
nor U23233 (N_23233,N_17939,N_19247);
and U23234 (N_23234,N_16336,N_19630);
and U23235 (N_23235,N_15056,N_16186);
and U23236 (N_23236,N_17581,N_15349);
and U23237 (N_23237,N_15442,N_17126);
xor U23238 (N_23238,N_18502,N_19713);
and U23239 (N_23239,N_16146,N_16238);
or U23240 (N_23240,N_18829,N_18293);
nand U23241 (N_23241,N_19523,N_15400);
xor U23242 (N_23242,N_15293,N_15290);
nor U23243 (N_23243,N_17284,N_16342);
or U23244 (N_23244,N_18468,N_17086);
and U23245 (N_23245,N_18728,N_18703);
nor U23246 (N_23246,N_17798,N_18752);
nand U23247 (N_23247,N_18546,N_15645);
nor U23248 (N_23248,N_18074,N_15097);
and U23249 (N_23249,N_18880,N_16905);
or U23250 (N_23250,N_15633,N_16804);
xnor U23251 (N_23251,N_15757,N_17960);
nor U23252 (N_23252,N_17687,N_17760);
nor U23253 (N_23253,N_16279,N_15462);
or U23254 (N_23254,N_19506,N_19355);
nand U23255 (N_23255,N_19351,N_16971);
and U23256 (N_23256,N_17998,N_17804);
nand U23257 (N_23257,N_17707,N_18504);
and U23258 (N_23258,N_18915,N_15450);
nand U23259 (N_23259,N_15743,N_19563);
or U23260 (N_23260,N_16698,N_15721);
xnor U23261 (N_23261,N_19805,N_19631);
nand U23262 (N_23262,N_19119,N_19595);
xor U23263 (N_23263,N_16995,N_18828);
or U23264 (N_23264,N_18024,N_19992);
or U23265 (N_23265,N_18543,N_19751);
nor U23266 (N_23266,N_18848,N_19755);
xor U23267 (N_23267,N_18917,N_18969);
nor U23268 (N_23268,N_15641,N_19572);
and U23269 (N_23269,N_17918,N_16351);
nand U23270 (N_23270,N_15655,N_19941);
or U23271 (N_23271,N_19971,N_18388);
nor U23272 (N_23272,N_15711,N_18096);
and U23273 (N_23273,N_15851,N_19820);
and U23274 (N_23274,N_19620,N_15964);
or U23275 (N_23275,N_17193,N_18918);
nand U23276 (N_23276,N_15965,N_19904);
and U23277 (N_23277,N_15143,N_15950);
nor U23278 (N_23278,N_17971,N_15623);
or U23279 (N_23279,N_15065,N_17232);
nor U23280 (N_23280,N_19622,N_16335);
nand U23281 (N_23281,N_16684,N_16163);
xnor U23282 (N_23282,N_15545,N_19313);
or U23283 (N_23283,N_17708,N_16275);
xor U23284 (N_23284,N_18809,N_18168);
xnor U23285 (N_23285,N_15589,N_17704);
nor U23286 (N_23286,N_19934,N_19168);
or U23287 (N_23287,N_19022,N_16354);
or U23288 (N_23288,N_18782,N_16804);
nor U23289 (N_23289,N_15169,N_16195);
or U23290 (N_23290,N_19378,N_19952);
or U23291 (N_23291,N_19610,N_17344);
and U23292 (N_23292,N_16237,N_19696);
and U23293 (N_23293,N_19514,N_19813);
nand U23294 (N_23294,N_17890,N_18259);
and U23295 (N_23295,N_16573,N_18760);
xnor U23296 (N_23296,N_16583,N_17823);
nor U23297 (N_23297,N_16120,N_18034);
nand U23298 (N_23298,N_19156,N_16741);
or U23299 (N_23299,N_17819,N_16446);
and U23300 (N_23300,N_17140,N_16399);
xor U23301 (N_23301,N_18625,N_16128);
or U23302 (N_23302,N_17072,N_17829);
and U23303 (N_23303,N_17714,N_16683);
or U23304 (N_23304,N_16309,N_17760);
nor U23305 (N_23305,N_15776,N_15497);
and U23306 (N_23306,N_18571,N_15132);
and U23307 (N_23307,N_19101,N_17169);
xor U23308 (N_23308,N_19954,N_18670);
and U23309 (N_23309,N_15372,N_16640);
nor U23310 (N_23310,N_17019,N_15179);
and U23311 (N_23311,N_19093,N_19600);
nor U23312 (N_23312,N_19709,N_17046);
or U23313 (N_23313,N_15203,N_16653);
nor U23314 (N_23314,N_18506,N_15701);
or U23315 (N_23315,N_15339,N_15728);
or U23316 (N_23316,N_18337,N_19878);
xor U23317 (N_23317,N_15104,N_16157);
and U23318 (N_23318,N_16377,N_18575);
and U23319 (N_23319,N_18744,N_18542);
and U23320 (N_23320,N_15775,N_16012);
and U23321 (N_23321,N_18997,N_17389);
and U23322 (N_23322,N_16512,N_19484);
nand U23323 (N_23323,N_18887,N_18357);
xor U23324 (N_23324,N_18449,N_16743);
nand U23325 (N_23325,N_15948,N_15671);
xnor U23326 (N_23326,N_19602,N_18118);
xor U23327 (N_23327,N_15709,N_19234);
xnor U23328 (N_23328,N_19509,N_19599);
or U23329 (N_23329,N_17325,N_18047);
nor U23330 (N_23330,N_18809,N_18949);
or U23331 (N_23331,N_18034,N_19259);
or U23332 (N_23332,N_18549,N_18529);
and U23333 (N_23333,N_15408,N_19860);
xor U23334 (N_23334,N_15427,N_18328);
nor U23335 (N_23335,N_19103,N_17220);
xnor U23336 (N_23336,N_15674,N_16563);
or U23337 (N_23337,N_15942,N_15278);
nor U23338 (N_23338,N_19569,N_18680);
xor U23339 (N_23339,N_18995,N_15897);
nor U23340 (N_23340,N_19290,N_18729);
xnor U23341 (N_23341,N_18989,N_19737);
and U23342 (N_23342,N_19501,N_16684);
and U23343 (N_23343,N_16627,N_16734);
nand U23344 (N_23344,N_19251,N_17088);
nand U23345 (N_23345,N_19352,N_16439);
nand U23346 (N_23346,N_16284,N_17660);
xnor U23347 (N_23347,N_15671,N_17890);
and U23348 (N_23348,N_19111,N_18723);
or U23349 (N_23349,N_17339,N_17312);
xnor U23350 (N_23350,N_15053,N_16112);
nand U23351 (N_23351,N_15526,N_15889);
and U23352 (N_23352,N_18941,N_18246);
nand U23353 (N_23353,N_17543,N_19655);
nor U23354 (N_23354,N_19790,N_17520);
and U23355 (N_23355,N_16310,N_19229);
xnor U23356 (N_23356,N_15768,N_17510);
xnor U23357 (N_23357,N_18362,N_18578);
nor U23358 (N_23358,N_16552,N_16934);
and U23359 (N_23359,N_15527,N_15490);
nand U23360 (N_23360,N_18629,N_15657);
and U23361 (N_23361,N_19557,N_17816);
nor U23362 (N_23362,N_19635,N_18612);
and U23363 (N_23363,N_16458,N_19919);
xor U23364 (N_23364,N_19817,N_16680);
xnor U23365 (N_23365,N_16177,N_15439);
nand U23366 (N_23366,N_18729,N_19716);
nor U23367 (N_23367,N_16922,N_17929);
nor U23368 (N_23368,N_18018,N_18399);
nand U23369 (N_23369,N_19061,N_18496);
nor U23370 (N_23370,N_18115,N_16127);
xnor U23371 (N_23371,N_15050,N_15041);
and U23372 (N_23372,N_18343,N_17506);
and U23373 (N_23373,N_16447,N_19125);
and U23374 (N_23374,N_16483,N_19150);
nor U23375 (N_23375,N_19906,N_17848);
xor U23376 (N_23376,N_17609,N_15703);
xnor U23377 (N_23377,N_17605,N_18812);
and U23378 (N_23378,N_15344,N_17561);
xor U23379 (N_23379,N_16859,N_17263);
nor U23380 (N_23380,N_17029,N_18710);
xor U23381 (N_23381,N_19554,N_19151);
xor U23382 (N_23382,N_19265,N_17677);
nand U23383 (N_23383,N_15058,N_15362);
nor U23384 (N_23384,N_16690,N_19928);
nand U23385 (N_23385,N_17644,N_18063);
xnor U23386 (N_23386,N_18966,N_17631);
xnor U23387 (N_23387,N_18332,N_19807);
xnor U23388 (N_23388,N_15552,N_19167);
nor U23389 (N_23389,N_16888,N_17447);
nand U23390 (N_23390,N_18278,N_16813);
xnor U23391 (N_23391,N_18864,N_17550);
nor U23392 (N_23392,N_15308,N_17015);
nand U23393 (N_23393,N_16997,N_17226);
nand U23394 (N_23394,N_17275,N_18013);
and U23395 (N_23395,N_16165,N_17380);
and U23396 (N_23396,N_18324,N_19271);
nand U23397 (N_23397,N_16636,N_18514);
xor U23398 (N_23398,N_16189,N_15768);
xnor U23399 (N_23399,N_19394,N_17984);
and U23400 (N_23400,N_15050,N_16533);
xor U23401 (N_23401,N_16177,N_15921);
xnor U23402 (N_23402,N_16877,N_16232);
and U23403 (N_23403,N_17057,N_18485);
or U23404 (N_23404,N_18129,N_16781);
nor U23405 (N_23405,N_17510,N_15689);
or U23406 (N_23406,N_17802,N_15389);
and U23407 (N_23407,N_16479,N_19676);
nand U23408 (N_23408,N_17455,N_15957);
nor U23409 (N_23409,N_15397,N_17874);
and U23410 (N_23410,N_16018,N_15739);
xnor U23411 (N_23411,N_16854,N_15859);
or U23412 (N_23412,N_17802,N_16627);
nor U23413 (N_23413,N_17603,N_16626);
nor U23414 (N_23414,N_17049,N_16880);
or U23415 (N_23415,N_19884,N_18883);
nor U23416 (N_23416,N_17853,N_16985);
or U23417 (N_23417,N_19161,N_19200);
or U23418 (N_23418,N_15251,N_16445);
or U23419 (N_23419,N_16247,N_19074);
nand U23420 (N_23420,N_19691,N_18773);
or U23421 (N_23421,N_15378,N_18173);
nor U23422 (N_23422,N_19759,N_17885);
and U23423 (N_23423,N_16146,N_15477);
or U23424 (N_23424,N_17320,N_15954);
nand U23425 (N_23425,N_16078,N_19322);
nand U23426 (N_23426,N_15350,N_18755);
nand U23427 (N_23427,N_17386,N_19751);
nor U23428 (N_23428,N_18484,N_16337);
xnor U23429 (N_23429,N_15440,N_16720);
and U23430 (N_23430,N_15377,N_18342);
or U23431 (N_23431,N_18187,N_16502);
xnor U23432 (N_23432,N_15643,N_19746);
or U23433 (N_23433,N_18048,N_17981);
xnor U23434 (N_23434,N_18172,N_17910);
and U23435 (N_23435,N_16149,N_15040);
nor U23436 (N_23436,N_19596,N_19015);
xor U23437 (N_23437,N_18029,N_15318);
and U23438 (N_23438,N_17685,N_15626);
nand U23439 (N_23439,N_16235,N_19338);
xor U23440 (N_23440,N_17017,N_19014);
nor U23441 (N_23441,N_19617,N_17709);
nor U23442 (N_23442,N_15609,N_19618);
xor U23443 (N_23443,N_15449,N_19683);
and U23444 (N_23444,N_15437,N_19893);
nand U23445 (N_23445,N_17502,N_16892);
and U23446 (N_23446,N_17875,N_16080);
nor U23447 (N_23447,N_18377,N_17603);
xor U23448 (N_23448,N_16877,N_15048);
nand U23449 (N_23449,N_15465,N_18614);
xnor U23450 (N_23450,N_15148,N_19666);
nand U23451 (N_23451,N_15475,N_15618);
and U23452 (N_23452,N_15018,N_17074);
and U23453 (N_23453,N_16069,N_16392);
and U23454 (N_23454,N_16922,N_18167);
or U23455 (N_23455,N_16996,N_15374);
nand U23456 (N_23456,N_15376,N_17864);
or U23457 (N_23457,N_18982,N_17409);
and U23458 (N_23458,N_15427,N_16264);
xor U23459 (N_23459,N_15273,N_15561);
nand U23460 (N_23460,N_17819,N_18790);
xnor U23461 (N_23461,N_17938,N_19167);
nand U23462 (N_23462,N_16827,N_16891);
nor U23463 (N_23463,N_19313,N_15888);
and U23464 (N_23464,N_18577,N_16026);
or U23465 (N_23465,N_19270,N_16724);
nor U23466 (N_23466,N_17221,N_19389);
or U23467 (N_23467,N_18153,N_18809);
xnor U23468 (N_23468,N_19366,N_16699);
and U23469 (N_23469,N_16648,N_17461);
xnor U23470 (N_23470,N_19196,N_15668);
nor U23471 (N_23471,N_18755,N_17566);
nor U23472 (N_23472,N_17640,N_17685);
or U23473 (N_23473,N_15105,N_16193);
or U23474 (N_23474,N_16184,N_18236);
xnor U23475 (N_23475,N_19619,N_18287);
and U23476 (N_23476,N_18041,N_18323);
xor U23477 (N_23477,N_16753,N_15336);
nor U23478 (N_23478,N_18218,N_15172);
xor U23479 (N_23479,N_16541,N_16414);
xor U23480 (N_23480,N_16500,N_16749);
nand U23481 (N_23481,N_15134,N_17419);
xor U23482 (N_23482,N_15776,N_15981);
and U23483 (N_23483,N_17376,N_16210);
nor U23484 (N_23484,N_19368,N_18318);
nor U23485 (N_23485,N_19310,N_17536);
and U23486 (N_23486,N_15386,N_18287);
nor U23487 (N_23487,N_17110,N_16949);
or U23488 (N_23488,N_16736,N_17112);
and U23489 (N_23489,N_17482,N_17824);
xnor U23490 (N_23490,N_17686,N_16550);
nand U23491 (N_23491,N_19462,N_19922);
nand U23492 (N_23492,N_18145,N_15180);
or U23493 (N_23493,N_17310,N_16445);
xor U23494 (N_23494,N_16824,N_15691);
and U23495 (N_23495,N_18246,N_16109);
nand U23496 (N_23496,N_17541,N_17893);
nand U23497 (N_23497,N_15195,N_18723);
and U23498 (N_23498,N_17566,N_15080);
nor U23499 (N_23499,N_19603,N_16336);
nand U23500 (N_23500,N_15750,N_18582);
or U23501 (N_23501,N_17345,N_17218);
nand U23502 (N_23502,N_16955,N_18525);
nor U23503 (N_23503,N_15475,N_17126);
or U23504 (N_23504,N_18262,N_17627);
nand U23505 (N_23505,N_17795,N_18353);
nor U23506 (N_23506,N_19564,N_17163);
nand U23507 (N_23507,N_19398,N_17946);
nor U23508 (N_23508,N_15925,N_19584);
nand U23509 (N_23509,N_19026,N_18710);
and U23510 (N_23510,N_16797,N_18484);
xor U23511 (N_23511,N_19960,N_15408);
and U23512 (N_23512,N_19885,N_19149);
nor U23513 (N_23513,N_15889,N_19602);
nand U23514 (N_23514,N_17169,N_16944);
xnor U23515 (N_23515,N_17949,N_19014);
xnor U23516 (N_23516,N_15730,N_18697);
and U23517 (N_23517,N_15399,N_19139);
or U23518 (N_23518,N_19941,N_16083);
and U23519 (N_23519,N_16838,N_15092);
or U23520 (N_23520,N_18319,N_15439);
and U23521 (N_23521,N_17904,N_15874);
or U23522 (N_23522,N_17707,N_16675);
nor U23523 (N_23523,N_18513,N_18953);
or U23524 (N_23524,N_16423,N_19365);
nor U23525 (N_23525,N_19335,N_19148);
nand U23526 (N_23526,N_18776,N_18270);
nor U23527 (N_23527,N_19152,N_17099);
and U23528 (N_23528,N_18632,N_15135);
nand U23529 (N_23529,N_17089,N_18291);
xor U23530 (N_23530,N_19242,N_18285);
and U23531 (N_23531,N_16070,N_18627);
nor U23532 (N_23532,N_15957,N_19544);
and U23533 (N_23533,N_19175,N_15621);
or U23534 (N_23534,N_19676,N_15485);
or U23535 (N_23535,N_17454,N_16795);
and U23536 (N_23536,N_19870,N_16052);
xnor U23537 (N_23537,N_15858,N_16952);
and U23538 (N_23538,N_15017,N_18049);
or U23539 (N_23539,N_16232,N_19871);
xnor U23540 (N_23540,N_15814,N_15223);
nand U23541 (N_23541,N_18918,N_16718);
nand U23542 (N_23542,N_17636,N_16702);
xnor U23543 (N_23543,N_15632,N_17592);
nor U23544 (N_23544,N_17747,N_17443);
and U23545 (N_23545,N_19184,N_15461);
nor U23546 (N_23546,N_15746,N_15141);
or U23547 (N_23547,N_18954,N_19964);
and U23548 (N_23548,N_18784,N_16158);
nand U23549 (N_23549,N_16814,N_18056);
nor U23550 (N_23550,N_15107,N_15633);
and U23551 (N_23551,N_18211,N_16618);
xnor U23552 (N_23552,N_15238,N_18178);
nand U23553 (N_23553,N_15036,N_17285);
nor U23554 (N_23554,N_18628,N_16859);
nor U23555 (N_23555,N_17954,N_16889);
xnor U23556 (N_23556,N_17905,N_19599);
nand U23557 (N_23557,N_17182,N_15890);
and U23558 (N_23558,N_19966,N_16090);
xnor U23559 (N_23559,N_19356,N_16979);
or U23560 (N_23560,N_16453,N_18388);
and U23561 (N_23561,N_17603,N_15415);
and U23562 (N_23562,N_18105,N_15376);
xor U23563 (N_23563,N_16633,N_17289);
or U23564 (N_23564,N_15093,N_15180);
nand U23565 (N_23565,N_19190,N_15931);
or U23566 (N_23566,N_17942,N_18031);
nor U23567 (N_23567,N_17413,N_19824);
or U23568 (N_23568,N_18989,N_19610);
or U23569 (N_23569,N_17475,N_16067);
nor U23570 (N_23570,N_19027,N_15078);
or U23571 (N_23571,N_18989,N_19548);
nand U23572 (N_23572,N_17401,N_17423);
nand U23573 (N_23573,N_17027,N_16213);
nor U23574 (N_23574,N_18152,N_19129);
nand U23575 (N_23575,N_16677,N_19383);
xor U23576 (N_23576,N_18228,N_19871);
nand U23577 (N_23577,N_15754,N_15357);
nand U23578 (N_23578,N_17341,N_16652);
and U23579 (N_23579,N_18425,N_19845);
or U23580 (N_23580,N_19030,N_15255);
or U23581 (N_23581,N_15585,N_18358);
or U23582 (N_23582,N_18669,N_19331);
nor U23583 (N_23583,N_19425,N_18302);
or U23584 (N_23584,N_15575,N_15428);
nor U23585 (N_23585,N_19614,N_18876);
xor U23586 (N_23586,N_17118,N_18207);
nor U23587 (N_23587,N_16735,N_15283);
xor U23588 (N_23588,N_16413,N_15677);
xnor U23589 (N_23589,N_16235,N_16820);
and U23590 (N_23590,N_16954,N_17756);
xor U23591 (N_23591,N_17249,N_16859);
xnor U23592 (N_23592,N_17905,N_17913);
or U23593 (N_23593,N_17904,N_17184);
or U23594 (N_23594,N_16638,N_16547);
and U23595 (N_23595,N_17800,N_16465);
nor U23596 (N_23596,N_16692,N_16766);
xor U23597 (N_23597,N_19739,N_17959);
and U23598 (N_23598,N_18593,N_19121);
and U23599 (N_23599,N_15701,N_17770);
and U23600 (N_23600,N_18323,N_18550);
and U23601 (N_23601,N_19664,N_16641);
nand U23602 (N_23602,N_17320,N_19125);
or U23603 (N_23603,N_17518,N_15677);
and U23604 (N_23604,N_16973,N_19838);
nand U23605 (N_23605,N_15762,N_15045);
and U23606 (N_23606,N_17216,N_17059);
nand U23607 (N_23607,N_15716,N_17695);
and U23608 (N_23608,N_19755,N_16101);
and U23609 (N_23609,N_18746,N_15785);
and U23610 (N_23610,N_19522,N_18768);
nor U23611 (N_23611,N_18919,N_18796);
or U23612 (N_23612,N_15977,N_15423);
nor U23613 (N_23613,N_16297,N_16108);
nor U23614 (N_23614,N_18748,N_18217);
nor U23615 (N_23615,N_15673,N_19208);
nand U23616 (N_23616,N_18660,N_17095);
and U23617 (N_23617,N_16664,N_16253);
xnor U23618 (N_23618,N_18910,N_15566);
or U23619 (N_23619,N_18314,N_15121);
or U23620 (N_23620,N_19867,N_16514);
nand U23621 (N_23621,N_15766,N_15634);
nand U23622 (N_23622,N_18199,N_16751);
nor U23623 (N_23623,N_17641,N_19705);
xor U23624 (N_23624,N_15478,N_15260);
nand U23625 (N_23625,N_18612,N_16067);
xor U23626 (N_23626,N_18962,N_17220);
nand U23627 (N_23627,N_16685,N_17882);
or U23628 (N_23628,N_15551,N_18816);
and U23629 (N_23629,N_16532,N_17069);
nor U23630 (N_23630,N_15217,N_15503);
and U23631 (N_23631,N_19074,N_18755);
or U23632 (N_23632,N_16900,N_16980);
nor U23633 (N_23633,N_15470,N_15032);
xor U23634 (N_23634,N_16701,N_19993);
nand U23635 (N_23635,N_18111,N_19268);
and U23636 (N_23636,N_15337,N_18251);
nand U23637 (N_23637,N_16583,N_18440);
and U23638 (N_23638,N_19409,N_17335);
nor U23639 (N_23639,N_16953,N_15870);
nor U23640 (N_23640,N_15681,N_15921);
nor U23641 (N_23641,N_17638,N_19158);
nor U23642 (N_23642,N_19834,N_15682);
nand U23643 (N_23643,N_19515,N_17161);
and U23644 (N_23644,N_15958,N_15465);
and U23645 (N_23645,N_19859,N_17769);
and U23646 (N_23646,N_18352,N_16857);
and U23647 (N_23647,N_19211,N_19322);
nand U23648 (N_23648,N_16643,N_15703);
nor U23649 (N_23649,N_15394,N_19426);
nor U23650 (N_23650,N_19584,N_16060);
or U23651 (N_23651,N_17096,N_18816);
and U23652 (N_23652,N_15179,N_17485);
xor U23653 (N_23653,N_15415,N_15791);
or U23654 (N_23654,N_17350,N_17897);
and U23655 (N_23655,N_18212,N_15401);
nand U23656 (N_23656,N_18508,N_18405);
xor U23657 (N_23657,N_18156,N_15699);
nand U23658 (N_23658,N_15510,N_17171);
and U23659 (N_23659,N_15681,N_17020);
nand U23660 (N_23660,N_17070,N_19064);
or U23661 (N_23661,N_18713,N_17978);
nand U23662 (N_23662,N_15605,N_18029);
or U23663 (N_23663,N_15507,N_17819);
nor U23664 (N_23664,N_17410,N_18211);
and U23665 (N_23665,N_17542,N_15671);
nand U23666 (N_23666,N_19907,N_17734);
xor U23667 (N_23667,N_19488,N_17844);
xor U23668 (N_23668,N_15814,N_19568);
nor U23669 (N_23669,N_17301,N_17146);
xnor U23670 (N_23670,N_17404,N_19567);
nor U23671 (N_23671,N_15317,N_19212);
xor U23672 (N_23672,N_19388,N_19865);
nor U23673 (N_23673,N_18131,N_15267);
and U23674 (N_23674,N_19457,N_16875);
xnor U23675 (N_23675,N_15186,N_17045);
nand U23676 (N_23676,N_15297,N_18572);
nor U23677 (N_23677,N_17124,N_16157);
and U23678 (N_23678,N_18999,N_15225);
or U23679 (N_23679,N_18200,N_17983);
and U23680 (N_23680,N_15174,N_17933);
xor U23681 (N_23681,N_17124,N_18871);
and U23682 (N_23682,N_17374,N_17347);
and U23683 (N_23683,N_16569,N_19666);
xor U23684 (N_23684,N_18869,N_18979);
xor U23685 (N_23685,N_17216,N_19239);
or U23686 (N_23686,N_15706,N_16767);
nand U23687 (N_23687,N_16160,N_15550);
or U23688 (N_23688,N_19226,N_19500);
and U23689 (N_23689,N_16460,N_19837);
nor U23690 (N_23690,N_15786,N_18228);
and U23691 (N_23691,N_15598,N_16033);
or U23692 (N_23692,N_16052,N_17169);
or U23693 (N_23693,N_16277,N_19223);
or U23694 (N_23694,N_19033,N_15948);
nor U23695 (N_23695,N_15437,N_19536);
nor U23696 (N_23696,N_17977,N_18506);
xor U23697 (N_23697,N_15339,N_19075);
nand U23698 (N_23698,N_18282,N_17300);
or U23699 (N_23699,N_18953,N_19996);
nand U23700 (N_23700,N_18763,N_19405);
and U23701 (N_23701,N_17498,N_15547);
nand U23702 (N_23702,N_15734,N_17764);
and U23703 (N_23703,N_17244,N_15230);
or U23704 (N_23704,N_16660,N_18379);
nand U23705 (N_23705,N_16043,N_19056);
xor U23706 (N_23706,N_15810,N_18415);
nand U23707 (N_23707,N_18869,N_15119);
or U23708 (N_23708,N_19812,N_17394);
nand U23709 (N_23709,N_16316,N_18764);
nor U23710 (N_23710,N_17597,N_15458);
and U23711 (N_23711,N_17288,N_15431);
nand U23712 (N_23712,N_15633,N_18148);
xnor U23713 (N_23713,N_16160,N_18734);
xnor U23714 (N_23714,N_19246,N_19309);
and U23715 (N_23715,N_19585,N_16891);
nor U23716 (N_23716,N_17565,N_17892);
nand U23717 (N_23717,N_19713,N_19841);
and U23718 (N_23718,N_15707,N_19020);
nand U23719 (N_23719,N_16992,N_19030);
and U23720 (N_23720,N_15102,N_16821);
or U23721 (N_23721,N_16080,N_19852);
xnor U23722 (N_23722,N_19329,N_16806);
and U23723 (N_23723,N_18758,N_16650);
or U23724 (N_23724,N_17662,N_16240);
or U23725 (N_23725,N_17540,N_16106);
nor U23726 (N_23726,N_15963,N_18350);
and U23727 (N_23727,N_17742,N_16266);
or U23728 (N_23728,N_16812,N_19445);
nand U23729 (N_23729,N_17539,N_16472);
nand U23730 (N_23730,N_19217,N_15092);
and U23731 (N_23731,N_18136,N_15887);
nand U23732 (N_23732,N_17057,N_16953);
nor U23733 (N_23733,N_17445,N_16999);
nor U23734 (N_23734,N_15171,N_16512);
xnor U23735 (N_23735,N_15351,N_16823);
or U23736 (N_23736,N_16427,N_18302);
xor U23737 (N_23737,N_16375,N_15951);
and U23738 (N_23738,N_19736,N_17222);
and U23739 (N_23739,N_18337,N_15516);
or U23740 (N_23740,N_16792,N_19802);
nand U23741 (N_23741,N_18614,N_19423);
or U23742 (N_23742,N_18663,N_17834);
nand U23743 (N_23743,N_16263,N_19252);
or U23744 (N_23744,N_18549,N_18049);
and U23745 (N_23745,N_15723,N_17267);
or U23746 (N_23746,N_18809,N_16313);
xnor U23747 (N_23747,N_17630,N_17916);
or U23748 (N_23748,N_15946,N_19567);
or U23749 (N_23749,N_17725,N_18088);
nor U23750 (N_23750,N_15401,N_19292);
xor U23751 (N_23751,N_19160,N_19208);
and U23752 (N_23752,N_15138,N_17095);
nor U23753 (N_23753,N_18511,N_19793);
and U23754 (N_23754,N_16797,N_15097);
nor U23755 (N_23755,N_18022,N_15592);
or U23756 (N_23756,N_15960,N_16503);
nand U23757 (N_23757,N_18450,N_17811);
or U23758 (N_23758,N_19264,N_15390);
and U23759 (N_23759,N_15548,N_19960);
or U23760 (N_23760,N_18656,N_19609);
and U23761 (N_23761,N_15546,N_18574);
or U23762 (N_23762,N_19873,N_15928);
or U23763 (N_23763,N_16251,N_15487);
xnor U23764 (N_23764,N_16839,N_18478);
nand U23765 (N_23765,N_18186,N_18614);
xor U23766 (N_23766,N_16553,N_17043);
xnor U23767 (N_23767,N_16993,N_18683);
nand U23768 (N_23768,N_15087,N_17033);
nand U23769 (N_23769,N_15449,N_17306);
or U23770 (N_23770,N_17458,N_17080);
or U23771 (N_23771,N_15186,N_18941);
xor U23772 (N_23772,N_19202,N_18678);
nor U23773 (N_23773,N_15763,N_18473);
xor U23774 (N_23774,N_18331,N_16019);
nand U23775 (N_23775,N_16753,N_15940);
or U23776 (N_23776,N_15435,N_16181);
and U23777 (N_23777,N_19704,N_19392);
and U23778 (N_23778,N_18173,N_16902);
or U23779 (N_23779,N_16477,N_19579);
or U23780 (N_23780,N_17998,N_16280);
xnor U23781 (N_23781,N_19726,N_19497);
or U23782 (N_23782,N_18740,N_19278);
and U23783 (N_23783,N_15646,N_15544);
or U23784 (N_23784,N_19359,N_18536);
and U23785 (N_23785,N_19864,N_16315);
nand U23786 (N_23786,N_18372,N_15505);
xnor U23787 (N_23787,N_17076,N_18597);
xnor U23788 (N_23788,N_19290,N_15566);
nand U23789 (N_23789,N_16941,N_19422);
nor U23790 (N_23790,N_16097,N_15926);
xnor U23791 (N_23791,N_17262,N_19636);
or U23792 (N_23792,N_19009,N_17074);
nand U23793 (N_23793,N_18321,N_19444);
xnor U23794 (N_23794,N_15942,N_19059);
nand U23795 (N_23795,N_19225,N_16854);
and U23796 (N_23796,N_17619,N_17076);
xor U23797 (N_23797,N_15847,N_15162);
nand U23798 (N_23798,N_17282,N_17734);
nand U23799 (N_23799,N_18803,N_18576);
and U23800 (N_23800,N_18445,N_19473);
or U23801 (N_23801,N_19544,N_16409);
nand U23802 (N_23802,N_18900,N_15425);
or U23803 (N_23803,N_18701,N_16249);
and U23804 (N_23804,N_16975,N_15888);
nand U23805 (N_23805,N_18484,N_15558);
nor U23806 (N_23806,N_16248,N_18763);
xor U23807 (N_23807,N_17526,N_17834);
or U23808 (N_23808,N_15299,N_19141);
xor U23809 (N_23809,N_16210,N_15442);
nand U23810 (N_23810,N_16052,N_18490);
nand U23811 (N_23811,N_17205,N_19860);
nand U23812 (N_23812,N_15668,N_18411);
or U23813 (N_23813,N_18133,N_19407);
or U23814 (N_23814,N_16919,N_17948);
and U23815 (N_23815,N_15475,N_16335);
or U23816 (N_23816,N_17018,N_19124);
nor U23817 (N_23817,N_16651,N_16197);
nand U23818 (N_23818,N_16515,N_17444);
xnor U23819 (N_23819,N_18588,N_18975);
nand U23820 (N_23820,N_16848,N_15571);
nand U23821 (N_23821,N_15516,N_16139);
and U23822 (N_23822,N_16085,N_18864);
nand U23823 (N_23823,N_15358,N_15030);
nor U23824 (N_23824,N_19550,N_17914);
nand U23825 (N_23825,N_18262,N_17808);
and U23826 (N_23826,N_18424,N_18288);
and U23827 (N_23827,N_15716,N_17153);
nand U23828 (N_23828,N_18540,N_15613);
or U23829 (N_23829,N_19573,N_16798);
or U23830 (N_23830,N_15866,N_15484);
nand U23831 (N_23831,N_17325,N_19865);
and U23832 (N_23832,N_19642,N_18053);
nor U23833 (N_23833,N_18763,N_16659);
or U23834 (N_23834,N_19227,N_19216);
and U23835 (N_23835,N_15293,N_15306);
or U23836 (N_23836,N_17404,N_17333);
nand U23837 (N_23837,N_19301,N_18400);
nand U23838 (N_23838,N_18002,N_16783);
or U23839 (N_23839,N_16990,N_16560);
nor U23840 (N_23840,N_18304,N_18290);
nor U23841 (N_23841,N_19431,N_17136);
or U23842 (N_23842,N_17792,N_17045);
nor U23843 (N_23843,N_16449,N_15355);
and U23844 (N_23844,N_18893,N_19772);
nor U23845 (N_23845,N_18657,N_16796);
or U23846 (N_23846,N_17586,N_15852);
nor U23847 (N_23847,N_16870,N_15499);
and U23848 (N_23848,N_16129,N_15498);
and U23849 (N_23849,N_18309,N_16885);
nand U23850 (N_23850,N_16537,N_15726);
nand U23851 (N_23851,N_16323,N_16783);
or U23852 (N_23852,N_18743,N_18680);
nor U23853 (N_23853,N_19895,N_19796);
nor U23854 (N_23854,N_17365,N_19356);
or U23855 (N_23855,N_16006,N_19011);
xor U23856 (N_23856,N_19139,N_17882);
or U23857 (N_23857,N_19504,N_19974);
nand U23858 (N_23858,N_19524,N_16296);
xnor U23859 (N_23859,N_15957,N_19419);
and U23860 (N_23860,N_15221,N_18019);
or U23861 (N_23861,N_16442,N_16625);
or U23862 (N_23862,N_19762,N_19400);
and U23863 (N_23863,N_19809,N_15452);
nand U23864 (N_23864,N_16210,N_18245);
nor U23865 (N_23865,N_18462,N_18346);
nor U23866 (N_23866,N_19273,N_18159);
or U23867 (N_23867,N_15028,N_15928);
nand U23868 (N_23868,N_18487,N_19782);
and U23869 (N_23869,N_16356,N_15309);
nand U23870 (N_23870,N_18686,N_16314);
nand U23871 (N_23871,N_17846,N_17120);
nor U23872 (N_23872,N_16066,N_17413);
nor U23873 (N_23873,N_15509,N_19502);
nand U23874 (N_23874,N_17901,N_16313);
or U23875 (N_23875,N_19622,N_19270);
or U23876 (N_23876,N_19678,N_15006);
and U23877 (N_23877,N_16639,N_19190);
xor U23878 (N_23878,N_16187,N_19184);
or U23879 (N_23879,N_19734,N_18391);
nor U23880 (N_23880,N_19916,N_19889);
and U23881 (N_23881,N_19496,N_19736);
xnor U23882 (N_23882,N_16357,N_17357);
nor U23883 (N_23883,N_19702,N_19641);
nor U23884 (N_23884,N_16882,N_16786);
or U23885 (N_23885,N_18341,N_16058);
and U23886 (N_23886,N_18804,N_17643);
xnor U23887 (N_23887,N_18218,N_18123);
xnor U23888 (N_23888,N_15340,N_15408);
or U23889 (N_23889,N_16239,N_16295);
nand U23890 (N_23890,N_15750,N_18152);
xnor U23891 (N_23891,N_16482,N_19355);
xor U23892 (N_23892,N_19562,N_19229);
nor U23893 (N_23893,N_17848,N_17593);
or U23894 (N_23894,N_18648,N_18464);
nand U23895 (N_23895,N_15494,N_16212);
and U23896 (N_23896,N_18210,N_16933);
nand U23897 (N_23897,N_16397,N_18496);
xor U23898 (N_23898,N_16043,N_18951);
and U23899 (N_23899,N_18268,N_16674);
or U23900 (N_23900,N_18657,N_19054);
xor U23901 (N_23901,N_16691,N_19483);
and U23902 (N_23902,N_17562,N_15731);
nand U23903 (N_23903,N_18834,N_15120);
xnor U23904 (N_23904,N_15109,N_17943);
and U23905 (N_23905,N_17642,N_18018);
and U23906 (N_23906,N_17765,N_15520);
or U23907 (N_23907,N_15524,N_15681);
or U23908 (N_23908,N_19615,N_15533);
xnor U23909 (N_23909,N_19865,N_15722);
xor U23910 (N_23910,N_17878,N_16629);
nand U23911 (N_23911,N_17687,N_15620);
nor U23912 (N_23912,N_17611,N_16285);
nand U23913 (N_23913,N_16109,N_18699);
nor U23914 (N_23914,N_17794,N_19749);
nor U23915 (N_23915,N_15447,N_17348);
and U23916 (N_23916,N_18524,N_16525);
xor U23917 (N_23917,N_19644,N_15316);
and U23918 (N_23918,N_17593,N_18721);
and U23919 (N_23919,N_19805,N_19143);
or U23920 (N_23920,N_16365,N_19722);
and U23921 (N_23921,N_17801,N_15499);
nor U23922 (N_23922,N_16222,N_18165);
nor U23923 (N_23923,N_16342,N_17434);
xnor U23924 (N_23924,N_17437,N_15885);
or U23925 (N_23925,N_17198,N_19095);
or U23926 (N_23926,N_17903,N_15439);
and U23927 (N_23927,N_16345,N_17417);
and U23928 (N_23928,N_18990,N_17162);
nor U23929 (N_23929,N_19355,N_18268);
and U23930 (N_23930,N_16985,N_19338);
or U23931 (N_23931,N_15840,N_17044);
and U23932 (N_23932,N_15215,N_18770);
xor U23933 (N_23933,N_15986,N_18661);
xnor U23934 (N_23934,N_17108,N_19381);
and U23935 (N_23935,N_19668,N_18261);
and U23936 (N_23936,N_19191,N_18814);
or U23937 (N_23937,N_15110,N_15133);
nand U23938 (N_23938,N_17183,N_16668);
and U23939 (N_23939,N_15375,N_18195);
nor U23940 (N_23940,N_19698,N_18681);
xor U23941 (N_23941,N_16610,N_15977);
nand U23942 (N_23942,N_18730,N_19685);
nor U23943 (N_23943,N_18863,N_18643);
xnor U23944 (N_23944,N_16929,N_19436);
or U23945 (N_23945,N_15875,N_16687);
nor U23946 (N_23946,N_19277,N_16785);
nand U23947 (N_23947,N_15797,N_17109);
nor U23948 (N_23948,N_16986,N_17648);
nand U23949 (N_23949,N_18295,N_18665);
xnor U23950 (N_23950,N_19359,N_16160);
nor U23951 (N_23951,N_18738,N_19720);
nor U23952 (N_23952,N_15987,N_18968);
xor U23953 (N_23953,N_19661,N_18005);
and U23954 (N_23954,N_16207,N_18022);
or U23955 (N_23955,N_15672,N_18415);
xnor U23956 (N_23956,N_15320,N_18101);
or U23957 (N_23957,N_16895,N_15767);
nand U23958 (N_23958,N_18078,N_18369);
nor U23959 (N_23959,N_15406,N_19872);
nor U23960 (N_23960,N_17925,N_18173);
xor U23961 (N_23961,N_15673,N_19156);
xor U23962 (N_23962,N_17957,N_19799);
nand U23963 (N_23963,N_19533,N_18816);
nand U23964 (N_23964,N_18140,N_15824);
and U23965 (N_23965,N_16602,N_18162);
and U23966 (N_23966,N_15018,N_18285);
nor U23967 (N_23967,N_15954,N_17863);
or U23968 (N_23968,N_15414,N_19333);
xnor U23969 (N_23969,N_15151,N_16154);
nand U23970 (N_23970,N_19477,N_17512);
or U23971 (N_23971,N_16695,N_17000);
or U23972 (N_23972,N_19540,N_15705);
nor U23973 (N_23973,N_19542,N_15722);
xnor U23974 (N_23974,N_16568,N_17174);
xor U23975 (N_23975,N_17764,N_16612);
and U23976 (N_23976,N_17536,N_16082);
or U23977 (N_23977,N_19098,N_15886);
or U23978 (N_23978,N_16103,N_16505);
and U23979 (N_23979,N_17900,N_18462);
nand U23980 (N_23980,N_15331,N_15190);
or U23981 (N_23981,N_18775,N_19604);
and U23982 (N_23982,N_15126,N_17585);
nor U23983 (N_23983,N_16224,N_18818);
nand U23984 (N_23984,N_15443,N_15338);
nor U23985 (N_23985,N_16971,N_18537);
nand U23986 (N_23986,N_16131,N_16875);
xor U23987 (N_23987,N_19815,N_17631);
or U23988 (N_23988,N_18822,N_17990);
nor U23989 (N_23989,N_17190,N_16216);
xnor U23990 (N_23990,N_17218,N_15604);
or U23991 (N_23991,N_19566,N_17051);
nand U23992 (N_23992,N_19917,N_15227);
nand U23993 (N_23993,N_15503,N_19213);
xnor U23994 (N_23994,N_18556,N_15018);
or U23995 (N_23995,N_19485,N_16370);
nor U23996 (N_23996,N_18100,N_15763);
and U23997 (N_23997,N_16179,N_19486);
nand U23998 (N_23998,N_18831,N_17763);
xor U23999 (N_23999,N_19487,N_19406);
and U24000 (N_24000,N_16173,N_15609);
and U24001 (N_24001,N_16701,N_17546);
nor U24002 (N_24002,N_19770,N_17980);
and U24003 (N_24003,N_15128,N_17039);
and U24004 (N_24004,N_17468,N_15370);
nor U24005 (N_24005,N_19607,N_19662);
nor U24006 (N_24006,N_17143,N_19055);
nor U24007 (N_24007,N_15224,N_16951);
nor U24008 (N_24008,N_16298,N_17461);
or U24009 (N_24009,N_18791,N_18230);
or U24010 (N_24010,N_19316,N_18339);
xnor U24011 (N_24011,N_17288,N_18820);
nand U24012 (N_24012,N_16412,N_15860);
nor U24013 (N_24013,N_18185,N_16917);
nand U24014 (N_24014,N_15472,N_17137);
nor U24015 (N_24015,N_15962,N_19531);
nand U24016 (N_24016,N_16407,N_18007);
and U24017 (N_24017,N_18341,N_19554);
nor U24018 (N_24018,N_15595,N_15980);
and U24019 (N_24019,N_17413,N_17941);
nor U24020 (N_24020,N_19235,N_19955);
nor U24021 (N_24021,N_19766,N_15311);
nand U24022 (N_24022,N_18960,N_19866);
nand U24023 (N_24023,N_15611,N_18977);
nand U24024 (N_24024,N_15298,N_19231);
or U24025 (N_24025,N_17912,N_19508);
xnor U24026 (N_24026,N_16527,N_17085);
xnor U24027 (N_24027,N_16109,N_16900);
xnor U24028 (N_24028,N_15512,N_19697);
xor U24029 (N_24029,N_18164,N_16849);
and U24030 (N_24030,N_18531,N_17981);
or U24031 (N_24031,N_15385,N_18303);
nor U24032 (N_24032,N_16061,N_17830);
nand U24033 (N_24033,N_17095,N_17647);
nand U24034 (N_24034,N_17898,N_19131);
nand U24035 (N_24035,N_18197,N_15639);
nand U24036 (N_24036,N_17742,N_18584);
and U24037 (N_24037,N_15637,N_15105);
or U24038 (N_24038,N_17138,N_16246);
nand U24039 (N_24039,N_15924,N_16476);
nor U24040 (N_24040,N_19294,N_18048);
nor U24041 (N_24041,N_19726,N_19941);
nor U24042 (N_24042,N_19574,N_15118);
xor U24043 (N_24043,N_18673,N_17446);
nand U24044 (N_24044,N_18572,N_19278);
and U24045 (N_24045,N_16483,N_16526);
xnor U24046 (N_24046,N_17281,N_18605);
and U24047 (N_24047,N_19244,N_17459);
or U24048 (N_24048,N_18871,N_15262);
or U24049 (N_24049,N_19163,N_16563);
and U24050 (N_24050,N_15976,N_18780);
or U24051 (N_24051,N_19469,N_17268);
nor U24052 (N_24052,N_19250,N_18939);
xor U24053 (N_24053,N_18227,N_15218);
nand U24054 (N_24054,N_17765,N_15776);
and U24055 (N_24055,N_17348,N_15000);
nor U24056 (N_24056,N_15810,N_15884);
and U24057 (N_24057,N_15989,N_15821);
nand U24058 (N_24058,N_16983,N_17249);
nor U24059 (N_24059,N_15466,N_18515);
nand U24060 (N_24060,N_16089,N_17848);
nand U24061 (N_24061,N_19114,N_16866);
xor U24062 (N_24062,N_16184,N_17997);
xor U24063 (N_24063,N_15517,N_15163);
and U24064 (N_24064,N_18823,N_18376);
and U24065 (N_24065,N_15202,N_17639);
and U24066 (N_24066,N_17743,N_18989);
nand U24067 (N_24067,N_17453,N_16473);
nand U24068 (N_24068,N_16933,N_18800);
nand U24069 (N_24069,N_16834,N_19451);
and U24070 (N_24070,N_19186,N_18031);
xnor U24071 (N_24071,N_18972,N_19312);
or U24072 (N_24072,N_17905,N_18935);
and U24073 (N_24073,N_16686,N_19830);
nand U24074 (N_24074,N_16360,N_15688);
nor U24075 (N_24075,N_16869,N_16505);
or U24076 (N_24076,N_15948,N_16256);
and U24077 (N_24077,N_16704,N_19645);
nand U24078 (N_24078,N_17894,N_16555);
and U24079 (N_24079,N_18178,N_15768);
and U24080 (N_24080,N_17316,N_15443);
or U24081 (N_24081,N_16535,N_15565);
and U24082 (N_24082,N_16230,N_19792);
nor U24083 (N_24083,N_17878,N_19338);
nor U24084 (N_24084,N_16241,N_19487);
and U24085 (N_24085,N_18548,N_18270);
nor U24086 (N_24086,N_15679,N_19227);
nor U24087 (N_24087,N_15295,N_17098);
nand U24088 (N_24088,N_16792,N_18195);
xnor U24089 (N_24089,N_17211,N_18297);
nand U24090 (N_24090,N_17468,N_19590);
nor U24091 (N_24091,N_16972,N_19443);
nand U24092 (N_24092,N_18345,N_18620);
or U24093 (N_24093,N_18747,N_15824);
nand U24094 (N_24094,N_18793,N_15150);
or U24095 (N_24095,N_18425,N_17681);
nor U24096 (N_24096,N_18014,N_17695);
nor U24097 (N_24097,N_15843,N_15887);
and U24098 (N_24098,N_16218,N_17088);
nand U24099 (N_24099,N_15587,N_19116);
and U24100 (N_24100,N_16442,N_17192);
or U24101 (N_24101,N_15192,N_16316);
xor U24102 (N_24102,N_19058,N_19946);
or U24103 (N_24103,N_16100,N_19733);
or U24104 (N_24104,N_19935,N_19901);
and U24105 (N_24105,N_19616,N_16209);
nand U24106 (N_24106,N_16296,N_15608);
nor U24107 (N_24107,N_19001,N_19166);
nand U24108 (N_24108,N_16823,N_15801);
and U24109 (N_24109,N_16698,N_19953);
and U24110 (N_24110,N_18854,N_18640);
or U24111 (N_24111,N_17265,N_19002);
nor U24112 (N_24112,N_16619,N_16605);
or U24113 (N_24113,N_15924,N_18695);
nor U24114 (N_24114,N_15100,N_18734);
nand U24115 (N_24115,N_19122,N_15472);
nand U24116 (N_24116,N_16576,N_17669);
nand U24117 (N_24117,N_19324,N_16318);
or U24118 (N_24118,N_16446,N_18826);
nand U24119 (N_24119,N_17457,N_18220);
xnor U24120 (N_24120,N_18109,N_19340);
nand U24121 (N_24121,N_18794,N_17763);
or U24122 (N_24122,N_19735,N_18406);
nor U24123 (N_24123,N_19294,N_17949);
xnor U24124 (N_24124,N_18834,N_18583);
nand U24125 (N_24125,N_15816,N_19711);
and U24126 (N_24126,N_15779,N_16487);
xor U24127 (N_24127,N_17019,N_15530);
nor U24128 (N_24128,N_17295,N_17062);
xor U24129 (N_24129,N_19267,N_18587);
or U24130 (N_24130,N_16698,N_17728);
nor U24131 (N_24131,N_15757,N_18714);
nor U24132 (N_24132,N_18469,N_16363);
xor U24133 (N_24133,N_15600,N_16494);
and U24134 (N_24134,N_17280,N_19686);
nand U24135 (N_24135,N_18991,N_17900);
nand U24136 (N_24136,N_15687,N_18826);
or U24137 (N_24137,N_17562,N_18540);
nor U24138 (N_24138,N_18971,N_19752);
and U24139 (N_24139,N_16636,N_17856);
xnor U24140 (N_24140,N_18931,N_19818);
and U24141 (N_24141,N_18491,N_17958);
or U24142 (N_24142,N_17790,N_17444);
and U24143 (N_24143,N_17031,N_19878);
nor U24144 (N_24144,N_19619,N_18126);
nor U24145 (N_24145,N_17598,N_19033);
or U24146 (N_24146,N_15227,N_17498);
nor U24147 (N_24147,N_17215,N_18229);
and U24148 (N_24148,N_19186,N_15906);
nor U24149 (N_24149,N_15498,N_19140);
or U24150 (N_24150,N_15100,N_15363);
or U24151 (N_24151,N_18872,N_18540);
nand U24152 (N_24152,N_19748,N_16741);
and U24153 (N_24153,N_15462,N_15373);
or U24154 (N_24154,N_18710,N_16136);
and U24155 (N_24155,N_18736,N_17686);
or U24156 (N_24156,N_17292,N_19285);
xnor U24157 (N_24157,N_18079,N_15351);
or U24158 (N_24158,N_17550,N_19097);
and U24159 (N_24159,N_16020,N_17906);
nor U24160 (N_24160,N_16513,N_19538);
and U24161 (N_24161,N_16169,N_19050);
or U24162 (N_24162,N_15007,N_15669);
or U24163 (N_24163,N_17140,N_19001);
xor U24164 (N_24164,N_17418,N_19918);
nand U24165 (N_24165,N_15466,N_15015);
xnor U24166 (N_24166,N_19439,N_16623);
and U24167 (N_24167,N_18314,N_19264);
or U24168 (N_24168,N_15009,N_15094);
xor U24169 (N_24169,N_15515,N_18397);
xnor U24170 (N_24170,N_17618,N_16479);
nor U24171 (N_24171,N_18982,N_19625);
nand U24172 (N_24172,N_15091,N_16972);
xnor U24173 (N_24173,N_17748,N_16344);
xor U24174 (N_24174,N_17197,N_19753);
and U24175 (N_24175,N_19036,N_16490);
nand U24176 (N_24176,N_16991,N_18691);
nor U24177 (N_24177,N_16778,N_15639);
nand U24178 (N_24178,N_15468,N_16047);
nor U24179 (N_24179,N_18861,N_18116);
nor U24180 (N_24180,N_15228,N_18450);
nand U24181 (N_24181,N_17697,N_18759);
nand U24182 (N_24182,N_16286,N_19740);
nand U24183 (N_24183,N_17993,N_18988);
nor U24184 (N_24184,N_18065,N_17235);
nand U24185 (N_24185,N_17609,N_16302);
and U24186 (N_24186,N_15244,N_18094);
and U24187 (N_24187,N_18376,N_16179);
xnor U24188 (N_24188,N_18054,N_17345);
or U24189 (N_24189,N_18971,N_17943);
or U24190 (N_24190,N_16689,N_16148);
nand U24191 (N_24191,N_17093,N_18105);
or U24192 (N_24192,N_15299,N_18053);
or U24193 (N_24193,N_17833,N_18902);
xnor U24194 (N_24194,N_18328,N_19602);
or U24195 (N_24195,N_16453,N_18224);
and U24196 (N_24196,N_16720,N_16870);
xor U24197 (N_24197,N_17697,N_16995);
nand U24198 (N_24198,N_18444,N_16438);
and U24199 (N_24199,N_17422,N_19982);
xor U24200 (N_24200,N_16215,N_19739);
xor U24201 (N_24201,N_15000,N_15682);
nor U24202 (N_24202,N_17016,N_18280);
xor U24203 (N_24203,N_15531,N_16657);
or U24204 (N_24204,N_15547,N_15999);
or U24205 (N_24205,N_16505,N_18545);
and U24206 (N_24206,N_17372,N_15887);
and U24207 (N_24207,N_15486,N_18084);
or U24208 (N_24208,N_18875,N_18477);
nand U24209 (N_24209,N_17283,N_19951);
xor U24210 (N_24210,N_16194,N_15557);
nand U24211 (N_24211,N_16168,N_16353);
nand U24212 (N_24212,N_17816,N_15179);
or U24213 (N_24213,N_15536,N_16892);
nand U24214 (N_24214,N_19993,N_19906);
xnor U24215 (N_24215,N_19845,N_19443);
or U24216 (N_24216,N_16007,N_16097);
or U24217 (N_24217,N_18343,N_15731);
xnor U24218 (N_24218,N_16139,N_15405);
nor U24219 (N_24219,N_18775,N_16038);
and U24220 (N_24220,N_19592,N_19072);
and U24221 (N_24221,N_19627,N_15020);
and U24222 (N_24222,N_15605,N_17000);
or U24223 (N_24223,N_17044,N_17400);
xnor U24224 (N_24224,N_19074,N_16613);
or U24225 (N_24225,N_15696,N_18879);
or U24226 (N_24226,N_19903,N_17962);
and U24227 (N_24227,N_18167,N_18163);
or U24228 (N_24228,N_16989,N_15467);
xnor U24229 (N_24229,N_18690,N_19757);
and U24230 (N_24230,N_19734,N_15405);
nor U24231 (N_24231,N_18164,N_18670);
and U24232 (N_24232,N_16811,N_17517);
nor U24233 (N_24233,N_17629,N_15550);
or U24234 (N_24234,N_16642,N_18223);
nand U24235 (N_24235,N_18880,N_18591);
nor U24236 (N_24236,N_17208,N_17394);
xor U24237 (N_24237,N_18409,N_18149);
or U24238 (N_24238,N_17271,N_16621);
and U24239 (N_24239,N_17161,N_15722);
or U24240 (N_24240,N_16121,N_19842);
xnor U24241 (N_24241,N_15275,N_15486);
and U24242 (N_24242,N_19822,N_17469);
xor U24243 (N_24243,N_16766,N_17400);
or U24244 (N_24244,N_16162,N_17115);
xor U24245 (N_24245,N_17663,N_18593);
nand U24246 (N_24246,N_17114,N_19900);
or U24247 (N_24247,N_16535,N_18355);
and U24248 (N_24248,N_18181,N_18309);
nand U24249 (N_24249,N_18521,N_18101);
nand U24250 (N_24250,N_16876,N_17887);
and U24251 (N_24251,N_17638,N_19854);
nand U24252 (N_24252,N_17024,N_16665);
or U24253 (N_24253,N_19586,N_16800);
and U24254 (N_24254,N_19129,N_17720);
or U24255 (N_24255,N_15635,N_19919);
nor U24256 (N_24256,N_19112,N_17760);
or U24257 (N_24257,N_17481,N_17581);
and U24258 (N_24258,N_15579,N_17519);
and U24259 (N_24259,N_18319,N_18276);
and U24260 (N_24260,N_18006,N_19421);
xor U24261 (N_24261,N_15782,N_16727);
or U24262 (N_24262,N_16806,N_16933);
nor U24263 (N_24263,N_18375,N_19917);
nand U24264 (N_24264,N_15717,N_18093);
or U24265 (N_24265,N_16670,N_18485);
or U24266 (N_24266,N_19651,N_19591);
xor U24267 (N_24267,N_15175,N_16705);
nand U24268 (N_24268,N_19445,N_15273);
nand U24269 (N_24269,N_16911,N_19453);
or U24270 (N_24270,N_15494,N_16477);
nand U24271 (N_24271,N_15271,N_16600);
or U24272 (N_24272,N_18748,N_18283);
nand U24273 (N_24273,N_18706,N_16070);
or U24274 (N_24274,N_19686,N_18776);
or U24275 (N_24275,N_19106,N_15842);
and U24276 (N_24276,N_15043,N_19129);
and U24277 (N_24277,N_19164,N_18653);
and U24278 (N_24278,N_15123,N_16837);
xnor U24279 (N_24279,N_18114,N_18496);
and U24280 (N_24280,N_16904,N_19091);
and U24281 (N_24281,N_15281,N_16427);
nand U24282 (N_24282,N_15853,N_18396);
or U24283 (N_24283,N_17422,N_15103);
xor U24284 (N_24284,N_17081,N_16800);
nand U24285 (N_24285,N_19270,N_15081);
xor U24286 (N_24286,N_19444,N_18206);
xor U24287 (N_24287,N_18005,N_16042);
nor U24288 (N_24288,N_16761,N_19336);
nor U24289 (N_24289,N_17197,N_19392);
nand U24290 (N_24290,N_16185,N_17440);
nor U24291 (N_24291,N_17572,N_16685);
or U24292 (N_24292,N_18467,N_19090);
xnor U24293 (N_24293,N_17531,N_16796);
or U24294 (N_24294,N_18247,N_16564);
or U24295 (N_24295,N_19095,N_15942);
and U24296 (N_24296,N_18961,N_16328);
nand U24297 (N_24297,N_16157,N_17012);
and U24298 (N_24298,N_16559,N_16491);
nand U24299 (N_24299,N_17092,N_16863);
or U24300 (N_24300,N_16968,N_15344);
nor U24301 (N_24301,N_16536,N_19170);
and U24302 (N_24302,N_16010,N_15400);
and U24303 (N_24303,N_19587,N_18342);
nor U24304 (N_24304,N_15064,N_17850);
nor U24305 (N_24305,N_17252,N_18733);
nor U24306 (N_24306,N_16139,N_17834);
xor U24307 (N_24307,N_18221,N_18939);
and U24308 (N_24308,N_17246,N_16740);
xor U24309 (N_24309,N_16565,N_19697);
or U24310 (N_24310,N_18200,N_19900);
and U24311 (N_24311,N_19234,N_17241);
nand U24312 (N_24312,N_15709,N_15860);
xor U24313 (N_24313,N_17327,N_17351);
xor U24314 (N_24314,N_19690,N_19746);
nor U24315 (N_24315,N_16456,N_19143);
nor U24316 (N_24316,N_17207,N_17424);
xor U24317 (N_24317,N_15443,N_16178);
and U24318 (N_24318,N_16970,N_18764);
nand U24319 (N_24319,N_15186,N_19645);
nand U24320 (N_24320,N_15578,N_17183);
and U24321 (N_24321,N_17723,N_19879);
nand U24322 (N_24322,N_19611,N_17946);
and U24323 (N_24323,N_19825,N_17287);
xnor U24324 (N_24324,N_17712,N_16620);
nand U24325 (N_24325,N_16998,N_16068);
xnor U24326 (N_24326,N_18472,N_19123);
nand U24327 (N_24327,N_15896,N_18841);
nor U24328 (N_24328,N_17035,N_18507);
xnor U24329 (N_24329,N_15221,N_15517);
xnor U24330 (N_24330,N_17596,N_16752);
or U24331 (N_24331,N_15958,N_17709);
nor U24332 (N_24332,N_16718,N_17149);
or U24333 (N_24333,N_15137,N_16315);
and U24334 (N_24334,N_15992,N_19308);
xor U24335 (N_24335,N_18041,N_17059);
nor U24336 (N_24336,N_17359,N_17311);
nor U24337 (N_24337,N_18365,N_15161);
xor U24338 (N_24338,N_15179,N_16385);
or U24339 (N_24339,N_15273,N_16480);
nand U24340 (N_24340,N_17673,N_19623);
nand U24341 (N_24341,N_15765,N_17675);
or U24342 (N_24342,N_16933,N_18548);
nor U24343 (N_24343,N_16486,N_18139);
and U24344 (N_24344,N_18316,N_18456);
and U24345 (N_24345,N_18701,N_16439);
nand U24346 (N_24346,N_17651,N_16261);
and U24347 (N_24347,N_18751,N_17855);
xnor U24348 (N_24348,N_16724,N_15612);
nand U24349 (N_24349,N_16564,N_16078);
and U24350 (N_24350,N_16853,N_18032);
or U24351 (N_24351,N_18679,N_16588);
nor U24352 (N_24352,N_18326,N_19947);
and U24353 (N_24353,N_16150,N_18906);
nand U24354 (N_24354,N_17530,N_19038);
nand U24355 (N_24355,N_16856,N_15745);
or U24356 (N_24356,N_18654,N_16388);
nand U24357 (N_24357,N_19002,N_19610);
or U24358 (N_24358,N_17219,N_15331);
nand U24359 (N_24359,N_16916,N_19211);
nand U24360 (N_24360,N_19875,N_18935);
and U24361 (N_24361,N_16105,N_19665);
xor U24362 (N_24362,N_18530,N_16463);
xor U24363 (N_24363,N_19896,N_17239);
nand U24364 (N_24364,N_19341,N_15940);
nor U24365 (N_24365,N_17574,N_19731);
and U24366 (N_24366,N_16696,N_19346);
and U24367 (N_24367,N_17355,N_15023);
xnor U24368 (N_24368,N_15419,N_19868);
or U24369 (N_24369,N_16884,N_19856);
nor U24370 (N_24370,N_16569,N_16799);
nor U24371 (N_24371,N_19267,N_18755);
and U24372 (N_24372,N_16480,N_17015);
nand U24373 (N_24373,N_18029,N_19451);
nor U24374 (N_24374,N_17437,N_18339);
and U24375 (N_24375,N_15784,N_18562);
and U24376 (N_24376,N_18491,N_18445);
and U24377 (N_24377,N_18832,N_17680);
nor U24378 (N_24378,N_18286,N_18090);
xnor U24379 (N_24379,N_15572,N_17455);
or U24380 (N_24380,N_15589,N_17817);
or U24381 (N_24381,N_15282,N_15918);
and U24382 (N_24382,N_17968,N_19595);
xor U24383 (N_24383,N_19072,N_15950);
and U24384 (N_24384,N_18726,N_16797);
or U24385 (N_24385,N_18029,N_19213);
or U24386 (N_24386,N_17856,N_17171);
xnor U24387 (N_24387,N_19223,N_15324);
and U24388 (N_24388,N_18817,N_19118);
nand U24389 (N_24389,N_16462,N_16962);
nor U24390 (N_24390,N_19180,N_17024);
and U24391 (N_24391,N_17363,N_16798);
or U24392 (N_24392,N_15691,N_17690);
nand U24393 (N_24393,N_16471,N_15676);
nand U24394 (N_24394,N_17535,N_19964);
xor U24395 (N_24395,N_17348,N_18287);
nor U24396 (N_24396,N_19269,N_17477);
nor U24397 (N_24397,N_15830,N_17967);
nand U24398 (N_24398,N_15903,N_17640);
nand U24399 (N_24399,N_19299,N_18866);
or U24400 (N_24400,N_15082,N_15590);
nand U24401 (N_24401,N_17144,N_16133);
nor U24402 (N_24402,N_17128,N_15623);
nand U24403 (N_24403,N_15136,N_18611);
nor U24404 (N_24404,N_19659,N_15902);
nand U24405 (N_24405,N_19813,N_15975);
xor U24406 (N_24406,N_18005,N_19937);
and U24407 (N_24407,N_16562,N_15142);
and U24408 (N_24408,N_18128,N_15075);
or U24409 (N_24409,N_19114,N_17059);
nor U24410 (N_24410,N_17987,N_19518);
nor U24411 (N_24411,N_17116,N_15991);
xor U24412 (N_24412,N_17781,N_15320);
xnor U24413 (N_24413,N_17821,N_16115);
xnor U24414 (N_24414,N_15729,N_19622);
or U24415 (N_24415,N_15675,N_16113);
or U24416 (N_24416,N_17854,N_19973);
xnor U24417 (N_24417,N_19418,N_17972);
nor U24418 (N_24418,N_17498,N_18892);
nand U24419 (N_24419,N_18529,N_18105);
nor U24420 (N_24420,N_18390,N_15594);
xnor U24421 (N_24421,N_17408,N_17994);
nand U24422 (N_24422,N_19770,N_15495);
nand U24423 (N_24423,N_16098,N_19825);
xnor U24424 (N_24424,N_17180,N_17637);
nor U24425 (N_24425,N_19176,N_15574);
and U24426 (N_24426,N_19094,N_15676);
nand U24427 (N_24427,N_16979,N_15524);
and U24428 (N_24428,N_15035,N_16439);
nor U24429 (N_24429,N_16922,N_18878);
nand U24430 (N_24430,N_19759,N_16621);
and U24431 (N_24431,N_15857,N_18870);
or U24432 (N_24432,N_18264,N_16839);
or U24433 (N_24433,N_17524,N_16689);
nor U24434 (N_24434,N_19167,N_17706);
and U24435 (N_24435,N_17249,N_16951);
and U24436 (N_24436,N_18932,N_17787);
or U24437 (N_24437,N_18749,N_16963);
and U24438 (N_24438,N_19831,N_15080);
and U24439 (N_24439,N_17464,N_15733);
xor U24440 (N_24440,N_15265,N_19255);
or U24441 (N_24441,N_16880,N_15716);
xor U24442 (N_24442,N_17953,N_17848);
nand U24443 (N_24443,N_18302,N_19434);
xor U24444 (N_24444,N_16427,N_16563);
nor U24445 (N_24445,N_16247,N_17907);
and U24446 (N_24446,N_18494,N_18358);
or U24447 (N_24447,N_16096,N_18427);
xor U24448 (N_24448,N_18223,N_15553);
nor U24449 (N_24449,N_16631,N_18963);
or U24450 (N_24450,N_16904,N_15422);
and U24451 (N_24451,N_17830,N_19362);
nand U24452 (N_24452,N_15319,N_16193);
nor U24453 (N_24453,N_15717,N_17887);
nor U24454 (N_24454,N_18082,N_19073);
xnor U24455 (N_24455,N_16726,N_19594);
nand U24456 (N_24456,N_15690,N_18470);
xnor U24457 (N_24457,N_18647,N_17683);
nand U24458 (N_24458,N_15272,N_17453);
or U24459 (N_24459,N_18141,N_16287);
or U24460 (N_24460,N_15947,N_15877);
nor U24461 (N_24461,N_18056,N_16331);
xor U24462 (N_24462,N_18048,N_18219);
or U24463 (N_24463,N_17642,N_15356);
xnor U24464 (N_24464,N_15244,N_19215);
nand U24465 (N_24465,N_19688,N_16331);
nor U24466 (N_24466,N_17338,N_18784);
nor U24467 (N_24467,N_15050,N_18558);
or U24468 (N_24468,N_16635,N_18353);
nor U24469 (N_24469,N_16248,N_16511);
nand U24470 (N_24470,N_19060,N_17570);
nor U24471 (N_24471,N_17999,N_18523);
nand U24472 (N_24472,N_19938,N_19836);
nand U24473 (N_24473,N_18237,N_17003);
nor U24474 (N_24474,N_19227,N_16053);
or U24475 (N_24475,N_19543,N_18170);
and U24476 (N_24476,N_15149,N_18618);
nand U24477 (N_24477,N_15383,N_17510);
or U24478 (N_24478,N_19269,N_15873);
nand U24479 (N_24479,N_18009,N_19550);
or U24480 (N_24480,N_19976,N_16205);
and U24481 (N_24481,N_18395,N_19011);
nor U24482 (N_24482,N_19275,N_15828);
nor U24483 (N_24483,N_16791,N_16819);
nor U24484 (N_24484,N_15459,N_15527);
and U24485 (N_24485,N_15457,N_18753);
nor U24486 (N_24486,N_16583,N_17644);
or U24487 (N_24487,N_18292,N_17869);
nor U24488 (N_24488,N_18084,N_19144);
xnor U24489 (N_24489,N_18825,N_17413);
or U24490 (N_24490,N_18493,N_18444);
and U24491 (N_24491,N_15505,N_17488);
xor U24492 (N_24492,N_17347,N_16521);
and U24493 (N_24493,N_15960,N_15500);
nor U24494 (N_24494,N_19275,N_15885);
xor U24495 (N_24495,N_15753,N_15673);
nor U24496 (N_24496,N_18742,N_17794);
or U24497 (N_24497,N_19244,N_17366);
nand U24498 (N_24498,N_18561,N_16293);
and U24499 (N_24499,N_17360,N_16029);
nor U24500 (N_24500,N_16296,N_15304);
nand U24501 (N_24501,N_17592,N_15935);
and U24502 (N_24502,N_16697,N_17381);
and U24503 (N_24503,N_18016,N_17844);
nand U24504 (N_24504,N_15996,N_15719);
nor U24505 (N_24505,N_15574,N_15310);
nand U24506 (N_24506,N_16206,N_19480);
or U24507 (N_24507,N_16446,N_15683);
or U24508 (N_24508,N_16409,N_19242);
and U24509 (N_24509,N_16049,N_17645);
and U24510 (N_24510,N_15704,N_17972);
and U24511 (N_24511,N_18324,N_16061);
or U24512 (N_24512,N_17700,N_19600);
or U24513 (N_24513,N_16665,N_18835);
nor U24514 (N_24514,N_15298,N_16358);
xnor U24515 (N_24515,N_18003,N_16985);
xor U24516 (N_24516,N_18037,N_15478);
or U24517 (N_24517,N_15439,N_15494);
nor U24518 (N_24518,N_15392,N_17334);
or U24519 (N_24519,N_16561,N_15373);
nand U24520 (N_24520,N_18477,N_17436);
nand U24521 (N_24521,N_19297,N_19162);
nor U24522 (N_24522,N_15328,N_17158);
and U24523 (N_24523,N_17699,N_15313);
or U24524 (N_24524,N_17802,N_18419);
and U24525 (N_24525,N_19666,N_15478);
nand U24526 (N_24526,N_16881,N_17603);
and U24527 (N_24527,N_18299,N_17256);
nor U24528 (N_24528,N_19200,N_16725);
and U24529 (N_24529,N_19731,N_16393);
xor U24530 (N_24530,N_18715,N_15166);
and U24531 (N_24531,N_15392,N_17219);
nand U24532 (N_24532,N_19063,N_15519);
nor U24533 (N_24533,N_19480,N_18429);
and U24534 (N_24534,N_18199,N_15882);
xnor U24535 (N_24535,N_17245,N_19873);
and U24536 (N_24536,N_15421,N_18975);
xor U24537 (N_24537,N_15310,N_19947);
nand U24538 (N_24538,N_17751,N_15241);
and U24539 (N_24539,N_16137,N_16204);
nand U24540 (N_24540,N_18767,N_18075);
nand U24541 (N_24541,N_17095,N_16007);
nor U24542 (N_24542,N_16044,N_16795);
xor U24543 (N_24543,N_18063,N_18591);
and U24544 (N_24544,N_17256,N_18393);
xor U24545 (N_24545,N_15253,N_18690);
and U24546 (N_24546,N_17159,N_15609);
and U24547 (N_24547,N_18171,N_15516);
or U24548 (N_24548,N_18515,N_16531);
nand U24549 (N_24549,N_17623,N_15078);
xnor U24550 (N_24550,N_15120,N_19801);
nand U24551 (N_24551,N_16617,N_15366);
nand U24552 (N_24552,N_19570,N_19964);
and U24553 (N_24553,N_18401,N_18177);
and U24554 (N_24554,N_18121,N_18283);
and U24555 (N_24555,N_15996,N_19389);
nor U24556 (N_24556,N_19414,N_18792);
nor U24557 (N_24557,N_16831,N_16926);
nor U24558 (N_24558,N_19340,N_17592);
and U24559 (N_24559,N_16879,N_15635);
or U24560 (N_24560,N_16833,N_16463);
nand U24561 (N_24561,N_19572,N_18878);
and U24562 (N_24562,N_15831,N_18297);
nand U24563 (N_24563,N_19446,N_16998);
and U24564 (N_24564,N_16685,N_15165);
xnor U24565 (N_24565,N_18000,N_19795);
nand U24566 (N_24566,N_19997,N_19495);
nor U24567 (N_24567,N_16892,N_17672);
nor U24568 (N_24568,N_18609,N_19414);
xnor U24569 (N_24569,N_17750,N_16962);
xnor U24570 (N_24570,N_18576,N_16067);
or U24571 (N_24571,N_16283,N_19003);
nand U24572 (N_24572,N_17085,N_17845);
and U24573 (N_24573,N_15129,N_18740);
nand U24574 (N_24574,N_19441,N_17885);
nor U24575 (N_24575,N_15306,N_19561);
or U24576 (N_24576,N_16341,N_19133);
and U24577 (N_24577,N_16942,N_16285);
and U24578 (N_24578,N_17467,N_19203);
or U24579 (N_24579,N_19826,N_19544);
or U24580 (N_24580,N_17768,N_19759);
nand U24581 (N_24581,N_17864,N_16460);
and U24582 (N_24582,N_18918,N_17749);
or U24583 (N_24583,N_17119,N_15139);
or U24584 (N_24584,N_19392,N_16768);
and U24585 (N_24585,N_17606,N_18212);
or U24586 (N_24586,N_19813,N_16845);
nand U24587 (N_24587,N_18383,N_19272);
and U24588 (N_24588,N_15176,N_15089);
and U24589 (N_24589,N_17612,N_15836);
and U24590 (N_24590,N_18303,N_19282);
and U24591 (N_24591,N_15722,N_16278);
nand U24592 (N_24592,N_17608,N_16410);
or U24593 (N_24593,N_16732,N_15447);
nand U24594 (N_24594,N_17616,N_17824);
nand U24595 (N_24595,N_19383,N_16041);
and U24596 (N_24596,N_18468,N_17893);
nand U24597 (N_24597,N_16784,N_19285);
or U24598 (N_24598,N_18938,N_18607);
and U24599 (N_24599,N_16640,N_16363);
or U24600 (N_24600,N_16890,N_16296);
or U24601 (N_24601,N_19084,N_16559);
nor U24602 (N_24602,N_18247,N_17960);
and U24603 (N_24603,N_17776,N_19490);
and U24604 (N_24604,N_16734,N_17926);
nor U24605 (N_24605,N_18168,N_17940);
or U24606 (N_24606,N_17399,N_17973);
and U24607 (N_24607,N_16935,N_19462);
and U24608 (N_24608,N_19054,N_16537);
nand U24609 (N_24609,N_17396,N_15815);
or U24610 (N_24610,N_19938,N_15576);
nor U24611 (N_24611,N_18249,N_17222);
nand U24612 (N_24612,N_17659,N_18243);
nor U24613 (N_24613,N_15993,N_17776);
and U24614 (N_24614,N_16900,N_19092);
nor U24615 (N_24615,N_15662,N_18107);
and U24616 (N_24616,N_19663,N_15418);
nor U24617 (N_24617,N_16805,N_17093);
nand U24618 (N_24618,N_18015,N_17415);
and U24619 (N_24619,N_15372,N_18718);
nand U24620 (N_24620,N_16568,N_17733);
nor U24621 (N_24621,N_15349,N_15931);
nand U24622 (N_24622,N_16755,N_19173);
nor U24623 (N_24623,N_17101,N_17803);
nand U24624 (N_24624,N_17282,N_15302);
or U24625 (N_24625,N_16946,N_19079);
or U24626 (N_24626,N_18404,N_15725);
nand U24627 (N_24627,N_17092,N_19715);
and U24628 (N_24628,N_19446,N_18970);
nor U24629 (N_24629,N_16574,N_15652);
nand U24630 (N_24630,N_15269,N_18044);
nor U24631 (N_24631,N_17600,N_16676);
nor U24632 (N_24632,N_17892,N_19975);
or U24633 (N_24633,N_19815,N_17291);
nor U24634 (N_24634,N_16395,N_19606);
nand U24635 (N_24635,N_15820,N_16591);
nor U24636 (N_24636,N_19801,N_19763);
nand U24637 (N_24637,N_16997,N_19521);
nand U24638 (N_24638,N_18176,N_18600);
or U24639 (N_24639,N_15625,N_17980);
and U24640 (N_24640,N_18667,N_18042);
nand U24641 (N_24641,N_15089,N_18462);
or U24642 (N_24642,N_17947,N_18906);
nor U24643 (N_24643,N_16943,N_19964);
xor U24644 (N_24644,N_17813,N_15588);
or U24645 (N_24645,N_18137,N_18633);
nor U24646 (N_24646,N_18966,N_17600);
nor U24647 (N_24647,N_15168,N_19833);
nand U24648 (N_24648,N_17626,N_18233);
or U24649 (N_24649,N_19595,N_17126);
nand U24650 (N_24650,N_19305,N_19648);
nor U24651 (N_24651,N_18851,N_16047);
nand U24652 (N_24652,N_16774,N_16778);
xnor U24653 (N_24653,N_16388,N_17671);
and U24654 (N_24654,N_18762,N_17865);
nand U24655 (N_24655,N_16660,N_17827);
xnor U24656 (N_24656,N_18243,N_19101);
xnor U24657 (N_24657,N_19772,N_17531);
nor U24658 (N_24658,N_15252,N_19664);
nand U24659 (N_24659,N_17995,N_17215);
nor U24660 (N_24660,N_15929,N_18128);
and U24661 (N_24661,N_19652,N_15729);
nor U24662 (N_24662,N_19123,N_19940);
nor U24663 (N_24663,N_16591,N_16921);
nand U24664 (N_24664,N_15811,N_19049);
xor U24665 (N_24665,N_17205,N_17185);
or U24666 (N_24666,N_19029,N_17732);
nand U24667 (N_24667,N_15151,N_18795);
or U24668 (N_24668,N_19825,N_18648);
nand U24669 (N_24669,N_16153,N_16819);
nor U24670 (N_24670,N_15684,N_16773);
nor U24671 (N_24671,N_18547,N_16507);
or U24672 (N_24672,N_18951,N_15848);
nor U24673 (N_24673,N_16758,N_17236);
and U24674 (N_24674,N_19289,N_18073);
nand U24675 (N_24675,N_17416,N_18918);
nor U24676 (N_24676,N_15472,N_16838);
nor U24677 (N_24677,N_17118,N_18259);
xor U24678 (N_24678,N_16394,N_19221);
or U24679 (N_24679,N_16097,N_15165);
nor U24680 (N_24680,N_16496,N_15611);
or U24681 (N_24681,N_17997,N_17751);
or U24682 (N_24682,N_15282,N_18797);
nand U24683 (N_24683,N_15195,N_18223);
nor U24684 (N_24684,N_17158,N_15944);
nor U24685 (N_24685,N_19139,N_15260);
and U24686 (N_24686,N_17323,N_18261);
and U24687 (N_24687,N_17633,N_18259);
nor U24688 (N_24688,N_19744,N_17035);
nand U24689 (N_24689,N_17722,N_17152);
nor U24690 (N_24690,N_18237,N_19415);
nand U24691 (N_24691,N_18509,N_15730);
or U24692 (N_24692,N_18667,N_18822);
and U24693 (N_24693,N_15304,N_15497);
or U24694 (N_24694,N_16356,N_18488);
nor U24695 (N_24695,N_19269,N_19365);
xnor U24696 (N_24696,N_17905,N_18636);
or U24697 (N_24697,N_17372,N_15402);
nand U24698 (N_24698,N_15589,N_19595);
xnor U24699 (N_24699,N_15258,N_16426);
nor U24700 (N_24700,N_16254,N_19140);
or U24701 (N_24701,N_19264,N_18658);
or U24702 (N_24702,N_19742,N_18946);
xnor U24703 (N_24703,N_16205,N_19428);
nand U24704 (N_24704,N_18333,N_18418);
nand U24705 (N_24705,N_19730,N_19209);
xor U24706 (N_24706,N_15906,N_18220);
xor U24707 (N_24707,N_15060,N_16608);
nor U24708 (N_24708,N_18887,N_18983);
or U24709 (N_24709,N_17060,N_16112);
and U24710 (N_24710,N_15024,N_17991);
or U24711 (N_24711,N_16850,N_18594);
nand U24712 (N_24712,N_17854,N_19633);
nor U24713 (N_24713,N_17770,N_18074);
nor U24714 (N_24714,N_17671,N_16106);
or U24715 (N_24715,N_18079,N_16213);
and U24716 (N_24716,N_18964,N_19421);
or U24717 (N_24717,N_15799,N_16054);
and U24718 (N_24718,N_17596,N_19043);
nand U24719 (N_24719,N_15648,N_16476);
and U24720 (N_24720,N_18954,N_18792);
xor U24721 (N_24721,N_19834,N_18565);
nor U24722 (N_24722,N_19241,N_19759);
xnor U24723 (N_24723,N_18814,N_19249);
xor U24724 (N_24724,N_15131,N_18835);
nand U24725 (N_24725,N_15726,N_17477);
nand U24726 (N_24726,N_19895,N_16565);
and U24727 (N_24727,N_17956,N_19511);
and U24728 (N_24728,N_18553,N_15993);
xnor U24729 (N_24729,N_18121,N_15565);
xnor U24730 (N_24730,N_18550,N_17514);
xnor U24731 (N_24731,N_19633,N_16769);
and U24732 (N_24732,N_19732,N_19367);
xor U24733 (N_24733,N_16673,N_18551);
and U24734 (N_24734,N_19227,N_17948);
or U24735 (N_24735,N_15330,N_19660);
xnor U24736 (N_24736,N_18000,N_17334);
or U24737 (N_24737,N_19922,N_16107);
and U24738 (N_24738,N_16195,N_16264);
xnor U24739 (N_24739,N_16099,N_16152);
nor U24740 (N_24740,N_19162,N_15007);
or U24741 (N_24741,N_15522,N_16581);
or U24742 (N_24742,N_17454,N_15351);
nor U24743 (N_24743,N_19644,N_19362);
xor U24744 (N_24744,N_15814,N_15402);
nand U24745 (N_24745,N_19215,N_17623);
nand U24746 (N_24746,N_16895,N_18033);
or U24747 (N_24747,N_15711,N_18541);
nand U24748 (N_24748,N_19084,N_18381);
and U24749 (N_24749,N_16178,N_18649);
nand U24750 (N_24750,N_15697,N_17301);
nand U24751 (N_24751,N_19548,N_17896);
or U24752 (N_24752,N_16112,N_17030);
and U24753 (N_24753,N_17778,N_17784);
nand U24754 (N_24754,N_17973,N_19176);
nor U24755 (N_24755,N_19713,N_17772);
nand U24756 (N_24756,N_16947,N_15982);
and U24757 (N_24757,N_18741,N_19285);
nor U24758 (N_24758,N_19837,N_18156);
or U24759 (N_24759,N_17364,N_16617);
nand U24760 (N_24760,N_17944,N_15813);
nor U24761 (N_24761,N_17662,N_15302);
and U24762 (N_24762,N_15265,N_18185);
nor U24763 (N_24763,N_19915,N_18059);
or U24764 (N_24764,N_16803,N_18871);
nor U24765 (N_24765,N_18533,N_18485);
nor U24766 (N_24766,N_15588,N_17592);
xnor U24767 (N_24767,N_16985,N_17947);
nor U24768 (N_24768,N_19044,N_16473);
nand U24769 (N_24769,N_18908,N_19881);
xor U24770 (N_24770,N_18998,N_16892);
and U24771 (N_24771,N_16985,N_18894);
or U24772 (N_24772,N_15220,N_18579);
nor U24773 (N_24773,N_19340,N_16009);
xor U24774 (N_24774,N_19019,N_15160);
xnor U24775 (N_24775,N_18524,N_18526);
nor U24776 (N_24776,N_19547,N_19744);
nor U24777 (N_24777,N_16203,N_16436);
or U24778 (N_24778,N_15766,N_15863);
nand U24779 (N_24779,N_16944,N_15150);
and U24780 (N_24780,N_15942,N_19146);
nor U24781 (N_24781,N_19619,N_19372);
nand U24782 (N_24782,N_19757,N_15390);
and U24783 (N_24783,N_19429,N_15682);
or U24784 (N_24784,N_17353,N_19748);
nand U24785 (N_24785,N_15927,N_17677);
nor U24786 (N_24786,N_15525,N_16451);
or U24787 (N_24787,N_16366,N_15347);
xor U24788 (N_24788,N_17193,N_19383);
or U24789 (N_24789,N_18974,N_18311);
xnor U24790 (N_24790,N_19902,N_17123);
xor U24791 (N_24791,N_17543,N_16812);
nand U24792 (N_24792,N_16773,N_19381);
nand U24793 (N_24793,N_17666,N_18590);
and U24794 (N_24794,N_17522,N_17735);
and U24795 (N_24795,N_17455,N_19837);
or U24796 (N_24796,N_17389,N_16679);
xnor U24797 (N_24797,N_16744,N_19006);
or U24798 (N_24798,N_18251,N_17704);
or U24799 (N_24799,N_19914,N_16005);
nand U24800 (N_24800,N_17698,N_17483);
xnor U24801 (N_24801,N_18799,N_15580);
and U24802 (N_24802,N_17836,N_15535);
xor U24803 (N_24803,N_19290,N_15528);
nor U24804 (N_24804,N_15942,N_18201);
and U24805 (N_24805,N_18533,N_15310);
nor U24806 (N_24806,N_15659,N_16558);
xnor U24807 (N_24807,N_17786,N_19637);
nand U24808 (N_24808,N_17000,N_15705);
and U24809 (N_24809,N_17188,N_18269);
nand U24810 (N_24810,N_19415,N_18187);
nand U24811 (N_24811,N_16885,N_17837);
xor U24812 (N_24812,N_18234,N_17853);
nand U24813 (N_24813,N_19642,N_19057);
nand U24814 (N_24814,N_17005,N_16454);
nand U24815 (N_24815,N_18081,N_16935);
nor U24816 (N_24816,N_16385,N_15914);
xor U24817 (N_24817,N_18325,N_19491);
or U24818 (N_24818,N_15432,N_15659);
or U24819 (N_24819,N_19081,N_19358);
and U24820 (N_24820,N_15664,N_16326);
nor U24821 (N_24821,N_15299,N_15533);
nand U24822 (N_24822,N_19223,N_18212);
xor U24823 (N_24823,N_19255,N_15797);
or U24824 (N_24824,N_15998,N_19361);
nand U24825 (N_24825,N_15670,N_17517);
or U24826 (N_24826,N_15677,N_17384);
and U24827 (N_24827,N_17571,N_15828);
or U24828 (N_24828,N_15916,N_18323);
and U24829 (N_24829,N_17071,N_16463);
xnor U24830 (N_24830,N_18134,N_15023);
nor U24831 (N_24831,N_15764,N_17819);
xor U24832 (N_24832,N_15400,N_18325);
nand U24833 (N_24833,N_16427,N_15446);
nor U24834 (N_24834,N_16239,N_19824);
xor U24835 (N_24835,N_16981,N_19720);
nand U24836 (N_24836,N_19281,N_16020);
nor U24837 (N_24837,N_16756,N_19235);
xnor U24838 (N_24838,N_19302,N_17175);
or U24839 (N_24839,N_19418,N_19909);
xnor U24840 (N_24840,N_17631,N_18439);
xnor U24841 (N_24841,N_17979,N_18206);
and U24842 (N_24842,N_17021,N_16682);
nand U24843 (N_24843,N_15495,N_18755);
xnor U24844 (N_24844,N_19047,N_17011);
xor U24845 (N_24845,N_17831,N_19436);
and U24846 (N_24846,N_18280,N_15335);
xor U24847 (N_24847,N_17825,N_18533);
or U24848 (N_24848,N_17718,N_17619);
nand U24849 (N_24849,N_17538,N_17894);
and U24850 (N_24850,N_17624,N_17256);
xor U24851 (N_24851,N_15846,N_17315);
nor U24852 (N_24852,N_16918,N_17492);
or U24853 (N_24853,N_19166,N_15053);
xnor U24854 (N_24854,N_18185,N_17542);
xnor U24855 (N_24855,N_17045,N_15899);
or U24856 (N_24856,N_19603,N_16779);
or U24857 (N_24857,N_19563,N_15605);
nand U24858 (N_24858,N_18430,N_15792);
nor U24859 (N_24859,N_17338,N_17631);
or U24860 (N_24860,N_16546,N_18028);
and U24861 (N_24861,N_16962,N_18670);
xnor U24862 (N_24862,N_19452,N_17077);
xnor U24863 (N_24863,N_18918,N_16396);
xnor U24864 (N_24864,N_18041,N_18481);
nand U24865 (N_24865,N_17180,N_18114);
xor U24866 (N_24866,N_18644,N_16519);
nor U24867 (N_24867,N_18649,N_19291);
and U24868 (N_24868,N_15879,N_15515);
or U24869 (N_24869,N_17041,N_19755);
nand U24870 (N_24870,N_18663,N_15933);
and U24871 (N_24871,N_18004,N_18858);
and U24872 (N_24872,N_18795,N_16719);
nand U24873 (N_24873,N_16676,N_17722);
or U24874 (N_24874,N_18703,N_19798);
xnor U24875 (N_24875,N_17053,N_17617);
xnor U24876 (N_24876,N_17616,N_19946);
or U24877 (N_24877,N_18000,N_16180);
xor U24878 (N_24878,N_17591,N_18183);
xor U24879 (N_24879,N_18761,N_16016);
nand U24880 (N_24880,N_19992,N_15044);
nor U24881 (N_24881,N_17449,N_17972);
and U24882 (N_24882,N_19682,N_16501);
or U24883 (N_24883,N_17847,N_15303);
nor U24884 (N_24884,N_15762,N_15363);
and U24885 (N_24885,N_18323,N_16776);
xor U24886 (N_24886,N_16862,N_17809);
and U24887 (N_24887,N_17819,N_15628);
nor U24888 (N_24888,N_16825,N_18925);
or U24889 (N_24889,N_16359,N_16252);
and U24890 (N_24890,N_16368,N_19615);
xnor U24891 (N_24891,N_18472,N_18348);
nand U24892 (N_24892,N_19922,N_17113);
nor U24893 (N_24893,N_15948,N_18891);
nand U24894 (N_24894,N_15601,N_17166);
nor U24895 (N_24895,N_15304,N_17484);
nor U24896 (N_24896,N_19329,N_19238);
and U24897 (N_24897,N_19453,N_16840);
nor U24898 (N_24898,N_17152,N_19700);
xnor U24899 (N_24899,N_19240,N_15046);
nor U24900 (N_24900,N_15836,N_15203);
xor U24901 (N_24901,N_15096,N_18485);
and U24902 (N_24902,N_18260,N_18369);
xor U24903 (N_24903,N_17400,N_16002);
and U24904 (N_24904,N_17040,N_18551);
nand U24905 (N_24905,N_18923,N_19129);
nor U24906 (N_24906,N_15240,N_16477);
xor U24907 (N_24907,N_17884,N_18158);
nand U24908 (N_24908,N_16653,N_19328);
or U24909 (N_24909,N_19024,N_17455);
nor U24910 (N_24910,N_18142,N_18690);
and U24911 (N_24911,N_16853,N_19587);
or U24912 (N_24912,N_19959,N_15272);
xnor U24913 (N_24913,N_15988,N_19730);
and U24914 (N_24914,N_18953,N_15319);
or U24915 (N_24915,N_18731,N_17931);
or U24916 (N_24916,N_18723,N_18526);
nand U24917 (N_24917,N_19346,N_17365);
nand U24918 (N_24918,N_19662,N_16137);
and U24919 (N_24919,N_19352,N_15157);
and U24920 (N_24920,N_19750,N_19463);
nor U24921 (N_24921,N_15899,N_19232);
or U24922 (N_24922,N_16546,N_19830);
xnor U24923 (N_24923,N_16644,N_18623);
or U24924 (N_24924,N_19428,N_17191);
nand U24925 (N_24925,N_17087,N_19752);
xor U24926 (N_24926,N_15156,N_16558);
nand U24927 (N_24927,N_15416,N_18802);
nor U24928 (N_24928,N_17905,N_17175);
nand U24929 (N_24929,N_15997,N_16351);
or U24930 (N_24930,N_18318,N_19746);
or U24931 (N_24931,N_18690,N_17357);
nor U24932 (N_24932,N_15713,N_17235);
nor U24933 (N_24933,N_17932,N_19232);
nand U24934 (N_24934,N_16706,N_17440);
nor U24935 (N_24935,N_19166,N_16790);
or U24936 (N_24936,N_18396,N_16075);
nor U24937 (N_24937,N_17762,N_19356);
and U24938 (N_24938,N_16389,N_15194);
nor U24939 (N_24939,N_15406,N_15901);
or U24940 (N_24940,N_17132,N_16704);
and U24941 (N_24941,N_19030,N_15109);
xor U24942 (N_24942,N_16179,N_15951);
xnor U24943 (N_24943,N_16270,N_15898);
xor U24944 (N_24944,N_17486,N_16308);
nor U24945 (N_24945,N_19242,N_15337);
nand U24946 (N_24946,N_18525,N_15288);
nor U24947 (N_24947,N_17035,N_18005);
nand U24948 (N_24948,N_16386,N_18231);
or U24949 (N_24949,N_15914,N_15985);
xor U24950 (N_24950,N_17976,N_16770);
or U24951 (N_24951,N_16357,N_15590);
xnor U24952 (N_24952,N_15945,N_19930);
and U24953 (N_24953,N_18770,N_15483);
xor U24954 (N_24954,N_16428,N_16273);
or U24955 (N_24955,N_19004,N_17161);
nand U24956 (N_24956,N_19124,N_16181);
xor U24957 (N_24957,N_16710,N_16476);
or U24958 (N_24958,N_18772,N_18367);
xor U24959 (N_24959,N_19133,N_17475);
or U24960 (N_24960,N_18014,N_15121);
nor U24961 (N_24961,N_15461,N_17483);
nor U24962 (N_24962,N_16982,N_15196);
xnor U24963 (N_24963,N_18904,N_19519);
or U24964 (N_24964,N_19254,N_16872);
nand U24965 (N_24965,N_16645,N_18774);
nor U24966 (N_24966,N_15962,N_19026);
xnor U24967 (N_24967,N_18168,N_16415);
and U24968 (N_24968,N_18845,N_17621);
xnor U24969 (N_24969,N_18983,N_16009);
nand U24970 (N_24970,N_18517,N_19216);
nand U24971 (N_24971,N_19249,N_17075);
xnor U24972 (N_24972,N_19432,N_19380);
nor U24973 (N_24973,N_18041,N_19508);
and U24974 (N_24974,N_15434,N_18536);
and U24975 (N_24975,N_16573,N_16951);
nand U24976 (N_24976,N_15919,N_19675);
and U24977 (N_24977,N_17196,N_18828);
nor U24978 (N_24978,N_18132,N_17220);
or U24979 (N_24979,N_17495,N_16812);
nand U24980 (N_24980,N_15751,N_16332);
and U24981 (N_24981,N_18257,N_19107);
nor U24982 (N_24982,N_17974,N_16107);
xnor U24983 (N_24983,N_15831,N_16807);
nor U24984 (N_24984,N_18345,N_19446);
nor U24985 (N_24985,N_19415,N_18565);
nand U24986 (N_24986,N_15658,N_19141);
nor U24987 (N_24987,N_18510,N_18651);
or U24988 (N_24988,N_19399,N_19173);
and U24989 (N_24989,N_18582,N_15707);
and U24990 (N_24990,N_17656,N_16125);
and U24991 (N_24991,N_16901,N_15373);
xor U24992 (N_24992,N_16345,N_15288);
nand U24993 (N_24993,N_18182,N_19056);
or U24994 (N_24994,N_19950,N_18275);
or U24995 (N_24995,N_15785,N_16056);
nand U24996 (N_24996,N_18441,N_18742);
or U24997 (N_24997,N_18311,N_15407);
nor U24998 (N_24998,N_15227,N_16208);
nand U24999 (N_24999,N_15638,N_16340);
nor U25000 (N_25000,N_20504,N_23235);
xnor U25001 (N_25001,N_22771,N_23834);
nand U25002 (N_25002,N_24480,N_20176);
nand U25003 (N_25003,N_22480,N_20101);
nor U25004 (N_25004,N_21741,N_23978);
xor U25005 (N_25005,N_22744,N_21284);
nor U25006 (N_25006,N_22093,N_24328);
xnor U25007 (N_25007,N_23273,N_23988);
and U25008 (N_25008,N_23347,N_24377);
or U25009 (N_25009,N_24993,N_21313);
nor U25010 (N_25010,N_23511,N_21645);
xor U25011 (N_25011,N_22784,N_22357);
and U25012 (N_25012,N_23109,N_21420);
and U25013 (N_25013,N_20384,N_24374);
nor U25014 (N_25014,N_23787,N_23086);
nand U25015 (N_25015,N_24369,N_22290);
xnor U25016 (N_25016,N_24709,N_20635);
nand U25017 (N_25017,N_22007,N_22871);
and U25018 (N_25018,N_23369,N_23823);
nor U25019 (N_25019,N_23845,N_23772);
xnor U25020 (N_25020,N_22176,N_20732);
nor U25021 (N_25021,N_23567,N_23015);
and U25022 (N_25022,N_22205,N_23091);
nand U25023 (N_25023,N_23625,N_23671);
xor U25024 (N_25024,N_23357,N_23316);
nor U25025 (N_25025,N_23938,N_22616);
and U25026 (N_25026,N_22360,N_21646);
xnor U25027 (N_25027,N_20116,N_20055);
nor U25028 (N_25028,N_21933,N_20302);
nand U25029 (N_25029,N_22502,N_22371);
nand U25030 (N_25030,N_22299,N_21263);
or U25031 (N_25031,N_21002,N_20427);
nand U25032 (N_25032,N_23519,N_24692);
nor U25033 (N_25033,N_24782,N_24247);
nand U25034 (N_25034,N_23844,N_21943);
xor U25035 (N_25035,N_23523,N_22722);
nand U25036 (N_25036,N_23463,N_20725);
nor U25037 (N_25037,N_22317,N_22970);
xor U25038 (N_25038,N_23001,N_21948);
nor U25039 (N_25039,N_22495,N_21049);
or U25040 (N_25040,N_24125,N_23478);
or U25041 (N_25041,N_24655,N_21044);
nor U25042 (N_25042,N_24508,N_24264);
xor U25043 (N_25043,N_22267,N_22258);
or U25044 (N_25044,N_22080,N_23635);
nand U25045 (N_25045,N_23547,N_24477);
nand U25046 (N_25046,N_20373,N_22174);
nand U25047 (N_25047,N_20202,N_21012);
xor U25048 (N_25048,N_24471,N_22570);
nor U25049 (N_25049,N_22583,N_22352);
and U25050 (N_25050,N_24585,N_21866);
or U25051 (N_25051,N_23422,N_22454);
xor U25052 (N_25052,N_24548,N_22433);
xnor U25053 (N_25053,N_20749,N_24953);
and U25054 (N_25054,N_22972,N_21843);
xor U25055 (N_25055,N_21615,N_21084);
or U25056 (N_25056,N_20014,N_22919);
or U25057 (N_25057,N_23892,N_20882);
nor U25058 (N_25058,N_21549,N_20412);
and U25059 (N_25059,N_21105,N_20807);
and U25060 (N_25060,N_24493,N_23609);
nor U25061 (N_25061,N_24600,N_21216);
or U25062 (N_25062,N_22119,N_23502);
nand U25063 (N_25063,N_22742,N_23954);
or U25064 (N_25064,N_24997,N_24140);
xnor U25065 (N_25065,N_21592,N_24873);
nand U25066 (N_25066,N_21042,N_22032);
xor U25067 (N_25067,N_21046,N_20716);
xor U25068 (N_25068,N_22941,N_21715);
or U25069 (N_25069,N_22719,N_22362);
xor U25070 (N_25070,N_20124,N_20416);
xnor U25071 (N_25071,N_20540,N_24014);
xor U25072 (N_25072,N_24973,N_21782);
or U25073 (N_25073,N_22144,N_21818);
xnor U25074 (N_25074,N_23971,N_22687);
and U25075 (N_25075,N_24724,N_22387);
nor U25076 (N_25076,N_22527,N_24384);
nor U25077 (N_25077,N_24142,N_21480);
or U25078 (N_25078,N_21725,N_24312);
nor U25079 (N_25079,N_24964,N_21026);
xnor U25080 (N_25080,N_21990,N_22667);
nand U25081 (N_25081,N_21637,N_24040);
nand U25082 (N_25082,N_20328,N_24778);
nor U25083 (N_25083,N_22643,N_23364);
nor U25084 (N_25084,N_22295,N_24892);
xnor U25085 (N_25085,N_20814,N_24875);
and U25086 (N_25086,N_21817,N_20399);
or U25087 (N_25087,N_21240,N_23754);
nor U25088 (N_25088,N_23883,N_21522);
nor U25089 (N_25089,N_20354,N_22228);
xnor U25090 (N_25090,N_23393,N_23918);
and U25091 (N_25091,N_23376,N_21217);
xor U25092 (N_25092,N_21078,N_21429);
nand U25093 (N_25093,N_22653,N_20080);
or U25094 (N_25094,N_22512,N_23919);
xnor U25095 (N_25095,N_23542,N_22861);
or U25096 (N_25096,N_23569,N_20349);
and U25097 (N_25097,N_22854,N_24888);
and U25098 (N_25098,N_24524,N_23668);
and U25099 (N_25099,N_21542,N_22876);
xnor U25100 (N_25100,N_21022,N_23072);
and U25101 (N_25101,N_24760,N_24042);
nor U25102 (N_25102,N_21041,N_20190);
and U25103 (N_25103,N_20403,N_22928);
nor U25104 (N_25104,N_21932,N_22005);
xor U25105 (N_25105,N_24478,N_21714);
nor U25106 (N_25106,N_20198,N_23512);
or U25107 (N_25107,N_22600,N_20062);
and U25108 (N_25108,N_24295,N_20338);
nor U25109 (N_25109,N_20441,N_22903);
and U25110 (N_25110,N_20479,N_23476);
nand U25111 (N_25111,N_24966,N_22549);
nor U25112 (N_25112,N_23417,N_23014);
nor U25113 (N_25113,N_21872,N_24206);
nor U25114 (N_25114,N_24425,N_20229);
nor U25115 (N_25115,N_22816,N_21811);
nand U25116 (N_25116,N_20144,N_24667);
xnor U25117 (N_25117,N_21917,N_21833);
xnor U25118 (N_25118,N_20396,N_21267);
or U25119 (N_25119,N_21381,N_22048);
nor U25120 (N_25120,N_20942,N_21836);
nand U25121 (N_25121,N_21772,N_22640);
nand U25122 (N_25122,N_24912,N_20858);
nand U25123 (N_25123,N_20836,N_21854);
nor U25124 (N_25124,N_24913,N_21861);
nand U25125 (N_25125,N_20787,N_20561);
xnor U25126 (N_25126,N_20761,N_22206);
nand U25127 (N_25127,N_23809,N_24194);
xor U25128 (N_25128,N_20555,N_21186);
and U25129 (N_25129,N_24470,N_21413);
and U25130 (N_25130,N_24451,N_21457);
nand U25131 (N_25131,N_23033,N_22444);
and U25132 (N_25132,N_23193,N_22723);
nand U25133 (N_25133,N_20805,N_20829);
and U25134 (N_25134,N_20015,N_24544);
nand U25135 (N_25135,N_21510,N_21193);
xor U25136 (N_25136,N_21979,N_22629);
xor U25137 (N_25137,N_23751,N_24057);
nand U25138 (N_25138,N_23020,N_20218);
nor U25139 (N_25139,N_22329,N_24924);
or U25140 (N_25140,N_21210,N_21226);
nand U25141 (N_25141,N_24276,N_22323);
nand U25142 (N_25142,N_24519,N_24530);
or U25143 (N_25143,N_21143,N_21517);
xor U25144 (N_25144,N_20030,N_24895);
or U25145 (N_25145,N_22756,N_24688);
xor U25146 (N_25146,N_20899,N_21058);
nand U25147 (N_25147,N_22171,N_24004);
xor U25148 (N_25148,N_20040,N_24539);
nor U25149 (N_25149,N_21898,N_21584);
and U25150 (N_25150,N_24996,N_21635);
xor U25151 (N_25151,N_24638,N_22960);
nand U25152 (N_25152,N_24754,N_21163);
and U25153 (N_25153,N_23113,N_21047);
nand U25154 (N_25154,N_24881,N_22259);
nor U25155 (N_25155,N_23474,N_23815);
nor U25156 (N_25156,N_24126,N_24624);
nor U25157 (N_25157,N_20099,N_24383);
and U25158 (N_25158,N_20126,N_21994);
or U25159 (N_25159,N_21737,N_21452);
or U25160 (N_25160,N_23669,N_23544);
nand U25161 (N_25161,N_21273,N_24682);
nor U25162 (N_25162,N_23793,N_22358);
nor U25163 (N_25163,N_22392,N_21529);
nor U25164 (N_25164,N_20081,N_21754);
and U25165 (N_25165,N_24923,N_23881);
and U25166 (N_25166,N_20930,N_23570);
and U25167 (N_25167,N_23025,N_21072);
and U25168 (N_25168,N_24424,N_21770);
nand U25169 (N_25169,N_22402,N_21339);
xor U25170 (N_25170,N_23945,N_21649);
nand U25171 (N_25171,N_21281,N_22375);
nor U25172 (N_25172,N_23348,N_23225);
xnor U25173 (N_25173,N_20944,N_23755);
or U25174 (N_25174,N_23308,N_20178);
nand U25175 (N_25175,N_21805,N_23377);
nand U25176 (N_25176,N_24339,N_23785);
or U25177 (N_25177,N_20020,N_24550);
or U25178 (N_25178,N_20448,N_20609);
and U25179 (N_25179,N_21519,N_24486);
and U25180 (N_25180,N_21242,N_21056);
and U25181 (N_25181,N_21853,N_22630);
or U25182 (N_25182,N_21513,N_20119);
and U25183 (N_25183,N_24664,N_23598);
and U25184 (N_25184,N_22904,N_22155);
nand U25185 (N_25185,N_24410,N_20627);
and U25186 (N_25186,N_20738,N_24442);
and U25187 (N_25187,N_24735,N_24504);
or U25188 (N_25188,N_23730,N_22597);
xnor U25189 (N_25189,N_20482,N_21369);
nor U25190 (N_25190,N_23638,N_20687);
nand U25191 (N_25191,N_24189,N_22364);
nand U25192 (N_25192,N_21241,N_22849);
xnor U25193 (N_25193,N_22445,N_24208);
xor U25194 (N_25194,N_24313,N_20951);
and U25195 (N_25195,N_24070,N_21254);
and U25196 (N_25196,N_21135,N_23155);
nor U25197 (N_25197,N_24498,N_22002);
nand U25198 (N_25198,N_22733,N_24263);
or U25199 (N_25199,N_20681,N_23851);
or U25200 (N_25200,N_21486,N_21523);
nand U25201 (N_25201,N_21015,N_22526);
nor U25202 (N_25202,N_22421,N_24644);
and U25203 (N_25203,N_20445,N_21613);
nand U25204 (N_25204,N_23263,N_24261);
nand U25205 (N_25205,N_22844,N_22031);
nand U25206 (N_25206,N_22846,N_24121);
nor U25207 (N_25207,N_24378,N_21891);
or U25208 (N_25208,N_20327,N_21655);
xnor U25209 (N_25209,N_20606,N_21699);
xor U25210 (N_25210,N_22054,N_21156);
or U25211 (N_25211,N_21100,N_20893);
nor U25212 (N_25212,N_20850,N_21051);
nand U25213 (N_25213,N_20250,N_23061);
nor U25214 (N_25214,N_23021,N_21200);
nand U25215 (N_25215,N_24526,N_22191);
or U25216 (N_25216,N_24691,N_23035);
nand U25217 (N_25217,N_24930,N_23739);
or U25218 (N_25218,N_20634,N_23990);
xnor U25219 (N_25219,N_21469,N_23993);
nand U25220 (N_25220,N_24491,N_22069);
or U25221 (N_25221,N_23734,N_22310);
nand U25222 (N_25222,N_23168,N_22948);
xnor U25223 (N_25223,N_23367,N_22099);
and U25224 (N_25224,N_21370,N_23160);
nand U25225 (N_25225,N_22927,N_20209);
or U25226 (N_25226,N_22049,N_20310);
xnor U25227 (N_25227,N_22661,N_23176);
nor U25228 (N_25228,N_20623,N_24641);
nor U25229 (N_25229,N_23584,N_24858);
xnor U25230 (N_25230,N_23071,N_24635);
nor U25231 (N_25231,N_20969,N_21676);
nand U25232 (N_25232,N_20484,N_24299);
nand U25233 (N_25233,N_24080,N_20923);
and U25234 (N_25234,N_22071,N_24262);
xor U25235 (N_25235,N_21427,N_24325);
nand U25236 (N_25236,N_24932,N_23447);
nor U25237 (N_25237,N_21619,N_24693);
and U25238 (N_25238,N_24010,N_22405);
and U25239 (N_25239,N_23283,N_24193);
nand U25240 (N_25240,N_22935,N_21177);
nor U25241 (N_25241,N_21985,N_21206);
xor U25242 (N_25242,N_23878,N_20877);
nor U25243 (N_25243,N_21142,N_22969);
xnor U25244 (N_25244,N_23178,N_23663);
and U25245 (N_25245,N_23788,N_24007);
xor U25246 (N_25246,N_22247,N_23192);
nand U25247 (N_25247,N_24429,N_24363);
and U25248 (N_25248,N_24173,N_20919);
nor U25249 (N_25249,N_20977,N_21577);
xnor U25250 (N_25250,N_22396,N_24686);
or U25251 (N_25251,N_23451,N_23023);
nand U25252 (N_25252,N_21773,N_24166);
nor U25253 (N_25253,N_20414,N_24707);
or U25254 (N_25254,N_22864,N_23218);
nor U25255 (N_25255,N_22254,N_24191);
xor U25256 (N_25256,N_22499,N_20108);
xnor U25257 (N_25257,N_23290,N_24153);
nor U25258 (N_25258,N_21280,N_22797);
xor U25259 (N_25259,N_21298,N_21272);
or U25260 (N_25260,N_23649,N_22209);
nand U25261 (N_25261,N_24000,N_22509);
xor U25262 (N_25262,N_23282,N_24331);
xor U25263 (N_25263,N_23477,N_23890);
or U25264 (N_25264,N_22645,N_22278);
nor U25265 (N_25265,N_24116,N_20968);
xor U25266 (N_25266,N_22465,N_20656);
nand U25267 (N_25267,N_23172,N_23572);
nor U25268 (N_25268,N_20910,N_23517);
or U25269 (N_25269,N_23041,N_23145);
and U25270 (N_25270,N_20762,N_21461);
nand U25271 (N_25271,N_21398,N_22143);
or U25272 (N_25272,N_20164,N_22218);
xor U25273 (N_25273,N_22442,N_21867);
nor U25274 (N_25274,N_20451,N_22335);
xor U25275 (N_25275,N_21809,N_21344);
nor U25276 (N_25276,N_24254,N_21875);
nor U25277 (N_25277,N_20402,N_21487);
nand U25278 (N_25278,N_23704,N_22452);
nor U25279 (N_25279,N_22417,N_21261);
or U25280 (N_25280,N_24500,N_24948);
nor U25281 (N_25281,N_21329,N_22468);
xnor U25282 (N_25282,N_20098,N_24001);
nand U25283 (N_25283,N_23827,N_23532);
xor U25284 (N_25284,N_23937,N_20652);
and U25285 (N_25285,N_21382,N_23317);
and U25286 (N_25286,N_22165,N_24677);
and U25287 (N_25287,N_24711,N_21746);
and U25288 (N_25288,N_20519,N_23770);
nand U25289 (N_25289,N_22727,N_20813);
and U25290 (N_25290,N_22072,N_21835);
xnor U25291 (N_25291,N_22710,N_22141);
nand U25292 (N_25292,N_22152,N_20068);
xnor U25293 (N_25293,N_20167,N_20881);
and U25294 (N_25294,N_21325,N_21279);
xnor U25295 (N_25295,N_21717,N_20425);
nor U25296 (N_25296,N_23483,N_20952);
nor U25297 (N_25297,N_23104,N_22656);
nor U25298 (N_25298,N_23498,N_24492);
and U25299 (N_25299,N_23245,N_22252);
nor U25300 (N_25300,N_20503,N_24083);
or U25301 (N_25301,N_21838,N_21219);
xnor U25302 (N_25302,N_20525,N_23833);
or U25303 (N_25303,N_24859,N_24386);
and U25304 (N_25304,N_22859,N_20802);
xnor U25305 (N_25305,N_21978,N_23154);
nor U25306 (N_25306,N_20689,N_22293);
nor U25307 (N_25307,N_21930,N_20215);
and U25308 (N_25308,N_23475,N_23301);
xnor U25309 (N_25309,N_24257,N_21019);
nor U25310 (N_25310,N_20397,N_21133);
nor U25311 (N_25311,N_20498,N_23051);
and U25312 (N_25312,N_22520,N_23431);
xnor U25313 (N_25313,N_21903,N_23928);
nand U25314 (N_25314,N_24808,N_22251);
or U25315 (N_25315,N_24370,N_20568);
nand U25316 (N_25316,N_21587,N_24931);
and U25317 (N_25317,N_20735,N_22697);
and U25318 (N_25318,N_23497,N_21724);
nand U25319 (N_25319,N_22325,N_22246);
and U25320 (N_25320,N_24949,N_23921);
xnor U25321 (N_25321,N_23875,N_21976);
and U25322 (N_25322,N_21851,N_21849);
and U25323 (N_25323,N_23070,N_21421);
nand U25324 (N_25324,N_21781,N_20960);
nand U25325 (N_25325,N_24285,N_20292);
and U25326 (N_25326,N_21060,N_20613);
nor U25327 (N_25327,N_22470,N_20758);
xor U25328 (N_25328,N_21463,N_22106);
nand U25329 (N_25329,N_21547,N_23737);
nand U25330 (N_25330,N_20905,N_24184);
nor U25331 (N_25331,N_21799,N_22937);
nor U25332 (N_25332,N_20010,N_21251);
and U25333 (N_25333,N_24183,N_21098);
xnor U25334 (N_25334,N_20494,N_22020);
xor U25335 (N_25335,N_24998,N_24666);
nor U25336 (N_25336,N_21119,N_23075);
xor U25337 (N_25337,N_24016,N_24460);
or U25338 (N_25338,N_23262,N_24834);
xor U25339 (N_25339,N_22166,N_24965);
and U25340 (N_25340,N_24514,N_21150);
xnor U25341 (N_25341,N_20457,N_22573);
nand U25342 (N_25342,N_23757,N_20261);
nand U25343 (N_25343,N_20563,N_22706);
nor U25344 (N_25344,N_23661,N_24642);
nand U25345 (N_25345,N_21684,N_23555);
xnor U25346 (N_25346,N_22092,N_21085);
xnor U25347 (N_25347,N_23637,N_22917);
and U25348 (N_25348,N_20665,N_24018);
nand U25349 (N_25349,N_23681,N_21199);
xnor U25350 (N_25350,N_21104,N_21407);
nor U25351 (N_25351,N_20811,N_24592);
and U25352 (N_25352,N_24303,N_21692);
or U25353 (N_25353,N_22493,N_22224);
nand U25354 (N_25354,N_23097,N_24758);
xnor U25355 (N_25355,N_23974,N_24154);
nor U25356 (N_25356,N_23471,N_20926);
or U25357 (N_25357,N_24110,N_21785);
nand U25358 (N_25358,N_20047,N_23366);
xnor U25359 (N_25359,N_23127,N_23198);
nand U25360 (N_25360,N_21195,N_21379);
or U25361 (N_25361,N_21550,N_21639);
nand U25362 (N_25362,N_20784,N_24269);
or U25363 (N_25363,N_24177,N_24708);
nand U25364 (N_25364,N_24938,N_23655);
and U25365 (N_25365,N_20175,N_21732);
xor U25366 (N_25366,N_24929,N_24444);
xnor U25367 (N_25367,N_24375,N_20468);
xor U25368 (N_25368,N_23931,N_23752);
nor U25369 (N_25369,N_23749,N_22262);
or U25370 (N_25370,N_23666,N_20203);
or U25371 (N_25371,N_21102,N_20793);
or U25372 (N_25372,N_24676,N_20490);
nand U25373 (N_25373,N_21146,N_22306);
xnor U25374 (N_25374,N_22632,N_23568);
nor U25375 (N_25375,N_24521,N_23210);
xnor U25376 (N_25376,N_20812,N_23191);
xor U25377 (N_25377,N_21360,N_22225);
and U25378 (N_25378,N_24174,N_20618);
nand U25379 (N_25379,N_22473,N_24487);
nor U25380 (N_25380,N_23406,N_22648);
or U25381 (N_25381,N_23966,N_22955);
and U25382 (N_25382,N_24773,N_20674);
nand U25383 (N_25383,N_22507,N_24237);
nand U25384 (N_25384,N_22750,N_20573);
or U25385 (N_25385,N_23370,N_20100);
xor U25386 (N_25386,N_22582,N_23100);
nor U25387 (N_25387,N_23571,N_21695);
xor U25388 (N_25388,N_22647,N_23505);
xor U25389 (N_25389,N_23839,N_23731);
nor U25390 (N_25390,N_21942,N_24739);
and U25391 (N_25391,N_22068,N_21808);
xor U25392 (N_25392,N_23373,N_23232);
xor U25393 (N_25393,N_23684,N_22595);
and U25394 (N_25394,N_20820,N_20360);
nand U25395 (N_25395,N_21634,N_21496);
nor U25396 (N_25396,N_22558,N_24265);
nor U25397 (N_25397,N_24823,N_20703);
nand U25398 (N_25398,N_24025,N_22688);
nor U25399 (N_25399,N_24430,N_24556);
nand U25400 (N_25400,N_22460,N_20326);
xor U25401 (N_25401,N_22250,N_22256);
and U25402 (N_25402,N_22212,N_24196);
nor U25403 (N_25403,N_20883,N_21905);
nor U25404 (N_25404,N_22944,N_22178);
or U25405 (N_25405,N_23284,N_20998);
nand U25406 (N_25406,N_21071,N_21077);
xor U25407 (N_25407,N_21266,N_22901);
nand U25408 (N_25408,N_23115,N_21340);
xor U25409 (N_25409,N_20174,N_22283);
nor U25410 (N_25410,N_22231,N_20273);
and U25411 (N_25411,N_20604,N_22279);
xnor U25412 (N_25412,N_21045,N_23083);
nor U25413 (N_25413,N_20120,N_23608);
xor U25414 (N_25414,N_20879,N_23820);
nand U25415 (N_25415,N_24417,N_22270);
and U25416 (N_25416,N_22192,N_24286);
and U25417 (N_25417,N_20632,N_21963);
nand U25418 (N_25418,N_22950,N_23953);
nor U25419 (N_25419,N_22019,N_21696);
nor U25420 (N_25420,N_20916,N_24910);
nand U25421 (N_25421,N_23190,N_20011);
nand U25422 (N_25422,N_22959,N_23619);
and U25423 (N_25423,N_22091,N_24171);
nor U25424 (N_25424,N_24988,N_24054);
or U25425 (N_25425,N_22631,N_22971);
nand U25426 (N_25426,N_20012,N_23234);
and U25427 (N_25427,N_24974,N_24715);
or U25428 (N_25428,N_23328,N_21239);
nand U25429 (N_25429,N_20059,N_22676);
nor U25430 (N_25430,N_20323,N_20630);
xor U25431 (N_25431,N_22947,N_24774);
nor U25432 (N_25432,N_20036,N_21134);
nor U25433 (N_25433,N_20386,N_24844);
and U25434 (N_25434,N_21434,N_20972);
nand U25435 (N_25435,N_24723,N_24879);
nand U25436 (N_25436,N_20230,N_21801);
nand U25437 (N_25437,N_23553,N_24227);
nand U25438 (N_25438,N_24185,N_24647);
and U25439 (N_25439,N_23963,N_20564);
xor U25440 (N_25440,N_21238,N_20316);
xor U25441 (N_25441,N_21007,N_20382);
or U25442 (N_25442,N_23425,N_22617);
nor U25443 (N_25443,N_21097,N_23900);
xnor U25444 (N_25444,N_20935,N_23808);
and U25445 (N_25445,N_21418,N_21593);
or U25446 (N_25446,N_23776,N_23428);
and U25447 (N_25447,N_24400,N_23501);
nor U25448 (N_25448,N_20868,N_20289);
nor U25449 (N_25449,N_20443,N_21445);
or U25450 (N_25450,N_24020,N_22496);
nand U25451 (N_25451,N_23107,N_21346);
or U25452 (N_25452,N_24978,N_20009);
and U25453 (N_25453,N_22765,N_22660);
or U25454 (N_25454,N_20056,N_23027);
nor U25455 (N_25455,N_24608,N_21659);
xor U25456 (N_25456,N_20431,N_22151);
and U25457 (N_25457,N_22413,N_22187);
nand U25458 (N_25458,N_24045,N_23006);
and U25459 (N_25459,N_24673,N_21511);
nand U25460 (N_25460,N_21387,N_24882);
xnor U25461 (N_25461,N_21493,N_21556);
nor U25462 (N_25462,N_22348,N_24800);
nor U25463 (N_25463,N_22888,N_21812);
nor U25464 (N_25464,N_23645,N_22052);
and U25465 (N_25465,N_21599,N_24373);
nand U25466 (N_25466,N_24914,N_24065);
nor U25467 (N_25467,N_23390,N_21814);
nand U25468 (N_25468,N_21920,N_23520);
xor U25469 (N_25469,N_23819,N_24230);
nor U25470 (N_25470,N_20305,N_24736);
nand U25471 (N_25471,N_22931,N_20515);
or U25472 (N_25472,N_21825,N_23134);
and U25473 (N_25473,N_20590,N_20086);
xnor U25474 (N_25474,N_23654,N_22389);
or U25475 (N_25475,N_22240,N_22945);
nand U25476 (N_25476,N_20611,N_23226);
nor U25477 (N_25477,N_20122,N_22728);
nor U25478 (N_25478,N_23246,N_21385);
and U25479 (N_25479,N_20194,N_20072);
nor U25480 (N_25480,N_22977,N_20123);
nor U25481 (N_25481,N_20508,N_22566);
nand U25482 (N_25482,N_21464,N_23882);
and U25483 (N_25483,N_23840,N_24679);
nor U25484 (N_25484,N_22369,N_24405);
nand U25485 (N_25485,N_20708,N_23458);
nor U25486 (N_25486,N_24032,N_24406);
xnor U25487 (N_25487,N_23067,N_23549);
xnor U25488 (N_25488,N_21941,N_23457);
nand U25489 (N_25489,N_24385,N_24130);
or U25490 (N_25490,N_23643,N_23574);
xor U25491 (N_25491,N_23494,N_20254);
nand U25492 (N_25492,N_22973,N_24084);
or U25493 (N_25493,N_23439,N_20922);
nor U25494 (N_25494,N_24991,N_22025);
or U25495 (N_25495,N_23632,N_23142);
nor U25496 (N_25496,N_24041,N_23556);
and U25497 (N_25497,N_21802,N_21089);
or U25498 (N_25498,N_23504,N_21479);
and U25499 (N_25499,N_22746,N_23054);
xnor U25500 (N_25500,N_21597,N_23618);
or U25501 (N_25501,N_24776,N_21000);
nand U25502 (N_25502,N_23206,N_21531);
and U25503 (N_25503,N_20650,N_23338);
nand U25504 (N_25504,N_20024,N_21130);
and U25505 (N_25505,N_23897,N_20529);
nand U25506 (N_25506,N_23123,N_21443);
nand U25507 (N_25507,N_23472,N_24352);
and U25508 (N_25508,N_22911,N_24076);
and U25509 (N_25509,N_24761,N_22916);
xor U25510 (N_25510,N_20981,N_23078);
or U25511 (N_25511,N_24807,N_24567);
nor U25512 (N_25512,N_23453,N_22594);
xnor U25513 (N_25513,N_24740,N_24743);
nand U25514 (N_25514,N_20105,N_24008);
nor U25515 (N_25515,N_22281,N_20557);
xor U25516 (N_25516,N_20688,N_24201);
nand U25517 (N_25517,N_21878,N_22918);
or U25518 (N_25518,N_21178,N_21157);
nor U25519 (N_25519,N_22965,N_23410);
or U25520 (N_25520,N_22772,N_23438);
nand U25521 (N_25521,N_23540,N_22836);
nor U25522 (N_25522,N_23415,N_22510);
and U25523 (N_25523,N_22110,N_22029);
or U25524 (N_25524,N_24427,N_23899);
nor U25525 (N_25525,N_20240,N_24553);
and U25526 (N_25526,N_23727,N_22312);
xor U25527 (N_25527,N_23697,N_20361);
and U25528 (N_25528,N_20092,N_20343);
and U25529 (N_25529,N_22770,N_22196);
or U25530 (N_25530,N_23509,N_22008);
or U25531 (N_25531,N_20740,N_21879);
nor U25532 (N_25532,N_22115,N_22451);
nor U25533 (N_25533,N_22921,N_21483);
or U25534 (N_25534,N_21612,N_20842);
and U25535 (N_25535,N_21620,N_24928);
nand U25536 (N_25536,N_22415,N_23872);
nor U25537 (N_25537,N_21630,N_21710);
and U25538 (N_25538,N_23660,N_22966);
nand U25539 (N_25539,N_22793,N_20364);
nor U25540 (N_25540,N_24283,N_24476);
nor U25541 (N_25541,N_20900,N_23389);
and U25542 (N_25542,N_23199,N_23345);
and U25543 (N_25543,N_20137,N_20659);
and U25544 (N_25544,N_20466,N_21912);
xnor U25545 (N_25545,N_21532,N_21682);
xor U25546 (N_25546,N_23830,N_21196);
and U25547 (N_25547,N_20710,N_24234);
xor U25548 (N_25548,N_24055,N_20408);
xor U25549 (N_25549,N_22015,N_20633);
nor U25550 (N_25550,N_24391,N_22519);
or U25551 (N_25551,N_22162,N_23744);
nor U25552 (N_25552,N_22650,N_21175);
nor U25553 (N_25553,N_21537,N_23750);
and U25554 (N_25554,N_23514,N_24846);
or U25555 (N_25555,N_24983,N_22277);
or U25556 (N_25556,N_22500,N_20260);
xor U25557 (N_25557,N_23583,N_24023);
or U25558 (N_25558,N_23984,N_21489);
nor U25559 (N_25559,N_20410,N_24672);
or U25560 (N_25560,N_20661,N_23853);
and U25561 (N_25561,N_20363,N_20134);
and U25562 (N_25562,N_24522,N_20411);
xnor U25563 (N_25563,N_24064,N_24050);
and U25564 (N_25564,N_24138,N_23383);
xnor U25565 (N_25565,N_24179,N_23331);
or U25566 (N_25566,N_22654,N_22156);
and U25567 (N_25567,N_20959,N_22998);
nand U25568 (N_25568,N_23264,N_21295);
nor U25569 (N_25569,N_22203,N_20608);
nand U25570 (N_25570,N_22073,N_20393);
and U25571 (N_25571,N_23161,N_20587);
nor U25572 (N_25572,N_21111,N_20578);
or U25573 (N_25573,N_22300,N_21282);
xnor U25574 (N_25574,N_22365,N_21957);
and U25575 (N_25575,N_22575,N_21552);
and U25576 (N_25576,N_22796,N_21271);
nand U25577 (N_25577,N_20160,N_23189);
nor U25578 (N_25578,N_21362,N_20992);
and U25579 (N_25579,N_22211,N_24750);
xor U25580 (N_25580,N_21910,N_23258);
or U25581 (N_25581,N_21160,N_21769);
nor U25582 (N_25582,N_20131,N_21909);
nand U25583 (N_25583,N_20132,N_22145);
nand U25584 (N_25584,N_24623,N_20104);
nand U25585 (N_25585,N_24720,N_20827);
nand U25586 (N_25586,N_21099,N_23735);
nor U25587 (N_25587,N_23073,N_22410);
or U25588 (N_25588,N_22789,N_23880);
or U25589 (N_25589,N_23150,N_23724);
nand U25590 (N_25590,N_20896,N_23257);
nor U25591 (N_25591,N_21306,N_23854);
xor U25592 (N_25592,N_23329,N_21694);
nand U25593 (N_25593,N_22568,N_21914);
xnor U25594 (N_25594,N_22555,N_23024);
xnor U25595 (N_25595,N_24804,N_23495);
nand U25596 (N_25596,N_21484,N_21989);
nor U25597 (N_25597,N_20937,N_21829);
nor U25598 (N_25598,N_22716,N_22319);
nand U25599 (N_25599,N_21345,N_22378);
nand U25600 (N_25600,N_21426,N_22328);
xor U25601 (N_25601,N_24395,N_22628);
nand U25602 (N_25602,N_24925,N_20541);
nand U25603 (N_25603,N_24863,N_22128);
xnor U25604 (N_25604,N_24315,N_23324);
xor U25605 (N_25605,N_23614,N_22377);
nor U25606 (N_25606,N_24318,N_21245);
xor U25607 (N_25607,N_23141,N_20085);
nand U25608 (N_25608,N_20864,N_21170);
nor U25609 (N_25609,N_22561,N_24232);
nor U25610 (N_25610,N_24815,N_21795);
nor U25611 (N_25611,N_23482,N_20987);
nand U25612 (N_25612,N_24026,N_23589);
nor U25613 (N_25613,N_22721,N_20810);
nand U25614 (N_25614,N_22724,N_20913);
and U25615 (N_25615,N_20884,N_21579);
nor U25616 (N_25616,N_20855,N_23048);
nor U25617 (N_25617,N_21703,N_23813);
nor U25618 (N_25618,N_22592,N_20161);
and U25619 (N_25619,N_20188,N_22804);
xor U25620 (N_25620,N_24255,N_23534);
or U25621 (N_25621,N_24095,N_23762);
or U25622 (N_25622,N_20547,N_24525);
nand U25623 (N_25623,N_23579,N_24481);
nor U25624 (N_25624,N_22609,N_21886);
or U25625 (N_25625,N_24379,N_23288);
nor U25626 (N_25626,N_21377,N_23894);
nand U25627 (N_25627,N_22523,N_20019);
and U25628 (N_25628,N_23162,N_24015);
xnor U25629 (N_25629,N_21459,N_23339);
nand U25630 (N_25630,N_23548,N_20005);
or U25631 (N_25631,N_22372,N_22939);
nand U25632 (N_25632,N_22714,N_22535);
xor U25633 (N_25633,N_20179,N_21775);
and U25634 (N_25634,N_24770,N_21503);
nor U25635 (N_25635,N_20329,N_23780);
and U25636 (N_25636,N_22453,N_20276);
nand U25637 (N_25637,N_20891,N_22620);
nor U25638 (N_25638,N_20701,N_24260);
nor U25639 (N_25639,N_24577,N_24511);
xor U25640 (N_25640,N_24485,N_24857);
xor U25641 (N_25641,N_23745,N_20789);
xnor U25642 (N_25642,N_24643,N_20620);
xor U25643 (N_25643,N_22210,N_21953);
or U25644 (N_25644,N_22016,N_23388);
xnor U25645 (N_25645,N_21997,N_21706);
and U25646 (N_25646,N_23241,N_20078);
xnor U25647 (N_25647,N_20377,N_23841);
nand U25648 (N_25648,N_23058,N_23319);
or U25649 (N_25649,N_23909,N_22508);
or U25650 (N_25650,N_21212,N_24684);
nor U25651 (N_25651,N_24217,N_21742);
and U25652 (N_25652,N_21499,N_21540);
xnor U25653 (N_25653,N_20031,N_22055);
xnor U25654 (N_25654,N_24066,N_21128);
or U25655 (N_25655,N_20157,N_21069);
nor U25656 (N_25656,N_23228,N_20359);
and U25657 (N_25657,N_23859,N_23889);
nor U25658 (N_25658,N_20544,N_21359);
nor U25659 (N_25659,N_21218,N_24102);
and U25660 (N_25660,N_24231,N_23886);
nor U25661 (N_25661,N_21482,N_21698);
xnor U25662 (N_25662,N_21736,N_21318);
nor U25663 (N_25663,N_24132,N_21380);
nor U25664 (N_25664,N_20763,N_20667);
or U25665 (N_25665,N_24239,N_20748);
and U25666 (N_25666,N_21462,N_20537);
xor U25667 (N_25667,N_21604,N_21600);
xor U25668 (N_25668,N_20697,N_21711);
or U25669 (N_25669,N_21411,N_20112);
xnor U25670 (N_25670,N_24789,N_22622);
nor U25671 (N_25671,N_24432,N_24322);
xnor U25672 (N_25672,N_20275,N_22331);
or U25673 (N_25673,N_20244,N_22428);
xnor U25674 (N_25674,N_24775,N_21631);
nand U25675 (N_25675,N_23658,N_23702);
xor U25676 (N_25676,N_20984,N_22983);
nor U25677 (N_25677,N_24330,N_20224);
or U25678 (N_25678,N_21870,N_22121);
or U25679 (N_25679,N_20830,N_22625);
xnor U25680 (N_25680,N_24887,N_23002);
nor U25681 (N_25681,N_22855,N_20401);
nor U25682 (N_25682,N_24768,N_24056);
or U25683 (N_25683,N_21308,N_23998);
or U25684 (N_25684,N_20769,N_20865);
nand U25685 (N_25685,N_22659,N_24212);
nand U25686 (N_25686,N_24072,N_21244);
or U25687 (N_25687,N_24058,N_23775);
and U25688 (N_25688,N_20997,N_24038);
xnor U25689 (N_25689,N_20640,N_23360);
nand U25690 (N_25690,N_24098,N_20670);
xor U25691 (N_25691,N_21166,N_23910);
nand U25692 (N_25692,N_23310,N_23354);
nor U25693 (N_25693,N_21184,N_22553);
and U25694 (N_25694,N_22457,N_24402);
nor U25695 (N_25695,N_22175,N_22168);
xor U25696 (N_25696,N_20339,N_22501);
nand U25697 (N_25697,N_24622,N_23479);
and U25698 (N_25698,N_21700,N_20474);
nor U25699 (N_25699,N_21068,N_21029);
or U25700 (N_25700,N_22248,N_20892);
nand U25701 (N_25701,N_23194,N_20299);
and U25702 (N_25702,N_20454,N_24663);
nor U25703 (N_25703,N_20724,N_22980);
nor U25704 (N_25704,N_23040,N_22336);
xor U25705 (N_25705,N_21153,N_20263);
nor U25706 (N_25706,N_20347,N_23565);
and U25707 (N_25707,N_22596,N_24490);
nor U25708 (N_25708,N_20872,N_22567);
xor U25709 (N_25709,N_20915,N_20385);
nand U25710 (N_25710,N_21303,N_23112);
nand U25711 (N_25711,N_22705,N_24075);
xor U25712 (N_25712,N_20989,N_24029);
nor U25713 (N_25713,N_23713,N_22541);
xor U25714 (N_25714,N_20073,N_22759);
nor U25715 (N_25715,N_22265,N_21324);
nand U25716 (N_25716,N_24005,N_24797);
or U25717 (N_25717,N_23602,N_23255);
or U25718 (N_25718,N_22001,N_21624);
nor U25719 (N_25719,N_21330,N_20619);
xnor U25720 (N_25720,N_22626,N_21882);
nor U25721 (N_25721,N_20567,N_20521);
or U25722 (N_25722,N_22780,N_23304);
or U25723 (N_25723,N_20469,N_24660);
and U25724 (N_25724,N_22326,N_22111);
nand U25725 (N_25725,N_23539,N_22537);
xor U25726 (N_25726,N_24680,N_20902);
nand U25727 (N_25727,N_22695,N_21425);
and U25728 (N_25728,N_20979,N_22067);
xor U25729 (N_25729,N_24351,N_21307);
xnor U25730 (N_25730,N_20449,N_20602);
or U25731 (N_25731,N_21771,N_21983);
nand U25732 (N_25732,N_23173,N_20423);
nor U25733 (N_25733,N_22275,N_22613);
nor U25734 (N_25734,N_23824,N_22062);
nor U25735 (N_25735,N_24467,N_23914);
nor U25736 (N_25736,N_20156,N_23761);
nand U25737 (N_25737,N_23013,N_20654);
nor U25738 (N_25738,N_23575,N_21412);
and U25739 (N_25739,N_20187,N_23911);
or U25740 (N_25740,N_21850,N_23271);
and U25741 (N_25741,N_24848,N_20777);
or U25742 (N_25742,N_22112,N_23219);
and U25743 (N_25743,N_21893,N_20622);
or U25744 (N_25744,N_23396,N_23079);
nor U25745 (N_25745,N_20723,N_21040);
or U25746 (N_25746,N_20840,N_21661);
and U25747 (N_25747,N_24967,N_22084);
xor U25748 (N_25748,N_24727,N_23462);
nand U25749 (N_25749,N_21763,N_22462);
and U25750 (N_25750,N_20133,N_23527);
or U25751 (N_25751,N_24971,N_24527);
and U25752 (N_25752,N_21830,N_22822);
nor U25753 (N_25753,N_24415,N_21557);
and U25754 (N_25754,N_20933,N_21117);
nor U25755 (N_25755,N_23783,N_24653);
and U25756 (N_25756,N_20087,N_24078);
nor U25757 (N_25757,N_22610,N_22416);
and U25758 (N_25758,N_24565,N_23979);
nand U25759 (N_25759,N_21666,N_22198);
or U25760 (N_25760,N_21846,N_24036);
and U25761 (N_25761,N_20415,N_24898);
nor U25762 (N_25762,N_23672,N_20874);
nor U25763 (N_25763,N_23076,N_21858);
xor U25764 (N_25764,N_21672,N_22736);
and U25765 (N_25765,N_22036,N_21844);
and U25766 (N_25766,N_23018,N_22584);
or U25767 (N_25767,N_24896,N_21567);
or U25768 (N_25768,N_23325,N_21039);
nor U25769 (N_25769,N_23361,N_24954);
xnor U25770 (N_25770,N_24621,N_20239);
xor U25771 (N_25771,N_24689,N_22397);
xnor U25772 (N_25772,N_20962,N_22936);
nand U25773 (N_25773,N_24678,N_23742);
nand U25774 (N_25774,N_20369,N_21969);
nor U25775 (N_25775,N_22051,N_23081);
or U25776 (N_25776,N_22702,N_24131);
and U25777 (N_25777,N_22671,N_23967);
or U25778 (N_25778,N_21402,N_23927);
xnor U25779 (N_25779,N_22872,N_23386);
xnor U25780 (N_25780,N_21815,N_24073);
nor U25781 (N_25781,N_24893,N_24507);
xor U25782 (N_25782,N_24419,N_24781);
xor U25783 (N_25783,N_22954,N_23022);
xor U25784 (N_25784,N_23667,N_24905);
or U25785 (N_25785,N_23616,N_20594);
or U25786 (N_25786,N_21662,N_20028);
nand U25787 (N_25787,N_24850,N_23876);
and U25788 (N_25788,N_21996,N_22887);
nand U25789 (N_25789,N_23986,N_20695);
and U25790 (N_25790,N_24135,N_22222);
nor U25791 (N_25791,N_22276,N_24300);
xor U25792 (N_25792,N_20006,N_20253);
nor U25793 (N_25793,N_24809,N_24701);
or U25794 (N_25794,N_22641,N_20265);
nand U25795 (N_25795,N_20579,N_22949);
or U25796 (N_25796,N_23445,N_20461);
nor U25797 (N_25797,N_22953,N_20043);
nor U25798 (N_25798,N_22652,N_21607);
and U25799 (N_25799,N_20846,N_20878);
nand U25800 (N_25800,N_20869,N_23664);
nand U25801 (N_25801,N_24982,N_21108);
or U25802 (N_25802,N_21628,N_21230);
or U25803 (N_25803,N_22824,N_24192);
and U25804 (N_25804,N_22226,N_24278);
nor U25805 (N_25805,N_22337,N_21632);
nor U25806 (N_25806,N_22464,N_20222);
nor U25807 (N_25807,N_21252,N_21083);
or U25808 (N_25808,N_23648,N_20436);
and U25809 (N_25809,N_23877,N_22233);
and U25810 (N_25810,N_24690,N_23309);
or U25811 (N_25811,N_23152,N_21509);
xnor U25812 (N_25812,N_20233,N_23700);
and U25813 (N_25813,N_21059,N_23487);
xor U25814 (N_25814,N_20381,N_22920);
or U25815 (N_25815,N_23677,N_20727);
or U25816 (N_25816,N_20707,N_22794);
or U25817 (N_25817,N_24650,N_24437);
or U25818 (N_25818,N_24947,N_20792);
nor U25819 (N_25819,N_22161,N_20728);
nor U25820 (N_25820,N_20121,N_23133);
xnor U25821 (N_25821,N_24916,N_24017);
nand U25822 (N_25822,N_22725,N_23034);
and U25823 (N_25823,N_20280,N_20785);
or U25824 (N_25824,N_23266,N_20595);
or U25825 (N_25825,N_20077,N_21713);
nand U25826 (N_25826,N_24367,N_23292);
and U25827 (N_25827,N_21121,N_22528);
nor U25828 (N_25828,N_22818,N_22202);
or U25829 (N_25829,N_22805,N_23507);
xnor U25830 (N_25830,N_24697,N_23102);
nor U25831 (N_25831,N_21526,N_21616);
xor U25832 (N_25832,N_22740,N_24314);
xnor U25833 (N_25833,N_20214,N_23885);
xnor U25834 (N_25834,N_20711,N_23867);
xnor U25835 (N_25835,N_22137,N_24394);
nand U25836 (N_25836,N_23493,N_23852);
nand U25837 (N_25837,N_22933,N_24915);
or U25838 (N_25838,N_23515,N_23518);
xnor U25839 (N_25839,N_22757,N_22763);
nor U25840 (N_25840,N_20616,N_20733);
nand U25841 (N_25841,N_23265,N_20934);
and U25842 (N_25842,N_24097,N_22425);
nand U25843 (N_25843,N_24091,N_24128);
or U25844 (N_25844,N_23491,N_21779);
nor U25845 (N_25845,N_23156,N_23720);
nor U25846 (N_25846,N_20539,N_21350);
nor U25847 (N_25847,N_22856,N_22838);
or U25848 (N_25848,N_22194,N_21762);
or U25849 (N_25849,N_20102,N_22136);
xor U25850 (N_25850,N_24291,N_21625);
or U25851 (N_25851,N_22715,N_23233);
xor U25852 (N_25852,N_22992,N_24092);
nor U25853 (N_25853,N_21902,N_23970);
nand U25854 (N_25854,N_24465,N_20257);
nand U25855 (N_25855,N_22868,N_23330);
nand U25856 (N_25856,N_21416,N_23363);
nand U25857 (N_25857,N_20141,N_21954);
nand U25858 (N_25858,N_21018,N_24995);
or U25859 (N_25859,N_23371,N_22436);
xnor U25860 (N_25860,N_24981,N_22589);
or U25861 (N_25861,N_21623,N_24909);
xnor U25862 (N_25862,N_22531,N_23804);
or U25863 (N_25863,N_23807,N_24802);
nand U25864 (N_25864,N_20452,N_23763);
nand U25865 (N_25865,N_24628,N_21096);
nor U25866 (N_25866,N_22355,N_22304);
xnor U25867 (N_25867,N_24551,N_20463);
nor U25868 (N_25868,N_23631,N_20168);
xnor U25869 (N_25869,N_23696,N_24052);
nand U25870 (N_25870,N_21035,N_21475);
nor U25871 (N_25871,N_20196,N_22012);
and U25872 (N_25872,N_24927,N_21823);
xnor U25873 (N_25873,N_23994,N_22429);
nor U25874 (N_25874,N_21573,N_23709);
xnor U25875 (N_25875,N_20390,N_23545);
nand U25876 (N_25876,N_20706,N_22424);
and U25877 (N_25877,N_22076,N_22427);
xnor U25878 (N_25878,N_21294,N_22082);
and U25879 (N_25879,N_23687,N_20398);
and U25880 (N_25880,N_20348,N_24785);
or U25881 (N_25881,N_20269,N_20199);
or U25882 (N_25882,N_24615,N_22882);
nand U25883 (N_25883,N_24618,N_23450);
or U25884 (N_25884,N_24440,N_20278);
or U25885 (N_25885,N_20434,N_22743);
and U25886 (N_25886,N_20293,N_21939);
and U25887 (N_25887,N_20447,N_21580);
nor U25888 (N_25888,N_21131,N_22522);
nand U25889 (N_25889,N_22905,N_22853);
and U25890 (N_25890,N_22874,N_24968);
nor U25891 (N_25891,N_24788,N_20429);
xnor U25892 (N_25892,N_20643,N_20246);
or U25893 (N_25893,N_24752,N_22316);
or U25894 (N_25894,N_20556,N_21435);
xor U25895 (N_25895,N_22320,N_23244);
and U25896 (N_25896,N_21353,N_20453);
xnor U25897 (N_25897,N_22146,N_22302);
or U25898 (N_25898,N_23973,N_20281);
or U25899 (N_25899,N_24421,N_21712);
and U25900 (N_25900,N_20669,N_20897);
nor U25901 (N_25901,N_24027,N_24917);
xnor U25902 (N_25902,N_20799,N_21906);
xor U25903 (N_25903,N_24068,N_23305);
nor U25904 (N_25904,N_23817,N_23578);
and U25905 (N_25905,N_23786,N_20971);
nor U25906 (N_25906,N_22734,N_23513);
xor U25907 (N_25907,N_23607,N_21126);
nand U25908 (N_25908,N_23049,N_22065);
xor U25909 (N_25909,N_22545,N_20392);
xor U25910 (N_25910,N_24168,N_24501);
and U25911 (N_25911,N_23759,N_24759);
xor U25912 (N_25912,N_22926,N_22043);
xor U25913 (N_25913,N_21365,N_24529);
nor U25914 (N_25914,N_24587,N_20581);
nor U25915 (N_25915,N_22190,N_23604);
or U25916 (N_25916,N_21438,N_24865);
nand U25917 (N_25917,N_22739,N_24251);
and U25918 (N_25918,N_24209,N_22547);
nand U25919 (N_25919,N_21918,N_24979);
nor U25920 (N_25920,N_22367,N_24767);
nor U25921 (N_25921,N_24292,N_21351);
or U25922 (N_25922,N_20542,N_24118);
xnor U25923 (N_25923,N_21168,N_21276);
xnor U25924 (N_25924,N_22621,N_24393);
and U25925 (N_25925,N_23434,N_24669);
nand U25926 (N_25926,N_20599,N_24108);
and U25927 (N_25927,N_23847,N_24822);
xnor U25928 (N_25928,N_20876,N_20404);
nand U25929 (N_25929,N_21368,N_20856);
nor U25930 (N_25930,N_24557,N_24479);
xor U25931 (N_25931,N_20497,N_23375);
nor U25932 (N_25932,N_24627,N_23293);
xor U25933 (N_25933,N_22173,N_24742);
or U25934 (N_25934,N_21705,N_20736);
and U25935 (N_25935,N_23530,N_20839);
or U25936 (N_25936,N_23551,N_24176);
nand U25937 (N_25937,N_21977,N_23250);
or U25938 (N_25938,N_20258,N_21738);
and U25939 (N_25939,N_23531,N_20844);
or U25940 (N_25940,N_22581,N_20271);
nor U25941 (N_25941,N_23976,N_21968);
nor U25942 (N_25942,N_22134,N_22914);
nor U25943 (N_25943,N_24107,N_23996);
and U25944 (N_25944,N_23741,N_21681);
or U25945 (N_25945,N_24323,N_23171);
xor U25946 (N_25946,N_21938,N_23215);
and U25947 (N_25947,N_20021,N_24728);
or U25948 (N_25948,N_23059,N_24279);
and U25949 (N_25949,N_24651,N_20346);
xnor U25950 (N_25950,N_23420,N_24349);
and U25951 (N_25951,N_24164,N_22243);
xnor U25952 (N_25952,N_22268,N_23975);
xnor U25953 (N_25953,N_20973,N_21506);
xnor U25954 (N_25954,N_23005,N_23119);
or U25955 (N_25955,N_22557,N_21422);
nor U25956 (N_25956,N_22673,N_20139);
nand U25957 (N_25957,N_22353,N_24143);
and U25958 (N_25958,N_24475,N_24170);
and U25959 (N_25959,N_24272,N_20655);
nand U25960 (N_25960,N_22735,N_22488);
xor U25961 (N_25961,N_21563,N_22604);
or U25962 (N_25962,N_20290,N_22274);
nand U25963 (N_25963,N_21877,N_23822);
xnor U25964 (N_25964,N_20140,N_24214);
xor U25965 (N_25965,N_20017,N_22768);
xnor U25966 (N_25966,N_23947,N_24972);
nand U25967 (N_25967,N_24751,N_21679);
nand U25968 (N_25968,N_24700,N_24584);
xnor U25969 (N_25969,N_22486,N_21289);
and U25970 (N_25970,N_24310,N_20895);
xnor U25971 (N_25971,N_20383,N_23821);
xnor U25972 (N_25972,N_23499,N_22552);
nand U25973 (N_25973,N_24517,N_22564);
nand U25974 (N_25974,N_24155,N_22184);
and U25975 (N_25975,N_20917,N_20806);
or U25976 (N_25976,N_22354,N_22598);
and U25977 (N_25977,N_24082,N_24271);
nor U25978 (N_25978,N_21256,N_21702);
nand U25979 (N_25979,N_21328,N_24186);
nor U25980 (N_25980,N_23708,N_21768);
and U25981 (N_25981,N_23503,N_23712);
or U25982 (N_25982,N_21743,N_22929);
and U25983 (N_25983,N_24610,N_23802);
and U25984 (N_25984,N_21819,N_21824);
xnor U25985 (N_25985,N_23065,N_24037);
nor U25986 (N_25986,N_20775,N_23591);
nand U25987 (N_25987,N_21678,N_20013);
and U25988 (N_25988,N_22023,N_24236);
or U25989 (N_25989,N_20191,N_21691);
nor U25990 (N_25990,N_24213,N_21562);
or U25991 (N_25991,N_22618,N_22058);
and U25992 (N_25992,N_20135,N_23989);
and U25993 (N_25993,N_21999,N_23043);
or U25994 (N_25994,N_22380,N_22761);
xnor U25995 (N_25995,N_21404,N_23766);
xor U25996 (N_25996,N_22754,N_22704);
xor U25997 (N_25997,N_21956,N_21708);
nand U25998 (N_25998,N_22199,N_21804);
and U25999 (N_25999,N_22779,N_23722);
nor U26000 (N_26000,N_20939,N_21430);
nor U26001 (N_26001,N_23860,N_22952);
nor U26002 (N_26002,N_24473,N_23898);
nand U26003 (N_26003,N_24307,N_20908);
and U26004 (N_26004,N_20887,N_23449);
and U26005 (N_26005,N_24870,N_24765);
and U26006 (N_26006,N_23871,N_20957);
and U26007 (N_26007,N_23796,N_20467);
nand U26008 (N_26008,N_20007,N_22150);
or U26009 (N_26009,N_24806,N_22646);
nor U26010 (N_26010,N_24124,N_21647);
or U26011 (N_26011,N_21590,N_23599);
xnor U26012 (N_26012,N_20136,N_21055);
xnor U26013 (N_26013,N_24620,N_23423);
or U26014 (N_26014,N_20514,N_24975);
or U26015 (N_26015,N_24958,N_21927);
nand U26016 (N_26016,N_24163,N_22638);
nand U26017 (N_26017,N_22961,N_20550);
nand U26018 (N_26018,N_24619,N_20378);
and U26019 (N_26019,N_24753,N_23960);
nor U26020 (N_26020,N_21936,N_23089);
nand U26021 (N_26021,N_24235,N_20746);
and U26022 (N_26022,N_21497,N_21050);
and U26023 (N_26023,N_21031,N_21568);
xor U26024 (N_26024,N_24134,N_22758);
xnor U26025 (N_26025,N_23209,N_21064);
xnor U26026 (N_26026,N_22327,N_20475);
and U26027 (N_26027,N_22050,N_20268);
or U26028 (N_26028,N_21481,N_22674);
and U26029 (N_26029,N_22841,N_20692);
nand U26030 (N_26030,N_22096,N_20002);
and U26031 (N_26031,N_24244,N_24407);
and U26032 (N_26032,N_23465,N_22477);
and U26033 (N_26033,N_23214,N_24365);
nor U26034 (N_26034,N_24354,N_22026);
nand U26035 (N_26035,N_22678,N_24090);
and U26036 (N_26036,N_20768,N_24268);
and U26037 (N_26037,N_21642,N_24648);
nor U26038 (N_26038,N_23506,N_20721);
xnor U26039 (N_26039,N_21589,N_23011);
nor U26040 (N_26040,N_23185,N_21950);
and U26041 (N_26041,N_23842,N_20334);
and U26042 (N_26042,N_20486,N_22562);
nor U26043 (N_26043,N_24051,N_23717);
nand U26044 (N_26044,N_20444,N_23334);
nor U26045 (N_26045,N_23733,N_21776);
or U26046 (N_26046,N_20950,N_22100);
nand U26047 (N_26047,N_24855,N_23118);
nand U26048 (N_26048,N_22412,N_21871);
nand U26049 (N_26049,N_24799,N_23208);
xor U26050 (N_26050,N_23541,N_22560);
nor U26051 (N_26051,N_22682,N_21685);
nand U26052 (N_26052,N_21285,N_24319);
or U26053 (N_26053,N_22297,N_23084);
and U26054 (N_26054,N_20225,N_21638);
xnor U26055 (N_26055,N_21154,N_24646);
nor U26056 (N_26056,N_20759,N_23995);
or U26057 (N_26057,N_24448,N_23341);
xor U26058 (N_26058,N_24408,N_21063);
and U26059 (N_26059,N_22532,N_22075);
nor U26060 (N_26060,N_24403,N_21960);
nand U26061 (N_26061,N_22775,N_22677);
nor U26062 (N_26062,N_20576,N_21118);
nand U26063 (N_26063,N_20217,N_23374);
xnor U26064 (N_26064,N_20825,N_24749);
xnor U26065 (N_26065,N_21492,N_24399);
and U26066 (N_26066,N_24445,N_23461);
and U26067 (N_26067,N_22964,N_22894);
and U26068 (N_26068,N_24901,N_23856);
or U26069 (N_26069,N_21439,N_21973);
and U26070 (N_26070,N_21965,N_22821);
or U26071 (N_26071,N_22282,N_24327);
and U26072 (N_26072,N_21578,N_23095);
nor U26073 (N_26073,N_22711,N_21928);
or U26074 (N_26074,N_22975,N_20337);
and U26075 (N_26075,N_24463,N_20610);
or U26076 (N_26076,N_20355,N_20888);
and U26077 (N_26077,N_20694,N_20353);
or U26078 (N_26078,N_24583,N_24943);
nand U26079 (N_26079,N_24649,N_23032);
nor U26080 (N_26080,N_21316,N_22154);
xnor U26081 (N_26081,N_24474,N_21507);
nand U26082 (N_26082,N_21831,N_20256);
and U26083 (N_26083,N_24136,N_23862);
nand U26084 (N_26084,N_20298,N_24849);
xnor U26085 (N_26085,N_21376,N_21658);
and U26086 (N_26086,N_20782,N_21923);
nor U26087 (N_26087,N_20804,N_22498);
or U26088 (N_26088,N_20534,N_22487);
nand U26089 (N_26089,N_21610,N_24945);
nand U26090 (N_26090,N_20666,N_22879);
nand U26091 (N_26091,N_21397,N_24002);
or U26092 (N_26092,N_24342,N_20920);
nor U26093 (N_26093,N_22546,N_20904);
nor U26094 (N_26094,N_22591,N_20238);
nand U26095 (N_26095,N_22373,N_24368);
nor U26096 (N_26096,N_21862,N_21467);
xor U26097 (N_26097,N_21752,N_24531);
or U26098 (N_26098,N_20958,N_22748);
nand U26099 (N_26099,N_20480,N_23381);
nor U26100 (N_26100,N_20201,N_22578);
or U26101 (N_26101,N_23398,N_22993);
xnor U26102 (N_26102,N_23351,N_23105);
nand U26103 (N_26103,N_24595,N_21149);
xnor U26104 (N_26104,N_22351,N_24218);
nand U26105 (N_26105,N_21151,N_23315);
or U26106 (N_26106,N_23401,N_23108);
and U26107 (N_26107,N_23444,N_24053);
nand U26108 (N_26108,N_22284,N_20629);
nand U26109 (N_26109,N_22577,N_24290);
and U26110 (N_26110,N_21777,N_21784);
or U26111 (N_26111,N_23533,N_22130);
nand U26112 (N_26112,N_20797,N_20270);
nand U26113 (N_26113,N_24497,N_24537);
and U26114 (N_26114,N_24216,N_23828);
and U26115 (N_26115,N_22418,N_23158);
nor U26116 (N_26116,N_21410,N_22515);
xor U26117 (N_26117,N_20924,N_24957);
and U26118 (N_26118,N_23728,N_22913);
xnor U26119 (N_26119,N_23448,N_21934);
xnor U26120 (N_26120,N_24878,N_21449);
and U26121 (N_26121,N_23469,N_21123);
nor U26122 (N_26122,N_24871,N_21061);
nor U26123 (N_26123,N_20313,N_24900);
nand U26124 (N_26124,N_21320,N_22717);
xor U26125 (N_26125,N_22635,N_22943);
nand U26126 (N_26126,N_22215,N_20153);
or U26127 (N_26127,N_20389,N_23818);
nor U26128 (N_26128,N_21911,N_23247);
or U26129 (N_26129,N_21221,N_21571);
or U26130 (N_26130,N_21856,N_21723);
xor U26131 (N_26131,N_22898,N_22957);
and U26132 (N_26132,N_22066,N_21312);
or U26133 (N_26133,N_20660,N_20715);
and U26134 (N_26134,N_24616,N_21640);
nor U26135 (N_26135,N_22946,N_20776);
or U26136 (N_26136,N_20584,N_22542);
xnor U26137 (N_26137,N_21792,N_24662);
xor U26138 (N_26138,N_23537,N_24157);
xor U26139 (N_26139,N_24614,N_22484);
xnor U26140 (N_26140,N_20491,N_20663);
xor U26141 (N_26141,N_22234,N_24028);
or U26142 (N_26142,N_20705,N_21260);
and U26143 (N_26143,N_21140,N_20995);
nand U26144 (N_26144,N_20319,N_24540);
or U26145 (N_26145,N_21395,N_22662);
xor U26146 (N_26146,N_21183,N_20255);
and U26147 (N_26147,N_20195,N_24658);
nand U26148 (N_26148,N_22346,N_22390);
or U26149 (N_26149,N_24324,N_21305);
or U26150 (N_26150,N_22808,N_20045);
or U26151 (N_26151,N_21232,N_21998);
xnor U26152 (N_26152,N_20702,N_22848);
nand U26153 (N_26153,N_22097,N_20662);
nand U26154 (N_26154,N_20653,N_22511);
and U26155 (N_26155,N_21310,N_22074);
and U26156 (N_26156,N_24335,N_23794);
xnor U26157 (N_26157,N_24190,N_23825);
nand U26158 (N_26158,N_23486,N_23612);
nor U26159 (N_26159,N_20272,N_23992);
or U26160 (N_26160,N_22221,N_22967);
xor U26161 (N_26161,N_23442,N_21652);
nand U26162 (N_26162,N_24617,N_22420);
and U26163 (N_26163,N_22741,N_22524);
nor U26164 (N_26164,N_23812,N_22590);
nand U26165 (N_26165,N_22514,N_22345);
and U26166 (N_26166,N_24270,N_24748);
nand U26167 (N_26167,N_22843,N_21331);
and U26168 (N_26168,N_24552,N_21406);
xnor U26169 (N_26169,N_20312,N_20476);
and U26170 (N_26170,N_20948,N_22504);
or U26171 (N_26171,N_20691,N_21176);
or U26172 (N_26172,N_22685,N_24306);
or U26173 (N_26173,N_23064,N_20675);
xnor U26174 (N_26174,N_22830,N_22434);
and U26175 (N_26175,N_24178,N_20471);
nor U26176 (N_26176,N_23777,N_22045);
nand U26177 (N_26177,N_20075,N_21894);
and U26178 (N_26178,N_21521,N_22463);
xor U26179 (N_26179,N_24181,N_20442);
nand U26180 (N_26180,N_24423,N_20211);
xnor U26181 (N_26181,N_21009,N_24994);
or U26182 (N_26182,N_21348,N_23920);
nor U26183 (N_26183,N_22393,N_21207);
nand U26184 (N_26184,N_24969,N_22408);
and U26185 (N_26185,N_24435,N_20315);
nor U26186 (N_26186,N_20696,N_20873);
xnor U26187 (N_26187,N_21124,N_22668);
xnor U26188 (N_26188,N_23411,N_23394);
nor U26189 (N_26189,N_24113,N_21548);
and U26190 (N_26190,N_22476,N_22764);
nor U26191 (N_26191,N_24311,N_22895);
and U26192 (N_26192,N_22242,N_24762);
or U26193 (N_26193,N_20745,N_22782);
or U26194 (N_26194,N_21554,N_20795);
and U26195 (N_26195,N_24911,N_24077);
and U26196 (N_26196,N_20982,N_23063);
and U26197 (N_26197,N_20862,N_23650);
or U26198 (N_26198,N_24877,N_24441);
or U26199 (N_26199,N_20324,N_24161);
or U26200 (N_26200,N_21863,N_24418);
nor U26201 (N_26201,N_21122,N_22521);
nand U26202 (N_26202,N_24035,N_24338);
or U26203 (N_26203,N_24590,N_20487);
nor U26204 (N_26204,N_21816,N_24683);
and U26205 (N_26205,N_21322,N_21137);
nor U26206 (N_26206,N_21536,N_22529);
xor U26207 (N_26207,N_21574,N_21220);
nor U26208 (N_26208,N_24734,N_20717);
nor U26209 (N_26209,N_23686,N_22403);
xnor U26210 (N_26210,N_24147,N_20183);
xnor U26211 (N_26211,N_22612,N_22506);
xnor U26212 (N_26212,N_23180,N_22907);
xnor U26213 (N_26213,N_22458,N_24468);
or U26214 (N_26214,N_20956,N_20282);
xnor U26215 (N_26215,N_21388,N_20034);
nor U26216 (N_26216,N_24992,N_20536);
and U26217 (N_26217,N_23675,N_24115);
or U26218 (N_26218,N_24361,N_24301);
nand U26219 (N_26219,N_20322,N_21793);
or U26220 (N_26220,N_24801,N_24358);
nor U26221 (N_26221,N_23336,N_20418);
xor U26222 (N_26222,N_22213,N_22359);
nor U26223 (N_26223,N_21657,N_20949);
or U26224 (N_26224,N_23901,N_24902);
xnor U26225 (N_26225,N_20849,N_22139);
nor U26226 (N_26226,N_23298,N_20286);
xnor U26227 (N_26227,N_20247,N_20834);
xor U26228 (N_26228,N_20350,N_24145);
xnor U26229 (N_26229,N_20052,N_20115);
and U26230 (N_26230,N_24357,N_23281);
and U26231 (N_26231,N_22586,N_21525);
and U26232 (N_26232,N_21321,N_24344);
xnor U26233 (N_26233,N_24694,N_20163);
nand U26234 (N_26234,N_21403,N_22469);
or U26235 (N_26235,N_20601,N_21356);
or U26236 (N_26236,N_22611,N_22795);
or U26237 (N_26237,N_20076,N_23803);
or U26238 (N_26238,N_24355,N_23610);
nand U26239 (N_26239,N_24831,N_20303);
and U26240 (N_26240,N_21860,N_20880);
and U26241 (N_26241,N_22296,N_24229);
nor U26242 (N_26242,N_24601,N_24946);
nand U26243 (N_26243,N_24861,N_21687);
nand U26244 (N_26244,N_22305,N_22516);
and U26245 (N_26245,N_22605,N_22694);
xnor U26246 (N_26246,N_22996,N_22987);
nand U26247 (N_26247,N_22229,N_24573);
nor U26248 (N_26248,N_24062,N_21139);
nand U26249 (N_26249,N_21651,N_21209);
nand U26250 (N_26250,N_20288,N_20061);
nand U26251 (N_26251,N_24578,N_22447);
or U26252 (N_26252,N_21336,N_20177);
nor U26253 (N_26253,N_24200,N_24656);
xor U26254 (N_26254,N_24277,N_21288);
nand U26255 (N_26255,N_24506,N_21534);
nand U26256 (N_26256,N_21614,N_22863);
and U26257 (N_26257,N_21821,N_23230);
or U26258 (N_26258,N_21384,N_24382);
or U26259 (N_26259,N_23416,N_22505);
or U26260 (N_26260,N_24825,N_20889);
or U26261 (N_26261,N_20375,N_20885);
and U26262 (N_26262,N_23368,N_24449);
and U26263 (N_26263,N_24872,N_23355);
nand U26264 (N_26264,N_23767,N_23850);
or U26265 (N_26265,N_24112,N_21883);
xor U26266 (N_26266,N_23707,N_23395);
xnor U26267 (N_26267,N_21915,N_20050);
xor U26268 (N_26268,N_20096,N_20374);
nand U26269 (N_26269,N_21755,N_21383);
and U26270 (N_26270,N_21488,N_23116);
or U26271 (N_26271,N_23087,N_20838);
xnor U26272 (N_26272,N_20356,N_23564);
xnor U26273 (N_26273,N_22636,N_23039);
and U26274 (N_26274,N_24842,N_24819);
nor U26275 (N_26275,N_21644,N_24744);
and U26276 (N_26276,N_22574,N_21453);
or U26277 (N_26277,N_23077,N_21066);
nor U26278 (N_26278,N_20221,N_22565);
or U26279 (N_26279,N_21629,N_24100);
nor U26280 (N_26280,N_21992,N_21796);
nor U26281 (N_26281,N_23036,N_23679);
or U26282 (N_26282,N_22261,N_23149);
or U26283 (N_26283,N_24757,N_20684);
nand U26284 (N_26284,N_22749,N_24006);
or U26285 (N_26285,N_23923,N_21501);
nand U26286 (N_26286,N_24659,N_22241);
xnor U26287 (N_26287,N_22655,N_21790);
xnor U26288 (N_26288,N_22244,N_22669);
nand U26289 (N_26289,N_22466,N_22285);
nand U26290 (N_26290,N_24304,N_23868);
xor U26291 (N_26291,N_23342,N_24908);
and U26292 (N_26292,N_20756,N_20833);
xor U26293 (N_26293,N_23550,N_20909);
nor U26294 (N_26294,N_24826,N_21275);
nand U26295 (N_26295,N_21553,N_23528);
and U26296 (N_26296,N_20614,N_22680);
or U26297 (N_26297,N_20990,N_24763);
xor U26298 (N_26298,N_23492,N_23044);
xnor U26299 (N_26299,N_22981,N_24990);
or U26300 (N_26300,N_20976,N_24096);
nand U26301 (N_26301,N_20766,N_22395);
or U26302 (N_26302,N_23748,N_22090);
and U26303 (N_26303,N_22382,N_23736);
nor U26304 (N_26304,N_22778,N_22003);
and U26305 (N_26305,N_20277,N_24220);
nand U26306 (N_26306,N_22614,N_22087);
and U26307 (N_26307,N_20821,N_21972);
and U26308 (N_26308,N_24847,N_21845);
xnor U26309 (N_26309,N_21473,N_24706);
or U26310 (N_26310,N_20455,N_21203);
nand U26311 (N_26311,N_24835,N_22245);
or U26312 (N_26312,N_23922,N_24392);
nor U26313 (N_26313,N_22906,N_23651);
nand U26314 (N_26314,N_21409,N_21606);
or U26315 (N_26315,N_23621,N_21287);
nand U26316 (N_26316,N_20234,N_23620);
nor U26317 (N_26317,N_20533,N_24505);
nor U26318 (N_26318,N_22149,N_22349);
nor U26319 (N_26319,N_20907,N_21229);
and U26320 (N_26320,N_23207,N_20700);
nor U26321 (N_26321,N_23980,N_21716);
xnor U26322 (N_26322,N_22021,N_22814);
nor U26323 (N_26323,N_20927,N_20488);
and U26324 (N_26324,N_21617,N_21865);
xnor U26325 (N_26325,N_21188,N_22891);
or U26326 (N_26326,N_22860,N_22172);
xor U26327 (N_26327,N_20344,N_21937);
or U26328 (N_26328,N_23678,N_24513);
xor U26329 (N_26329,N_24962,N_24899);
xnor U26330 (N_26330,N_21735,N_24564);
nor U26331 (N_26331,N_22193,N_23012);
or U26332 (N_26332,N_24816,N_23276);
or U26333 (N_26333,N_20848,N_22404);
or U26334 (N_26334,N_20064,N_22448);
and U26335 (N_26335,N_23756,N_23313);
and U26336 (N_26336,N_20679,N_21962);
nand U26337 (N_26337,N_21690,N_22986);
xor U26338 (N_26338,N_22334,N_21159);
nor U26339 (N_26339,N_24150,N_23464);
nand U26340 (N_26340,N_22730,N_20376);
or U26341 (N_26341,N_23323,N_20033);
xor U26342 (N_26342,N_24798,N_22799);
or U26343 (N_26343,N_23790,N_24716);
and U26344 (N_26344,N_21400,N_23714);
and U26345 (N_26345,N_21237,N_24137);
and U26346 (N_26346,N_21669,N_22033);
nand U26347 (N_26347,N_24837,N_22249);
or U26348 (N_26348,N_23295,N_21485);
nand U26349 (N_26349,N_21265,N_20794);
nor U26350 (N_26350,N_21302,N_20931);
nand U26351 (N_26351,N_22046,N_22922);
nand U26352 (N_26352,N_22422,N_20851);
and U26353 (N_26353,N_22745,N_21611);
or U26354 (N_26354,N_21474,N_21067);
nand U26355 (N_26355,N_23597,N_20181);
and U26356 (N_26356,N_21165,N_23484);
nor U26357 (N_26357,N_23443,N_24520);
nor U26358 (N_26358,N_24611,N_21357);
nor U26359 (N_26359,N_21355,N_21107);
nor U26360 (N_26360,N_23344,N_24593);
nand U26361 (N_26361,N_23222,N_20553);
nor U26362 (N_26362,N_20621,N_20495);
xnor U26363 (N_26363,N_21508,N_22170);
xor U26364 (N_26364,N_21608,N_24105);
xor U26365 (N_26365,N_20870,N_24939);
nand U26366 (N_26366,N_21158,N_24199);
nand U26367 (N_26367,N_22280,N_20859);
and U26368 (N_26368,N_20673,N_23307);
nor U26369 (N_26369,N_22138,N_22157);
nor U26370 (N_26370,N_22083,N_23585);
nor U26371 (N_26371,N_20803,N_21564);
or U26372 (N_26372,N_23624,N_24152);
or U26373 (N_26373,N_21949,N_24321);
nand U26374 (N_26374,N_22238,N_24198);
or U26375 (N_26375,N_24746,N_22414);
or U26376 (N_26376,N_21734,N_23120);
nand U26377 (N_26377,N_21921,N_23516);
nor U26378 (N_26378,N_20545,N_23452);
nor U26379 (N_26379,N_24503,N_22828);
xnor U26380 (N_26380,N_21292,N_22979);
or U26381 (N_26381,N_23811,N_21053);
and U26382 (N_26382,N_20575,N_21450);
nor U26383 (N_26383,N_23958,N_20185);
and U26384 (N_26384,N_21582,N_22271);
xor U26385 (N_26385,N_22430,N_22204);
and U26386 (N_26386,N_20420,N_20638);
xor U26387 (N_26387,N_23261,N_24772);
xor U26388 (N_26388,N_23874,N_20193);
xor U26389 (N_26389,N_20237,N_22047);
xor U26390 (N_26390,N_21466,N_21144);
nor U26391 (N_26391,N_20965,N_22803);
and U26392 (N_26392,N_21297,N_20554);
or U26393 (N_26393,N_20500,N_22318);
nor U26394 (N_26394,N_22588,N_21446);
nand U26395 (N_26395,N_22344,N_21739);
xor U26396 (N_26396,N_21211,N_24443);
xor U26397 (N_26397,N_22135,N_20559);
nand U26398 (N_26398,N_22379,N_23769);
nor U26399 (N_26399,N_23007,N_21465);
or U26400 (N_26400,N_21803,N_22700);
and U26401 (N_26401,N_20095,N_24977);
xnor U26402 (N_26402,N_20817,N_23552);
nand U26403 (N_26403,N_21189,N_20336);
nand U26404 (N_26404,N_24455,N_20481);
xnor U26405 (N_26405,N_24362,N_23269);
xnor U26406 (N_26406,N_20947,N_23488);
nor U26407 (N_26407,N_21358,N_21704);
nand U26408 (N_26408,N_22140,N_20593);
xor U26409 (N_26409,N_23327,N_21745);
nor U26410 (N_26410,N_22117,N_23466);
nor U26411 (N_26411,N_22053,N_20252);
and U26412 (N_26412,N_23930,N_23170);
and U26413 (N_26413,N_22314,N_22909);
or U26414 (N_26414,N_21733,N_24360);
nand U26415 (N_26415,N_24079,N_20685);
or U26416 (N_26416,N_23346,N_21436);
nor U26417 (N_26417,N_24308,N_22394);
or U26418 (N_26418,N_22056,N_21249);
xnor U26419 (N_26419,N_20946,N_23267);
and U26420 (N_26420,N_20974,N_23508);
nor U26421 (N_26421,N_22976,N_21797);
xnor U26422 (N_26422,N_20430,N_20304);
xor U26423 (N_26423,N_24259,N_23446);
nand U26424 (N_26424,N_24862,N_22890);
nor U26425 (N_26425,N_23831,N_20042);
and U26426 (N_26426,N_21857,N_24297);
xnor U26427 (N_26427,N_20816,N_22767);
xor U26428 (N_26428,N_24867,N_24094);
nand U26429 (N_26429,N_22088,N_21471);
or U26430 (N_26430,N_22307,N_24755);
or U26431 (N_26431,N_22309,N_23187);
xnor U26432 (N_26432,N_21798,N_24305);
xor U26433 (N_26433,N_22544,N_21304);
xor U26434 (N_26434,N_22865,N_24536);
xnor U26435 (N_26435,N_20615,N_24681);
nor U26436 (N_26436,N_24454,N_20367);
or U26437 (N_26437,N_22160,N_22449);
and U26438 (N_26438,N_21551,N_24547);
nor U26439 (N_26439,N_24830,N_21787);
and U26440 (N_26440,N_23056,N_24984);
nand U26441 (N_26441,N_23455,N_22361);
and U26442 (N_26442,N_21688,N_23964);
xor U26443 (N_26443,N_22712,N_22991);
nand U26444 (N_26444,N_21940,N_23365);
or U26445 (N_26445,N_23836,N_20358);
nor U26446 (N_26446,N_21765,N_21442);
xnor U26447 (N_26447,N_23887,N_24812);
or U26448 (N_26448,N_20770,N_23561);
and U26449 (N_26449,N_21500,N_22356);
nor U26450 (N_26450,N_24811,N_20709);
nor U26451 (N_26451,N_22342,N_21558);
or U26452 (N_26452,N_22024,N_24366);
nand U26453 (N_26453,N_20200,N_20901);
xnor U26454 (N_26454,N_24884,N_21964);
and U26455 (N_26455,N_20088,N_21751);
or U26456 (N_26456,N_21037,N_24221);
xor U26457 (N_26457,N_23546,N_24249);
or U26458 (N_26458,N_22873,N_23016);
xor U26459 (N_26459,N_22958,N_22875);
or U26460 (N_26460,N_24582,N_20435);
xnor U26461 (N_26461,N_24287,N_23706);
or U26462 (N_26462,N_21491,N_22148);
nor U26463 (N_26463,N_21065,N_21654);
or U26464 (N_26464,N_20648,N_24484);
nand U26465 (N_26465,N_21726,N_20165);
nor U26466 (N_26466,N_23969,N_23536);
and U26467 (N_26467,N_21586,N_24515);
nand U26468 (N_26468,N_21208,N_24195);
and U26469 (N_26469,N_24545,N_23082);
and U26470 (N_26470,N_23030,N_21456);
nand U26471 (N_26471,N_20279,N_20357);
or U26472 (N_26472,N_22321,N_20586);
nand U26473 (N_26473,N_23924,N_20118);
and U26474 (N_26474,N_20591,N_22009);
and U26475 (N_26475,N_21744,N_21428);
nand U26476 (N_26476,N_24696,N_21660);
and U26477 (N_26477,N_21030,N_20788);
and U26478 (N_26478,N_22580,N_24745);
xor U26479 (N_26479,N_24562,N_21874);
nor U26480 (N_26480,N_20790,N_20413);
nand U26481 (N_26481,N_22164,N_20066);
and U26482 (N_26482,N_24941,N_20128);
and U26483 (N_26483,N_21419,N_24856);
nor U26484 (N_26484,N_22550,N_21650);
xnor U26485 (N_26485,N_21399,N_24541);
or U26486 (N_26486,N_23124,N_24654);
and U26487 (N_26487,N_20342,N_24891);
nor U26488 (N_26488,N_22340,N_21837);
or U26489 (N_26489,N_22236,N_22459);
or U26490 (N_26490,N_24936,N_23052);
nand U26491 (N_26491,N_24223,N_20038);
nand U26492 (N_26492,N_21070,N_24483);
nor U26493 (N_26493,N_20127,N_22572);
and U26494 (N_26494,N_21757,N_22399);
nor U26495 (N_26495,N_23038,N_21155);
or U26496 (N_26496,N_20528,N_20297);
nand U26497 (N_26497,N_20251,N_24389);
nand U26498 (N_26498,N_20664,N_22889);
xnor U26499 (N_26499,N_20345,N_21904);
nand U26500 (N_26500,N_21375,N_20600);
nor U26501 (N_26501,N_23595,N_20626);
nor U26502 (N_26502,N_20668,N_22900);
or U26503 (N_26503,N_24569,N_24555);
nor U26504 (N_26504,N_21225,N_23543);
nor U26505 (N_26505,N_22409,N_20069);
nor U26506 (N_26506,N_24636,N_23197);
and U26507 (N_26507,N_23403,N_22908);
and U26508 (N_26508,N_21114,N_20117);
nand U26509 (N_26509,N_21054,N_20628);
nor U26510 (N_26510,N_21003,N_20372);
xor U26511 (N_26511,N_23279,N_22990);
and U26512 (N_26512,N_21794,N_23306);
xor U26513 (N_26513,N_24832,N_24886);
and U26514 (N_26514,N_23220,N_22472);
xor U26515 (N_26515,N_21335,N_23949);
and U26516 (N_26516,N_22034,N_21269);
and U26517 (N_26517,N_21301,N_21668);
nor U26518 (N_26518,N_24652,N_24959);
xnor U26519 (N_26519,N_20906,N_21363);
nor U26520 (N_26520,N_22398,N_24922);
and U26521 (N_26521,N_21300,N_24289);
and U26522 (N_26522,N_20301,N_21113);
xor U26523 (N_26523,N_24089,N_20734);
and U26524 (N_26524,N_22665,N_21683);
nor U26525 (N_26525,N_24242,N_24187);
or U26526 (N_26526,N_24952,N_20520);
nand U26527 (N_26527,N_23430,N_24428);
nand U26528 (N_26528,N_23068,N_20067);
nor U26529 (N_26529,N_24284,N_22608);
nand U26530 (N_26530,N_22018,N_21214);
xor U26531 (N_26531,N_21258,N_21347);
and U26532 (N_26532,N_20035,N_23908);
or U26533 (N_26533,N_21945,N_22997);
nor U26534 (N_26534,N_23773,N_20996);
nor U26535 (N_26535,N_23685,N_24149);
nand U26536 (N_26536,N_20417,N_21017);
nor U26537 (N_26537,N_22840,N_21062);
nand U26538 (N_26538,N_23204,N_22388);
nand U26539 (N_26539,N_20094,N_23904);
or U26540 (N_26540,N_20925,N_24818);
and U26541 (N_26541,N_23047,N_20368);
nor U26542 (N_26542,N_21576,N_22810);
nand U26543 (N_26543,N_23753,N_21544);
and U26544 (N_26544,N_24298,N_23946);
xnor U26545 (N_26545,N_20262,N_23662);
nor U26546 (N_26546,N_23441,N_21626);
nand U26547 (N_26547,N_20053,N_23760);
nand U26548 (N_26548,N_23093,N_23522);
and U26549 (N_26549,N_23805,N_24240);
nor U26550 (N_26550,N_22207,N_23053);
nand U26551 (N_26551,N_24874,N_20432);
xor U26552 (N_26552,N_20857,N_24671);
xor U26553 (N_26553,N_23201,N_22670);
and U26554 (N_26554,N_22956,N_22481);
xnor U26555 (N_26555,N_23835,N_20798);
xor U26556 (N_26556,N_24532,N_23432);
nand U26557 (N_26557,N_23665,N_23962);
or U26558 (N_26558,N_20171,N_21032);
nand U26559 (N_26559,N_23628,N_21748);
and U26560 (N_26560,N_21756,N_21202);
nor U26561 (N_26561,N_21975,N_24162);
nor U26562 (N_26562,N_22441,N_21674);
or U26563 (N_26563,N_23747,N_23581);
nand U26564 (N_26564,N_21440,N_24747);
or U26565 (N_26565,N_22027,N_22127);
and U26566 (N_26566,N_24345,N_21730);
nor U26567 (N_26567,N_21091,N_24067);
and U26568 (N_26568,N_22384,N_24604);
xor U26569 (N_26569,N_20771,N_23296);
nand U26570 (N_26570,N_20472,N_22752);
xnor U26571 (N_26571,N_22497,N_23725);
xnor U26572 (N_26572,N_22266,N_24633);
nand U26573 (N_26573,N_24274,N_20220);
xnor U26574 (N_26574,N_20267,N_24840);
or U26575 (N_26575,N_23412,N_20232);
and U26576 (N_26576,N_20970,N_20180);
nand U26577 (N_26577,N_24817,N_23873);
and U26578 (N_26578,N_24637,N_21006);
xor U26579 (N_26579,N_23916,N_24685);
nor U26580 (N_26580,N_20450,N_20460);
nor U26581 (N_26581,N_20658,N_24792);
and U26582 (N_26582,N_24412,N_23349);
and U26583 (N_26583,N_20589,N_24059);
or U26584 (N_26584,N_21393,N_21038);
nand U26585 (N_26585,N_22994,N_21869);
nand U26586 (N_26586,N_24160,N_20824);
xnor U26587 (N_26587,N_23701,N_22623);
and U26588 (N_26588,N_20741,N_21109);
or U26589 (N_26589,N_21946,N_24609);
and U26590 (N_26590,N_21194,N_20583);
nand U26591 (N_26591,N_22880,N_21283);
xnor U26592 (N_26592,N_21433,N_24868);
nand U26593 (N_26593,N_21986,N_23400);
nor U26594 (N_26594,N_22108,N_22664);
and U26595 (N_26595,N_22079,N_20341);
and U26596 (N_26596,N_21317,N_24814);
or U26597 (N_26597,N_20228,N_24317);
and U26598 (N_26598,N_20894,N_20223);
nand U26599 (N_26599,N_20103,N_23711);
or U26600 (N_26600,N_24495,N_23397);
nor U26601 (N_26601,N_22788,N_20818);
or U26602 (N_26602,N_20433,N_23223);
or U26603 (N_26603,N_21367,N_24326);
or U26604 (N_26604,N_20003,N_22663);
and U26605 (N_26605,N_22781,N_23322);
nor U26606 (N_26606,N_21476,N_22847);
nand U26607 (N_26607,N_24009,N_20835);
or U26608 (N_26608,N_20722,N_23132);
and U26609 (N_26609,N_23302,N_23865);
and U26610 (N_26610,N_24518,N_24275);
and U26611 (N_26611,N_24579,N_21760);
or U26612 (N_26612,N_22709,N_22437);
or U26613 (N_26613,N_23917,N_23771);
xor U26614 (N_26614,N_20646,N_22200);
or U26615 (N_26615,N_24081,N_23000);
and U26616 (N_26616,N_20985,N_20637);
or U26617 (N_26617,N_20060,N_20405);
and U26618 (N_26618,N_20631,N_24534);
or U26619 (N_26619,N_22819,N_23332);
or U26620 (N_26620,N_24099,N_22607);
nand U26621 (N_26621,N_24880,N_24581);
or U26622 (N_26622,N_23157,N_21545);
xor U26623 (N_26623,N_20184,N_20932);
or U26624 (N_26624,N_23849,N_21311);
or U26625 (N_26625,N_21832,N_22370);
nand U26626 (N_26626,N_22800,N_21028);
xor U26627 (N_26627,N_23562,N_21243);
and U26628 (N_26628,N_22942,N_24340);
nand U26629 (N_26629,N_23240,N_23588);
xnor U26630 (N_26630,N_24182,N_24756);
or U26631 (N_26631,N_23694,N_23582);
xor U26632 (N_26632,N_23985,N_21535);
nor U26633 (N_26633,N_23216,N_23159);
or U26634 (N_26634,N_24794,N_23045);
nand U26635 (N_26635,N_23999,N_23740);
nand U26636 (N_26636,N_23982,N_24704);
nand U26637 (N_26637,N_20582,N_22554);
and U26638 (N_26638,N_22101,N_20090);
nor U26639 (N_26639,N_24127,N_22726);
or U26640 (N_26640,N_21680,N_22078);
and U26641 (N_26641,N_22601,N_21826);
nor U26642 (N_26642,N_22787,N_24469);
and U26643 (N_26643,N_22513,N_20861);
or U26644 (N_26644,N_23436,N_22707);
xor U26645 (N_26645,N_24935,N_21641);
xor U26646 (N_26646,N_23285,N_23203);
or U26647 (N_26647,N_23636,N_20867);
nor U26648 (N_26648,N_20125,N_20778);
or U26649 (N_26649,N_24371,N_20379);
nand U26650 (N_26650,N_23580,N_23468);
or U26651 (N_26651,N_24726,N_20155);
xor U26652 (N_26652,N_20552,N_21697);
nand U26653 (N_26653,N_22538,N_23144);
nor U26654 (N_26654,N_23419,N_24087);
nor U26655 (N_26655,N_22103,N_21810);
nor U26656 (N_26656,N_22322,N_23151);
nor U26657 (N_26657,N_20914,N_20677);
nor U26658 (N_26658,N_24572,N_23405);
and U26659 (N_26659,N_24598,N_24864);
nor U26660 (N_26660,N_21848,N_20753);
nand U26661 (N_26661,N_22017,N_23138);
and U26662 (N_26662,N_23277,N_22040);
xor U26663 (N_26663,N_20871,N_20236);
and U26664 (N_26664,N_21840,N_23689);
and U26665 (N_26665,N_24456,N_21201);
nor U26666 (N_26666,N_23943,N_23721);
nor U26667 (N_26667,N_22189,N_21947);
nand U26668 (N_26668,N_21315,N_21010);
xor U26669 (N_26669,N_22829,N_24433);
or U26670 (N_26670,N_21179,N_22208);
or U26671 (N_26671,N_23163,N_22627);
nand U26672 (N_26672,N_24411,N_22038);
and U26673 (N_26673,N_23765,N_23587);
xor U26674 (N_26674,N_21800,N_20988);
nor U26675 (N_26675,N_20624,N_21309);
or U26676 (N_26676,N_21827,N_22214);
xor U26677 (N_26677,N_22491,N_24907);
nor U26678 (N_26678,N_23473,N_22835);
nor U26679 (N_26679,N_20351,N_22186);
xor U26680 (N_26680,N_24203,N_20983);
nand U26681 (N_26681,N_21408,N_23633);
and U26682 (N_26682,N_22540,N_22809);
nand U26683 (N_26683,N_24320,N_20464);
nor U26684 (N_26684,N_21895,N_21885);
and U26685 (N_26685,N_20243,N_22658);
or U26686 (N_26686,N_20216,N_20438);
nor U26687 (N_26687,N_22832,N_22534);
nor U26688 (N_26688,N_20757,N_20781);
or U26689 (N_26689,N_22366,N_23603);
or U26690 (N_26690,N_23294,N_20577);
and U26691 (N_26691,N_21591,N_22802);
or U26692 (N_26692,N_21235,N_22751);
and U26693 (N_26693,N_23948,N_20750);
and U26694 (N_26694,N_20084,N_22490);
nor U26695 (N_26695,N_20478,N_23080);
and U26696 (N_26696,N_23252,N_23593);
and U26697 (N_26697,N_22381,N_22450);
xor U26698 (N_26698,N_20213,N_20241);
nor U26699 (N_26699,N_23639,N_24921);
nor U26700 (N_26700,N_22886,N_23312);
and U26701 (N_26701,N_21378,N_21864);
and U26702 (N_26702,N_24489,N_24903);
xor U26703 (N_26703,N_20082,N_22169);
nor U26704 (N_26704,N_22938,N_21648);
xor U26705 (N_26705,N_24836,N_23026);
and U26706 (N_26706,N_21707,N_22923);
and U26707 (N_26707,N_22755,N_20928);
and U26708 (N_26708,N_22866,N_21374);
and U26709 (N_26709,N_21337,N_23950);
xor U26710 (N_26710,N_23485,N_24388);
nor U26711 (N_26711,N_20138,N_23715);
or U26712 (N_26712,N_21559,N_23239);
nand U26713 (N_26713,N_24793,N_22769);
and U26714 (N_26714,N_24906,N_21036);
nand U26715 (N_26715,N_22785,N_24766);
nor U26716 (N_26716,N_21967,N_23774);
nor U26717 (N_26717,N_21880,N_21516);
nor U26718 (N_26718,N_21533,N_22713);
nand U26719 (N_26719,N_20518,N_24252);
nor U26720 (N_26720,N_23798,N_21228);
and U26721 (N_26721,N_23270,N_21115);
nor U26722 (N_26722,N_20569,N_20592);
nor U26723 (N_26723,N_23321,N_21277);
nor U26724 (N_26724,N_24796,N_20309);
xor U26725 (N_26725,N_23941,N_23017);
xor U26726 (N_26726,N_24559,N_23644);
nand U26727 (N_26727,N_22185,N_21468);
and U26728 (N_26728,N_22492,N_24904);
nand U26729 (N_26729,N_24591,N_22932);
and U26730 (N_26730,N_21596,N_23879);
nor U26731 (N_26731,N_23718,N_20395);
nor U26732 (N_26732,N_24926,N_24554);
or U26733 (N_26733,N_21101,N_21120);
nor U26734 (N_26734,N_23577,N_24934);
or U26735 (N_26735,N_23454,N_20320);
and U26736 (N_26736,N_20712,N_23174);
or U26737 (N_26737,N_22383,N_24828);
nor U26738 (N_26738,N_24710,N_21414);
and U26739 (N_26739,N_21859,N_24612);
and U26740 (N_26740,N_21127,N_23259);
and U26741 (N_26741,N_23893,N_22217);
and U26742 (N_26742,N_20154,N_24122);
xnor U26743 (N_26743,N_21602,N_23538);
nand U26744 (N_26744,N_23074,N_23940);
nand U26745 (N_26745,N_20129,N_22438);
and U26746 (N_26746,N_24472,N_23594);
xnor U26747 (N_26747,N_23188,N_22257);
xor U26748 (N_26748,N_23983,N_21490);
and U26749 (N_26749,N_24273,N_20113);
nand U26750 (N_26750,N_21498,N_22530);
xnor U26751 (N_26751,N_22116,N_21148);
or U26752 (N_26752,N_21152,N_20760);
nor U26753 (N_26753,N_24606,N_24717);
nand U26754 (N_26754,N_23554,N_22057);
or U26755 (N_26755,N_21901,N_24820);
xnor U26756 (N_26756,N_23905,N_23435);
or U26757 (N_26757,N_23600,N_24764);
nand U26758 (N_26758,N_23129,N_20832);
nor U26759 (N_26759,N_21538,N_23352);
nand U26760 (N_26760,N_24937,N_20819);
nor U26761 (N_26761,N_20321,N_20380);
nand U26762 (N_26762,N_23489,N_23858);
xnor U26763 (N_26763,N_23143,N_20729);
xnor U26764 (N_26764,N_21389,N_22684);
nand U26765 (N_26765,N_23695,N_20004);
and U26766 (N_26766,N_24674,N_20532);
nor U26767 (N_26767,N_22385,N_21341);
xnor U26768 (N_26768,N_23299,N_20422);
or U26769 (N_26769,N_24063,N_20617);
nor U26770 (N_26770,N_23340,N_24024);
xnor U26771 (N_26771,N_20331,N_22807);
nand U26772 (N_26772,N_22615,N_23103);
or U26773 (N_26773,N_24348,N_21332);
nand U26774 (N_26774,N_24568,N_22338);
nand U26775 (N_26775,N_24980,N_24109);
nor U26776 (N_26776,N_23782,N_24048);
and U26777 (N_26777,N_20955,N_20048);
nand U26778 (N_26778,N_21900,N_20543);
xnor U26779 (N_26779,N_23470,N_24769);
xor U26780 (N_26780,N_22798,N_21246);
nor U26781 (N_26781,N_23814,N_22237);
nand U26782 (N_26782,N_22133,N_20676);
or U26783 (N_26783,N_23286,N_21424);
nand U26784 (N_26784,N_22870,N_22030);
or U26785 (N_26785,N_20737,N_23238);
nor U26786 (N_26786,N_21951,N_21916);
nand U26787 (N_26787,N_21270,N_24039);
nand U26788 (N_26788,N_21001,N_21255);
xor U26789 (N_26789,N_20407,N_24401);
nand U26790 (N_26790,N_22823,N_22826);
and U26791 (N_26791,N_20208,N_21366);
or U26792 (N_26792,N_20366,N_22129);
or U26793 (N_26793,N_20325,N_20259);
nand U26794 (N_26794,N_21514,N_21721);
nand U26795 (N_26795,N_20294,N_21008);
nand U26796 (N_26796,N_22400,N_20485);
nand U26797 (N_26797,N_20274,N_23164);
and U26798 (N_26798,N_22995,N_20162);
and U26799 (N_26799,N_23195,N_23408);
and U26800 (N_26800,N_21852,N_24457);
and U26801 (N_26801,N_24703,N_24238);
xor U26802 (N_26802,N_22791,N_20535);
or U26803 (N_26803,N_21460,N_23601);
and U26804 (N_26804,N_22988,N_22984);
and U26805 (N_26805,N_21145,N_22109);
nor U26806 (N_26806,N_21386,N_23955);
nand U26807 (N_26807,N_24942,N_24165);
xnor U26808 (N_26808,N_21224,N_21132);
nand U26809 (N_26809,N_23275,N_22813);
or U26810 (N_26810,N_23196,N_21264);
or U26811 (N_26811,N_20558,N_21187);
and U26812 (N_26812,N_23683,N_21530);
nand U26813 (N_26813,N_20406,N_24337);
nand U26814 (N_26814,N_21024,N_23935);
and U26815 (N_26815,N_23165,N_21173);
nand U26816 (N_26816,N_20400,N_21478);
xor U26817 (N_26817,N_20151,N_22489);
xnor U26818 (N_26818,N_22690,N_23884);
or U26819 (N_26819,N_21338,N_20898);
and U26820 (N_26820,N_23213,N_24438);
and U26821 (N_26821,N_22619,N_23622);
xnor U26822 (N_26822,N_23140,N_20284);
nor U26823 (N_26823,N_20704,N_21447);
nand U26824 (N_26824,N_20510,N_24436);
and U26825 (N_26825,N_23525,N_22801);
or U26826 (N_26826,N_22899,N_22089);
nor U26827 (N_26827,N_22760,N_24159);
nand U26828 (N_26828,N_20300,N_23682);
nor U26829 (N_26829,N_21627,N_20875);
nor U26830 (N_26830,N_23848,N_22461);
or U26831 (N_26831,N_22783,N_20172);
xor U26832 (N_26832,N_20683,N_22478);
nor U26833 (N_26833,N_24783,N_23179);
xnor U26834 (N_26834,N_20645,N_20826);
xor U26835 (N_26835,N_24207,N_23121);
or U26836 (N_26836,N_21364,N_22693);
xor U26837 (N_26837,N_24434,N_20526);
nor U26838 (N_26838,N_23670,N_23066);
nor U26839 (N_26839,N_23521,N_24447);
or U26840 (N_26840,N_24488,N_24228);
and U26841 (N_26841,N_21052,N_22439);
nor U26842 (N_26842,N_22294,N_23680);
nor U26843 (N_26843,N_24603,N_20731);
nor U26844 (N_26844,N_23907,N_21747);
nand U26845 (N_26845,N_22303,N_22766);
xor U26846 (N_26846,N_20765,N_22820);
nor U26847 (N_26847,N_24019,N_24211);
and U26848 (N_26848,N_20018,N_24563);
nand U26849 (N_26849,N_22485,N_21952);
nor U26850 (N_26850,N_23009,N_23652);
nor U26851 (N_26851,N_21502,N_21925);
or U26852 (N_26852,N_21926,N_21401);
and U26853 (N_26853,N_22731,N_20863);
or U26854 (N_26854,N_23705,N_21931);
xnor U26855 (N_26855,N_20308,N_23254);
xor U26856 (N_26856,N_24245,N_21437);
or U26857 (N_26857,N_23957,N_22333);
and U26858 (N_26858,N_22579,N_22011);
nand U26859 (N_26859,N_20682,N_23128);
nor U26860 (N_26860,N_20714,N_24061);
and U26861 (N_26861,N_24205,N_21783);
xnor U26862 (N_26862,N_21079,N_23997);
nand U26863 (N_26863,N_24043,N_21991);
nor U26864 (N_26864,N_20505,N_24341);
nand U26865 (N_26865,N_22812,N_20065);
or U26866 (N_26866,N_23110,N_22376);
nor U26867 (N_26867,N_21075,N_20170);
xnor U26868 (N_26868,N_22363,N_20847);
nand U26869 (N_26869,N_23384,N_23402);
nor U26870 (N_26870,N_24634,N_21454);
or U26871 (N_26871,N_22637,N_20828);
nand U26872 (N_26872,N_21959,N_22064);
and U26873 (N_26873,N_22182,N_22475);
xnor U26874 (N_26874,N_22884,N_24426);
nand U26875 (N_26875,N_22006,N_24738);
nor U26876 (N_26876,N_24461,N_21319);
xnor U26877 (N_26877,N_21970,N_21174);
xor U26878 (N_26878,N_24141,N_24940);
nand U26879 (N_26879,N_22776,N_24626);
or U26880 (N_26880,N_22181,N_24596);
and U26881 (N_26881,N_22272,N_21527);
nand U26882 (N_26882,N_23688,N_24960);
or U26883 (N_26883,N_22881,N_22132);
and U26884 (N_26884,N_21213,N_20698);
xor U26885 (N_26885,N_23251,N_20426);
nor U26886 (N_26886,N_22291,N_24833);
or U26887 (N_26887,N_20054,N_21944);
nor U26888 (N_26888,N_21372,N_22081);
nand U26889 (N_26889,N_21291,N_21086);
and U26890 (N_26890,N_22839,N_23729);
xor U26891 (N_26891,N_23560,N_23460);
xnor U26892 (N_26892,N_21094,N_24336);
xor U26893 (N_26893,N_22825,N_21171);
and U26894 (N_26894,N_22857,N_21982);
nor U26895 (N_26895,N_24387,N_21569);
nand U26896 (N_26896,N_22474,N_20772);
or U26897 (N_26897,N_23779,N_21740);
nor U26898 (N_26898,N_21633,N_20752);
and U26899 (N_26899,N_20462,N_20764);
nand U26900 (N_26900,N_20029,N_23253);
and U26901 (N_26901,N_20159,N_21922);
nor U26902 (N_26902,N_24022,N_21955);
or U26903 (N_26903,N_20639,N_22774);
and U26904 (N_26904,N_22587,N_22885);
nor U26905 (N_26905,N_21129,N_24266);
and U26906 (N_26906,N_23698,N_24944);
and U26907 (N_26907,N_20186,N_23912);
and U26908 (N_26908,N_20929,N_20823);
xnor U26909 (N_26909,N_21204,N_20106);
xor U26910 (N_26910,N_24699,N_24482);
nor U26911 (N_26911,N_23287,N_20083);
nor U26912 (N_26912,N_23716,N_24737);
xnor U26913 (N_26913,N_24172,N_23148);
nand U26914 (N_26914,N_24897,N_21913);
and U26915 (N_26915,N_23832,N_21257);
and U26916 (N_26916,N_22633,N_24730);
and U26917 (N_26917,N_22188,N_24919);
nand U26918 (N_26918,N_21890,N_22877);
nand U26919 (N_26919,N_21594,N_21494);
nor U26920 (N_26920,N_21720,N_23229);
and U26921 (N_26921,N_22142,N_23659);
nand U26922 (N_26922,N_22114,N_22347);
and U26923 (N_26923,N_24086,N_23606);
xor U26924 (N_26924,N_20560,N_22411);
nand U26925 (N_26925,N_21774,N_24657);
or U26926 (N_26926,N_23676,N_22696);
or U26927 (N_26927,N_23320,N_21561);
or U26928 (N_26928,N_22963,N_22042);
and U26929 (N_26929,N_21405,N_22014);
and U26930 (N_26930,N_24791,N_20853);
xnor U26931 (N_26931,N_20571,N_23710);
and U26932 (N_26932,N_23385,N_23166);
nor U26933 (N_26933,N_21873,N_20000);
nor U26934 (N_26934,N_22426,N_21057);
or U26935 (N_26935,N_21185,N_24117);
and U26936 (N_26936,N_23135,N_20227);
nand U26937 (N_26937,N_22482,N_24496);
and U26938 (N_26938,N_21834,N_21234);
and U26939 (N_26939,N_21899,N_21731);
or U26940 (N_26940,N_20938,N_23640);
nor U26941 (N_26941,N_20231,N_22041);
nand U26942 (N_26942,N_21847,N_23221);
or U26943 (N_26943,N_24013,N_20686);
and U26944 (N_26944,N_22230,N_21693);
or U26945 (N_26945,N_21924,N_24560);
nand U26946 (N_26946,N_23915,N_24509);
nor U26947 (N_26947,N_22292,N_23300);
and U26948 (N_26948,N_24111,N_21841);
or U26949 (N_26949,N_22902,N_24466);
xor U26950 (N_26950,N_20307,N_20551);
nand U26951 (N_26951,N_22471,N_21198);
and U26952 (N_26952,N_22951,N_23042);
or U26953 (N_26953,N_23139,N_21106);
and U26954 (N_26954,N_21138,N_22407);
and U26955 (N_26955,N_21727,N_21581);
and U26956 (N_26956,N_22273,N_23231);
nor U26957 (N_26957,N_23902,N_22332);
xor U26958 (N_26958,N_20921,N_21908);
nor U26959 (N_26959,N_20911,N_24502);
or U26960 (N_26960,N_24687,N_20963);
and U26961 (N_26961,N_21572,N_23169);
or U26962 (N_26962,N_24729,N_24714);
nand U26963 (N_26963,N_24538,N_20726);
and U26964 (N_26964,N_20978,N_23260);
nand U26965 (N_26965,N_22817,N_20808);
xor U26966 (N_26966,N_23674,N_21231);
nor U26967 (N_26967,N_24599,N_20049);
nor U26968 (N_26968,N_20391,N_21004);
xor U26969 (N_26969,N_23693,N_20097);
nor U26970 (N_26970,N_22070,N_20477);
nor U26971 (N_26971,N_23092,N_23314);
and U26972 (N_26972,N_24786,N_21689);
or U26973 (N_26973,N_20918,N_21618);
xor U26974 (N_26974,N_23019,N_21323);
nand U26975 (N_26975,N_22850,N_23183);
nand U26976 (N_26976,N_20783,N_21981);
xor U26977 (N_26977,N_22539,N_24074);
nand U26978 (N_26978,N_23167,N_21653);
nand U26979 (N_26979,N_24071,N_22028);
xor U26980 (N_26980,N_20538,N_23630);
xnor U26981 (N_26981,N_21820,N_22896);
nor U26982 (N_26982,N_20791,N_24044);
nor U26983 (N_26983,N_22163,N_24003);
xor U26984 (N_26984,N_20235,N_22831);
or U26985 (N_26985,N_23399,N_20936);
nand U26986 (N_26986,N_21415,N_21299);
nor U26987 (N_26987,N_23806,N_21233);
xor U26988 (N_26988,N_22639,N_22313);
xnor U26989 (N_26989,N_20954,N_24933);
or U26990 (N_26990,N_24033,N_23387);
xnor U26991 (N_26991,N_20837,N_23634);
and U26992 (N_26992,N_22288,N_20598);
and U26993 (N_26993,N_21749,N_21664);
xnor U26994 (N_26994,N_23864,N_22666);
xor U26995 (N_26995,N_22311,N_22435);
nand U26996 (N_26996,N_23289,N_20210);
nor U26997 (N_26997,N_24120,N_24151);
nand U26998 (N_26998,N_22708,N_24060);
nor U26999 (N_26999,N_23816,N_23723);
and U27000 (N_27000,N_20786,N_24146);
or U27001 (N_27001,N_23427,N_22105);
nand U27002 (N_27002,N_21136,N_22147);
nand U27003 (N_27003,N_21842,N_23490);
nand U27004 (N_27004,N_23421,N_22701);
nand U27005 (N_27005,N_23526,N_23956);
and U27006 (N_27006,N_22985,N_23318);
nor U27007 (N_27007,N_21868,N_23131);
nand U27008 (N_27008,N_22934,N_24129);
and U27009 (N_27009,N_22000,N_21512);
and U27010 (N_27010,N_23186,N_24282);
or U27011 (N_27011,N_21686,N_22035);
xor U27012 (N_27012,N_21248,N_22432);
nand U27013 (N_27013,N_20531,N_20548);
xor U27014 (N_27014,N_22683,N_20026);
nand U27015 (N_27015,N_20755,N_24597);
or U27016 (N_27016,N_23981,N_23965);
nand U27017 (N_27017,N_23111,N_24034);
and U27018 (N_27018,N_21585,N_24346);
nand U27019 (N_27019,N_20690,N_23944);
nand U27020 (N_27020,N_23335,N_21789);
or U27021 (N_27021,N_20459,N_24645);
or U27022 (N_27022,N_23781,N_22286);
and U27023 (N_27023,N_24805,N_23175);
nand U27024 (N_27024,N_20943,N_24458);
and U27025 (N_27025,N_22260,N_24280);
or U27026 (N_27026,N_24224,N_21093);
xnor U27027 (N_27027,N_23799,N_22925);
or U27028 (N_27028,N_24741,N_21349);
nand U27029 (N_27029,N_22235,N_24566);
nor U27030 (N_27030,N_23050,N_24987);
nand U27031 (N_27031,N_20142,N_22339);
or U27032 (N_27032,N_24787,N_23181);
or U27033 (N_27033,N_20249,N_23467);
nor U27034 (N_27034,N_24613,N_21470);
or U27035 (N_27035,N_23857,N_24309);
nor U27036 (N_27036,N_23414,N_22834);
nor U27037 (N_27037,N_20473,N_24372);
nand U27038 (N_27038,N_20647,N_21758);
nand U27039 (N_27039,N_23942,N_20522);
nand U27040 (N_27040,N_24350,N_20492);
or U27041 (N_27041,N_23605,N_22897);
nor U27042 (N_27042,N_20071,N_21441);
nor U27043 (N_27043,N_22456,N_23846);
xnor U27044 (N_27044,N_22343,N_23409);
nor U27045 (N_27045,N_23951,N_20340);
xor U27046 (N_27046,N_20801,N_23932);
xnor U27047 (N_27047,N_20512,N_20754);
and U27048 (N_27048,N_23611,N_23372);
nand U27049 (N_27049,N_21518,N_24713);
xor U27050 (N_27050,N_23122,N_20114);
and U27051 (N_27051,N_22974,N_22571);
nor U27052 (N_27052,N_24986,N_20605);
or U27053 (N_27053,N_21432,N_22308);
and U27054 (N_27054,N_21588,N_21892);
and U27055 (N_27055,N_20428,N_23896);
and U27056 (N_27056,N_24512,N_22159);
xnor U27057 (N_27057,N_24885,N_24588);
nor U27058 (N_27058,N_20150,N_21605);
nor U27059 (N_27059,N_23212,N_21728);
nor U27060 (N_27060,N_22851,N_23855);
or U27061 (N_27061,N_21278,N_21887);
or U27062 (N_27062,N_22624,N_23202);
nand U27063 (N_27063,N_24510,N_20975);
and U27064 (N_27064,N_22642,N_20780);
xor U27065 (N_27065,N_22962,N_24380);
xnor U27066 (N_27066,N_20607,N_24630);
xnor U27067 (N_27067,N_22675,N_20058);
xor U27068 (N_27068,N_24546,N_24533);
nand U27069 (N_27069,N_23237,N_23350);
xor U27070 (N_27070,N_20458,N_20219);
or U27071 (N_27071,N_23037,N_23952);
nand U27072 (N_27072,N_22063,N_22060);
nor U27073 (N_27073,N_22910,N_23459);
or U27074 (N_27074,N_23062,N_23959);
nor U27075 (N_27075,N_24790,N_23177);
or U27076 (N_27076,N_23278,N_24985);
xor U27077 (N_27077,N_20089,N_20999);
or U27078 (N_27078,N_23297,N_24158);
nand U27079 (N_27079,N_21253,N_24827);
xor U27080 (N_27080,N_22124,N_20699);
nor U27081 (N_27081,N_23861,N_22153);
and U27082 (N_27082,N_21172,N_22777);
nor U27083 (N_27083,N_21670,N_23699);
or U27084 (N_27084,N_21729,N_21528);
nand U27085 (N_27085,N_21889,N_21354);
and U27086 (N_27086,N_21164,N_20008);
nand U27087 (N_27087,N_21296,N_21455);
nand U27088 (N_27088,N_24364,N_23837);
or U27089 (N_27089,N_21822,N_24732);
nand U27090 (N_27090,N_23069,N_22220);
nor U27091 (N_27091,N_20517,N_23563);
or U27092 (N_27092,N_22517,N_20649);
or U27093 (N_27093,N_23433,N_20317);
nor U27094 (N_27094,N_23653,N_22219);
xnor U27095 (N_27095,N_20890,N_23153);
nor U27096 (N_27096,N_20079,N_24889);
nand U27097 (N_27097,N_21566,N_20527);
and U27098 (N_27098,N_24248,N_24839);
nand U27099 (N_27099,N_23429,N_21896);
xor U27100 (N_27100,N_22634,N_24780);
nor U27101 (N_27101,N_23248,N_22298);
nor U27102 (N_27102,N_24824,N_22837);
xnor U27103 (N_27103,N_24640,N_24258);
nor U27104 (N_27104,N_22269,N_22729);
nand U27105 (N_27105,N_20192,N_20860);
nand U27106 (N_27106,N_20961,N_20796);
xor U27107 (N_27107,N_21609,N_20713);
nor U27108 (N_27108,N_23903,N_20530);
or U27109 (N_27109,N_22738,N_23784);
and U27110 (N_27110,N_23791,N_20016);
or U27111 (N_27111,N_23101,N_22037);
nor U27112 (N_27112,N_24576,N_23843);
nand U27113 (N_27113,N_21247,N_21520);
xor U27114 (N_27114,N_21371,N_23972);
nor U27115 (N_27115,N_23703,N_23137);
nand U27116 (N_27116,N_23268,N_23311);
nor U27117 (N_27117,N_20866,N_24446);
or U27118 (N_27118,N_21543,N_21342);
or U27119 (N_27119,N_21663,N_23936);
nand U27120 (N_27120,N_22446,N_21431);
or U27121 (N_27121,N_21813,N_24668);
xnor U27122 (N_27122,N_21090,N_23590);
and U27123 (N_27123,N_22982,N_20182);
and U27124 (N_27124,N_21565,N_24876);
or U27125 (N_27125,N_21081,N_20822);
nor U27126 (N_27126,N_23358,N_21391);
xnor U27127 (N_27127,N_24580,N_23913);
or U27128 (N_27128,N_20953,N_21125);
and U27129 (N_27129,N_20446,N_20562);
nand U27130 (N_27130,N_21343,N_20041);
nand U27131 (N_27131,N_20352,N_22602);
or U27132 (N_27132,N_24359,N_21048);
and U27133 (N_27133,N_20111,N_20644);
or U27134 (N_27134,N_24989,N_24920);
nand U27135 (N_27135,N_21675,N_22672);
nand U27136 (N_27136,N_22893,N_21180);
or U27137 (N_27137,N_24139,N_21334);
nor U27138 (N_27138,N_22223,N_22686);
xor U27139 (N_27139,N_24675,N_23333);
or U27140 (N_27140,N_21919,N_20751);
xor U27141 (N_27141,N_22113,N_20966);
nand U27142 (N_27142,N_22179,N_24589);
xor U27143 (N_27143,N_20580,N_24549);
nand U27144 (N_27144,N_23353,N_20093);
or U27145 (N_27145,N_23797,N_24570);
nor U27146 (N_27146,N_24390,N_24413);
or U27147 (N_27147,N_21541,N_24810);
or U27148 (N_27148,N_22569,N_23641);
or U27149 (N_27149,N_24586,N_22747);
and U27150 (N_27150,N_22341,N_24106);
nand U27151 (N_27151,N_20291,N_21980);
nand U27152 (N_27152,N_21274,N_22718);
nand U27153 (N_27153,N_22107,N_23359);
and U27154 (N_27154,N_23094,N_23003);
nand U27155 (N_27155,N_20671,N_21073);
and U27156 (N_27156,N_22576,N_20335);
and U27157 (N_27157,N_20266,N_24101);
nand U27158 (N_27158,N_23657,N_22104);
or U27159 (N_27159,N_20439,N_24777);
and U27160 (N_27160,N_23573,N_23906);
nand U27161 (N_27161,N_23626,N_21076);
or U27162 (N_27162,N_21555,N_23615);
nor U27163 (N_27163,N_23236,N_20523);
and U27164 (N_27164,N_20815,N_20566);
xor U27165 (N_27165,N_22599,N_22044);
and U27166 (N_27166,N_22858,N_23424);
or U27167 (N_27167,N_23217,N_20642);
nand U27168 (N_27168,N_21286,N_23939);
and U27169 (N_27169,N_20025,N_21621);
nor U27170 (N_27170,N_21504,N_20964);
nand U27171 (N_27171,N_24719,N_20730);
and U27172 (N_27172,N_21262,N_24281);
nor U27173 (N_27173,N_23496,N_20332);
xnor U27174 (N_27174,N_21601,N_23392);
or U27175 (N_27175,N_21603,N_24695);
xor U27176 (N_27176,N_24829,N_22842);
or U27177 (N_27177,N_21884,N_24499);
or U27178 (N_27178,N_24012,N_20032);
and U27179 (N_27179,N_24021,N_23146);
xnor U27180 (N_27180,N_21191,N_23184);
nor U27181 (N_27181,N_21807,N_20107);
nor U27182 (N_27182,N_24334,N_21112);
and U27183 (N_27183,N_24288,N_24329);
nand U27184 (N_27184,N_21570,N_21250);
nand U27185 (N_27185,N_24347,N_20149);
xor U27186 (N_27186,N_22806,N_21665);
nand U27187 (N_27187,N_20226,N_22315);
nor U27188 (N_27188,N_24404,N_24088);
nand U27189 (N_27189,N_20993,N_20800);
and U27190 (N_27190,N_24119,N_23576);
nand U27191 (N_27191,N_23792,N_23566);
and U27192 (N_27192,N_23404,N_20678);
nor U27193 (N_27193,N_23617,N_20169);
nor U27194 (N_27194,N_22431,N_22330);
and U27195 (N_27195,N_21082,N_21828);
or U27196 (N_27196,N_22368,N_20744);
or U27197 (N_27197,N_23096,N_20456);
nor U27198 (N_27198,N_21396,N_20039);
nand U27199 (N_27199,N_23743,N_23764);
nor U27200 (N_27200,N_23613,N_23646);
nor U27201 (N_27201,N_22692,N_21722);
or U27202 (N_27202,N_24422,N_24316);
or U27203 (N_27203,N_20507,N_21656);
and U27204 (N_27204,N_20421,N_20242);
xor U27205 (N_27205,N_23136,N_22773);
nor U27206 (N_27206,N_22924,N_22195);
xnor U27207 (N_27207,N_21025,N_21888);
and U27208 (N_27208,N_20424,N_23558);
nor U27209 (N_27209,N_24169,N_22585);
and U27210 (N_27210,N_24381,N_22253);
xor U27211 (N_27211,N_23343,N_24219);
nor U27212 (N_27212,N_24114,N_24241);
or U27213 (N_27213,N_20742,N_22098);
nand U27214 (N_27214,N_21881,N_24148);
or U27215 (N_27215,N_23055,N_21595);
nand U27216 (N_27216,N_20506,N_20511);
nor U27217 (N_27217,N_23800,N_20546);
and U27218 (N_27218,N_22467,N_20570);
or U27219 (N_27219,N_23456,N_21259);
nand U27220 (N_27220,N_21033,N_24803);
nand U27221 (N_27221,N_22374,N_23929);
and U27222 (N_27222,N_20549,N_21929);
xnor U27223 (N_27223,N_20739,N_23726);
nand U27224 (N_27224,N_21205,N_20845);
nor U27225 (N_27225,N_23481,N_24602);
xor U27226 (N_27226,N_22232,N_20146);
nor U27227 (N_27227,N_20371,N_20572);
xor U27228 (N_27228,N_20720,N_22651);
or U27229 (N_27229,N_23147,N_22177);
xnor U27230 (N_27230,N_20212,N_23719);
nor U27231 (N_27231,N_22059,N_23961);
nor U27232 (N_27232,N_21268,N_23866);
and U27233 (N_27233,N_20657,N_22559);
xor U27234 (N_27234,N_20680,N_22762);
nor U27235 (N_27235,N_21390,N_24854);
and U27236 (N_27236,N_20779,N_23088);
nor U27237 (N_27237,N_22440,N_24718);
xnor U27238 (N_27238,N_21092,N_20941);
or U27239 (N_27239,N_21223,N_24665);
nand U27240 (N_27240,N_20205,N_22556);
or U27241 (N_27241,N_24093,N_24180);
xor U27242 (N_27242,N_23413,N_21643);
nand U27243 (N_27243,N_22999,N_20524);
nand U27244 (N_27244,N_21333,N_20370);
and U27245 (N_27245,N_20311,N_23592);
and U27246 (N_27246,N_24561,N_24226);
nand U27247 (N_27247,N_24103,N_20001);
nor U27248 (N_27248,N_23863,N_21116);
and U27249 (N_27249,N_20173,N_20440);
nor U27250 (N_27250,N_24156,N_20365);
nor U27251 (N_27251,N_24414,N_24398);
and U27252 (N_27252,N_23829,N_23795);
and U27253 (N_27253,N_20206,N_21182);
xnor U27254 (N_27254,N_23510,N_22324);
xnor U27255 (N_27255,N_20499,N_21750);
nand U27256 (N_27256,N_24133,N_24356);
and U27257 (N_27257,N_21472,N_23028);
and U27258 (N_27258,N_24452,N_24670);
xor U27259 (N_27259,N_20565,N_20283);
nand U27260 (N_27260,N_24733,N_21326);
nor U27261 (N_27261,N_22978,N_23440);
nor U27262 (N_27262,N_23732,N_24523);
or U27263 (N_27263,N_23130,N_24771);
or U27264 (N_27264,N_20245,N_20625);
nand U27265 (N_27265,N_23291,N_24571);
xnor U27266 (N_27266,N_24784,N_21897);
nand U27267 (N_27267,N_20903,N_21190);
nand U27268 (N_27268,N_20747,N_20130);
nor U27269 (N_27269,N_21515,N_23629);
xor U27270 (N_27270,N_22811,N_22753);
xnor U27271 (N_27271,N_24843,N_21110);
nand U27272 (N_27272,N_22167,N_21839);
nor U27273 (N_27273,N_24853,N_23888);
nor U27274 (N_27274,N_23968,N_21907);
and U27275 (N_27275,N_24420,N_21719);
nand U27276 (N_27276,N_20502,N_22419);
and U27277 (N_27277,N_21088,N_20314);
or U27278 (N_27278,N_22681,N_20603);
xnor U27279 (N_27279,N_22391,N_23926);
or U27280 (N_27280,N_20672,N_21361);
and U27281 (N_27281,N_24353,N_20046);
nand U27282 (N_27282,N_20070,N_23768);
nor U27283 (N_27283,N_24661,N_20148);
xnor U27284 (N_27284,N_21855,N_24409);
xnor U27285 (N_27285,N_22551,N_22479);
xnor U27286 (N_27286,N_20509,N_20513);
xor U27287 (N_27287,N_21417,N_23623);
or U27288 (N_27288,N_22852,N_20285);
nand U27289 (N_27289,N_24222,N_24197);
or U27290 (N_27290,N_22423,N_22494);
and U27291 (N_27291,N_21709,N_20945);
nor U27292 (N_27292,N_23243,N_21477);
nor U27293 (N_27293,N_23690,N_22989);
xor U27294 (N_27294,N_20091,N_24632);
and U27295 (N_27295,N_24431,N_23826);
nor U27296 (N_27296,N_23480,N_24333);
and U27297 (N_27297,N_20023,N_20991);
xnor U27298 (N_27298,N_20719,N_24516);
or U27299 (N_27299,N_24821,N_20409);
nor U27300 (N_27300,N_23242,N_20318);
xor U27301 (N_27301,N_23801,N_22536);
or U27302 (N_27302,N_20419,N_24594);
or U27303 (N_27303,N_23692,N_24869);
xnor U27304 (N_27304,N_22878,N_23362);
or U27305 (N_27305,N_22548,N_21394);
nand U27306 (N_27306,N_22833,N_20718);
xor U27307 (N_27307,N_21701,N_21215);
nand U27308 (N_27308,N_21876,N_23380);
nand U27309 (N_27309,N_20362,N_23337);
nand U27310 (N_27310,N_22301,N_23117);
nor U27311 (N_27311,N_20597,N_23098);
and U27312 (N_27312,N_23125,N_20516);
nand U27313 (N_27313,N_20641,N_21169);
xnor U27314 (N_27314,N_22720,N_21546);
nand U27315 (N_27315,N_21290,N_21167);
xor U27316 (N_27316,N_24296,N_23031);
or U27317 (N_27317,N_23303,N_22689);
nor U27318 (N_27318,N_21458,N_22061);
and U27319 (N_27319,N_24956,N_23382);
xor U27320 (N_27320,N_24343,N_22095);
or U27321 (N_27321,N_20027,N_23060);
xor U27322 (N_27322,N_24698,N_21448);
and U27323 (N_27323,N_24204,N_23004);
and U27324 (N_27324,N_23227,N_23326);
nor U27325 (N_27325,N_20074,N_22264);
nor U27326 (N_27326,N_21236,N_23114);
or U27327 (N_27327,N_20204,N_24253);
nand U27328 (N_27328,N_22443,N_24961);
and U27329 (N_27329,N_24631,N_24607);
and U27330 (N_27330,N_21181,N_22180);
or U27331 (N_27331,N_24464,N_24813);
nand U27332 (N_27332,N_22867,N_23933);
and U27333 (N_27333,N_23934,N_21764);
or U27334 (N_27334,N_21780,N_24725);
xnor U27335 (N_27335,N_24639,N_22350);
nand U27336 (N_27336,N_24963,N_24605);
nor U27337 (N_27337,N_22649,N_24841);
nand U27338 (N_27338,N_24795,N_24528);
and U27339 (N_27339,N_21147,N_20831);
or U27340 (N_27340,N_20166,N_24396);
xnor U27341 (N_27341,N_20465,N_23586);
or U27342 (N_27342,N_23378,N_20306);
or U27343 (N_27343,N_23656,N_24031);
xor U27344 (N_27344,N_23673,N_24542);
nand U27345 (N_27345,N_20197,N_24955);
nor U27346 (N_27346,N_24851,N_21958);
nor U27347 (N_27347,N_23596,N_22483);
or U27348 (N_27348,N_21677,N_21005);
xnor U27349 (N_27349,N_22603,N_24225);
nand U27350 (N_27350,N_21043,N_22039);
or U27351 (N_27351,N_22118,N_20330);
nand U27352 (N_27352,N_22010,N_24376);
and U27353 (N_27353,N_20248,N_20287);
and U27354 (N_27354,N_22732,N_22085);
and U27355 (N_27355,N_20588,N_24030);
nand U27356 (N_27356,N_20585,N_21583);
nand U27357 (N_27357,N_23869,N_23559);
xor U27358 (N_27358,N_24999,N_23758);
and U27359 (N_27359,N_22287,N_22940);
xnor U27360 (N_27360,N_20152,N_21753);
or U27361 (N_27361,N_23249,N_22968);
or U27362 (N_27362,N_21598,N_24011);
nand U27363 (N_27363,N_21971,N_23272);
xnor U27364 (N_27364,N_20693,N_24574);
and U27365 (N_27365,N_20022,N_24416);
nor U27366 (N_27366,N_21080,N_24459);
nor U27367 (N_27367,N_20912,N_24883);
xor U27368 (N_27368,N_23010,N_22869);
and U27369 (N_27369,N_24845,N_23789);
or U27370 (N_27370,N_22094,N_20189);
nor U27371 (N_27371,N_23418,N_22593);
or U27372 (N_27372,N_20854,N_24246);
xnor U27373 (N_27373,N_24069,N_22125);
nor U27374 (N_27374,N_21791,N_22915);
nand U27375 (N_27375,N_22892,N_24722);
xnor U27376 (N_27376,N_23057,N_20940);
xor U27377 (N_27377,N_20063,N_20207);
nand U27378 (N_27378,N_22525,N_20388);
or U27379 (N_27379,N_22102,N_23891);
and U27380 (N_27380,N_21524,N_21192);
nand U27381 (N_27381,N_20037,N_22122);
nand U27382 (N_27382,N_23126,N_21023);
xor U27383 (N_27383,N_23738,N_20295);
nor U27384 (N_27384,N_20809,N_22123);
nand U27385 (N_27385,N_22120,N_24838);
or U27386 (N_27386,N_24243,N_20986);
and U27387 (N_27387,N_21034,N_22086);
xor U27388 (N_27388,N_20483,N_23838);
nand U27389 (N_27389,N_21197,N_24575);
or U27390 (N_27390,N_21718,N_21423);
xnor U27391 (N_27391,N_24397,N_20057);
or U27392 (N_27392,N_20651,N_21667);
and U27393 (N_27393,N_20143,N_24951);
nor U27394 (N_27394,N_21352,N_23182);
and U27395 (N_27395,N_21995,N_24167);
nand U27396 (N_27396,N_23535,N_24629);
xor U27397 (N_27397,N_24453,N_21087);
nand U27398 (N_27398,N_24721,N_22657);
or U27399 (N_27399,N_24712,N_22703);
or U27400 (N_27400,N_23529,N_22077);
nand U27401 (N_27401,N_24302,N_24123);
nor U27402 (N_27402,N_20470,N_22815);
nand U27403 (N_27403,N_24215,N_22386);
nand U27404 (N_27404,N_20852,N_23437);
or U27405 (N_27405,N_23870,N_23224);
nand U27406 (N_27406,N_21505,N_20967);
and U27407 (N_27407,N_21014,N_21778);
and U27408 (N_27408,N_21636,N_22862);
nor U27409 (N_27409,N_23391,N_21539);
or U27410 (N_27410,N_24918,N_23925);
and U27411 (N_27411,N_20501,N_22533);
xnor U27412 (N_27412,N_20496,N_23256);
nand U27413 (N_27413,N_21327,N_23977);
nand U27414 (N_27414,N_22737,N_23379);
nand U27415 (N_27415,N_20612,N_21966);
and U27416 (N_27416,N_24188,N_21013);
nand U27417 (N_27417,N_22518,N_21161);
xnor U27418 (N_27418,N_23200,N_23046);
nor U27419 (N_27419,N_21222,N_22004);
nor U27420 (N_27420,N_23895,N_22563);
and U27421 (N_27421,N_24175,N_20574);
and U27422 (N_27422,N_21761,N_24144);
xor U27423 (N_27423,N_24970,N_20051);
xor U27424 (N_27424,N_20596,N_21575);
or U27425 (N_27425,N_22227,N_20109);
xnor U27426 (N_27426,N_24233,N_21961);
xor U27427 (N_27427,N_22239,N_22845);
or U27428 (N_27428,N_21162,N_21759);
or U27429 (N_27429,N_22022,N_20158);
and U27430 (N_27430,N_22263,N_21020);
xor U27431 (N_27431,N_20044,N_23008);
or U27432 (N_27432,N_23426,N_20437);
and U27433 (N_27433,N_24294,N_21671);
nand U27434 (N_27434,N_22401,N_22158);
xnor U27435 (N_27435,N_24558,N_24462);
nor U27436 (N_27436,N_21074,N_23557);
xor U27437 (N_27437,N_21673,N_22126);
xnor U27438 (N_27438,N_24625,N_23211);
or U27439 (N_27439,N_21392,N_20110);
nand U27440 (N_27440,N_23205,N_20843);
nor U27441 (N_27441,N_21788,N_23778);
or U27442 (N_27442,N_24543,N_22183);
xor U27443 (N_27443,N_24535,N_21987);
nor U27444 (N_27444,N_21103,N_20333);
or U27445 (N_27445,N_23642,N_21011);
or U27446 (N_27446,N_24852,N_24450);
or U27447 (N_27447,N_23647,N_23029);
nor U27448 (N_27448,N_20886,N_24866);
xnor U27449 (N_27449,N_22255,N_21974);
xnor U27450 (N_27450,N_20145,N_20841);
or U27451 (N_27451,N_20147,N_21806);
xor U27452 (N_27452,N_21451,N_24439);
nor U27453 (N_27453,N_23524,N_22013);
or U27454 (N_27454,N_23274,N_20636);
and U27455 (N_27455,N_22455,N_22289);
xnor U27456 (N_27456,N_24779,N_22699);
xnor U27457 (N_27457,N_22679,N_24250);
or U27458 (N_27458,N_20296,N_20743);
and U27459 (N_27459,N_22201,N_20980);
or U27460 (N_27460,N_20994,N_21935);
xnor U27461 (N_27461,N_20493,N_23691);
or U27462 (N_27462,N_22930,N_24046);
nand U27463 (N_27463,N_20774,N_23500);
nor U27464 (N_27464,N_24705,N_22691);
nor U27465 (N_27465,N_23407,N_24293);
nand U27466 (N_27466,N_21993,N_21141);
and U27467 (N_27467,N_22883,N_22406);
and U27468 (N_27468,N_24267,N_24731);
or U27469 (N_27469,N_22131,N_23987);
nand U27470 (N_27470,N_21444,N_23810);
nand U27471 (N_27471,N_24494,N_21027);
nand U27472 (N_27472,N_21016,N_21984);
nand U27473 (N_27473,N_20387,N_21314);
nand U27474 (N_27474,N_24890,N_23085);
and U27475 (N_27475,N_22912,N_22698);
nor U27476 (N_27476,N_20489,N_23280);
xnor U27477 (N_27477,N_22197,N_24049);
xor U27478 (N_27478,N_21495,N_21988);
nor U27479 (N_27479,N_22543,N_24332);
and U27480 (N_27480,N_24950,N_23090);
nand U27481 (N_27481,N_22606,N_22644);
or U27482 (N_27482,N_22790,N_21021);
and U27483 (N_27483,N_22792,N_21786);
nand U27484 (N_27484,N_24860,N_21767);
xnor U27485 (N_27485,N_24202,N_22216);
nor U27486 (N_27486,N_21766,N_23099);
and U27487 (N_27487,N_23991,N_21293);
nand U27488 (N_27488,N_24702,N_22827);
nand U27489 (N_27489,N_21622,N_23627);
xnor U27490 (N_27490,N_24047,N_22503);
xnor U27491 (N_27491,N_24210,N_20773);
nor U27492 (N_27492,N_21560,N_24976);
nand U27493 (N_27493,N_20264,N_24894);
and U27494 (N_27494,N_23356,N_21227);
nand U27495 (N_27495,N_21095,N_24104);
or U27496 (N_27496,N_20767,N_23746);
or U27497 (N_27497,N_20394,N_23106);
nand U27498 (N_27498,N_21373,N_24085);
and U27499 (N_27499,N_24256,N_22786);
nand U27500 (N_27500,N_20622,N_22599);
nand U27501 (N_27501,N_21636,N_21343);
and U27502 (N_27502,N_20329,N_21428);
and U27503 (N_27503,N_20747,N_20334);
nand U27504 (N_27504,N_24038,N_23532);
or U27505 (N_27505,N_23859,N_20046);
and U27506 (N_27506,N_24892,N_23197);
xnor U27507 (N_27507,N_24185,N_20945);
xnor U27508 (N_27508,N_21041,N_21752);
nor U27509 (N_27509,N_20867,N_24989);
and U27510 (N_27510,N_24801,N_20027);
nor U27511 (N_27511,N_24778,N_23019);
and U27512 (N_27512,N_21445,N_20884);
nand U27513 (N_27513,N_20308,N_21305);
or U27514 (N_27514,N_23924,N_22556);
xnor U27515 (N_27515,N_22494,N_23552);
and U27516 (N_27516,N_23003,N_22398);
and U27517 (N_27517,N_22702,N_24938);
and U27518 (N_27518,N_21822,N_21649);
xnor U27519 (N_27519,N_23033,N_23632);
or U27520 (N_27520,N_24269,N_21341);
xor U27521 (N_27521,N_23407,N_21860);
nor U27522 (N_27522,N_22329,N_24923);
or U27523 (N_27523,N_24319,N_24264);
xnor U27524 (N_27524,N_21524,N_20859);
or U27525 (N_27525,N_23522,N_22909);
and U27526 (N_27526,N_24552,N_23450);
nor U27527 (N_27527,N_24925,N_20648);
or U27528 (N_27528,N_24870,N_22590);
nor U27529 (N_27529,N_22236,N_24361);
and U27530 (N_27530,N_20921,N_20182);
and U27531 (N_27531,N_20268,N_23533);
xor U27532 (N_27532,N_23391,N_24905);
xnor U27533 (N_27533,N_20547,N_24595);
nor U27534 (N_27534,N_24885,N_22798);
and U27535 (N_27535,N_20164,N_21480);
or U27536 (N_27536,N_20640,N_22859);
nand U27537 (N_27537,N_24719,N_20566);
or U27538 (N_27538,N_21522,N_20082);
and U27539 (N_27539,N_20508,N_20495);
nand U27540 (N_27540,N_20009,N_22161);
nand U27541 (N_27541,N_24014,N_21778);
and U27542 (N_27542,N_20850,N_22074);
nor U27543 (N_27543,N_24164,N_20669);
nand U27544 (N_27544,N_20462,N_22382);
nand U27545 (N_27545,N_23992,N_21259);
and U27546 (N_27546,N_20311,N_20954);
or U27547 (N_27547,N_23578,N_23022);
nand U27548 (N_27548,N_23449,N_22434);
and U27549 (N_27549,N_20391,N_21481);
and U27550 (N_27550,N_23098,N_21196);
nor U27551 (N_27551,N_24041,N_23603);
or U27552 (N_27552,N_21357,N_20161);
xnor U27553 (N_27553,N_20249,N_24981);
or U27554 (N_27554,N_23527,N_20688);
xnor U27555 (N_27555,N_21798,N_24197);
or U27556 (N_27556,N_21067,N_21396);
xor U27557 (N_27557,N_21941,N_21322);
and U27558 (N_27558,N_21569,N_21994);
nand U27559 (N_27559,N_24192,N_24744);
nand U27560 (N_27560,N_23189,N_23605);
and U27561 (N_27561,N_21801,N_21360);
and U27562 (N_27562,N_23127,N_24813);
or U27563 (N_27563,N_21632,N_22585);
and U27564 (N_27564,N_23644,N_23816);
and U27565 (N_27565,N_23143,N_21400);
xor U27566 (N_27566,N_21809,N_24602);
or U27567 (N_27567,N_22063,N_21674);
and U27568 (N_27568,N_20490,N_21504);
xor U27569 (N_27569,N_23912,N_23973);
or U27570 (N_27570,N_23368,N_21467);
nor U27571 (N_27571,N_24107,N_22523);
or U27572 (N_27572,N_23225,N_22165);
or U27573 (N_27573,N_23785,N_21053);
nand U27574 (N_27574,N_20946,N_22987);
and U27575 (N_27575,N_24396,N_20257);
nand U27576 (N_27576,N_22786,N_24138);
xnor U27577 (N_27577,N_21721,N_23524);
xor U27578 (N_27578,N_23555,N_23647);
and U27579 (N_27579,N_23564,N_22781);
or U27580 (N_27580,N_24105,N_24603);
and U27581 (N_27581,N_23195,N_22097);
and U27582 (N_27582,N_22846,N_22657);
xor U27583 (N_27583,N_21591,N_21389);
nand U27584 (N_27584,N_23208,N_24545);
nor U27585 (N_27585,N_21279,N_21352);
xnor U27586 (N_27586,N_20500,N_24319);
nand U27587 (N_27587,N_22329,N_23415);
xnor U27588 (N_27588,N_21700,N_20293);
and U27589 (N_27589,N_24631,N_22110);
or U27590 (N_27590,N_21169,N_20646);
nand U27591 (N_27591,N_20918,N_21502);
and U27592 (N_27592,N_21339,N_22634);
nor U27593 (N_27593,N_22487,N_21368);
xor U27594 (N_27594,N_20864,N_20359);
xnor U27595 (N_27595,N_20446,N_20410);
nor U27596 (N_27596,N_23546,N_22768);
and U27597 (N_27597,N_20495,N_20922);
nor U27598 (N_27598,N_23267,N_20107);
or U27599 (N_27599,N_24051,N_20843);
xnor U27600 (N_27600,N_24620,N_24828);
nor U27601 (N_27601,N_21870,N_22037);
nor U27602 (N_27602,N_22268,N_20804);
or U27603 (N_27603,N_21519,N_21963);
and U27604 (N_27604,N_20017,N_24871);
or U27605 (N_27605,N_23817,N_23073);
nor U27606 (N_27606,N_22926,N_23373);
nor U27607 (N_27607,N_22507,N_20320);
or U27608 (N_27608,N_23126,N_22783);
xnor U27609 (N_27609,N_24167,N_23995);
nor U27610 (N_27610,N_22123,N_24185);
nand U27611 (N_27611,N_22594,N_22785);
and U27612 (N_27612,N_22851,N_20798);
and U27613 (N_27613,N_23067,N_22768);
and U27614 (N_27614,N_22340,N_22519);
xnor U27615 (N_27615,N_23502,N_24348);
xnor U27616 (N_27616,N_21555,N_23809);
or U27617 (N_27617,N_23713,N_24302);
and U27618 (N_27618,N_24441,N_22454);
or U27619 (N_27619,N_24974,N_20206);
nand U27620 (N_27620,N_20601,N_22736);
and U27621 (N_27621,N_24510,N_21134);
nor U27622 (N_27622,N_23916,N_22107);
or U27623 (N_27623,N_21405,N_21069);
xnor U27624 (N_27624,N_24513,N_24566);
nor U27625 (N_27625,N_23883,N_21744);
and U27626 (N_27626,N_21421,N_24247);
nor U27627 (N_27627,N_21849,N_24991);
or U27628 (N_27628,N_22632,N_23249);
nand U27629 (N_27629,N_24701,N_22755);
nand U27630 (N_27630,N_22705,N_23054);
nor U27631 (N_27631,N_21176,N_21863);
nand U27632 (N_27632,N_23993,N_22250);
or U27633 (N_27633,N_22987,N_21050);
nand U27634 (N_27634,N_24886,N_20497);
nor U27635 (N_27635,N_23089,N_24810);
or U27636 (N_27636,N_22715,N_24194);
nand U27637 (N_27637,N_23169,N_23617);
nand U27638 (N_27638,N_20532,N_21874);
nand U27639 (N_27639,N_24327,N_24667);
and U27640 (N_27640,N_20936,N_21895);
and U27641 (N_27641,N_23061,N_23344);
nor U27642 (N_27642,N_23055,N_20902);
nand U27643 (N_27643,N_20608,N_21307);
nor U27644 (N_27644,N_24142,N_24065);
nor U27645 (N_27645,N_20664,N_24029);
nor U27646 (N_27646,N_21136,N_22170);
and U27647 (N_27647,N_21707,N_20191);
and U27648 (N_27648,N_21465,N_20494);
and U27649 (N_27649,N_20118,N_21627);
and U27650 (N_27650,N_22332,N_21405);
and U27651 (N_27651,N_23272,N_24598);
xor U27652 (N_27652,N_20253,N_20169);
nor U27653 (N_27653,N_22074,N_20575);
nand U27654 (N_27654,N_20846,N_23816);
and U27655 (N_27655,N_20518,N_24284);
xor U27656 (N_27656,N_22300,N_22043);
nor U27657 (N_27657,N_23326,N_22163);
nand U27658 (N_27658,N_22152,N_23751);
or U27659 (N_27659,N_22543,N_23118);
or U27660 (N_27660,N_20308,N_21043);
nor U27661 (N_27661,N_21135,N_20635);
or U27662 (N_27662,N_20448,N_23230);
nand U27663 (N_27663,N_24010,N_20639);
nand U27664 (N_27664,N_21923,N_20827);
nand U27665 (N_27665,N_22499,N_20865);
xor U27666 (N_27666,N_22067,N_23764);
nor U27667 (N_27667,N_21065,N_20590);
nand U27668 (N_27668,N_20914,N_21636);
and U27669 (N_27669,N_23047,N_22648);
xor U27670 (N_27670,N_21431,N_22497);
nand U27671 (N_27671,N_20518,N_20146);
nor U27672 (N_27672,N_22575,N_21634);
nand U27673 (N_27673,N_20414,N_22258);
and U27674 (N_27674,N_23530,N_21316);
nor U27675 (N_27675,N_23288,N_20804);
xnor U27676 (N_27676,N_23396,N_23032);
nand U27677 (N_27677,N_22736,N_22034);
or U27678 (N_27678,N_22671,N_21934);
nor U27679 (N_27679,N_20865,N_23168);
xnor U27680 (N_27680,N_22615,N_23572);
xnor U27681 (N_27681,N_22113,N_24796);
and U27682 (N_27682,N_24570,N_22967);
nor U27683 (N_27683,N_23542,N_22785);
and U27684 (N_27684,N_21800,N_21761);
or U27685 (N_27685,N_24988,N_20302);
or U27686 (N_27686,N_20056,N_21922);
nand U27687 (N_27687,N_20942,N_22561);
xor U27688 (N_27688,N_22660,N_22746);
or U27689 (N_27689,N_23812,N_23951);
nand U27690 (N_27690,N_21707,N_23858);
or U27691 (N_27691,N_21346,N_20724);
nand U27692 (N_27692,N_24695,N_20910);
and U27693 (N_27693,N_21359,N_23705);
nand U27694 (N_27694,N_24470,N_20305);
nand U27695 (N_27695,N_21884,N_23386);
or U27696 (N_27696,N_22225,N_21868);
nor U27697 (N_27697,N_23599,N_21975);
nand U27698 (N_27698,N_22050,N_22028);
and U27699 (N_27699,N_24635,N_23770);
nor U27700 (N_27700,N_21003,N_20288);
nor U27701 (N_27701,N_23778,N_24186);
and U27702 (N_27702,N_23357,N_22805);
nor U27703 (N_27703,N_20935,N_22659);
nor U27704 (N_27704,N_20625,N_20085);
xnor U27705 (N_27705,N_20021,N_23391);
nand U27706 (N_27706,N_24580,N_22922);
xnor U27707 (N_27707,N_23992,N_24290);
nor U27708 (N_27708,N_24916,N_22991);
nor U27709 (N_27709,N_20856,N_23205);
and U27710 (N_27710,N_21321,N_22383);
nor U27711 (N_27711,N_24294,N_20863);
nor U27712 (N_27712,N_24907,N_22324);
nand U27713 (N_27713,N_21510,N_23323);
nor U27714 (N_27714,N_23294,N_20347);
nand U27715 (N_27715,N_23779,N_21632);
and U27716 (N_27716,N_22104,N_21474);
and U27717 (N_27717,N_22690,N_21466);
and U27718 (N_27718,N_22376,N_23913);
nor U27719 (N_27719,N_23675,N_23958);
xnor U27720 (N_27720,N_20563,N_20004);
nand U27721 (N_27721,N_24361,N_20040);
or U27722 (N_27722,N_23759,N_22740);
and U27723 (N_27723,N_23689,N_22476);
xnor U27724 (N_27724,N_20711,N_24686);
and U27725 (N_27725,N_22488,N_21685);
nand U27726 (N_27726,N_24718,N_20605);
or U27727 (N_27727,N_20546,N_22440);
nand U27728 (N_27728,N_24859,N_22709);
nor U27729 (N_27729,N_20453,N_22056);
nand U27730 (N_27730,N_20267,N_23602);
and U27731 (N_27731,N_24099,N_24491);
nor U27732 (N_27732,N_22300,N_24338);
and U27733 (N_27733,N_23939,N_23619);
and U27734 (N_27734,N_21281,N_23410);
nor U27735 (N_27735,N_23090,N_22365);
xor U27736 (N_27736,N_20194,N_21674);
or U27737 (N_27737,N_21828,N_20815);
xnor U27738 (N_27738,N_21464,N_21499);
xor U27739 (N_27739,N_23069,N_21117);
or U27740 (N_27740,N_21567,N_21248);
nor U27741 (N_27741,N_22277,N_23748);
nor U27742 (N_27742,N_22809,N_21616);
and U27743 (N_27743,N_22157,N_20865);
nand U27744 (N_27744,N_24140,N_21749);
and U27745 (N_27745,N_23164,N_20719);
or U27746 (N_27746,N_21703,N_23752);
and U27747 (N_27747,N_21657,N_23274);
nor U27748 (N_27748,N_23446,N_22478);
xnor U27749 (N_27749,N_24799,N_22785);
xnor U27750 (N_27750,N_24633,N_20841);
nand U27751 (N_27751,N_24879,N_24769);
nor U27752 (N_27752,N_24867,N_23340);
or U27753 (N_27753,N_24103,N_21404);
xor U27754 (N_27754,N_20105,N_23466);
xnor U27755 (N_27755,N_21452,N_22612);
nand U27756 (N_27756,N_24726,N_20676);
xnor U27757 (N_27757,N_24219,N_21409);
nand U27758 (N_27758,N_21254,N_24343);
nor U27759 (N_27759,N_21751,N_22831);
nand U27760 (N_27760,N_23248,N_23368);
xnor U27761 (N_27761,N_22099,N_21180);
nand U27762 (N_27762,N_21896,N_21592);
xnor U27763 (N_27763,N_24469,N_23289);
nand U27764 (N_27764,N_22395,N_23259);
or U27765 (N_27765,N_21390,N_21235);
nor U27766 (N_27766,N_23804,N_21915);
nor U27767 (N_27767,N_23791,N_20821);
and U27768 (N_27768,N_23502,N_23341);
nor U27769 (N_27769,N_24205,N_20806);
or U27770 (N_27770,N_23317,N_23649);
and U27771 (N_27771,N_24339,N_20746);
nor U27772 (N_27772,N_23604,N_23188);
and U27773 (N_27773,N_22148,N_23832);
nor U27774 (N_27774,N_21844,N_20843);
nand U27775 (N_27775,N_22496,N_24060);
nand U27776 (N_27776,N_21391,N_21779);
xor U27777 (N_27777,N_23041,N_22124);
nand U27778 (N_27778,N_20199,N_20158);
and U27779 (N_27779,N_21764,N_21549);
xnor U27780 (N_27780,N_21511,N_24311);
and U27781 (N_27781,N_22525,N_20137);
and U27782 (N_27782,N_24072,N_24107);
nor U27783 (N_27783,N_20222,N_23735);
nor U27784 (N_27784,N_21254,N_23153);
or U27785 (N_27785,N_20543,N_21494);
nor U27786 (N_27786,N_21828,N_24289);
nand U27787 (N_27787,N_20932,N_20276);
xor U27788 (N_27788,N_20251,N_21501);
or U27789 (N_27789,N_22777,N_23879);
nor U27790 (N_27790,N_24418,N_24775);
and U27791 (N_27791,N_24170,N_24240);
xor U27792 (N_27792,N_21706,N_22691);
nor U27793 (N_27793,N_24741,N_20849);
and U27794 (N_27794,N_21090,N_22824);
nor U27795 (N_27795,N_23210,N_24440);
and U27796 (N_27796,N_22549,N_24663);
and U27797 (N_27797,N_20601,N_23256);
nor U27798 (N_27798,N_24621,N_21296);
xnor U27799 (N_27799,N_20939,N_23791);
nor U27800 (N_27800,N_20843,N_22680);
or U27801 (N_27801,N_22518,N_24588);
and U27802 (N_27802,N_24152,N_23363);
or U27803 (N_27803,N_24191,N_24363);
xnor U27804 (N_27804,N_23433,N_20674);
or U27805 (N_27805,N_24960,N_22028);
xnor U27806 (N_27806,N_22984,N_24452);
xor U27807 (N_27807,N_21503,N_22272);
xor U27808 (N_27808,N_24460,N_23760);
xnor U27809 (N_27809,N_22280,N_21976);
nand U27810 (N_27810,N_24631,N_21659);
nor U27811 (N_27811,N_23151,N_23076);
and U27812 (N_27812,N_20290,N_21941);
or U27813 (N_27813,N_21371,N_21460);
xnor U27814 (N_27814,N_20796,N_24476);
or U27815 (N_27815,N_21093,N_24759);
nor U27816 (N_27816,N_21335,N_20815);
nand U27817 (N_27817,N_23800,N_23963);
nor U27818 (N_27818,N_24320,N_23885);
or U27819 (N_27819,N_24805,N_24744);
nand U27820 (N_27820,N_22512,N_24609);
nor U27821 (N_27821,N_24399,N_20319);
nand U27822 (N_27822,N_21703,N_21660);
xnor U27823 (N_27823,N_21852,N_24628);
nand U27824 (N_27824,N_22365,N_24591);
xor U27825 (N_27825,N_20083,N_23713);
nand U27826 (N_27826,N_21720,N_24582);
or U27827 (N_27827,N_20898,N_22093);
or U27828 (N_27828,N_22241,N_23427);
nand U27829 (N_27829,N_21033,N_24044);
and U27830 (N_27830,N_20273,N_20293);
nand U27831 (N_27831,N_20598,N_23981);
nor U27832 (N_27832,N_21023,N_23065);
xor U27833 (N_27833,N_23696,N_22046);
or U27834 (N_27834,N_22195,N_21269);
and U27835 (N_27835,N_21212,N_23779);
and U27836 (N_27836,N_24325,N_23865);
and U27837 (N_27837,N_21319,N_24447);
or U27838 (N_27838,N_22208,N_20797);
xor U27839 (N_27839,N_23170,N_22729);
xor U27840 (N_27840,N_23622,N_20513);
or U27841 (N_27841,N_20327,N_24297);
xnor U27842 (N_27842,N_20774,N_23389);
and U27843 (N_27843,N_23388,N_21512);
xor U27844 (N_27844,N_20183,N_21997);
xnor U27845 (N_27845,N_20268,N_24275);
nor U27846 (N_27846,N_24511,N_22600);
nand U27847 (N_27847,N_23020,N_23811);
and U27848 (N_27848,N_24781,N_23003);
and U27849 (N_27849,N_21827,N_22162);
nor U27850 (N_27850,N_21047,N_22827);
xor U27851 (N_27851,N_24597,N_21341);
nand U27852 (N_27852,N_22504,N_24885);
xnor U27853 (N_27853,N_21235,N_20408);
nor U27854 (N_27854,N_20454,N_22166);
xnor U27855 (N_27855,N_20750,N_22556);
and U27856 (N_27856,N_20825,N_23322);
nand U27857 (N_27857,N_22446,N_20501);
xor U27858 (N_27858,N_22759,N_23408);
nand U27859 (N_27859,N_20535,N_20689);
xnor U27860 (N_27860,N_23978,N_20813);
nor U27861 (N_27861,N_23501,N_22328);
nor U27862 (N_27862,N_22414,N_23036);
and U27863 (N_27863,N_22902,N_22753);
nand U27864 (N_27864,N_24318,N_23208);
nor U27865 (N_27865,N_22822,N_21969);
xnor U27866 (N_27866,N_21934,N_22041);
or U27867 (N_27867,N_23011,N_21877);
or U27868 (N_27868,N_24719,N_22654);
xor U27869 (N_27869,N_23476,N_21318);
or U27870 (N_27870,N_22786,N_20213);
or U27871 (N_27871,N_20577,N_22451);
nand U27872 (N_27872,N_23940,N_22432);
xnor U27873 (N_27873,N_21620,N_24005);
nor U27874 (N_27874,N_23741,N_22057);
or U27875 (N_27875,N_23238,N_23929);
xnor U27876 (N_27876,N_22003,N_21488);
nor U27877 (N_27877,N_21351,N_23352);
xor U27878 (N_27878,N_20422,N_22591);
xnor U27879 (N_27879,N_24903,N_22723);
xnor U27880 (N_27880,N_20296,N_20397);
nor U27881 (N_27881,N_20222,N_22593);
and U27882 (N_27882,N_20408,N_23140);
or U27883 (N_27883,N_22622,N_20632);
xnor U27884 (N_27884,N_20004,N_21720);
or U27885 (N_27885,N_21232,N_21287);
or U27886 (N_27886,N_23672,N_22029);
nand U27887 (N_27887,N_21549,N_23750);
nand U27888 (N_27888,N_24969,N_22212);
and U27889 (N_27889,N_21865,N_20731);
nor U27890 (N_27890,N_23519,N_24130);
nor U27891 (N_27891,N_24786,N_24510);
nor U27892 (N_27892,N_20624,N_24578);
or U27893 (N_27893,N_22395,N_21951);
or U27894 (N_27894,N_21343,N_20184);
nand U27895 (N_27895,N_22184,N_22846);
xor U27896 (N_27896,N_21642,N_24780);
nand U27897 (N_27897,N_23593,N_23948);
nand U27898 (N_27898,N_22705,N_20967);
or U27899 (N_27899,N_24598,N_22842);
nor U27900 (N_27900,N_23283,N_23605);
or U27901 (N_27901,N_24146,N_20972);
or U27902 (N_27902,N_22264,N_21546);
xor U27903 (N_27903,N_22850,N_20087);
nand U27904 (N_27904,N_21732,N_21629);
or U27905 (N_27905,N_24870,N_21336);
nand U27906 (N_27906,N_22521,N_21104);
xor U27907 (N_27907,N_23047,N_22787);
nor U27908 (N_27908,N_24319,N_20289);
xor U27909 (N_27909,N_20366,N_20018);
and U27910 (N_27910,N_21332,N_23035);
xor U27911 (N_27911,N_21933,N_20889);
xnor U27912 (N_27912,N_23490,N_21628);
nor U27913 (N_27913,N_21295,N_20156);
nand U27914 (N_27914,N_24885,N_20084);
xnor U27915 (N_27915,N_21412,N_20847);
or U27916 (N_27916,N_22592,N_23888);
nor U27917 (N_27917,N_24213,N_22890);
xnor U27918 (N_27918,N_20608,N_20854);
xor U27919 (N_27919,N_23807,N_22138);
and U27920 (N_27920,N_22374,N_20507);
nand U27921 (N_27921,N_20863,N_24322);
nand U27922 (N_27922,N_24422,N_24447);
nand U27923 (N_27923,N_22884,N_24345);
nor U27924 (N_27924,N_24237,N_23586);
xnor U27925 (N_27925,N_22505,N_24771);
nand U27926 (N_27926,N_24072,N_21850);
or U27927 (N_27927,N_21642,N_20256);
or U27928 (N_27928,N_23644,N_21946);
or U27929 (N_27929,N_23740,N_20706);
or U27930 (N_27930,N_23366,N_22256);
nand U27931 (N_27931,N_21524,N_21949);
and U27932 (N_27932,N_21303,N_22685);
and U27933 (N_27933,N_21624,N_23582);
and U27934 (N_27934,N_20210,N_24914);
nand U27935 (N_27935,N_24298,N_21729);
and U27936 (N_27936,N_22950,N_24864);
nand U27937 (N_27937,N_20332,N_23303);
nor U27938 (N_27938,N_24904,N_23693);
nor U27939 (N_27939,N_22855,N_23717);
nor U27940 (N_27940,N_24068,N_23425);
nor U27941 (N_27941,N_24350,N_21683);
or U27942 (N_27942,N_20927,N_20973);
xnor U27943 (N_27943,N_20690,N_20487);
xor U27944 (N_27944,N_21169,N_20699);
nand U27945 (N_27945,N_24203,N_22666);
and U27946 (N_27946,N_21663,N_21409);
nor U27947 (N_27947,N_24468,N_21442);
and U27948 (N_27948,N_23763,N_24081);
nand U27949 (N_27949,N_22397,N_21168);
xor U27950 (N_27950,N_22995,N_21112);
and U27951 (N_27951,N_24349,N_21250);
xor U27952 (N_27952,N_21445,N_23502);
nand U27953 (N_27953,N_22749,N_21938);
xor U27954 (N_27954,N_23171,N_24572);
and U27955 (N_27955,N_20576,N_24202);
nor U27956 (N_27956,N_21972,N_24639);
xnor U27957 (N_27957,N_20349,N_23707);
nand U27958 (N_27958,N_23576,N_24470);
nand U27959 (N_27959,N_22371,N_23957);
or U27960 (N_27960,N_22556,N_21469);
xor U27961 (N_27961,N_21389,N_24011);
xnor U27962 (N_27962,N_23219,N_21396);
nand U27963 (N_27963,N_24299,N_21407);
and U27964 (N_27964,N_21059,N_21842);
nor U27965 (N_27965,N_20698,N_20138);
nand U27966 (N_27966,N_23926,N_24628);
nor U27967 (N_27967,N_24567,N_22343);
and U27968 (N_27968,N_24879,N_20156);
nor U27969 (N_27969,N_24856,N_21330);
xnor U27970 (N_27970,N_20100,N_21155);
and U27971 (N_27971,N_22761,N_20438);
xnor U27972 (N_27972,N_22834,N_22670);
or U27973 (N_27973,N_24129,N_24939);
nand U27974 (N_27974,N_22081,N_21119);
nand U27975 (N_27975,N_22668,N_24055);
nor U27976 (N_27976,N_23965,N_22015);
and U27977 (N_27977,N_22724,N_20503);
or U27978 (N_27978,N_21988,N_22836);
or U27979 (N_27979,N_23388,N_24278);
nand U27980 (N_27980,N_22700,N_22617);
and U27981 (N_27981,N_21315,N_22691);
nor U27982 (N_27982,N_24876,N_23231);
xnor U27983 (N_27983,N_23759,N_23308);
nor U27984 (N_27984,N_21799,N_21457);
nand U27985 (N_27985,N_20577,N_23776);
and U27986 (N_27986,N_21625,N_21500);
nor U27987 (N_27987,N_24447,N_22052);
nand U27988 (N_27988,N_22554,N_22544);
xnor U27989 (N_27989,N_24536,N_23540);
and U27990 (N_27990,N_21078,N_22918);
and U27991 (N_27991,N_23796,N_20226);
nor U27992 (N_27992,N_21216,N_22358);
nor U27993 (N_27993,N_21044,N_20804);
xor U27994 (N_27994,N_22838,N_22346);
and U27995 (N_27995,N_20014,N_22883);
nand U27996 (N_27996,N_22006,N_22375);
and U27997 (N_27997,N_22752,N_22095);
and U27998 (N_27998,N_22243,N_24954);
or U27999 (N_27999,N_22905,N_24598);
nor U28000 (N_28000,N_20408,N_20965);
nor U28001 (N_28001,N_21643,N_22825);
nor U28002 (N_28002,N_21594,N_23479);
and U28003 (N_28003,N_24586,N_24308);
nor U28004 (N_28004,N_21377,N_21506);
and U28005 (N_28005,N_21925,N_23551);
nor U28006 (N_28006,N_24208,N_24313);
and U28007 (N_28007,N_20751,N_22170);
nor U28008 (N_28008,N_21283,N_24546);
nor U28009 (N_28009,N_24778,N_22563);
and U28010 (N_28010,N_24861,N_23797);
xor U28011 (N_28011,N_22353,N_24608);
nand U28012 (N_28012,N_22852,N_22675);
xor U28013 (N_28013,N_21527,N_23015);
xnor U28014 (N_28014,N_21522,N_20148);
nand U28015 (N_28015,N_20310,N_22025);
and U28016 (N_28016,N_24768,N_20113);
or U28017 (N_28017,N_22802,N_23010);
xor U28018 (N_28018,N_23990,N_20514);
xor U28019 (N_28019,N_24705,N_24633);
and U28020 (N_28020,N_20666,N_22951);
nor U28021 (N_28021,N_21981,N_24250);
nand U28022 (N_28022,N_22713,N_22866);
and U28023 (N_28023,N_24859,N_24105);
and U28024 (N_28024,N_23558,N_24194);
nand U28025 (N_28025,N_23132,N_21990);
xor U28026 (N_28026,N_22596,N_20754);
xor U28027 (N_28027,N_20903,N_21152);
nand U28028 (N_28028,N_21443,N_23453);
or U28029 (N_28029,N_20946,N_21200);
nand U28030 (N_28030,N_24033,N_21035);
xnor U28031 (N_28031,N_24711,N_20986);
nand U28032 (N_28032,N_23164,N_21000);
nand U28033 (N_28033,N_21215,N_21668);
nand U28034 (N_28034,N_20036,N_23799);
or U28035 (N_28035,N_20863,N_23960);
xor U28036 (N_28036,N_22548,N_24769);
and U28037 (N_28037,N_23032,N_21723);
nor U28038 (N_28038,N_21492,N_24524);
and U28039 (N_28039,N_24191,N_20029);
and U28040 (N_28040,N_23585,N_22679);
or U28041 (N_28041,N_21859,N_23167);
or U28042 (N_28042,N_21521,N_20523);
and U28043 (N_28043,N_21539,N_20025);
or U28044 (N_28044,N_22542,N_20336);
nor U28045 (N_28045,N_23975,N_24513);
or U28046 (N_28046,N_21665,N_20075);
nand U28047 (N_28047,N_21807,N_21888);
or U28048 (N_28048,N_24658,N_20556);
nor U28049 (N_28049,N_24609,N_24472);
or U28050 (N_28050,N_20442,N_24979);
nand U28051 (N_28051,N_24036,N_23814);
xor U28052 (N_28052,N_22356,N_24372);
and U28053 (N_28053,N_23527,N_20478);
xnor U28054 (N_28054,N_21962,N_22894);
nand U28055 (N_28055,N_22118,N_23870);
xor U28056 (N_28056,N_24307,N_21462);
and U28057 (N_28057,N_24474,N_21902);
nor U28058 (N_28058,N_20126,N_24681);
and U28059 (N_28059,N_20524,N_22941);
or U28060 (N_28060,N_23624,N_22304);
xnor U28061 (N_28061,N_21928,N_22072);
and U28062 (N_28062,N_20228,N_21043);
nand U28063 (N_28063,N_23057,N_24651);
or U28064 (N_28064,N_22359,N_24035);
nand U28065 (N_28065,N_24672,N_21678);
nor U28066 (N_28066,N_21919,N_24713);
xor U28067 (N_28067,N_20482,N_20305);
xnor U28068 (N_28068,N_21152,N_24617);
nor U28069 (N_28069,N_23636,N_21035);
nand U28070 (N_28070,N_23743,N_22731);
xnor U28071 (N_28071,N_20863,N_20438);
xor U28072 (N_28072,N_24813,N_21456);
and U28073 (N_28073,N_20024,N_23072);
and U28074 (N_28074,N_21453,N_22606);
and U28075 (N_28075,N_22394,N_20689);
and U28076 (N_28076,N_22985,N_22916);
nand U28077 (N_28077,N_20258,N_24207);
or U28078 (N_28078,N_22577,N_21084);
xnor U28079 (N_28079,N_20093,N_21136);
or U28080 (N_28080,N_22105,N_24797);
nor U28081 (N_28081,N_24463,N_22679);
or U28082 (N_28082,N_23684,N_21495);
nand U28083 (N_28083,N_24498,N_21739);
nor U28084 (N_28084,N_24340,N_20207);
nor U28085 (N_28085,N_21662,N_20172);
or U28086 (N_28086,N_21969,N_20826);
and U28087 (N_28087,N_21712,N_20957);
xnor U28088 (N_28088,N_22834,N_21830);
nor U28089 (N_28089,N_22789,N_24336);
xor U28090 (N_28090,N_20979,N_22254);
nand U28091 (N_28091,N_20993,N_22820);
or U28092 (N_28092,N_23554,N_21336);
nor U28093 (N_28093,N_21701,N_20736);
xnor U28094 (N_28094,N_22487,N_24811);
or U28095 (N_28095,N_24650,N_21676);
xor U28096 (N_28096,N_21460,N_20636);
nand U28097 (N_28097,N_24173,N_23103);
and U28098 (N_28098,N_23007,N_23860);
nor U28099 (N_28099,N_21474,N_24217);
and U28100 (N_28100,N_21707,N_21994);
or U28101 (N_28101,N_23918,N_20051);
nand U28102 (N_28102,N_22265,N_20610);
nand U28103 (N_28103,N_21505,N_23404);
xnor U28104 (N_28104,N_22809,N_21581);
and U28105 (N_28105,N_21429,N_22874);
nand U28106 (N_28106,N_22050,N_23967);
nand U28107 (N_28107,N_21482,N_20746);
nor U28108 (N_28108,N_21424,N_21466);
xor U28109 (N_28109,N_22552,N_20849);
xor U28110 (N_28110,N_20064,N_24751);
and U28111 (N_28111,N_22872,N_24101);
and U28112 (N_28112,N_21834,N_20737);
nand U28113 (N_28113,N_20521,N_24928);
and U28114 (N_28114,N_24436,N_20665);
nor U28115 (N_28115,N_23668,N_23502);
xnor U28116 (N_28116,N_23926,N_23020);
and U28117 (N_28117,N_22657,N_20354);
xnor U28118 (N_28118,N_22133,N_22201);
nand U28119 (N_28119,N_22299,N_23114);
nand U28120 (N_28120,N_24022,N_21152);
nand U28121 (N_28121,N_21799,N_23506);
xor U28122 (N_28122,N_23810,N_22989);
nor U28123 (N_28123,N_23452,N_24910);
or U28124 (N_28124,N_24112,N_21049);
nor U28125 (N_28125,N_20054,N_20636);
xor U28126 (N_28126,N_21780,N_22015);
nand U28127 (N_28127,N_20114,N_23985);
nand U28128 (N_28128,N_21365,N_24474);
or U28129 (N_28129,N_20290,N_23737);
xnor U28130 (N_28130,N_20973,N_23571);
xor U28131 (N_28131,N_20311,N_24061);
nand U28132 (N_28132,N_24583,N_23616);
nor U28133 (N_28133,N_20228,N_23499);
nand U28134 (N_28134,N_21231,N_23532);
nor U28135 (N_28135,N_20002,N_20886);
nor U28136 (N_28136,N_23377,N_21689);
nand U28137 (N_28137,N_21245,N_22159);
or U28138 (N_28138,N_20167,N_24985);
or U28139 (N_28139,N_20207,N_23792);
xor U28140 (N_28140,N_24687,N_21513);
nor U28141 (N_28141,N_20596,N_23461);
or U28142 (N_28142,N_23832,N_24076);
xor U28143 (N_28143,N_24633,N_24645);
or U28144 (N_28144,N_20696,N_21584);
nor U28145 (N_28145,N_22651,N_21886);
and U28146 (N_28146,N_23682,N_21123);
nor U28147 (N_28147,N_20040,N_20609);
xor U28148 (N_28148,N_21559,N_23203);
xnor U28149 (N_28149,N_24669,N_21789);
or U28150 (N_28150,N_23155,N_24737);
or U28151 (N_28151,N_22143,N_20475);
xnor U28152 (N_28152,N_23011,N_20765);
or U28153 (N_28153,N_20128,N_22643);
nand U28154 (N_28154,N_20349,N_21969);
nor U28155 (N_28155,N_22868,N_21956);
or U28156 (N_28156,N_23935,N_20754);
nor U28157 (N_28157,N_22528,N_24134);
or U28158 (N_28158,N_23657,N_20852);
or U28159 (N_28159,N_21938,N_20803);
xor U28160 (N_28160,N_23716,N_22928);
nand U28161 (N_28161,N_23290,N_20552);
nor U28162 (N_28162,N_24305,N_24800);
xor U28163 (N_28163,N_22704,N_24030);
xnor U28164 (N_28164,N_23291,N_22634);
nand U28165 (N_28165,N_24329,N_23426);
nand U28166 (N_28166,N_21627,N_22042);
nor U28167 (N_28167,N_20057,N_24340);
xnor U28168 (N_28168,N_22293,N_23289);
nor U28169 (N_28169,N_24380,N_21278);
nand U28170 (N_28170,N_21659,N_23425);
or U28171 (N_28171,N_22749,N_20094);
and U28172 (N_28172,N_23346,N_22292);
nor U28173 (N_28173,N_20451,N_20448);
nand U28174 (N_28174,N_23272,N_21818);
and U28175 (N_28175,N_24139,N_23489);
nor U28176 (N_28176,N_20367,N_23883);
or U28177 (N_28177,N_22958,N_23675);
nand U28178 (N_28178,N_20634,N_22113);
nand U28179 (N_28179,N_22190,N_23096);
xnor U28180 (N_28180,N_23549,N_20254);
nand U28181 (N_28181,N_22611,N_23877);
nor U28182 (N_28182,N_23313,N_24533);
nand U28183 (N_28183,N_24323,N_21223);
nor U28184 (N_28184,N_20186,N_22608);
or U28185 (N_28185,N_24788,N_23065);
xnor U28186 (N_28186,N_20488,N_23248);
xnor U28187 (N_28187,N_21405,N_23591);
xor U28188 (N_28188,N_22215,N_20568);
xnor U28189 (N_28189,N_22705,N_20381);
nand U28190 (N_28190,N_23442,N_21401);
nor U28191 (N_28191,N_21624,N_20866);
xor U28192 (N_28192,N_23954,N_23496);
xnor U28193 (N_28193,N_22352,N_22730);
and U28194 (N_28194,N_20645,N_21697);
or U28195 (N_28195,N_23605,N_22571);
or U28196 (N_28196,N_23166,N_20802);
nand U28197 (N_28197,N_20931,N_22674);
and U28198 (N_28198,N_20339,N_21508);
nand U28199 (N_28199,N_24766,N_21389);
or U28200 (N_28200,N_20803,N_23254);
xnor U28201 (N_28201,N_21204,N_23176);
and U28202 (N_28202,N_24151,N_22422);
nand U28203 (N_28203,N_24909,N_20085);
xnor U28204 (N_28204,N_24795,N_21884);
nand U28205 (N_28205,N_22719,N_22814);
nor U28206 (N_28206,N_22103,N_20425);
and U28207 (N_28207,N_21625,N_22200);
nand U28208 (N_28208,N_20771,N_22511);
nor U28209 (N_28209,N_24215,N_22483);
xnor U28210 (N_28210,N_23725,N_20181);
xnor U28211 (N_28211,N_23616,N_21070);
and U28212 (N_28212,N_22254,N_21242);
nor U28213 (N_28213,N_24845,N_23576);
xnor U28214 (N_28214,N_22931,N_21089);
xnor U28215 (N_28215,N_24393,N_21979);
nand U28216 (N_28216,N_21853,N_20576);
xnor U28217 (N_28217,N_22479,N_23104);
nand U28218 (N_28218,N_24245,N_20908);
and U28219 (N_28219,N_23070,N_21237);
and U28220 (N_28220,N_22458,N_23781);
and U28221 (N_28221,N_23017,N_21458);
nand U28222 (N_28222,N_23028,N_24623);
and U28223 (N_28223,N_21164,N_20044);
xnor U28224 (N_28224,N_21535,N_23126);
nor U28225 (N_28225,N_23756,N_20749);
xnor U28226 (N_28226,N_20959,N_20895);
nand U28227 (N_28227,N_22761,N_24429);
xnor U28228 (N_28228,N_22876,N_21662);
xor U28229 (N_28229,N_21271,N_23037);
or U28230 (N_28230,N_23000,N_20353);
nor U28231 (N_28231,N_22232,N_22513);
and U28232 (N_28232,N_21422,N_20239);
nand U28233 (N_28233,N_21978,N_23996);
xor U28234 (N_28234,N_22087,N_21386);
and U28235 (N_28235,N_22082,N_22213);
and U28236 (N_28236,N_22295,N_23176);
and U28237 (N_28237,N_20957,N_22923);
and U28238 (N_28238,N_20104,N_24206);
nor U28239 (N_28239,N_23286,N_23692);
nor U28240 (N_28240,N_20832,N_23547);
or U28241 (N_28241,N_24951,N_21855);
and U28242 (N_28242,N_20929,N_22272);
nor U28243 (N_28243,N_21817,N_24132);
nor U28244 (N_28244,N_23275,N_20526);
xnor U28245 (N_28245,N_20972,N_24689);
nand U28246 (N_28246,N_20338,N_22649);
nor U28247 (N_28247,N_23750,N_21304);
nand U28248 (N_28248,N_23619,N_21665);
nor U28249 (N_28249,N_23849,N_21574);
xor U28250 (N_28250,N_24137,N_21154);
nor U28251 (N_28251,N_20166,N_21746);
xnor U28252 (N_28252,N_20543,N_22998);
nor U28253 (N_28253,N_20333,N_21403);
nand U28254 (N_28254,N_20627,N_21523);
and U28255 (N_28255,N_20431,N_23127);
or U28256 (N_28256,N_20657,N_22639);
or U28257 (N_28257,N_22430,N_23309);
or U28258 (N_28258,N_21020,N_22156);
and U28259 (N_28259,N_24450,N_21591);
nand U28260 (N_28260,N_21635,N_23961);
nor U28261 (N_28261,N_20013,N_23986);
or U28262 (N_28262,N_22153,N_21890);
and U28263 (N_28263,N_21749,N_20993);
or U28264 (N_28264,N_21064,N_22228);
nand U28265 (N_28265,N_21844,N_23403);
and U28266 (N_28266,N_24392,N_24479);
or U28267 (N_28267,N_20155,N_20818);
nor U28268 (N_28268,N_23969,N_20825);
nand U28269 (N_28269,N_20390,N_20249);
nor U28270 (N_28270,N_20272,N_20774);
nand U28271 (N_28271,N_22176,N_20589);
nor U28272 (N_28272,N_24580,N_22060);
or U28273 (N_28273,N_21654,N_21277);
or U28274 (N_28274,N_20833,N_23077);
and U28275 (N_28275,N_20465,N_21733);
and U28276 (N_28276,N_20019,N_21853);
nor U28277 (N_28277,N_22307,N_24975);
xnor U28278 (N_28278,N_23873,N_22176);
or U28279 (N_28279,N_21043,N_21665);
and U28280 (N_28280,N_21483,N_23754);
nor U28281 (N_28281,N_23308,N_20667);
or U28282 (N_28282,N_23354,N_20034);
nand U28283 (N_28283,N_21363,N_21012);
and U28284 (N_28284,N_21977,N_22579);
nand U28285 (N_28285,N_21071,N_24808);
and U28286 (N_28286,N_23572,N_20262);
or U28287 (N_28287,N_20401,N_21175);
or U28288 (N_28288,N_22213,N_21630);
xor U28289 (N_28289,N_23780,N_23225);
or U28290 (N_28290,N_23366,N_20721);
nand U28291 (N_28291,N_20238,N_21765);
xnor U28292 (N_28292,N_22503,N_24247);
xnor U28293 (N_28293,N_21933,N_20597);
and U28294 (N_28294,N_21909,N_23541);
or U28295 (N_28295,N_22245,N_22097);
xnor U28296 (N_28296,N_20226,N_21087);
nor U28297 (N_28297,N_20843,N_24686);
nand U28298 (N_28298,N_23868,N_20746);
nor U28299 (N_28299,N_23832,N_24244);
and U28300 (N_28300,N_21884,N_21529);
nor U28301 (N_28301,N_20134,N_20769);
xnor U28302 (N_28302,N_21311,N_20080);
nor U28303 (N_28303,N_21779,N_21301);
nor U28304 (N_28304,N_21397,N_24370);
xor U28305 (N_28305,N_22876,N_20209);
xnor U28306 (N_28306,N_24716,N_22418);
or U28307 (N_28307,N_21736,N_22217);
or U28308 (N_28308,N_20445,N_24761);
and U28309 (N_28309,N_23969,N_22389);
or U28310 (N_28310,N_22717,N_23546);
or U28311 (N_28311,N_20635,N_22351);
nor U28312 (N_28312,N_24975,N_21692);
nor U28313 (N_28313,N_23840,N_23590);
xor U28314 (N_28314,N_22598,N_20364);
xnor U28315 (N_28315,N_21827,N_24849);
and U28316 (N_28316,N_24573,N_21526);
nor U28317 (N_28317,N_21576,N_24872);
xor U28318 (N_28318,N_21712,N_23043);
nor U28319 (N_28319,N_21532,N_24602);
nor U28320 (N_28320,N_23590,N_20241);
xnor U28321 (N_28321,N_20826,N_24738);
nand U28322 (N_28322,N_23761,N_22253);
xnor U28323 (N_28323,N_22531,N_21537);
or U28324 (N_28324,N_22721,N_21591);
nor U28325 (N_28325,N_22523,N_23175);
xor U28326 (N_28326,N_20828,N_24631);
or U28327 (N_28327,N_21696,N_24044);
nor U28328 (N_28328,N_24061,N_23718);
or U28329 (N_28329,N_24656,N_24467);
and U28330 (N_28330,N_20338,N_23988);
and U28331 (N_28331,N_23886,N_22076);
nor U28332 (N_28332,N_22459,N_21488);
xor U28333 (N_28333,N_21360,N_22450);
and U28334 (N_28334,N_24780,N_24976);
and U28335 (N_28335,N_20572,N_22892);
or U28336 (N_28336,N_24776,N_21087);
nor U28337 (N_28337,N_21674,N_23775);
nor U28338 (N_28338,N_20868,N_22553);
and U28339 (N_28339,N_24440,N_20921);
or U28340 (N_28340,N_24688,N_23966);
nor U28341 (N_28341,N_23897,N_23112);
nand U28342 (N_28342,N_20655,N_24855);
xnor U28343 (N_28343,N_22896,N_23163);
xnor U28344 (N_28344,N_21404,N_21660);
xor U28345 (N_28345,N_24828,N_23902);
and U28346 (N_28346,N_23677,N_24943);
nand U28347 (N_28347,N_21628,N_21663);
and U28348 (N_28348,N_23229,N_23179);
nand U28349 (N_28349,N_20331,N_20125);
xnor U28350 (N_28350,N_23849,N_23075);
nand U28351 (N_28351,N_24704,N_23882);
nor U28352 (N_28352,N_23757,N_21625);
or U28353 (N_28353,N_22328,N_23891);
or U28354 (N_28354,N_20513,N_22107);
xnor U28355 (N_28355,N_20266,N_22474);
nor U28356 (N_28356,N_24045,N_22719);
or U28357 (N_28357,N_20100,N_23790);
or U28358 (N_28358,N_22421,N_22869);
nor U28359 (N_28359,N_24577,N_21358);
or U28360 (N_28360,N_22482,N_20668);
nor U28361 (N_28361,N_23362,N_21001);
or U28362 (N_28362,N_24590,N_21566);
xor U28363 (N_28363,N_22940,N_21016);
or U28364 (N_28364,N_23468,N_21479);
nand U28365 (N_28365,N_24582,N_21327);
and U28366 (N_28366,N_22402,N_24696);
or U28367 (N_28367,N_20235,N_22293);
nor U28368 (N_28368,N_23482,N_22542);
or U28369 (N_28369,N_22541,N_22091);
nand U28370 (N_28370,N_22105,N_24342);
and U28371 (N_28371,N_20691,N_24166);
and U28372 (N_28372,N_22736,N_24768);
and U28373 (N_28373,N_24982,N_21569);
xor U28374 (N_28374,N_24858,N_23315);
and U28375 (N_28375,N_24767,N_24148);
nor U28376 (N_28376,N_22947,N_20338);
xor U28377 (N_28377,N_21346,N_23592);
nand U28378 (N_28378,N_23739,N_23194);
xnor U28379 (N_28379,N_21332,N_21996);
nor U28380 (N_28380,N_20967,N_20398);
nor U28381 (N_28381,N_24715,N_24034);
nand U28382 (N_28382,N_24461,N_20043);
nand U28383 (N_28383,N_21042,N_22220);
nand U28384 (N_28384,N_20627,N_23251);
xnor U28385 (N_28385,N_22742,N_24285);
xnor U28386 (N_28386,N_20823,N_20666);
or U28387 (N_28387,N_21083,N_23576);
and U28388 (N_28388,N_22717,N_23756);
or U28389 (N_28389,N_22523,N_24911);
and U28390 (N_28390,N_20165,N_20892);
or U28391 (N_28391,N_24311,N_23801);
nand U28392 (N_28392,N_23613,N_21180);
or U28393 (N_28393,N_21924,N_20634);
xor U28394 (N_28394,N_21877,N_20862);
and U28395 (N_28395,N_24860,N_23836);
nand U28396 (N_28396,N_23748,N_21722);
xor U28397 (N_28397,N_22626,N_24928);
nand U28398 (N_28398,N_23334,N_22037);
nor U28399 (N_28399,N_24199,N_22035);
or U28400 (N_28400,N_20720,N_21824);
and U28401 (N_28401,N_20474,N_21095);
and U28402 (N_28402,N_20157,N_24804);
and U28403 (N_28403,N_23410,N_24385);
and U28404 (N_28404,N_24085,N_21583);
and U28405 (N_28405,N_24865,N_22712);
nor U28406 (N_28406,N_23790,N_23897);
and U28407 (N_28407,N_21883,N_20919);
nor U28408 (N_28408,N_23792,N_24752);
or U28409 (N_28409,N_24452,N_20860);
nor U28410 (N_28410,N_20876,N_21290);
xor U28411 (N_28411,N_22844,N_20475);
nand U28412 (N_28412,N_21144,N_22563);
nor U28413 (N_28413,N_20620,N_23646);
and U28414 (N_28414,N_24916,N_23330);
xor U28415 (N_28415,N_22826,N_20974);
or U28416 (N_28416,N_23150,N_24136);
nor U28417 (N_28417,N_20703,N_21488);
or U28418 (N_28418,N_23430,N_21677);
nor U28419 (N_28419,N_24425,N_20673);
and U28420 (N_28420,N_20687,N_23364);
xor U28421 (N_28421,N_23072,N_20716);
or U28422 (N_28422,N_21804,N_23522);
nand U28423 (N_28423,N_20531,N_20808);
or U28424 (N_28424,N_23609,N_22962);
nand U28425 (N_28425,N_20127,N_22216);
nand U28426 (N_28426,N_23596,N_21659);
nor U28427 (N_28427,N_22251,N_21678);
and U28428 (N_28428,N_20228,N_21172);
xnor U28429 (N_28429,N_23789,N_23450);
and U28430 (N_28430,N_24695,N_20187);
and U28431 (N_28431,N_24284,N_22101);
nor U28432 (N_28432,N_23849,N_24616);
xnor U28433 (N_28433,N_20599,N_23444);
nand U28434 (N_28434,N_22077,N_20429);
or U28435 (N_28435,N_21062,N_23459);
nand U28436 (N_28436,N_20672,N_20490);
nand U28437 (N_28437,N_24922,N_24923);
nor U28438 (N_28438,N_24855,N_20803);
nor U28439 (N_28439,N_21402,N_21489);
nand U28440 (N_28440,N_24103,N_22363);
or U28441 (N_28441,N_20150,N_22407);
and U28442 (N_28442,N_23053,N_20258);
xor U28443 (N_28443,N_23711,N_23094);
xnor U28444 (N_28444,N_24585,N_20549);
nand U28445 (N_28445,N_24583,N_22386);
nor U28446 (N_28446,N_20383,N_22091);
nor U28447 (N_28447,N_20202,N_21888);
and U28448 (N_28448,N_23741,N_20192);
nor U28449 (N_28449,N_23455,N_22708);
nor U28450 (N_28450,N_24620,N_21215);
nand U28451 (N_28451,N_21404,N_22031);
and U28452 (N_28452,N_21145,N_21859);
and U28453 (N_28453,N_23856,N_22779);
nand U28454 (N_28454,N_21563,N_24659);
or U28455 (N_28455,N_24760,N_21835);
or U28456 (N_28456,N_22780,N_24278);
nor U28457 (N_28457,N_21723,N_24221);
and U28458 (N_28458,N_24074,N_24598);
xnor U28459 (N_28459,N_24258,N_23941);
xnor U28460 (N_28460,N_20571,N_22374);
and U28461 (N_28461,N_23091,N_22187);
or U28462 (N_28462,N_23864,N_23741);
and U28463 (N_28463,N_21774,N_20426);
or U28464 (N_28464,N_20733,N_20963);
nor U28465 (N_28465,N_21004,N_21164);
xnor U28466 (N_28466,N_20617,N_24384);
and U28467 (N_28467,N_24282,N_23712);
and U28468 (N_28468,N_24012,N_22010);
or U28469 (N_28469,N_22150,N_24611);
and U28470 (N_28470,N_24526,N_24844);
or U28471 (N_28471,N_24775,N_22638);
xor U28472 (N_28472,N_20185,N_20346);
nand U28473 (N_28473,N_20060,N_24820);
and U28474 (N_28474,N_22735,N_20818);
nand U28475 (N_28475,N_23152,N_21779);
or U28476 (N_28476,N_23022,N_22649);
nor U28477 (N_28477,N_20884,N_21356);
nor U28478 (N_28478,N_24723,N_24150);
nor U28479 (N_28479,N_22060,N_23617);
and U28480 (N_28480,N_20817,N_22420);
nor U28481 (N_28481,N_20350,N_23089);
xor U28482 (N_28482,N_23738,N_23788);
and U28483 (N_28483,N_22818,N_20962);
xor U28484 (N_28484,N_24689,N_23491);
nand U28485 (N_28485,N_23495,N_21230);
and U28486 (N_28486,N_21944,N_23825);
nor U28487 (N_28487,N_24710,N_24081);
nor U28488 (N_28488,N_24538,N_23123);
xnor U28489 (N_28489,N_24602,N_20439);
nand U28490 (N_28490,N_24463,N_24046);
and U28491 (N_28491,N_24416,N_22763);
or U28492 (N_28492,N_22068,N_23214);
xnor U28493 (N_28493,N_21630,N_22746);
nand U28494 (N_28494,N_23177,N_23934);
xor U28495 (N_28495,N_23979,N_24057);
or U28496 (N_28496,N_23425,N_20769);
or U28497 (N_28497,N_21461,N_21215);
nor U28498 (N_28498,N_23426,N_24571);
nor U28499 (N_28499,N_24079,N_22042);
or U28500 (N_28500,N_22770,N_23647);
and U28501 (N_28501,N_22410,N_22924);
nand U28502 (N_28502,N_23645,N_21247);
nor U28503 (N_28503,N_22267,N_24505);
nand U28504 (N_28504,N_20975,N_23439);
xnor U28505 (N_28505,N_22822,N_20099);
nor U28506 (N_28506,N_22075,N_22015);
and U28507 (N_28507,N_20970,N_23293);
or U28508 (N_28508,N_23026,N_24028);
and U28509 (N_28509,N_23336,N_23575);
xnor U28510 (N_28510,N_24381,N_21545);
nand U28511 (N_28511,N_22547,N_20639);
and U28512 (N_28512,N_22614,N_23423);
nor U28513 (N_28513,N_21021,N_20881);
xor U28514 (N_28514,N_22780,N_23324);
xor U28515 (N_28515,N_21900,N_21137);
xor U28516 (N_28516,N_23953,N_23873);
nand U28517 (N_28517,N_22576,N_22772);
xor U28518 (N_28518,N_21961,N_20240);
nand U28519 (N_28519,N_23514,N_24920);
and U28520 (N_28520,N_21048,N_21265);
nor U28521 (N_28521,N_22960,N_20970);
or U28522 (N_28522,N_23439,N_20772);
nand U28523 (N_28523,N_20613,N_24600);
nor U28524 (N_28524,N_23674,N_24805);
xor U28525 (N_28525,N_21708,N_20568);
or U28526 (N_28526,N_23365,N_21027);
nand U28527 (N_28527,N_21974,N_22990);
or U28528 (N_28528,N_22619,N_24217);
xnor U28529 (N_28529,N_21924,N_23226);
nor U28530 (N_28530,N_24338,N_21540);
nor U28531 (N_28531,N_20063,N_21712);
and U28532 (N_28532,N_23070,N_24905);
and U28533 (N_28533,N_23536,N_21410);
nor U28534 (N_28534,N_21916,N_23730);
or U28535 (N_28535,N_24784,N_24218);
xor U28536 (N_28536,N_21430,N_24369);
xor U28537 (N_28537,N_23258,N_20384);
nor U28538 (N_28538,N_23885,N_22972);
or U28539 (N_28539,N_20231,N_20388);
nand U28540 (N_28540,N_23747,N_22739);
xnor U28541 (N_28541,N_24317,N_21182);
nor U28542 (N_28542,N_24643,N_22681);
or U28543 (N_28543,N_23126,N_21382);
nand U28544 (N_28544,N_22170,N_20727);
xor U28545 (N_28545,N_21658,N_20679);
xor U28546 (N_28546,N_22310,N_23420);
xnor U28547 (N_28547,N_21854,N_23320);
and U28548 (N_28548,N_21210,N_24179);
and U28549 (N_28549,N_22531,N_20175);
nand U28550 (N_28550,N_20602,N_22701);
xnor U28551 (N_28551,N_23878,N_20412);
or U28552 (N_28552,N_22801,N_20655);
or U28553 (N_28553,N_21502,N_24948);
xor U28554 (N_28554,N_23222,N_23469);
xnor U28555 (N_28555,N_23224,N_20009);
nand U28556 (N_28556,N_20736,N_24700);
nand U28557 (N_28557,N_24282,N_20811);
xnor U28558 (N_28558,N_23236,N_21008);
or U28559 (N_28559,N_20384,N_21529);
xnor U28560 (N_28560,N_20917,N_22439);
and U28561 (N_28561,N_24342,N_23126);
or U28562 (N_28562,N_22016,N_22738);
nor U28563 (N_28563,N_22079,N_21876);
nand U28564 (N_28564,N_22911,N_22660);
nand U28565 (N_28565,N_22008,N_22237);
or U28566 (N_28566,N_22056,N_22666);
or U28567 (N_28567,N_23959,N_23106);
or U28568 (N_28568,N_21158,N_20139);
xor U28569 (N_28569,N_20116,N_24953);
nor U28570 (N_28570,N_23146,N_22555);
and U28571 (N_28571,N_20041,N_21486);
and U28572 (N_28572,N_24914,N_20050);
or U28573 (N_28573,N_21435,N_24023);
nor U28574 (N_28574,N_22240,N_21651);
nand U28575 (N_28575,N_21443,N_22605);
nand U28576 (N_28576,N_22953,N_20013);
nor U28577 (N_28577,N_24372,N_23191);
nor U28578 (N_28578,N_22837,N_22362);
or U28579 (N_28579,N_21196,N_20127);
xnor U28580 (N_28580,N_24327,N_24186);
and U28581 (N_28581,N_21452,N_23152);
or U28582 (N_28582,N_23870,N_22412);
nand U28583 (N_28583,N_24549,N_20089);
xnor U28584 (N_28584,N_20117,N_20917);
xor U28585 (N_28585,N_21681,N_22848);
nor U28586 (N_28586,N_21628,N_23790);
xor U28587 (N_28587,N_22477,N_21064);
or U28588 (N_28588,N_21416,N_24292);
nor U28589 (N_28589,N_20231,N_20210);
nor U28590 (N_28590,N_20707,N_21151);
and U28591 (N_28591,N_20869,N_24215);
and U28592 (N_28592,N_21074,N_20388);
nand U28593 (N_28593,N_20002,N_21457);
xor U28594 (N_28594,N_20722,N_24530);
and U28595 (N_28595,N_22185,N_21544);
nor U28596 (N_28596,N_20338,N_23304);
nor U28597 (N_28597,N_22279,N_20064);
nand U28598 (N_28598,N_21205,N_21691);
nand U28599 (N_28599,N_22435,N_20693);
or U28600 (N_28600,N_24077,N_22307);
or U28601 (N_28601,N_22172,N_23114);
xnor U28602 (N_28602,N_22746,N_21977);
and U28603 (N_28603,N_22958,N_22266);
nor U28604 (N_28604,N_21910,N_22856);
xnor U28605 (N_28605,N_24902,N_22670);
or U28606 (N_28606,N_21009,N_23317);
or U28607 (N_28607,N_21735,N_21191);
or U28608 (N_28608,N_22065,N_20141);
nand U28609 (N_28609,N_22911,N_23909);
and U28610 (N_28610,N_22849,N_22469);
nand U28611 (N_28611,N_21970,N_22894);
and U28612 (N_28612,N_20133,N_24672);
and U28613 (N_28613,N_24363,N_24485);
nor U28614 (N_28614,N_20768,N_23725);
or U28615 (N_28615,N_22800,N_24261);
nand U28616 (N_28616,N_23549,N_22639);
and U28617 (N_28617,N_20420,N_20997);
xnor U28618 (N_28618,N_20698,N_20728);
nor U28619 (N_28619,N_21837,N_24122);
and U28620 (N_28620,N_20681,N_20976);
nand U28621 (N_28621,N_22313,N_21503);
nor U28622 (N_28622,N_24824,N_21915);
and U28623 (N_28623,N_23015,N_21948);
nor U28624 (N_28624,N_22150,N_24830);
nor U28625 (N_28625,N_21190,N_24634);
nor U28626 (N_28626,N_20896,N_24083);
or U28627 (N_28627,N_21558,N_24294);
and U28628 (N_28628,N_21004,N_21897);
or U28629 (N_28629,N_23612,N_23427);
or U28630 (N_28630,N_23415,N_22039);
or U28631 (N_28631,N_21121,N_20763);
xnor U28632 (N_28632,N_21833,N_23635);
nor U28633 (N_28633,N_21686,N_23186);
or U28634 (N_28634,N_22531,N_20188);
and U28635 (N_28635,N_20305,N_20771);
nor U28636 (N_28636,N_23813,N_23852);
nor U28637 (N_28637,N_21210,N_23568);
or U28638 (N_28638,N_21083,N_20813);
nor U28639 (N_28639,N_24002,N_23491);
xnor U28640 (N_28640,N_23190,N_22432);
xnor U28641 (N_28641,N_22378,N_22316);
xor U28642 (N_28642,N_20317,N_21512);
nand U28643 (N_28643,N_22893,N_24576);
xor U28644 (N_28644,N_24187,N_23832);
nand U28645 (N_28645,N_20830,N_23084);
nand U28646 (N_28646,N_21035,N_20941);
or U28647 (N_28647,N_22035,N_20281);
nor U28648 (N_28648,N_23858,N_21138);
xor U28649 (N_28649,N_20964,N_23692);
nand U28650 (N_28650,N_23132,N_23626);
nor U28651 (N_28651,N_20672,N_24429);
xor U28652 (N_28652,N_24507,N_22817);
nor U28653 (N_28653,N_24159,N_23283);
nor U28654 (N_28654,N_20161,N_21769);
nand U28655 (N_28655,N_23706,N_22749);
nand U28656 (N_28656,N_23599,N_22240);
nand U28657 (N_28657,N_23186,N_20469);
and U28658 (N_28658,N_24569,N_21501);
or U28659 (N_28659,N_24535,N_22725);
nor U28660 (N_28660,N_22513,N_24587);
or U28661 (N_28661,N_23982,N_21643);
nand U28662 (N_28662,N_21659,N_21557);
nand U28663 (N_28663,N_22681,N_21370);
or U28664 (N_28664,N_23857,N_22072);
nand U28665 (N_28665,N_20343,N_22263);
nand U28666 (N_28666,N_22955,N_21319);
xor U28667 (N_28667,N_24590,N_22252);
xnor U28668 (N_28668,N_24435,N_23408);
nor U28669 (N_28669,N_23305,N_22512);
xnor U28670 (N_28670,N_20558,N_22130);
or U28671 (N_28671,N_23650,N_23870);
nand U28672 (N_28672,N_20057,N_24058);
and U28673 (N_28673,N_21249,N_24587);
xnor U28674 (N_28674,N_23289,N_22598);
xnor U28675 (N_28675,N_21639,N_23812);
and U28676 (N_28676,N_24672,N_21395);
nand U28677 (N_28677,N_23052,N_22789);
xnor U28678 (N_28678,N_21635,N_22955);
and U28679 (N_28679,N_22058,N_23375);
nand U28680 (N_28680,N_20426,N_22406);
and U28681 (N_28681,N_20893,N_24273);
xor U28682 (N_28682,N_23049,N_20090);
xor U28683 (N_28683,N_21145,N_20036);
and U28684 (N_28684,N_21539,N_22367);
or U28685 (N_28685,N_21477,N_21023);
nand U28686 (N_28686,N_23220,N_22421);
or U28687 (N_28687,N_22026,N_21632);
nor U28688 (N_28688,N_24127,N_23205);
and U28689 (N_28689,N_22114,N_22320);
xor U28690 (N_28690,N_23296,N_23080);
xor U28691 (N_28691,N_23441,N_21431);
nand U28692 (N_28692,N_20561,N_22576);
and U28693 (N_28693,N_20103,N_20316);
xor U28694 (N_28694,N_23632,N_22886);
nor U28695 (N_28695,N_24312,N_24612);
nor U28696 (N_28696,N_20715,N_20185);
or U28697 (N_28697,N_22557,N_22486);
nand U28698 (N_28698,N_22156,N_24202);
or U28699 (N_28699,N_21440,N_24358);
nor U28700 (N_28700,N_24093,N_21589);
and U28701 (N_28701,N_20872,N_22713);
and U28702 (N_28702,N_23508,N_20128);
xnor U28703 (N_28703,N_23456,N_20772);
and U28704 (N_28704,N_23466,N_21982);
xnor U28705 (N_28705,N_23915,N_22709);
nand U28706 (N_28706,N_22177,N_21311);
or U28707 (N_28707,N_23320,N_22100);
xor U28708 (N_28708,N_24117,N_24435);
and U28709 (N_28709,N_21848,N_23806);
or U28710 (N_28710,N_21163,N_20932);
or U28711 (N_28711,N_23444,N_21629);
or U28712 (N_28712,N_22133,N_23144);
or U28713 (N_28713,N_21052,N_24249);
nor U28714 (N_28714,N_23551,N_21094);
nor U28715 (N_28715,N_22981,N_22719);
or U28716 (N_28716,N_20554,N_20895);
xnor U28717 (N_28717,N_22475,N_24527);
nor U28718 (N_28718,N_24370,N_23828);
nor U28719 (N_28719,N_20788,N_22479);
and U28720 (N_28720,N_24222,N_23136);
nand U28721 (N_28721,N_23831,N_21880);
or U28722 (N_28722,N_24956,N_22434);
nand U28723 (N_28723,N_24531,N_23584);
nor U28724 (N_28724,N_24848,N_24633);
nor U28725 (N_28725,N_23729,N_24028);
nor U28726 (N_28726,N_22520,N_21133);
nor U28727 (N_28727,N_24396,N_22128);
nor U28728 (N_28728,N_21701,N_23894);
nor U28729 (N_28729,N_24390,N_24428);
or U28730 (N_28730,N_22385,N_22817);
xnor U28731 (N_28731,N_24142,N_22078);
or U28732 (N_28732,N_21373,N_23877);
nand U28733 (N_28733,N_22143,N_22399);
nand U28734 (N_28734,N_24847,N_22667);
and U28735 (N_28735,N_20280,N_24594);
or U28736 (N_28736,N_20167,N_22201);
xor U28737 (N_28737,N_23229,N_21288);
xor U28738 (N_28738,N_22365,N_24663);
nand U28739 (N_28739,N_21073,N_21586);
nor U28740 (N_28740,N_23493,N_21763);
and U28741 (N_28741,N_22794,N_23583);
nand U28742 (N_28742,N_24638,N_20045);
xor U28743 (N_28743,N_24680,N_24741);
nor U28744 (N_28744,N_24478,N_22858);
nand U28745 (N_28745,N_24232,N_22791);
or U28746 (N_28746,N_24801,N_20708);
nor U28747 (N_28747,N_21337,N_21292);
xnor U28748 (N_28748,N_24066,N_24359);
or U28749 (N_28749,N_23130,N_22097);
xnor U28750 (N_28750,N_23093,N_22988);
and U28751 (N_28751,N_22803,N_23866);
or U28752 (N_28752,N_23097,N_22598);
nor U28753 (N_28753,N_22286,N_21140);
nand U28754 (N_28754,N_23036,N_22169);
xor U28755 (N_28755,N_21497,N_20234);
nor U28756 (N_28756,N_21148,N_21814);
nand U28757 (N_28757,N_22945,N_20965);
nand U28758 (N_28758,N_21871,N_22537);
xor U28759 (N_28759,N_20630,N_21258);
xor U28760 (N_28760,N_22362,N_23658);
nand U28761 (N_28761,N_24069,N_24016);
or U28762 (N_28762,N_20149,N_20099);
nand U28763 (N_28763,N_20895,N_24527);
nor U28764 (N_28764,N_22839,N_21522);
nor U28765 (N_28765,N_23995,N_22670);
or U28766 (N_28766,N_20794,N_21296);
nor U28767 (N_28767,N_21629,N_20237);
xnor U28768 (N_28768,N_22647,N_23381);
and U28769 (N_28769,N_24035,N_21051);
and U28770 (N_28770,N_24387,N_21631);
and U28771 (N_28771,N_22681,N_20691);
or U28772 (N_28772,N_22168,N_24367);
nand U28773 (N_28773,N_23208,N_22217);
nor U28774 (N_28774,N_24064,N_23488);
nor U28775 (N_28775,N_23910,N_24703);
and U28776 (N_28776,N_24185,N_24261);
xnor U28777 (N_28777,N_23884,N_20604);
nand U28778 (N_28778,N_22010,N_24379);
nor U28779 (N_28779,N_24806,N_24100);
or U28780 (N_28780,N_20753,N_20631);
nand U28781 (N_28781,N_24245,N_22815);
nand U28782 (N_28782,N_21399,N_21439);
nor U28783 (N_28783,N_23610,N_20180);
or U28784 (N_28784,N_20282,N_22037);
nor U28785 (N_28785,N_23149,N_20119);
and U28786 (N_28786,N_21999,N_21677);
nor U28787 (N_28787,N_21225,N_24785);
or U28788 (N_28788,N_20609,N_22524);
and U28789 (N_28789,N_22770,N_21216);
and U28790 (N_28790,N_24750,N_20147);
or U28791 (N_28791,N_21370,N_23232);
and U28792 (N_28792,N_23685,N_23374);
nor U28793 (N_28793,N_24390,N_22615);
nor U28794 (N_28794,N_23276,N_23823);
and U28795 (N_28795,N_21055,N_23264);
and U28796 (N_28796,N_23470,N_23119);
or U28797 (N_28797,N_24281,N_23561);
or U28798 (N_28798,N_22863,N_21885);
nor U28799 (N_28799,N_22219,N_20414);
xnor U28800 (N_28800,N_24743,N_23440);
or U28801 (N_28801,N_22469,N_21781);
or U28802 (N_28802,N_23718,N_23867);
and U28803 (N_28803,N_24832,N_20078);
nand U28804 (N_28804,N_21878,N_21238);
nor U28805 (N_28805,N_20450,N_20953);
or U28806 (N_28806,N_23174,N_23646);
and U28807 (N_28807,N_21652,N_23708);
or U28808 (N_28808,N_24809,N_22485);
xnor U28809 (N_28809,N_24664,N_23508);
nor U28810 (N_28810,N_24742,N_21736);
or U28811 (N_28811,N_23828,N_22483);
and U28812 (N_28812,N_23951,N_22399);
and U28813 (N_28813,N_21048,N_23283);
and U28814 (N_28814,N_22182,N_22121);
and U28815 (N_28815,N_22679,N_22769);
and U28816 (N_28816,N_24674,N_22740);
nor U28817 (N_28817,N_23851,N_20831);
xnor U28818 (N_28818,N_23653,N_21952);
or U28819 (N_28819,N_22351,N_22250);
or U28820 (N_28820,N_20285,N_21993);
and U28821 (N_28821,N_20531,N_20556);
and U28822 (N_28822,N_23022,N_22275);
nand U28823 (N_28823,N_24816,N_23029);
or U28824 (N_28824,N_24802,N_21234);
or U28825 (N_28825,N_23177,N_22719);
nand U28826 (N_28826,N_21446,N_22875);
and U28827 (N_28827,N_20283,N_22819);
or U28828 (N_28828,N_20068,N_21103);
nand U28829 (N_28829,N_22464,N_22898);
or U28830 (N_28830,N_24349,N_21843);
or U28831 (N_28831,N_20102,N_21212);
or U28832 (N_28832,N_20110,N_20448);
nand U28833 (N_28833,N_20166,N_21415);
nand U28834 (N_28834,N_23394,N_23319);
or U28835 (N_28835,N_20692,N_20218);
and U28836 (N_28836,N_22525,N_22361);
and U28837 (N_28837,N_23317,N_23827);
nor U28838 (N_28838,N_20849,N_24028);
and U28839 (N_28839,N_24468,N_22117);
or U28840 (N_28840,N_21251,N_20914);
xnor U28841 (N_28841,N_24018,N_20918);
xor U28842 (N_28842,N_21739,N_22656);
xor U28843 (N_28843,N_22665,N_23030);
nand U28844 (N_28844,N_21107,N_21794);
xnor U28845 (N_28845,N_22647,N_22677);
xor U28846 (N_28846,N_23790,N_22425);
nand U28847 (N_28847,N_24950,N_20125);
nor U28848 (N_28848,N_20190,N_20917);
nand U28849 (N_28849,N_24260,N_21832);
xor U28850 (N_28850,N_21928,N_20409);
or U28851 (N_28851,N_21381,N_20817);
and U28852 (N_28852,N_24116,N_21231);
nor U28853 (N_28853,N_22438,N_24976);
nand U28854 (N_28854,N_24457,N_23444);
and U28855 (N_28855,N_21789,N_24418);
and U28856 (N_28856,N_22519,N_24129);
or U28857 (N_28857,N_22969,N_20839);
or U28858 (N_28858,N_21018,N_22523);
and U28859 (N_28859,N_22527,N_24692);
and U28860 (N_28860,N_21277,N_22835);
and U28861 (N_28861,N_24075,N_23783);
nand U28862 (N_28862,N_20802,N_22682);
nor U28863 (N_28863,N_22695,N_20704);
nor U28864 (N_28864,N_21177,N_20089);
and U28865 (N_28865,N_21360,N_22580);
and U28866 (N_28866,N_22260,N_23028);
xnor U28867 (N_28867,N_24701,N_23384);
or U28868 (N_28868,N_23621,N_20836);
xnor U28869 (N_28869,N_23627,N_24585);
nor U28870 (N_28870,N_22719,N_23525);
xnor U28871 (N_28871,N_20405,N_20511);
nor U28872 (N_28872,N_21183,N_20949);
or U28873 (N_28873,N_24277,N_24562);
and U28874 (N_28874,N_20969,N_23467);
and U28875 (N_28875,N_20925,N_24437);
or U28876 (N_28876,N_22895,N_21234);
nand U28877 (N_28877,N_24463,N_21803);
xnor U28878 (N_28878,N_24935,N_21639);
and U28879 (N_28879,N_24245,N_23584);
and U28880 (N_28880,N_20042,N_22105);
or U28881 (N_28881,N_20426,N_21868);
and U28882 (N_28882,N_21703,N_23534);
or U28883 (N_28883,N_22818,N_22909);
nor U28884 (N_28884,N_22024,N_21408);
and U28885 (N_28885,N_22212,N_22411);
nor U28886 (N_28886,N_22213,N_23735);
or U28887 (N_28887,N_22178,N_20819);
xor U28888 (N_28888,N_21094,N_22778);
or U28889 (N_28889,N_24079,N_20711);
nand U28890 (N_28890,N_24305,N_21964);
xor U28891 (N_28891,N_22995,N_24321);
nand U28892 (N_28892,N_23681,N_20636);
or U28893 (N_28893,N_23982,N_20527);
nand U28894 (N_28894,N_22602,N_24032);
and U28895 (N_28895,N_20589,N_22364);
xnor U28896 (N_28896,N_22019,N_22012);
and U28897 (N_28897,N_22841,N_22275);
nor U28898 (N_28898,N_22669,N_21289);
and U28899 (N_28899,N_21834,N_24056);
and U28900 (N_28900,N_22432,N_20943);
nor U28901 (N_28901,N_23212,N_22310);
and U28902 (N_28902,N_24004,N_23656);
nand U28903 (N_28903,N_21668,N_22798);
nor U28904 (N_28904,N_22487,N_24498);
and U28905 (N_28905,N_23949,N_24191);
and U28906 (N_28906,N_24562,N_21392);
or U28907 (N_28907,N_20741,N_23224);
nand U28908 (N_28908,N_23338,N_23962);
xor U28909 (N_28909,N_24761,N_24575);
nand U28910 (N_28910,N_23498,N_22610);
xnor U28911 (N_28911,N_24501,N_21184);
or U28912 (N_28912,N_20963,N_24412);
nand U28913 (N_28913,N_23156,N_24294);
nand U28914 (N_28914,N_22131,N_23048);
nor U28915 (N_28915,N_22828,N_22866);
nor U28916 (N_28916,N_22702,N_24967);
nand U28917 (N_28917,N_24112,N_20571);
nor U28918 (N_28918,N_23395,N_24496);
and U28919 (N_28919,N_21175,N_23458);
xor U28920 (N_28920,N_24107,N_24282);
nor U28921 (N_28921,N_21941,N_21414);
xnor U28922 (N_28922,N_20278,N_21071);
nor U28923 (N_28923,N_21784,N_21907);
or U28924 (N_28924,N_22957,N_20782);
xnor U28925 (N_28925,N_20519,N_23876);
or U28926 (N_28926,N_22642,N_22212);
and U28927 (N_28927,N_20922,N_23371);
and U28928 (N_28928,N_22197,N_21792);
nand U28929 (N_28929,N_23836,N_20165);
and U28930 (N_28930,N_24488,N_23847);
nor U28931 (N_28931,N_22455,N_20305);
and U28932 (N_28932,N_23244,N_20278);
and U28933 (N_28933,N_24088,N_22072);
or U28934 (N_28934,N_21261,N_21941);
xnor U28935 (N_28935,N_23060,N_20488);
and U28936 (N_28936,N_20571,N_23483);
or U28937 (N_28937,N_23341,N_24877);
or U28938 (N_28938,N_24689,N_22583);
nor U28939 (N_28939,N_22603,N_23342);
nand U28940 (N_28940,N_24996,N_21146);
xnor U28941 (N_28941,N_21692,N_20805);
nor U28942 (N_28942,N_22538,N_20595);
or U28943 (N_28943,N_23843,N_20328);
nand U28944 (N_28944,N_22872,N_21663);
nor U28945 (N_28945,N_24353,N_23136);
and U28946 (N_28946,N_22473,N_21805);
xnor U28947 (N_28947,N_21144,N_21446);
and U28948 (N_28948,N_21913,N_20537);
or U28949 (N_28949,N_24121,N_21360);
xor U28950 (N_28950,N_20644,N_20785);
nor U28951 (N_28951,N_21237,N_24503);
nor U28952 (N_28952,N_23205,N_23008);
xor U28953 (N_28953,N_24846,N_21160);
or U28954 (N_28954,N_23417,N_21550);
nor U28955 (N_28955,N_20542,N_24100);
or U28956 (N_28956,N_23645,N_21083);
nor U28957 (N_28957,N_21719,N_21818);
nor U28958 (N_28958,N_20755,N_21881);
nor U28959 (N_28959,N_22387,N_20933);
nand U28960 (N_28960,N_21192,N_20820);
xnor U28961 (N_28961,N_21216,N_21149);
nor U28962 (N_28962,N_20541,N_24317);
and U28963 (N_28963,N_24593,N_24759);
nand U28964 (N_28964,N_24509,N_22587);
nor U28965 (N_28965,N_21611,N_20864);
nor U28966 (N_28966,N_21099,N_21287);
xor U28967 (N_28967,N_24938,N_23019);
nand U28968 (N_28968,N_22090,N_21710);
and U28969 (N_28969,N_24826,N_22980);
and U28970 (N_28970,N_20541,N_20211);
nor U28971 (N_28971,N_24440,N_22098);
nand U28972 (N_28972,N_21287,N_23959);
nand U28973 (N_28973,N_23762,N_21835);
nand U28974 (N_28974,N_23192,N_20757);
nor U28975 (N_28975,N_23798,N_21031);
nor U28976 (N_28976,N_21066,N_21189);
nor U28977 (N_28977,N_22155,N_21436);
or U28978 (N_28978,N_20761,N_23901);
nor U28979 (N_28979,N_21096,N_21609);
xnor U28980 (N_28980,N_22946,N_24905);
and U28981 (N_28981,N_21304,N_22945);
nor U28982 (N_28982,N_24344,N_22677);
or U28983 (N_28983,N_22250,N_24701);
or U28984 (N_28984,N_24473,N_21007);
or U28985 (N_28985,N_24974,N_24175);
or U28986 (N_28986,N_20010,N_21493);
or U28987 (N_28987,N_22038,N_22656);
and U28988 (N_28988,N_22588,N_21807);
or U28989 (N_28989,N_22003,N_21620);
nand U28990 (N_28990,N_20837,N_21917);
xnor U28991 (N_28991,N_20016,N_24250);
or U28992 (N_28992,N_23087,N_22564);
nor U28993 (N_28993,N_21565,N_22490);
and U28994 (N_28994,N_20854,N_21652);
and U28995 (N_28995,N_24325,N_21114);
nor U28996 (N_28996,N_20940,N_20387);
xnor U28997 (N_28997,N_24868,N_22225);
or U28998 (N_28998,N_22775,N_24761);
or U28999 (N_28999,N_20156,N_22678);
xnor U29000 (N_29000,N_23535,N_23010);
and U29001 (N_29001,N_20106,N_23882);
and U29002 (N_29002,N_21986,N_23367);
xnor U29003 (N_29003,N_23639,N_23560);
nand U29004 (N_29004,N_21482,N_23736);
xor U29005 (N_29005,N_22865,N_23922);
or U29006 (N_29006,N_24073,N_24051);
nand U29007 (N_29007,N_22577,N_24150);
nand U29008 (N_29008,N_21423,N_20087);
or U29009 (N_29009,N_23027,N_24524);
or U29010 (N_29010,N_22200,N_22078);
or U29011 (N_29011,N_20484,N_21923);
nand U29012 (N_29012,N_21569,N_23756);
nand U29013 (N_29013,N_22626,N_21720);
or U29014 (N_29014,N_20037,N_21178);
and U29015 (N_29015,N_22989,N_21899);
or U29016 (N_29016,N_21755,N_24317);
or U29017 (N_29017,N_21502,N_24026);
nand U29018 (N_29018,N_21313,N_21875);
nor U29019 (N_29019,N_24192,N_20612);
xnor U29020 (N_29020,N_22050,N_23836);
nand U29021 (N_29021,N_24235,N_24754);
xnor U29022 (N_29022,N_22045,N_21207);
and U29023 (N_29023,N_24846,N_23048);
nand U29024 (N_29024,N_20216,N_22517);
or U29025 (N_29025,N_24343,N_21836);
nor U29026 (N_29026,N_22084,N_22194);
xor U29027 (N_29027,N_23848,N_20550);
nand U29028 (N_29028,N_24149,N_24746);
nor U29029 (N_29029,N_20017,N_21300);
and U29030 (N_29030,N_23637,N_21218);
nor U29031 (N_29031,N_24463,N_21059);
xor U29032 (N_29032,N_22329,N_24031);
and U29033 (N_29033,N_21452,N_22083);
nor U29034 (N_29034,N_22438,N_23606);
or U29035 (N_29035,N_23338,N_23619);
nand U29036 (N_29036,N_20968,N_22888);
nor U29037 (N_29037,N_20695,N_23507);
xor U29038 (N_29038,N_20882,N_21949);
xnor U29039 (N_29039,N_21540,N_22838);
and U29040 (N_29040,N_23647,N_24064);
nor U29041 (N_29041,N_20686,N_24964);
xor U29042 (N_29042,N_23046,N_22915);
nor U29043 (N_29043,N_22477,N_24534);
or U29044 (N_29044,N_21482,N_22685);
or U29045 (N_29045,N_23572,N_22793);
and U29046 (N_29046,N_23017,N_20773);
nor U29047 (N_29047,N_24218,N_21479);
xnor U29048 (N_29048,N_21987,N_24234);
nor U29049 (N_29049,N_23763,N_24519);
nor U29050 (N_29050,N_21082,N_22577);
nand U29051 (N_29051,N_21054,N_22422);
nand U29052 (N_29052,N_21042,N_24509);
nor U29053 (N_29053,N_24084,N_22845);
and U29054 (N_29054,N_23197,N_20965);
xnor U29055 (N_29055,N_21674,N_24386);
nand U29056 (N_29056,N_21694,N_23057);
nor U29057 (N_29057,N_23476,N_20232);
nor U29058 (N_29058,N_23356,N_24122);
xnor U29059 (N_29059,N_22061,N_24547);
or U29060 (N_29060,N_24628,N_22988);
xor U29061 (N_29061,N_23910,N_20239);
xor U29062 (N_29062,N_21785,N_20610);
xor U29063 (N_29063,N_21316,N_21169);
or U29064 (N_29064,N_21007,N_23598);
or U29065 (N_29065,N_21346,N_21810);
nand U29066 (N_29066,N_21465,N_22678);
and U29067 (N_29067,N_21538,N_22970);
xor U29068 (N_29068,N_23802,N_22574);
and U29069 (N_29069,N_21097,N_22076);
or U29070 (N_29070,N_24011,N_23678);
and U29071 (N_29071,N_24319,N_24635);
and U29072 (N_29072,N_21534,N_24761);
or U29073 (N_29073,N_20491,N_22336);
xor U29074 (N_29074,N_23387,N_20466);
nor U29075 (N_29075,N_21722,N_23971);
nand U29076 (N_29076,N_20485,N_23846);
nor U29077 (N_29077,N_21301,N_20485);
nand U29078 (N_29078,N_24354,N_21118);
nor U29079 (N_29079,N_24431,N_24314);
nor U29080 (N_29080,N_20569,N_24150);
and U29081 (N_29081,N_24269,N_22279);
or U29082 (N_29082,N_21013,N_21176);
or U29083 (N_29083,N_20127,N_22574);
and U29084 (N_29084,N_23883,N_24749);
nor U29085 (N_29085,N_21442,N_24623);
nand U29086 (N_29086,N_20664,N_24491);
xnor U29087 (N_29087,N_21003,N_21347);
xnor U29088 (N_29088,N_20841,N_23197);
xnor U29089 (N_29089,N_23464,N_20229);
or U29090 (N_29090,N_24534,N_24698);
nand U29091 (N_29091,N_22808,N_24227);
nand U29092 (N_29092,N_21441,N_21258);
xnor U29093 (N_29093,N_21331,N_24958);
nand U29094 (N_29094,N_23518,N_23966);
or U29095 (N_29095,N_21190,N_24916);
or U29096 (N_29096,N_21999,N_20405);
nor U29097 (N_29097,N_22723,N_21998);
nand U29098 (N_29098,N_22184,N_21160);
or U29099 (N_29099,N_24577,N_23132);
xnor U29100 (N_29100,N_24101,N_22183);
xor U29101 (N_29101,N_23837,N_20738);
nor U29102 (N_29102,N_20127,N_24919);
nor U29103 (N_29103,N_24495,N_24933);
or U29104 (N_29104,N_20940,N_24918);
xor U29105 (N_29105,N_24389,N_23769);
nor U29106 (N_29106,N_24271,N_22084);
or U29107 (N_29107,N_23724,N_24495);
or U29108 (N_29108,N_21764,N_21544);
xor U29109 (N_29109,N_23454,N_20146);
xnor U29110 (N_29110,N_20574,N_24975);
nor U29111 (N_29111,N_22881,N_23049);
and U29112 (N_29112,N_24018,N_24953);
xor U29113 (N_29113,N_20116,N_23367);
nor U29114 (N_29114,N_21379,N_24004);
xor U29115 (N_29115,N_20091,N_23721);
or U29116 (N_29116,N_20819,N_20632);
nand U29117 (N_29117,N_20349,N_23027);
nor U29118 (N_29118,N_24491,N_24257);
or U29119 (N_29119,N_20586,N_23246);
nor U29120 (N_29120,N_24083,N_20242);
nand U29121 (N_29121,N_21162,N_24752);
and U29122 (N_29122,N_23679,N_22588);
xor U29123 (N_29123,N_23950,N_20956);
nand U29124 (N_29124,N_24971,N_24871);
nand U29125 (N_29125,N_20195,N_23300);
nand U29126 (N_29126,N_20149,N_21124);
nand U29127 (N_29127,N_23799,N_23153);
nand U29128 (N_29128,N_20131,N_23893);
and U29129 (N_29129,N_21800,N_20384);
nor U29130 (N_29130,N_23330,N_21671);
nor U29131 (N_29131,N_21180,N_21249);
xor U29132 (N_29132,N_21705,N_23272);
or U29133 (N_29133,N_23025,N_22793);
or U29134 (N_29134,N_20965,N_22899);
nor U29135 (N_29135,N_21978,N_22769);
and U29136 (N_29136,N_20138,N_20750);
and U29137 (N_29137,N_24331,N_22463);
and U29138 (N_29138,N_22392,N_20967);
nand U29139 (N_29139,N_21367,N_20566);
nor U29140 (N_29140,N_22112,N_23734);
and U29141 (N_29141,N_24151,N_24769);
and U29142 (N_29142,N_22268,N_22702);
nor U29143 (N_29143,N_23294,N_20832);
or U29144 (N_29144,N_21655,N_22882);
or U29145 (N_29145,N_21300,N_20496);
xnor U29146 (N_29146,N_22967,N_21580);
and U29147 (N_29147,N_21469,N_22277);
or U29148 (N_29148,N_23718,N_22420);
xnor U29149 (N_29149,N_21408,N_21606);
nor U29150 (N_29150,N_24973,N_21671);
and U29151 (N_29151,N_23139,N_23202);
and U29152 (N_29152,N_21060,N_20286);
and U29153 (N_29153,N_24494,N_20680);
and U29154 (N_29154,N_23581,N_22746);
xnor U29155 (N_29155,N_22401,N_21641);
and U29156 (N_29156,N_22197,N_23028);
nand U29157 (N_29157,N_23887,N_24845);
nand U29158 (N_29158,N_22434,N_22886);
and U29159 (N_29159,N_21838,N_21060);
nor U29160 (N_29160,N_21118,N_23997);
nand U29161 (N_29161,N_22987,N_20899);
nand U29162 (N_29162,N_24315,N_22085);
nor U29163 (N_29163,N_21632,N_22121);
or U29164 (N_29164,N_23254,N_23218);
nor U29165 (N_29165,N_22401,N_24728);
or U29166 (N_29166,N_21818,N_21585);
or U29167 (N_29167,N_20072,N_23648);
nor U29168 (N_29168,N_21103,N_23933);
nor U29169 (N_29169,N_21172,N_24257);
nor U29170 (N_29170,N_22867,N_24348);
nor U29171 (N_29171,N_21059,N_20483);
or U29172 (N_29172,N_23854,N_20938);
and U29173 (N_29173,N_23796,N_24068);
nor U29174 (N_29174,N_23463,N_21237);
nor U29175 (N_29175,N_22668,N_22154);
and U29176 (N_29176,N_22740,N_24200);
xor U29177 (N_29177,N_20997,N_21127);
nand U29178 (N_29178,N_20481,N_23778);
and U29179 (N_29179,N_24139,N_23597);
or U29180 (N_29180,N_24829,N_24115);
or U29181 (N_29181,N_21136,N_22894);
or U29182 (N_29182,N_21234,N_23534);
and U29183 (N_29183,N_21088,N_22489);
or U29184 (N_29184,N_23936,N_21374);
xnor U29185 (N_29185,N_23970,N_20076);
or U29186 (N_29186,N_21930,N_23139);
or U29187 (N_29187,N_24420,N_22594);
nor U29188 (N_29188,N_23046,N_20503);
nor U29189 (N_29189,N_22505,N_24047);
nand U29190 (N_29190,N_21936,N_21384);
or U29191 (N_29191,N_23488,N_20842);
nand U29192 (N_29192,N_23690,N_23789);
nand U29193 (N_29193,N_20610,N_23871);
xnor U29194 (N_29194,N_21883,N_21513);
nand U29195 (N_29195,N_20838,N_20484);
and U29196 (N_29196,N_21985,N_23451);
nor U29197 (N_29197,N_20749,N_24786);
nand U29198 (N_29198,N_24077,N_22716);
nor U29199 (N_29199,N_20280,N_20572);
nand U29200 (N_29200,N_21076,N_20158);
and U29201 (N_29201,N_21299,N_21183);
or U29202 (N_29202,N_21949,N_24700);
xnor U29203 (N_29203,N_23889,N_23021);
nor U29204 (N_29204,N_23017,N_22932);
xnor U29205 (N_29205,N_22813,N_23976);
nor U29206 (N_29206,N_24288,N_22096);
xnor U29207 (N_29207,N_23239,N_21570);
nand U29208 (N_29208,N_22291,N_21282);
xor U29209 (N_29209,N_20719,N_24281);
xor U29210 (N_29210,N_23385,N_24702);
and U29211 (N_29211,N_22203,N_23115);
and U29212 (N_29212,N_22715,N_21054);
nand U29213 (N_29213,N_21320,N_20741);
nand U29214 (N_29214,N_21173,N_24231);
and U29215 (N_29215,N_23521,N_24467);
nand U29216 (N_29216,N_23900,N_22908);
and U29217 (N_29217,N_21397,N_20966);
and U29218 (N_29218,N_23009,N_20044);
nor U29219 (N_29219,N_24509,N_23865);
nor U29220 (N_29220,N_20046,N_24908);
or U29221 (N_29221,N_23303,N_21191);
nor U29222 (N_29222,N_23996,N_20069);
xor U29223 (N_29223,N_23327,N_24805);
nand U29224 (N_29224,N_24027,N_24583);
and U29225 (N_29225,N_21470,N_23537);
or U29226 (N_29226,N_24943,N_21228);
and U29227 (N_29227,N_20166,N_21627);
nor U29228 (N_29228,N_24042,N_21044);
nor U29229 (N_29229,N_23975,N_23022);
or U29230 (N_29230,N_23569,N_22260);
xor U29231 (N_29231,N_23283,N_21996);
xnor U29232 (N_29232,N_20238,N_22503);
nor U29233 (N_29233,N_20622,N_24218);
nor U29234 (N_29234,N_21060,N_20980);
nor U29235 (N_29235,N_22694,N_22501);
and U29236 (N_29236,N_21094,N_24514);
and U29237 (N_29237,N_21008,N_22908);
nand U29238 (N_29238,N_24967,N_23573);
nand U29239 (N_29239,N_20296,N_20056);
xnor U29240 (N_29240,N_23244,N_20713);
nand U29241 (N_29241,N_23710,N_23457);
xnor U29242 (N_29242,N_21114,N_22243);
xor U29243 (N_29243,N_23327,N_21516);
or U29244 (N_29244,N_23568,N_23072);
xor U29245 (N_29245,N_20999,N_22646);
and U29246 (N_29246,N_24689,N_20060);
nor U29247 (N_29247,N_21964,N_24738);
nand U29248 (N_29248,N_20959,N_22476);
xor U29249 (N_29249,N_24416,N_21268);
xor U29250 (N_29250,N_20512,N_22134);
and U29251 (N_29251,N_22034,N_21605);
nand U29252 (N_29252,N_22976,N_22492);
nand U29253 (N_29253,N_21277,N_24456);
or U29254 (N_29254,N_21550,N_24868);
and U29255 (N_29255,N_21731,N_24808);
nor U29256 (N_29256,N_21662,N_22558);
or U29257 (N_29257,N_20480,N_20357);
or U29258 (N_29258,N_22048,N_23124);
and U29259 (N_29259,N_20911,N_21784);
or U29260 (N_29260,N_24707,N_22480);
nor U29261 (N_29261,N_23156,N_23488);
nor U29262 (N_29262,N_23642,N_21257);
nand U29263 (N_29263,N_23008,N_21340);
and U29264 (N_29264,N_21473,N_24081);
nor U29265 (N_29265,N_20422,N_21467);
and U29266 (N_29266,N_22524,N_24021);
and U29267 (N_29267,N_21439,N_21080);
nor U29268 (N_29268,N_24923,N_22933);
nor U29269 (N_29269,N_22360,N_20763);
and U29270 (N_29270,N_21336,N_21851);
nand U29271 (N_29271,N_22466,N_20081);
nand U29272 (N_29272,N_24422,N_21241);
or U29273 (N_29273,N_20736,N_23205);
xnor U29274 (N_29274,N_21859,N_22378);
and U29275 (N_29275,N_21649,N_20409);
nor U29276 (N_29276,N_23992,N_21938);
nor U29277 (N_29277,N_20060,N_20901);
xnor U29278 (N_29278,N_24627,N_22121);
or U29279 (N_29279,N_21915,N_20210);
and U29280 (N_29280,N_22377,N_23971);
nand U29281 (N_29281,N_22240,N_22770);
nand U29282 (N_29282,N_23741,N_23913);
xor U29283 (N_29283,N_24176,N_24803);
and U29284 (N_29284,N_24105,N_24069);
or U29285 (N_29285,N_20957,N_22822);
nor U29286 (N_29286,N_24216,N_22391);
nand U29287 (N_29287,N_21180,N_23600);
and U29288 (N_29288,N_20782,N_24426);
nor U29289 (N_29289,N_24132,N_23741);
xnor U29290 (N_29290,N_20089,N_24505);
nor U29291 (N_29291,N_23649,N_23510);
nand U29292 (N_29292,N_23986,N_20082);
or U29293 (N_29293,N_24044,N_22297);
and U29294 (N_29294,N_22754,N_22190);
or U29295 (N_29295,N_24822,N_22243);
nand U29296 (N_29296,N_20785,N_24602);
and U29297 (N_29297,N_20398,N_21448);
or U29298 (N_29298,N_24147,N_24953);
nand U29299 (N_29299,N_24177,N_22652);
xnor U29300 (N_29300,N_21417,N_20238);
xor U29301 (N_29301,N_20474,N_22580);
nand U29302 (N_29302,N_20688,N_23569);
nand U29303 (N_29303,N_23168,N_20490);
nor U29304 (N_29304,N_21790,N_24195);
nand U29305 (N_29305,N_20686,N_24762);
nor U29306 (N_29306,N_21176,N_24474);
or U29307 (N_29307,N_20744,N_23805);
or U29308 (N_29308,N_24952,N_23157);
and U29309 (N_29309,N_23409,N_23122);
or U29310 (N_29310,N_21520,N_22294);
nor U29311 (N_29311,N_21256,N_21142);
nand U29312 (N_29312,N_21250,N_24078);
and U29313 (N_29313,N_22642,N_23321);
nand U29314 (N_29314,N_23136,N_22277);
and U29315 (N_29315,N_21124,N_22272);
or U29316 (N_29316,N_22653,N_23673);
xnor U29317 (N_29317,N_20364,N_22636);
nand U29318 (N_29318,N_24979,N_22629);
nor U29319 (N_29319,N_24560,N_22624);
xor U29320 (N_29320,N_21404,N_23556);
or U29321 (N_29321,N_20898,N_20790);
and U29322 (N_29322,N_20183,N_23408);
xor U29323 (N_29323,N_23439,N_20996);
and U29324 (N_29324,N_22796,N_24718);
and U29325 (N_29325,N_20377,N_22275);
xnor U29326 (N_29326,N_24980,N_22353);
and U29327 (N_29327,N_22576,N_24180);
xnor U29328 (N_29328,N_21972,N_20144);
or U29329 (N_29329,N_23052,N_24383);
and U29330 (N_29330,N_20503,N_24761);
nor U29331 (N_29331,N_21345,N_22548);
nor U29332 (N_29332,N_20175,N_20379);
or U29333 (N_29333,N_24179,N_20759);
nor U29334 (N_29334,N_21613,N_24731);
or U29335 (N_29335,N_24504,N_21759);
nand U29336 (N_29336,N_20773,N_20551);
xor U29337 (N_29337,N_20831,N_22196);
xor U29338 (N_29338,N_22229,N_24181);
xnor U29339 (N_29339,N_22142,N_22925);
xor U29340 (N_29340,N_22433,N_24272);
xnor U29341 (N_29341,N_23697,N_23575);
xnor U29342 (N_29342,N_20969,N_21721);
nor U29343 (N_29343,N_22242,N_23635);
xor U29344 (N_29344,N_24461,N_24519);
nor U29345 (N_29345,N_20136,N_20222);
nand U29346 (N_29346,N_20458,N_24666);
and U29347 (N_29347,N_21887,N_21808);
xnor U29348 (N_29348,N_23351,N_23416);
or U29349 (N_29349,N_23913,N_20292);
xnor U29350 (N_29350,N_20282,N_23508);
nor U29351 (N_29351,N_20152,N_23416);
or U29352 (N_29352,N_22546,N_20567);
nand U29353 (N_29353,N_20434,N_24131);
or U29354 (N_29354,N_22869,N_23583);
or U29355 (N_29355,N_24771,N_20634);
nand U29356 (N_29356,N_23043,N_21921);
nor U29357 (N_29357,N_24249,N_22626);
or U29358 (N_29358,N_23556,N_20791);
and U29359 (N_29359,N_20563,N_21232);
xor U29360 (N_29360,N_23333,N_20169);
nor U29361 (N_29361,N_22076,N_24307);
nor U29362 (N_29362,N_20083,N_24379);
and U29363 (N_29363,N_20481,N_22081);
xor U29364 (N_29364,N_23392,N_20232);
nor U29365 (N_29365,N_21131,N_24285);
xor U29366 (N_29366,N_20286,N_20592);
nor U29367 (N_29367,N_23339,N_24700);
xor U29368 (N_29368,N_20345,N_20898);
nand U29369 (N_29369,N_24731,N_21850);
nand U29370 (N_29370,N_20343,N_22291);
and U29371 (N_29371,N_21168,N_23121);
nand U29372 (N_29372,N_21624,N_23748);
xor U29373 (N_29373,N_22906,N_21021);
and U29374 (N_29374,N_23648,N_22004);
xor U29375 (N_29375,N_22747,N_20879);
and U29376 (N_29376,N_24477,N_20567);
or U29377 (N_29377,N_24667,N_24093);
nand U29378 (N_29378,N_23291,N_22712);
nand U29379 (N_29379,N_22758,N_20581);
and U29380 (N_29380,N_21063,N_22236);
xnor U29381 (N_29381,N_22363,N_22795);
or U29382 (N_29382,N_24713,N_20020);
xor U29383 (N_29383,N_20294,N_23754);
or U29384 (N_29384,N_20432,N_21957);
nand U29385 (N_29385,N_22320,N_23016);
nor U29386 (N_29386,N_20559,N_20119);
nor U29387 (N_29387,N_21429,N_23972);
and U29388 (N_29388,N_24234,N_20084);
or U29389 (N_29389,N_24641,N_24489);
nor U29390 (N_29390,N_22040,N_21567);
nor U29391 (N_29391,N_20731,N_23893);
nor U29392 (N_29392,N_23641,N_20959);
nor U29393 (N_29393,N_22687,N_20648);
nand U29394 (N_29394,N_22065,N_21191);
xnor U29395 (N_29395,N_20798,N_24623);
or U29396 (N_29396,N_20196,N_21137);
nand U29397 (N_29397,N_24253,N_22130);
nor U29398 (N_29398,N_22087,N_24913);
nor U29399 (N_29399,N_20347,N_22414);
xnor U29400 (N_29400,N_23268,N_21922);
xnor U29401 (N_29401,N_23075,N_23759);
nand U29402 (N_29402,N_24444,N_23534);
nand U29403 (N_29403,N_23849,N_20830);
or U29404 (N_29404,N_23084,N_20066);
xnor U29405 (N_29405,N_24920,N_20019);
or U29406 (N_29406,N_22551,N_24478);
or U29407 (N_29407,N_22151,N_20475);
nand U29408 (N_29408,N_24773,N_23929);
and U29409 (N_29409,N_23488,N_24859);
or U29410 (N_29410,N_22135,N_20445);
xor U29411 (N_29411,N_22280,N_21706);
or U29412 (N_29412,N_23391,N_23531);
nand U29413 (N_29413,N_24032,N_22386);
xnor U29414 (N_29414,N_22912,N_23787);
nand U29415 (N_29415,N_20723,N_24089);
nor U29416 (N_29416,N_21077,N_23465);
nand U29417 (N_29417,N_21525,N_20241);
and U29418 (N_29418,N_20031,N_21632);
or U29419 (N_29419,N_21265,N_24428);
or U29420 (N_29420,N_22714,N_24501);
xnor U29421 (N_29421,N_20358,N_22345);
and U29422 (N_29422,N_21873,N_24545);
nand U29423 (N_29423,N_23210,N_20595);
and U29424 (N_29424,N_21344,N_22409);
nor U29425 (N_29425,N_22576,N_24272);
nor U29426 (N_29426,N_21560,N_21763);
nand U29427 (N_29427,N_23510,N_20858);
and U29428 (N_29428,N_24505,N_24133);
nand U29429 (N_29429,N_22225,N_24032);
nand U29430 (N_29430,N_20195,N_20987);
nand U29431 (N_29431,N_24876,N_24487);
and U29432 (N_29432,N_22608,N_21233);
nand U29433 (N_29433,N_24051,N_21290);
xnor U29434 (N_29434,N_21819,N_20699);
and U29435 (N_29435,N_20439,N_22263);
nor U29436 (N_29436,N_20841,N_22501);
and U29437 (N_29437,N_24859,N_20419);
nor U29438 (N_29438,N_20165,N_24639);
nor U29439 (N_29439,N_24657,N_22634);
nand U29440 (N_29440,N_24924,N_21728);
or U29441 (N_29441,N_20740,N_20034);
or U29442 (N_29442,N_23543,N_22241);
nor U29443 (N_29443,N_21185,N_21364);
xnor U29444 (N_29444,N_21765,N_23788);
xnor U29445 (N_29445,N_24543,N_24605);
or U29446 (N_29446,N_24272,N_21760);
nand U29447 (N_29447,N_21527,N_22855);
nand U29448 (N_29448,N_23597,N_23696);
nor U29449 (N_29449,N_22097,N_21917);
nand U29450 (N_29450,N_22702,N_24062);
or U29451 (N_29451,N_23318,N_23511);
nor U29452 (N_29452,N_20836,N_20931);
xnor U29453 (N_29453,N_21494,N_23542);
xor U29454 (N_29454,N_24644,N_23335);
nor U29455 (N_29455,N_22174,N_22217);
nor U29456 (N_29456,N_22723,N_24308);
nor U29457 (N_29457,N_20346,N_21478);
nand U29458 (N_29458,N_22975,N_20546);
nor U29459 (N_29459,N_22099,N_22646);
or U29460 (N_29460,N_24134,N_23046);
or U29461 (N_29461,N_22723,N_21810);
xor U29462 (N_29462,N_20085,N_24595);
nor U29463 (N_29463,N_20572,N_22008);
nor U29464 (N_29464,N_23431,N_24952);
xor U29465 (N_29465,N_20882,N_23460);
nor U29466 (N_29466,N_22043,N_23396);
and U29467 (N_29467,N_24380,N_23008);
nand U29468 (N_29468,N_23674,N_20440);
nand U29469 (N_29469,N_21050,N_22186);
and U29470 (N_29470,N_22881,N_20413);
nor U29471 (N_29471,N_20873,N_20034);
xor U29472 (N_29472,N_22041,N_20980);
xnor U29473 (N_29473,N_20116,N_21460);
and U29474 (N_29474,N_22673,N_22643);
nand U29475 (N_29475,N_21328,N_21120);
and U29476 (N_29476,N_21735,N_20890);
xor U29477 (N_29477,N_20430,N_22256);
nand U29478 (N_29478,N_21719,N_22180);
or U29479 (N_29479,N_22729,N_20071);
or U29480 (N_29480,N_24903,N_20618);
nand U29481 (N_29481,N_20124,N_22331);
and U29482 (N_29482,N_24535,N_20659);
and U29483 (N_29483,N_21270,N_24482);
and U29484 (N_29484,N_22663,N_21139);
nand U29485 (N_29485,N_20994,N_20324);
or U29486 (N_29486,N_20919,N_23739);
xnor U29487 (N_29487,N_21150,N_21790);
xor U29488 (N_29488,N_20527,N_24635);
xnor U29489 (N_29489,N_21649,N_21040);
or U29490 (N_29490,N_23291,N_21648);
nor U29491 (N_29491,N_22045,N_23697);
or U29492 (N_29492,N_23199,N_23256);
nand U29493 (N_29493,N_23367,N_21506);
and U29494 (N_29494,N_22829,N_22751);
or U29495 (N_29495,N_20348,N_21125);
or U29496 (N_29496,N_20107,N_24716);
xor U29497 (N_29497,N_21083,N_20678);
or U29498 (N_29498,N_20617,N_24335);
or U29499 (N_29499,N_22086,N_22589);
nor U29500 (N_29500,N_22841,N_22287);
xnor U29501 (N_29501,N_24443,N_24027);
nor U29502 (N_29502,N_21817,N_24207);
and U29503 (N_29503,N_24328,N_21863);
nand U29504 (N_29504,N_21178,N_24878);
or U29505 (N_29505,N_24004,N_20163);
nand U29506 (N_29506,N_24479,N_24677);
nor U29507 (N_29507,N_20102,N_20487);
or U29508 (N_29508,N_24596,N_23025);
xnor U29509 (N_29509,N_23558,N_21191);
and U29510 (N_29510,N_23593,N_21896);
xnor U29511 (N_29511,N_24001,N_22132);
nor U29512 (N_29512,N_21303,N_22512);
and U29513 (N_29513,N_22431,N_21127);
and U29514 (N_29514,N_23094,N_22032);
nor U29515 (N_29515,N_21386,N_21785);
nand U29516 (N_29516,N_24437,N_21528);
nand U29517 (N_29517,N_24965,N_21498);
and U29518 (N_29518,N_22904,N_21152);
nor U29519 (N_29519,N_22814,N_23186);
and U29520 (N_29520,N_20666,N_23831);
nand U29521 (N_29521,N_22319,N_20246);
and U29522 (N_29522,N_20193,N_21505);
and U29523 (N_29523,N_20179,N_20212);
nor U29524 (N_29524,N_24958,N_20396);
nand U29525 (N_29525,N_20300,N_24355);
nand U29526 (N_29526,N_20611,N_24788);
nor U29527 (N_29527,N_24580,N_24538);
nand U29528 (N_29528,N_24405,N_23656);
or U29529 (N_29529,N_20279,N_24479);
nand U29530 (N_29530,N_22590,N_24983);
nor U29531 (N_29531,N_22514,N_21612);
nor U29532 (N_29532,N_23513,N_21036);
nand U29533 (N_29533,N_22550,N_24095);
nor U29534 (N_29534,N_24582,N_21129);
or U29535 (N_29535,N_20506,N_21908);
xor U29536 (N_29536,N_23790,N_21014);
nor U29537 (N_29537,N_20850,N_20451);
nand U29538 (N_29538,N_20542,N_23353);
nor U29539 (N_29539,N_22273,N_24520);
or U29540 (N_29540,N_20666,N_23947);
nor U29541 (N_29541,N_21454,N_20765);
and U29542 (N_29542,N_24850,N_20200);
or U29543 (N_29543,N_24780,N_23627);
nor U29544 (N_29544,N_23690,N_22995);
and U29545 (N_29545,N_23154,N_22073);
and U29546 (N_29546,N_23407,N_21084);
or U29547 (N_29547,N_21819,N_22310);
xnor U29548 (N_29548,N_22644,N_20349);
nor U29549 (N_29549,N_22113,N_21819);
nor U29550 (N_29550,N_21646,N_21184);
or U29551 (N_29551,N_24932,N_21436);
and U29552 (N_29552,N_20122,N_23571);
and U29553 (N_29553,N_22875,N_20389);
xnor U29554 (N_29554,N_23182,N_23745);
nand U29555 (N_29555,N_24901,N_21814);
nand U29556 (N_29556,N_23491,N_23205);
xor U29557 (N_29557,N_23463,N_20151);
nand U29558 (N_29558,N_21373,N_24540);
nand U29559 (N_29559,N_22174,N_23180);
nor U29560 (N_29560,N_21922,N_22039);
xnor U29561 (N_29561,N_20809,N_23540);
nand U29562 (N_29562,N_24367,N_22527);
or U29563 (N_29563,N_24601,N_23768);
nor U29564 (N_29564,N_23866,N_20104);
or U29565 (N_29565,N_20022,N_22293);
or U29566 (N_29566,N_23908,N_20210);
nor U29567 (N_29567,N_20696,N_23556);
and U29568 (N_29568,N_23723,N_24582);
and U29569 (N_29569,N_23129,N_24920);
nand U29570 (N_29570,N_24935,N_22709);
nand U29571 (N_29571,N_23722,N_22493);
nand U29572 (N_29572,N_22848,N_22576);
or U29573 (N_29573,N_20525,N_24380);
and U29574 (N_29574,N_21677,N_24183);
and U29575 (N_29575,N_22483,N_23330);
nor U29576 (N_29576,N_21494,N_21820);
or U29577 (N_29577,N_20053,N_24575);
nand U29578 (N_29578,N_22441,N_22407);
xor U29579 (N_29579,N_22614,N_22267);
or U29580 (N_29580,N_20603,N_21932);
or U29581 (N_29581,N_23929,N_22965);
or U29582 (N_29582,N_23631,N_24454);
nand U29583 (N_29583,N_20545,N_21308);
nand U29584 (N_29584,N_22043,N_24616);
xnor U29585 (N_29585,N_23647,N_20407);
nor U29586 (N_29586,N_20968,N_20237);
xor U29587 (N_29587,N_21172,N_22792);
or U29588 (N_29588,N_21672,N_21739);
xor U29589 (N_29589,N_21694,N_23575);
xnor U29590 (N_29590,N_23348,N_23854);
xor U29591 (N_29591,N_21009,N_24773);
and U29592 (N_29592,N_20316,N_21660);
or U29593 (N_29593,N_22052,N_20862);
and U29594 (N_29594,N_20781,N_23521);
nor U29595 (N_29595,N_23200,N_20940);
nor U29596 (N_29596,N_23140,N_20173);
or U29597 (N_29597,N_23648,N_23125);
nand U29598 (N_29598,N_23359,N_20776);
nand U29599 (N_29599,N_24458,N_21526);
nor U29600 (N_29600,N_23946,N_23487);
xor U29601 (N_29601,N_21807,N_24410);
nor U29602 (N_29602,N_23340,N_23604);
nand U29603 (N_29603,N_22363,N_24146);
or U29604 (N_29604,N_23157,N_24434);
and U29605 (N_29605,N_24685,N_24613);
or U29606 (N_29606,N_20753,N_23584);
nor U29607 (N_29607,N_21140,N_22166);
or U29608 (N_29608,N_24459,N_24533);
or U29609 (N_29609,N_24188,N_20945);
nand U29610 (N_29610,N_20401,N_20788);
xor U29611 (N_29611,N_23190,N_23269);
nor U29612 (N_29612,N_24676,N_23757);
nand U29613 (N_29613,N_20866,N_23580);
and U29614 (N_29614,N_21160,N_21593);
xnor U29615 (N_29615,N_24328,N_23249);
or U29616 (N_29616,N_20573,N_20532);
and U29617 (N_29617,N_20583,N_23459);
or U29618 (N_29618,N_24227,N_22183);
or U29619 (N_29619,N_22668,N_21338);
nand U29620 (N_29620,N_20025,N_24889);
nor U29621 (N_29621,N_21539,N_23598);
nor U29622 (N_29622,N_23276,N_20667);
nor U29623 (N_29623,N_21653,N_24430);
or U29624 (N_29624,N_24769,N_22630);
or U29625 (N_29625,N_20597,N_23944);
nor U29626 (N_29626,N_22781,N_22913);
xor U29627 (N_29627,N_22581,N_21914);
nor U29628 (N_29628,N_22102,N_21576);
nand U29629 (N_29629,N_20778,N_20948);
and U29630 (N_29630,N_23495,N_24891);
or U29631 (N_29631,N_23152,N_22151);
xnor U29632 (N_29632,N_21317,N_23879);
or U29633 (N_29633,N_23608,N_24609);
and U29634 (N_29634,N_21954,N_21560);
xnor U29635 (N_29635,N_24516,N_23038);
nand U29636 (N_29636,N_22826,N_22223);
nand U29637 (N_29637,N_23133,N_20051);
and U29638 (N_29638,N_20198,N_23802);
or U29639 (N_29639,N_23469,N_23997);
or U29640 (N_29640,N_20848,N_21620);
nor U29641 (N_29641,N_22278,N_21544);
nand U29642 (N_29642,N_24802,N_21152);
nand U29643 (N_29643,N_23161,N_24575);
nand U29644 (N_29644,N_23182,N_22576);
nor U29645 (N_29645,N_20166,N_24133);
or U29646 (N_29646,N_24748,N_23127);
nand U29647 (N_29647,N_23088,N_22583);
and U29648 (N_29648,N_22553,N_23928);
and U29649 (N_29649,N_21205,N_21798);
and U29650 (N_29650,N_21021,N_23243);
and U29651 (N_29651,N_20278,N_22282);
or U29652 (N_29652,N_21163,N_21761);
nand U29653 (N_29653,N_23235,N_22202);
nor U29654 (N_29654,N_20566,N_22883);
or U29655 (N_29655,N_22138,N_24398);
and U29656 (N_29656,N_21971,N_22697);
or U29657 (N_29657,N_21402,N_20955);
or U29658 (N_29658,N_20040,N_21101);
nand U29659 (N_29659,N_20646,N_22104);
xor U29660 (N_29660,N_24991,N_21691);
nor U29661 (N_29661,N_22532,N_23865);
nor U29662 (N_29662,N_23461,N_23504);
nand U29663 (N_29663,N_23823,N_20105);
xor U29664 (N_29664,N_22284,N_20395);
and U29665 (N_29665,N_20217,N_22042);
nand U29666 (N_29666,N_22595,N_20415);
nand U29667 (N_29667,N_24672,N_22124);
or U29668 (N_29668,N_22060,N_21447);
xnor U29669 (N_29669,N_20596,N_20501);
nand U29670 (N_29670,N_22503,N_22806);
and U29671 (N_29671,N_23231,N_22217);
and U29672 (N_29672,N_20991,N_21440);
nor U29673 (N_29673,N_22073,N_23984);
nor U29674 (N_29674,N_23014,N_21999);
or U29675 (N_29675,N_21686,N_24215);
nor U29676 (N_29676,N_23797,N_21245);
and U29677 (N_29677,N_21123,N_20269);
or U29678 (N_29678,N_21238,N_23153);
xor U29679 (N_29679,N_22696,N_21992);
and U29680 (N_29680,N_22978,N_20748);
and U29681 (N_29681,N_24371,N_22543);
and U29682 (N_29682,N_21024,N_21004);
and U29683 (N_29683,N_22030,N_22970);
or U29684 (N_29684,N_23713,N_21919);
and U29685 (N_29685,N_24532,N_23245);
or U29686 (N_29686,N_20720,N_20716);
nand U29687 (N_29687,N_21719,N_20891);
or U29688 (N_29688,N_21449,N_20804);
and U29689 (N_29689,N_22767,N_20854);
nand U29690 (N_29690,N_21433,N_21368);
and U29691 (N_29691,N_24113,N_24760);
nand U29692 (N_29692,N_23969,N_22719);
xor U29693 (N_29693,N_22848,N_20902);
nand U29694 (N_29694,N_24406,N_22342);
or U29695 (N_29695,N_20572,N_20901);
and U29696 (N_29696,N_20834,N_20753);
nand U29697 (N_29697,N_21477,N_20297);
nor U29698 (N_29698,N_21846,N_24863);
or U29699 (N_29699,N_22031,N_24195);
and U29700 (N_29700,N_24465,N_23503);
and U29701 (N_29701,N_24336,N_24835);
xnor U29702 (N_29702,N_22869,N_20540);
nor U29703 (N_29703,N_21090,N_21451);
xor U29704 (N_29704,N_22857,N_20490);
or U29705 (N_29705,N_21651,N_22606);
nand U29706 (N_29706,N_20540,N_22967);
and U29707 (N_29707,N_21137,N_22621);
nor U29708 (N_29708,N_20215,N_21381);
and U29709 (N_29709,N_23105,N_20227);
nor U29710 (N_29710,N_22160,N_20305);
nand U29711 (N_29711,N_24294,N_22571);
and U29712 (N_29712,N_23436,N_22367);
nor U29713 (N_29713,N_20906,N_24684);
xor U29714 (N_29714,N_22854,N_22160);
nand U29715 (N_29715,N_23274,N_21792);
xor U29716 (N_29716,N_21600,N_21941);
nor U29717 (N_29717,N_24277,N_23432);
xnor U29718 (N_29718,N_24344,N_22095);
xor U29719 (N_29719,N_23046,N_22912);
nor U29720 (N_29720,N_23734,N_24562);
nand U29721 (N_29721,N_21969,N_21456);
xor U29722 (N_29722,N_21035,N_20505);
and U29723 (N_29723,N_20098,N_24465);
xor U29724 (N_29724,N_21807,N_20355);
nor U29725 (N_29725,N_22286,N_20948);
and U29726 (N_29726,N_20934,N_22188);
nand U29727 (N_29727,N_20199,N_22075);
or U29728 (N_29728,N_21137,N_20903);
xor U29729 (N_29729,N_21863,N_23419);
or U29730 (N_29730,N_22454,N_23952);
and U29731 (N_29731,N_21779,N_22640);
nand U29732 (N_29732,N_23515,N_23344);
and U29733 (N_29733,N_23832,N_23262);
or U29734 (N_29734,N_24670,N_21312);
or U29735 (N_29735,N_21135,N_23843);
nor U29736 (N_29736,N_22066,N_20559);
and U29737 (N_29737,N_20889,N_24849);
nand U29738 (N_29738,N_23370,N_20169);
and U29739 (N_29739,N_24293,N_20897);
nand U29740 (N_29740,N_21040,N_24870);
and U29741 (N_29741,N_24622,N_20412);
or U29742 (N_29742,N_24962,N_22869);
and U29743 (N_29743,N_21102,N_24506);
or U29744 (N_29744,N_22766,N_20285);
or U29745 (N_29745,N_21627,N_21580);
nor U29746 (N_29746,N_23741,N_24600);
and U29747 (N_29747,N_20108,N_21225);
or U29748 (N_29748,N_21278,N_23178);
and U29749 (N_29749,N_22356,N_21974);
nand U29750 (N_29750,N_20544,N_21936);
or U29751 (N_29751,N_20786,N_21532);
and U29752 (N_29752,N_24299,N_22608);
nor U29753 (N_29753,N_23788,N_23777);
xor U29754 (N_29754,N_20429,N_22326);
nand U29755 (N_29755,N_21084,N_23234);
nand U29756 (N_29756,N_23178,N_23855);
or U29757 (N_29757,N_21175,N_21403);
nand U29758 (N_29758,N_20184,N_21641);
xnor U29759 (N_29759,N_24247,N_21915);
nor U29760 (N_29760,N_20844,N_24141);
or U29761 (N_29761,N_24544,N_20037);
or U29762 (N_29762,N_24136,N_22805);
xnor U29763 (N_29763,N_21916,N_22221);
nand U29764 (N_29764,N_20525,N_24124);
nor U29765 (N_29765,N_20887,N_24556);
xnor U29766 (N_29766,N_23750,N_20300);
and U29767 (N_29767,N_23578,N_22968);
nor U29768 (N_29768,N_23485,N_24805);
nand U29769 (N_29769,N_21932,N_22749);
xnor U29770 (N_29770,N_22501,N_20319);
and U29771 (N_29771,N_24482,N_24900);
and U29772 (N_29772,N_22336,N_20469);
nand U29773 (N_29773,N_21615,N_24132);
nand U29774 (N_29774,N_22790,N_23366);
nand U29775 (N_29775,N_20254,N_23012);
or U29776 (N_29776,N_24176,N_21965);
nor U29777 (N_29777,N_21644,N_22898);
or U29778 (N_29778,N_21639,N_23124);
xor U29779 (N_29779,N_22982,N_22289);
and U29780 (N_29780,N_22846,N_22647);
or U29781 (N_29781,N_24227,N_20834);
or U29782 (N_29782,N_23462,N_22935);
xor U29783 (N_29783,N_24612,N_21998);
and U29784 (N_29784,N_20998,N_24147);
nor U29785 (N_29785,N_20046,N_21924);
or U29786 (N_29786,N_21256,N_20632);
or U29787 (N_29787,N_20332,N_20752);
nor U29788 (N_29788,N_24985,N_20816);
nor U29789 (N_29789,N_21025,N_23070);
xnor U29790 (N_29790,N_23252,N_20101);
nor U29791 (N_29791,N_20229,N_23518);
nor U29792 (N_29792,N_21264,N_22210);
nor U29793 (N_29793,N_20646,N_22058);
xnor U29794 (N_29794,N_21655,N_20728);
xor U29795 (N_29795,N_21621,N_23001);
and U29796 (N_29796,N_23753,N_24846);
or U29797 (N_29797,N_24458,N_23725);
nand U29798 (N_29798,N_21441,N_21526);
nor U29799 (N_29799,N_21417,N_24013);
xor U29800 (N_29800,N_21064,N_20770);
and U29801 (N_29801,N_21353,N_24692);
and U29802 (N_29802,N_20243,N_21922);
nand U29803 (N_29803,N_24420,N_20403);
nand U29804 (N_29804,N_20352,N_21725);
or U29805 (N_29805,N_20434,N_22235);
nand U29806 (N_29806,N_21055,N_22727);
xnor U29807 (N_29807,N_20505,N_24873);
nor U29808 (N_29808,N_22518,N_24109);
xor U29809 (N_29809,N_23957,N_23589);
nand U29810 (N_29810,N_22390,N_24417);
nand U29811 (N_29811,N_21220,N_22390);
or U29812 (N_29812,N_20575,N_22595);
or U29813 (N_29813,N_23583,N_24568);
and U29814 (N_29814,N_23228,N_20997);
nor U29815 (N_29815,N_22848,N_22238);
xnor U29816 (N_29816,N_20548,N_23045);
xor U29817 (N_29817,N_23991,N_24726);
nor U29818 (N_29818,N_23495,N_24257);
and U29819 (N_29819,N_21640,N_21074);
xor U29820 (N_29820,N_23268,N_21865);
and U29821 (N_29821,N_24869,N_21095);
xor U29822 (N_29822,N_20805,N_21581);
or U29823 (N_29823,N_20432,N_21374);
and U29824 (N_29824,N_23376,N_20149);
nand U29825 (N_29825,N_22354,N_24499);
xor U29826 (N_29826,N_23505,N_21940);
or U29827 (N_29827,N_24199,N_21944);
or U29828 (N_29828,N_20778,N_24626);
and U29829 (N_29829,N_22619,N_22811);
or U29830 (N_29830,N_23664,N_22732);
nand U29831 (N_29831,N_23973,N_20088);
nor U29832 (N_29832,N_21262,N_21935);
xnor U29833 (N_29833,N_21858,N_20541);
nor U29834 (N_29834,N_23329,N_20419);
xor U29835 (N_29835,N_22313,N_24839);
nand U29836 (N_29836,N_21518,N_21235);
xnor U29837 (N_29837,N_24788,N_21958);
xnor U29838 (N_29838,N_24569,N_20388);
xor U29839 (N_29839,N_24819,N_21051);
nor U29840 (N_29840,N_21800,N_20621);
or U29841 (N_29841,N_23172,N_22022);
nand U29842 (N_29842,N_23393,N_23165);
xnor U29843 (N_29843,N_21838,N_22908);
or U29844 (N_29844,N_21947,N_20890);
or U29845 (N_29845,N_24402,N_24424);
xnor U29846 (N_29846,N_20916,N_21356);
nor U29847 (N_29847,N_22380,N_21467);
or U29848 (N_29848,N_23958,N_23606);
nand U29849 (N_29849,N_24576,N_22982);
xor U29850 (N_29850,N_24671,N_24572);
xnor U29851 (N_29851,N_23959,N_23495);
nor U29852 (N_29852,N_23023,N_21998);
xor U29853 (N_29853,N_21145,N_21519);
xor U29854 (N_29854,N_20981,N_23640);
and U29855 (N_29855,N_23149,N_23054);
or U29856 (N_29856,N_22020,N_22479);
or U29857 (N_29857,N_20541,N_20754);
and U29858 (N_29858,N_20436,N_20968);
xor U29859 (N_29859,N_21142,N_22343);
nor U29860 (N_29860,N_24615,N_20549);
nand U29861 (N_29861,N_24194,N_23322);
nand U29862 (N_29862,N_21631,N_22219);
and U29863 (N_29863,N_22653,N_24190);
nand U29864 (N_29864,N_24491,N_21026);
or U29865 (N_29865,N_23149,N_22974);
and U29866 (N_29866,N_22415,N_24337);
nand U29867 (N_29867,N_24554,N_20832);
nand U29868 (N_29868,N_20130,N_22463);
xor U29869 (N_29869,N_23588,N_22866);
nand U29870 (N_29870,N_21590,N_23817);
xor U29871 (N_29871,N_21023,N_21367);
or U29872 (N_29872,N_21163,N_22063);
or U29873 (N_29873,N_24446,N_20778);
nand U29874 (N_29874,N_23887,N_23656);
nor U29875 (N_29875,N_23673,N_23574);
or U29876 (N_29876,N_20070,N_21858);
xnor U29877 (N_29877,N_21358,N_20295);
nor U29878 (N_29878,N_23918,N_22367);
or U29879 (N_29879,N_21352,N_20474);
xnor U29880 (N_29880,N_21297,N_22216);
xnor U29881 (N_29881,N_23833,N_21166);
or U29882 (N_29882,N_22303,N_22142);
xor U29883 (N_29883,N_24232,N_22313);
and U29884 (N_29884,N_24231,N_22881);
and U29885 (N_29885,N_21585,N_21522);
nand U29886 (N_29886,N_22963,N_23262);
xnor U29887 (N_29887,N_23819,N_23063);
and U29888 (N_29888,N_23940,N_21918);
and U29889 (N_29889,N_21708,N_23525);
nand U29890 (N_29890,N_21178,N_23566);
xor U29891 (N_29891,N_23306,N_23928);
nor U29892 (N_29892,N_21758,N_24640);
and U29893 (N_29893,N_21646,N_23599);
nor U29894 (N_29894,N_23743,N_23496);
nor U29895 (N_29895,N_23904,N_21899);
nand U29896 (N_29896,N_20508,N_22448);
nand U29897 (N_29897,N_23354,N_20756);
and U29898 (N_29898,N_24831,N_24943);
xnor U29899 (N_29899,N_23368,N_20185);
nand U29900 (N_29900,N_20124,N_23331);
nor U29901 (N_29901,N_22071,N_23270);
or U29902 (N_29902,N_20019,N_24159);
and U29903 (N_29903,N_20196,N_21323);
or U29904 (N_29904,N_24117,N_24273);
nor U29905 (N_29905,N_23001,N_22614);
or U29906 (N_29906,N_20681,N_22822);
or U29907 (N_29907,N_20585,N_23217);
and U29908 (N_29908,N_23010,N_20626);
and U29909 (N_29909,N_23116,N_20832);
and U29910 (N_29910,N_24117,N_22368);
nand U29911 (N_29911,N_23346,N_21470);
nor U29912 (N_29912,N_24836,N_22278);
or U29913 (N_29913,N_21192,N_22795);
xor U29914 (N_29914,N_21119,N_23980);
or U29915 (N_29915,N_23962,N_24157);
nand U29916 (N_29916,N_21601,N_22989);
nor U29917 (N_29917,N_22366,N_20584);
nor U29918 (N_29918,N_24171,N_24806);
nor U29919 (N_29919,N_21684,N_22204);
and U29920 (N_29920,N_24642,N_20613);
nand U29921 (N_29921,N_21540,N_22201);
or U29922 (N_29922,N_24496,N_21446);
xnor U29923 (N_29923,N_24654,N_20699);
and U29924 (N_29924,N_24596,N_20365);
xnor U29925 (N_29925,N_20502,N_22301);
nor U29926 (N_29926,N_24404,N_24123);
and U29927 (N_29927,N_23442,N_23580);
nor U29928 (N_29928,N_23086,N_24004);
and U29929 (N_29929,N_21921,N_23107);
or U29930 (N_29930,N_21379,N_21745);
nor U29931 (N_29931,N_23502,N_22223);
nor U29932 (N_29932,N_20611,N_23383);
nand U29933 (N_29933,N_23592,N_20819);
xnor U29934 (N_29934,N_22512,N_22932);
nor U29935 (N_29935,N_23393,N_20327);
xnor U29936 (N_29936,N_21649,N_20754);
or U29937 (N_29937,N_22558,N_23803);
xor U29938 (N_29938,N_22329,N_21318);
and U29939 (N_29939,N_22744,N_24805);
nor U29940 (N_29940,N_23691,N_20119);
nor U29941 (N_29941,N_21168,N_23853);
xnor U29942 (N_29942,N_23445,N_22057);
or U29943 (N_29943,N_23034,N_24294);
xor U29944 (N_29944,N_23665,N_22907);
nor U29945 (N_29945,N_23301,N_24585);
or U29946 (N_29946,N_24777,N_22214);
xnor U29947 (N_29947,N_23448,N_23821);
nor U29948 (N_29948,N_21628,N_23141);
nand U29949 (N_29949,N_24318,N_23014);
or U29950 (N_29950,N_24493,N_24858);
nor U29951 (N_29951,N_22418,N_24413);
and U29952 (N_29952,N_21235,N_23835);
and U29953 (N_29953,N_21507,N_23808);
or U29954 (N_29954,N_20225,N_20529);
xor U29955 (N_29955,N_23842,N_23346);
or U29956 (N_29956,N_20222,N_23952);
and U29957 (N_29957,N_23898,N_24909);
nor U29958 (N_29958,N_23386,N_21343);
nor U29959 (N_29959,N_24480,N_21657);
nor U29960 (N_29960,N_22417,N_22024);
or U29961 (N_29961,N_24322,N_20033);
and U29962 (N_29962,N_23419,N_20097);
or U29963 (N_29963,N_20971,N_22830);
or U29964 (N_29964,N_21127,N_20286);
xor U29965 (N_29965,N_23247,N_21688);
nand U29966 (N_29966,N_24628,N_23309);
or U29967 (N_29967,N_24874,N_23615);
or U29968 (N_29968,N_20121,N_21185);
xor U29969 (N_29969,N_21444,N_21860);
and U29970 (N_29970,N_21201,N_21118);
nor U29971 (N_29971,N_24826,N_21052);
nand U29972 (N_29972,N_23017,N_24238);
nor U29973 (N_29973,N_20781,N_20027);
xor U29974 (N_29974,N_20643,N_20223);
xor U29975 (N_29975,N_22711,N_20353);
and U29976 (N_29976,N_23685,N_20832);
nor U29977 (N_29977,N_23328,N_24649);
and U29978 (N_29978,N_24934,N_21870);
nor U29979 (N_29979,N_21914,N_20343);
nor U29980 (N_29980,N_21943,N_20585);
nor U29981 (N_29981,N_20741,N_23024);
and U29982 (N_29982,N_21164,N_23106);
xor U29983 (N_29983,N_21705,N_23989);
or U29984 (N_29984,N_23971,N_22061);
or U29985 (N_29985,N_20312,N_22170);
or U29986 (N_29986,N_21539,N_21102);
nand U29987 (N_29987,N_21012,N_24220);
and U29988 (N_29988,N_24425,N_20593);
nand U29989 (N_29989,N_23239,N_20792);
xor U29990 (N_29990,N_20245,N_20856);
xor U29991 (N_29991,N_22007,N_20174);
or U29992 (N_29992,N_24152,N_23344);
nand U29993 (N_29993,N_20016,N_21371);
nor U29994 (N_29994,N_20518,N_20763);
xor U29995 (N_29995,N_21143,N_24869);
and U29996 (N_29996,N_21219,N_20106);
nand U29997 (N_29997,N_22049,N_22401);
and U29998 (N_29998,N_20965,N_24367);
and U29999 (N_29999,N_23235,N_22701);
nor UO_0 (O_0,N_29925,N_28701);
and UO_1 (O_1,N_27473,N_26799);
xnor UO_2 (O_2,N_26526,N_27936);
nor UO_3 (O_3,N_25984,N_26516);
xor UO_4 (O_4,N_29545,N_27318);
and UO_5 (O_5,N_29717,N_25847);
nand UO_6 (O_6,N_25795,N_25176);
nor UO_7 (O_7,N_28871,N_29492);
xnor UO_8 (O_8,N_28860,N_29824);
nand UO_9 (O_9,N_29100,N_25724);
xnor UO_10 (O_10,N_27345,N_29738);
or UO_11 (O_11,N_29047,N_25899);
nor UO_12 (O_12,N_25565,N_28094);
nor UO_13 (O_13,N_28543,N_28633);
nor UO_14 (O_14,N_25946,N_27464);
nor UO_15 (O_15,N_26333,N_29860);
or UO_16 (O_16,N_26861,N_26590);
and UO_17 (O_17,N_27928,N_29064);
nor UO_18 (O_18,N_28341,N_27064);
nor UO_19 (O_19,N_25287,N_25369);
nor UO_20 (O_20,N_26462,N_29097);
nor UO_21 (O_21,N_28625,N_26910);
nand UO_22 (O_22,N_26903,N_28529);
and UO_23 (O_23,N_25943,N_26334);
and UO_24 (O_24,N_26427,N_26052);
nor UO_25 (O_25,N_26351,N_27522);
xnor UO_26 (O_26,N_27149,N_27783);
xor UO_27 (O_27,N_25342,N_26500);
nand UO_28 (O_28,N_28746,N_25221);
nand UO_29 (O_29,N_26827,N_29179);
nor UO_30 (O_30,N_29940,N_26814);
and UO_31 (O_31,N_25508,N_26485);
nor UO_32 (O_32,N_25306,N_28904);
nand UO_33 (O_33,N_26089,N_28219);
nor UO_34 (O_34,N_29266,N_29536);
nor UO_35 (O_35,N_26320,N_28009);
or UO_36 (O_36,N_27301,N_27240);
nand UO_37 (O_37,N_27135,N_29283);
nor UO_38 (O_38,N_29051,N_25875);
or UO_39 (O_39,N_29389,N_28263);
nand UO_40 (O_40,N_28235,N_25307);
nand UO_41 (O_41,N_26640,N_29515);
nor UO_42 (O_42,N_29714,N_25750);
and UO_43 (O_43,N_25643,N_29092);
or UO_44 (O_44,N_27644,N_28544);
nand UO_45 (O_45,N_25671,N_29247);
nor UO_46 (O_46,N_27577,N_28195);
and UO_47 (O_47,N_29629,N_26624);
xor UO_48 (O_48,N_25297,N_28878);
nor UO_49 (O_49,N_28946,N_25664);
and UO_50 (O_50,N_28022,N_26115);
or UO_51 (O_51,N_29317,N_28705);
nor UO_52 (O_52,N_28634,N_25361);
or UO_53 (O_53,N_25553,N_29391);
and UO_54 (O_54,N_25790,N_29954);
xnor UO_55 (O_55,N_25957,N_27799);
or UO_56 (O_56,N_25350,N_25763);
nor UO_57 (O_57,N_29110,N_29405);
or UO_58 (O_58,N_27435,N_25362);
and UO_59 (O_59,N_27333,N_28355);
and UO_60 (O_60,N_27676,N_28794);
nand UO_61 (O_61,N_26033,N_28314);
xnor UO_62 (O_62,N_25700,N_29964);
nand UO_63 (O_63,N_27172,N_28295);
nor UO_64 (O_64,N_29140,N_26917);
or UO_65 (O_65,N_25405,N_27935);
nor UO_66 (O_66,N_26387,N_29206);
nand UO_67 (O_67,N_27750,N_27263);
xor UO_68 (O_68,N_29382,N_25239);
xnor UO_69 (O_69,N_25961,N_29188);
nor UO_70 (O_70,N_26330,N_26482);
xnor UO_71 (O_71,N_29335,N_29586);
nand UO_72 (O_72,N_27985,N_29640);
or UO_73 (O_73,N_25107,N_28498);
nand UO_74 (O_74,N_27252,N_26449);
xnor UO_75 (O_75,N_28863,N_29300);
nand UO_76 (O_76,N_26815,N_27698);
nand UO_77 (O_77,N_25608,N_29618);
nor UO_78 (O_78,N_26847,N_28364);
nor UO_79 (O_79,N_26786,N_29584);
nand UO_80 (O_80,N_28218,N_28367);
nand UO_81 (O_81,N_29921,N_26931);
nand UO_82 (O_82,N_29692,N_27626);
or UO_83 (O_83,N_26353,N_26593);
nand UO_84 (O_84,N_27290,N_28286);
and UO_85 (O_85,N_28053,N_29856);
nor UO_86 (O_86,N_27036,N_29022);
or UO_87 (O_87,N_27083,N_25662);
nand UO_88 (O_88,N_25436,N_25948);
or UO_89 (O_89,N_26774,N_25432);
and UO_90 (O_90,N_29747,N_29647);
and UO_91 (O_91,N_25916,N_29839);
or UO_92 (O_92,N_25595,N_27885);
xor UO_93 (O_93,N_28587,N_26388);
xor UO_94 (O_94,N_27631,N_26906);
xor UO_95 (O_95,N_26182,N_27490);
and UO_96 (O_96,N_29712,N_27023);
or UO_97 (O_97,N_25484,N_26397);
nor UO_98 (O_98,N_28636,N_28256);
and UO_99 (O_99,N_26629,N_27098);
or UO_100 (O_100,N_27510,N_28621);
or UO_101 (O_101,N_27743,N_28249);
nand UO_102 (O_102,N_29253,N_27923);
nand UO_103 (O_103,N_27168,N_28120);
nand UO_104 (O_104,N_27525,N_28895);
and UO_105 (O_105,N_26378,N_27071);
xor UO_106 (O_106,N_27370,N_29204);
or UO_107 (O_107,N_26776,N_26288);
or UO_108 (O_108,N_25157,N_27181);
and UO_109 (O_109,N_28958,N_26240);
nand UO_110 (O_110,N_28668,N_29819);
nand UO_111 (O_111,N_27331,N_25938);
nand UO_112 (O_112,N_27592,N_28266);
nand UO_113 (O_113,N_25618,N_26818);
and UO_114 (O_114,N_29522,N_29780);
and UO_115 (O_115,N_25151,N_25936);
nor UO_116 (O_116,N_28905,N_25966);
nand UO_117 (O_117,N_29018,N_29592);
and UO_118 (O_118,N_28005,N_28574);
or UO_119 (O_119,N_26015,N_25537);
xnor UO_120 (O_120,N_29828,N_28464);
xnor UO_121 (O_121,N_26731,N_28875);
nor UO_122 (O_122,N_26233,N_27894);
and UO_123 (O_123,N_25598,N_27983);
xnor UO_124 (O_124,N_27756,N_25979);
and UO_125 (O_125,N_28706,N_25744);
and UO_126 (O_126,N_28319,N_25516);
nor UO_127 (O_127,N_27237,N_27108);
and UO_128 (O_128,N_28399,N_25972);
and UO_129 (O_129,N_28952,N_28748);
xor UO_130 (O_130,N_29699,N_27326);
and UO_131 (O_131,N_26179,N_27578);
nand UO_132 (O_132,N_25403,N_25101);
nand UO_133 (O_133,N_25762,N_29128);
and UO_134 (O_134,N_25893,N_27657);
nor UO_135 (O_135,N_28615,N_25849);
xnor UO_136 (O_136,N_29636,N_27223);
and UO_137 (O_137,N_28977,N_27542);
nand UO_138 (O_138,N_29899,N_28043);
or UO_139 (O_139,N_27646,N_25100);
nand UO_140 (O_140,N_26669,N_29910);
nand UO_141 (O_141,N_26777,N_29285);
or UO_142 (O_142,N_29667,N_28788);
and UO_143 (O_143,N_29804,N_25329);
nor UO_144 (O_144,N_25973,N_25761);
xnor UO_145 (O_145,N_25850,N_29173);
and UO_146 (O_146,N_27161,N_27496);
xor UO_147 (O_147,N_26144,N_27664);
nand UO_148 (O_148,N_27685,N_29834);
and UO_149 (O_149,N_26087,N_27002);
and UO_150 (O_150,N_28530,N_28107);
nor UO_151 (O_151,N_25771,N_27014);
and UO_152 (O_152,N_27532,N_25816);
nand UO_153 (O_153,N_28976,N_26920);
nand UO_154 (O_154,N_27378,N_26783);
nand UO_155 (O_155,N_28929,N_26772);
xnor UO_156 (O_156,N_25424,N_29280);
and UO_157 (O_157,N_27017,N_29872);
nand UO_158 (O_158,N_25240,N_28606);
nand UO_159 (O_159,N_25788,N_25123);
or UO_160 (O_160,N_26909,N_25241);
nand UO_161 (O_161,N_26114,N_27896);
or UO_162 (O_162,N_25488,N_25862);
nor UO_163 (O_163,N_26242,N_25879);
nor UO_164 (O_164,N_28209,N_27277);
nand UO_165 (O_165,N_26996,N_26922);
xnor UO_166 (O_166,N_29024,N_28560);
and UO_167 (O_167,N_29124,N_29634);
or UO_168 (O_168,N_27294,N_28435);
xor UO_169 (O_169,N_28987,N_26307);
nor UO_170 (O_170,N_27786,N_28893);
xnor UO_171 (O_171,N_29044,N_26189);
nand UO_172 (O_172,N_28001,N_27120);
xor UO_173 (O_173,N_28371,N_27361);
nor UO_174 (O_174,N_27844,N_28911);
and UO_175 (O_175,N_25732,N_29996);
and UO_176 (O_176,N_29324,N_28801);
xnor UO_177 (O_177,N_25471,N_28690);
or UO_178 (O_178,N_27348,N_28796);
nor UO_179 (O_179,N_29086,N_28541);
nand UO_180 (O_180,N_27874,N_27125);
nand UO_181 (O_181,N_26675,N_25058);
nor UO_182 (O_182,N_27551,N_29531);
nand UO_183 (O_183,N_28052,N_28717);
or UO_184 (O_184,N_27570,N_29381);
nor UO_185 (O_185,N_25996,N_25854);
or UO_186 (O_186,N_29109,N_25443);
or UO_187 (O_187,N_25235,N_25170);
and UO_188 (O_188,N_25922,N_29347);
nor UO_189 (O_189,N_28630,N_29939);
or UO_190 (O_190,N_28756,N_27257);
and UO_191 (O_191,N_27797,N_25668);
nand UO_192 (O_192,N_28450,N_27207);
nand UO_193 (O_193,N_25346,N_25981);
nor UO_194 (O_194,N_27174,N_25060);
xnor UO_195 (O_195,N_29426,N_29526);
and UO_196 (O_196,N_25500,N_25962);
nor UO_197 (O_197,N_25498,N_29387);
and UO_198 (O_198,N_29552,N_26983);
or UO_199 (O_199,N_29931,N_28260);
nor UO_200 (O_200,N_29858,N_26444);
xnor UO_201 (O_201,N_29376,N_29581);
xor UO_202 (O_202,N_28859,N_26746);
or UO_203 (O_203,N_29924,N_28240);
or UO_204 (O_204,N_25428,N_29567);
or UO_205 (O_205,N_25673,N_28161);
and UO_206 (O_206,N_29183,N_25645);
nand UO_207 (O_207,N_25985,N_27085);
nand UO_208 (O_208,N_29811,N_28927);
nor UO_209 (O_209,N_25913,N_29332);
and UO_210 (O_210,N_26150,N_25928);
and UO_211 (O_211,N_28211,N_27892);
nor UO_212 (O_212,N_26941,N_25637);
xor UO_213 (O_213,N_26862,N_27735);
and UO_214 (O_214,N_25220,N_27443);
or UO_215 (O_215,N_29896,N_28106);
nor UO_216 (O_216,N_26030,N_28289);
or UO_217 (O_217,N_27600,N_25253);
or UO_218 (O_218,N_25709,N_29198);
and UO_219 (O_219,N_27933,N_28358);
nor UO_220 (O_220,N_25509,N_27792);
xnor UO_221 (O_221,N_28771,N_26771);
or UO_222 (O_222,N_28338,N_27707);
and UO_223 (O_223,N_28578,N_29455);
nand UO_224 (O_224,N_27654,N_29185);
and UO_225 (O_225,N_29609,N_26392);
and UO_226 (O_226,N_27506,N_26181);
nand UO_227 (O_227,N_26073,N_26788);
or UO_228 (O_228,N_26327,N_28956);
nand UO_229 (O_229,N_27701,N_27454);
and UO_230 (O_230,N_26702,N_26977);
xor UO_231 (O_231,N_25642,N_29123);
and UO_232 (O_232,N_29705,N_26391);
or UO_233 (O_233,N_27018,N_27068);
xnor UO_234 (O_234,N_27472,N_26721);
nand UO_235 (O_235,N_29637,N_27777);
nor UO_236 (O_236,N_27693,N_27813);
or UO_237 (O_237,N_27079,N_28718);
and UO_238 (O_238,N_26718,N_25791);
nand UO_239 (O_239,N_28309,N_25571);
and UO_240 (O_240,N_26328,N_26790);
xor UO_241 (O_241,N_26620,N_29386);
and UO_242 (O_242,N_27006,N_27820);
xor UO_243 (O_243,N_26113,N_27119);
nor UO_244 (O_244,N_28847,N_28590);
xnor UO_245 (O_245,N_26838,N_26231);
or UO_246 (O_246,N_28128,N_26987);
nand UO_247 (O_247,N_27480,N_28042);
xnor UO_248 (O_248,N_28000,N_29554);
and UO_249 (O_249,N_26681,N_28817);
or UO_250 (O_250,N_25734,N_25782);
nand UO_251 (O_251,N_29416,N_27846);
nor UO_252 (O_252,N_28025,N_29434);
and UO_253 (O_253,N_26876,N_26321);
xnor UO_254 (O_254,N_27711,N_27779);
nor UO_255 (O_255,N_27200,N_27955);
or UO_256 (O_256,N_25908,N_29116);
nor UO_257 (O_257,N_26759,N_27359);
nand UO_258 (O_258,N_28168,N_26365);
nand UO_259 (O_259,N_29762,N_25356);
and UO_260 (O_260,N_25939,N_27310);
and UO_261 (O_261,N_25841,N_29080);
and UO_262 (O_262,N_29916,N_25259);
and UO_263 (O_263,N_28045,N_29686);
nand UO_264 (O_264,N_29431,N_26588);
nand UO_265 (O_265,N_27791,N_26745);
xor UO_266 (O_266,N_26550,N_26125);
nand UO_267 (O_267,N_25703,N_25682);
nand UO_268 (O_268,N_26456,N_25839);
nor UO_269 (O_269,N_29418,N_29849);
nand UO_270 (O_270,N_28248,N_28844);
nor UO_271 (O_271,N_25396,N_27233);
nand UO_272 (O_272,N_28620,N_26698);
nor UO_273 (O_273,N_28509,N_29457);
xor UO_274 (O_274,N_25217,N_29749);
xnor UO_275 (O_275,N_27030,N_28599);
nand UO_276 (O_276,N_26200,N_25942);
nand UO_277 (O_277,N_28992,N_29730);
xor UO_278 (O_278,N_29371,N_26896);
nor UO_279 (O_279,N_25872,N_26578);
nand UO_280 (O_280,N_28826,N_26592);
nor UO_281 (O_281,N_27478,N_25360);
nand UO_282 (O_282,N_26406,N_27145);
nand UO_283 (O_283,N_28692,N_28362);
or UO_284 (O_284,N_28466,N_27548);
nand UO_285 (O_285,N_26763,N_27970);
nand UO_286 (O_286,N_25310,N_27619);
or UO_287 (O_287,N_25583,N_25377);
and UO_288 (O_288,N_26558,N_26540);
and UO_289 (O_289,N_25502,N_28051);
and UO_290 (O_290,N_26897,N_27497);
nor UO_291 (O_291,N_29721,N_26341);
nor UO_292 (O_292,N_28215,N_26061);
nand UO_293 (O_293,N_28657,N_26800);
nor UO_294 (O_294,N_25937,N_28184);
xor UO_295 (O_295,N_27856,N_27109);
or UO_296 (O_296,N_28872,N_25345);
or UO_297 (O_297,N_26904,N_26178);
nand UO_298 (O_298,N_25274,N_27298);
nor UO_299 (O_299,N_27710,N_28262);
and UO_300 (O_300,N_29467,N_27516);
nor UO_301 (O_301,N_27765,N_26562);
xor UO_302 (O_302,N_29241,N_25006);
and UO_303 (O_303,N_29155,N_25089);
or UO_304 (O_304,N_29299,N_25601);
and UO_305 (O_305,N_27709,N_26632);
xor UO_306 (O_306,N_27772,N_29569);
or UO_307 (O_307,N_28583,N_27686);
or UO_308 (O_308,N_26945,N_26937);
and UO_309 (O_309,N_28789,N_25534);
and UO_310 (O_310,N_25906,N_25786);
and UO_311 (O_311,N_29069,N_27342);
or UO_312 (O_312,N_26149,N_29913);
xor UO_313 (O_313,N_27214,N_29950);
xor UO_314 (O_314,N_29139,N_28959);
and UO_315 (O_315,N_27533,N_28348);
nor UO_316 (O_316,N_26374,N_28743);
xor UO_317 (O_317,N_27261,N_29679);
nor UO_318 (O_318,N_28004,N_26158);
or UO_319 (O_319,N_26175,N_28516);
xor UO_320 (O_320,N_29665,N_28199);
xnor UO_321 (O_321,N_29559,N_27192);
and UO_322 (O_322,N_28158,N_27862);
xor UO_323 (O_323,N_27387,N_29703);
and UO_324 (O_324,N_29876,N_26968);
nor UO_325 (O_325,N_28834,N_29658);
nand UO_326 (O_326,N_28963,N_29760);
xnor UO_327 (O_327,N_25382,N_28152);
xor UO_328 (O_328,N_27891,N_27875);
nand UO_329 (O_329,N_28499,N_25320);
nor UO_330 (O_330,N_28444,N_27971);
xor UO_331 (O_331,N_25232,N_26532);
or UO_332 (O_332,N_27332,N_25808);
and UO_333 (O_333,N_25557,N_29713);
nand UO_334 (O_334,N_28515,N_29944);
or UO_335 (O_335,N_27226,N_28588);
nor UO_336 (O_336,N_28411,N_28994);
nand UO_337 (O_337,N_27211,N_28085);
and UO_338 (O_338,N_26657,N_29566);
and UO_339 (O_339,N_26311,N_29011);
nor UO_340 (O_340,N_29904,N_26964);
nand UO_341 (O_341,N_27315,N_28949);
and UO_342 (O_342,N_25202,N_28484);
and UO_343 (O_343,N_27637,N_29920);
nor UO_344 (O_344,N_28334,N_25506);
nor UO_345 (O_345,N_26697,N_25820);
nand UO_346 (O_346,N_26716,N_27058);
xnor UO_347 (O_347,N_26643,N_26118);
or UO_348 (O_348,N_26907,N_29898);
nand UO_349 (O_349,N_28374,N_28637);
and UO_350 (O_350,N_27782,N_25780);
or UO_351 (O_351,N_25331,N_26618);
nand UO_352 (O_352,N_29257,N_28781);
nand UO_353 (O_353,N_26614,N_28137);
or UO_354 (O_354,N_29893,N_25366);
or UO_355 (O_355,N_26544,N_25125);
or UO_356 (O_356,N_25723,N_29107);
and UO_357 (O_357,N_25332,N_28275);
xnor UO_358 (O_358,N_25927,N_29114);
or UO_359 (O_359,N_27501,N_26025);
nand UO_360 (O_360,N_29468,N_27405);
nand UO_361 (O_361,N_27817,N_26266);
nand UO_362 (O_362,N_28500,N_25929);
nand UO_363 (O_363,N_26993,N_27680);
and UO_364 (O_364,N_29082,N_29776);
nor UO_365 (O_365,N_27216,N_26963);
nor UO_366 (O_366,N_28505,N_25654);
nand UO_367 (O_367,N_28322,N_29883);
nor UO_368 (O_368,N_26258,N_25002);
or UO_369 (O_369,N_28386,N_27751);
and UO_370 (O_370,N_29422,N_29682);
nor UO_371 (O_371,N_25691,N_26841);
nor UO_372 (O_372,N_27809,N_26802);
and UO_373 (O_373,N_28127,N_25144);
nor UO_374 (O_374,N_29981,N_27430);
xnor UO_375 (O_375,N_26140,N_27982);
and UO_376 (O_376,N_27581,N_25683);
and UO_377 (O_377,N_27273,N_28501);
xor UO_378 (O_378,N_25080,N_25930);
xnor UO_379 (O_379,N_26076,N_29252);
xnor UO_380 (O_380,N_29025,N_27732);
nand UO_381 (O_381,N_29725,N_26913);
nor UO_382 (O_382,N_25475,N_28869);
nor UO_383 (O_383,N_25309,N_27544);
xor UO_384 (O_384,N_27001,N_26713);
and UO_385 (O_385,N_27645,N_28575);
nor UO_386 (O_386,N_28613,N_27402);
or UO_387 (O_387,N_28317,N_29163);
or UO_388 (O_388,N_26335,N_28017);
and UO_389 (O_389,N_27814,N_27700);
nor UO_390 (O_390,N_28084,N_29167);
or UO_391 (O_391,N_28713,N_25255);
nand UO_392 (O_392,N_26092,N_25900);
nand UO_393 (O_393,N_29187,N_29953);
nor UO_394 (O_394,N_26960,N_27024);
xnor UO_395 (O_395,N_26433,N_27804);
and UO_396 (O_396,N_26944,N_25798);
nand UO_397 (O_397,N_29164,N_29832);
or UO_398 (O_398,N_28397,N_27563);
or UO_399 (O_399,N_26574,N_25825);
xor UO_400 (O_400,N_26429,N_27139);
xor UO_401 (O_401,N_26217,N_26357);
nor UO_402 (O_402,N_27433,N_29678);
or UO_403 (O_403,N_29708,N_29957);
and UO_404 (O_404,N_25234,N_26974);
or UO_405 (O_405,N_25019,N_27962);
or UO_406 (O_406,N_28350,N_28193);
nand UO_407 (O_407,N_28721,N_27111);
xnor UO_408 (O_408,N_26020,N_25884);
nand UO_409 (O_409,N_27748,N_27746);
and UO_410 (O_410,N_28975,N_25053);
and UO_411 (O_411,N_25237,N_29835);
nand UO_412 (O_412,N_29030,N_27587);
and UO_413 (O_413,N_27228,N_28594);
xor UO_414 (O_414,N_27594,N_28178);
or UO_415 (O_415,N_29734,N_29494);
and UO_416 (O_416,N_27458,N_25215);
or UO_417 (O_417,N_27210,N_26770);
nand UO_418 (O_418,N_26890,N_27288);
xor UO_419 (O_419,N_27988,N_26642);
nand UO_420 (O_420,N_26637,N_25914);
xor UO_421 (O_421,N_27633,N_29937);
nand UO_422 (O_422,N_25200,N_27967);
nor UO_423 (O_423,N_28420,N_27486);
or UO_424 (O_424,N_25415,N_27133);
or UO_425 (O_425,N_25052,N_27287);
or UO_426 (O_426,N_26159,N_25719);
or UO_427 (O_427,N_26256,N_27042);
nor UO_428 (O_428,N_25421,N_28308);
and UO_429 (O_429,N_25013,N_27840);
and UO_430 (O_430,N_25869,N_25273);
and UO_431 (O_431,N_29764,N_27218);
nand UO_432 (O_432,N_28778,N_28654);
or UO_433 (O_433,N_26893,N_27137);
nand UO_434 (O_434,N_25477,N_25667);
xor UO_435 (O_435,N_25876,N_29414);
and UO_436 (O_436,N_27423,N_26443);
nor UO_437 (O_437,N_25585,N_27785);
and UO_438 (O_438,N_27491,N_29960);
nand UO_439 (O_439,N_29877,N_29349);
nor UO_440 (O_440,N_25544,N_25931);
or UO_441 (O_441,N_26878,N_29604);
or UO_442 (O_442,N_26967,N_25828);
nor UO_443 (O_443,N_25755,N_27994);
and UO_444 (O_444,N_25041,N_26819);
or UO_445 (O_445,N_28730,N_29660);
or UO_446 (O_446,N_26916,N_26942);
or UO_447 (O_447,N_26930,N_25057);
and UO_448 (O_448,N_29078,N_29902);
xnor UO_449 (O_449,N_25472,N_28261);
or UO_450 (O_450,N_26650,N_28327);
nand UO_451 (O_451,N_29830,N_27078);
and UO_452 (O_452,N_27770,N_27830);
xor UO_453 (O_453,N_26739,N_28047);
nand UO_454 (O_454,N_25478,N_29650);
xor UO_455 (O_455,N_28431,N_27901);
xnor UO_456 (O_456,N_25017,N_29962);
or UO_457 (O_457,N_28907,N_25169);
and UO_458 (O_458,N_26290,N_28586);
or UO_459 (O_459,N_26733,N_27377);
xor UO_460 (O_460,N_26314,N_27417);
nand UO_461 (O_461,N_27066,N_27639);
or UO_462 (O_462,N_27759,N_29268);
nand UO_463 (O_463,N_29029,N_26728);
and UO_464 (O_464,N_26549,N_25614);
nand UO_465 (O_465,N_27324,N_27368);
nor UO_466 (O_466,N_29676,N_26091);
and UO_467 (O_467,N_28884,N_26660);
nand UO_468 (O_468,N_26059,N_27474);
nand UO_469 (O_469,N_25532,N_27255);
nor UO_470 (O_470,N_27169,N_28183);
nor UO_471 (O_471,N_26299,N_28091);
and UO_472 (O_472,N_25264,N_27725);
and UO_473 (O_473,N_25090,N_26938);
nand UO_474 (O_474,N_29499,N_29966);
nor UO_475 (O_475,N_28102,N_25247);
nand UO_476 (O_476,N_28438,N_27366);
nand UO_477 (O_477,N_25868,N_25395);
or UO_478 (O_478,N_28993,N_29008);
or UO_479 (O_479,N_26701,N_29793);
nand UO_480 (O_480,N_26208,N_26530);
or UO_481 (O_481,N_25848,N_29453);
nand UO_482 (O_482,N_26021,N_28745);
or UO_483 (O_483,N_29580,N_27339);
and UO_484 (O_484,N_29006,N_26292);
nand UO_485 (O_485,N_25865,N_26405);
or UO_486 (O_486,N_27268,N_27179);
and UO_487 (O_487,N_26889,N_29033);
or UO_488 (O_488,N_25552,N_26428);
xnor UO_489 (O_489,N_29224,N_25231);
xnor UO_490 (O_490,N_26738,N_29571);
nor UO_491 (O_491,N_28377,N_27566);
nand UO_492 (O_492,N_28930,N_29873);
nand UO_493 (O_493,N_27924,N_29974);
xor UO_494 (O_494,N_29121,N_26366);
or UO_495 (O_495,N_29067,N_28003);
or UO_496 (O_496,N_28873,N_28820);
nand UO_497 (O_497,N_25044,N_26204);
and UO_498 (O_498,N_28618,N_27107);
or UO_499 (O_499,N_26685,N_26817);
nor UO_500 (O_500,N_26779,N_29449);
nor UO_501 (O_501,N_29770,N_27527);
or UO_502 (O_502,N_28395,N_27100);
nand UO_503 (O_503,N_29134,N_26541);
xor UO_504 (O_504,N_29313,N_28252);
xnor UO_505 (O_505,N_26780,N_28156);
nand UO_506 (O_506,N_25097,N_25685);
xnor UO_507 (O_507,N_28551,N_29917);
or UO_508 (O_508,N_25684,N_28453);
and UO_509 (O_509,N_25735,N_27020);
or UO_510 (O_510,N_25610,N_29683);
xnor UO_511 (O_511,N_28809,N_28616);
or UO_512 (O_512,N_28276,N_27112);
nand UO_513 (O_513,N_29271,N_25776);
xnor UO_514 (O_514,N_28925,N_28101);
or UO_515 (O_515,N_26418,N_25263);
nor UO_516 (O_516,N_26582,N_29341);
or UO_517 (O_517,N_27457,N_27937);
nor UO_518 (O_518,N_27514,N_29845);
or UO_519 (O_519,N_26633,N_25246);
xor UO_520 (O_520,N_27302,N_27195);
and UO_521 (O_521,N_28458,N_27561);
nand UO_522 (O_522,N_29298,N_29942);
or UO_523 (O_523,N_25955,N_27056);
xor UO_524 (O_524,N_28130,N_27740);
xnor UO_525 (O_525,N_27659,N_26811);
and UO_526 (O_526,N_29918,N_26623);
xor UO_527 (O_527,N_28342,N_28422);
or UO_528 (O_528,N_27910,N_27373);
and UO_529 (O_529,N_27479,N_29158);
xnor UO_530 (O_530,N_28418,N_28175);
and UO_531 (O_531,N_28840,N_27934);
nand UO_532 (O_532,N_27309,N_26106);
xor UO_533 (O_533,N_29737,N_25450);
nor UO_534 (O_534,N_25286,N_28121);
nand UO_535 (O_535,N_29999,N_28092);
xnor UO_536 (O_536,N_27031,N_25122);
nor UO_537 (O_537,N_27374,N_27677);
and UO_538 (O_538,N_28792,N_26737);
and UO_539 (O_539,N_29000,N_27864);
or UO_540 (O_540,N_27199,N_25644);
nor UO_541 (O_541,N_25082,N_25034);
or UO_542 (O_542,N_27340,N_28080);
and UO_543 (O_543,N_26509,N_25406);
nor UO_544 (O_544,N_26111,N_29216);
xor UO_545 (O_545,N_26807,N_28361);
nor UO_546 (O_546,N_25230,N_26542);
nor UO_547 (O_547,N_27234,N_27666);
and UO_548 (O_548,N_27146,N_27660);
nor UO_549 (O_549,N_28177,N_25487);
nand UO_550 (O_550,N_25646,N_29277);
nand UO_551 (O_551,N_26611,N_25410);
nand UO_552 (O_552,N_28147,N_28716);
nor UO_553 (O_553,N_25726,N_27027);
and UO_554 (O_554,N_26035,N_27140);
xor UO_555 (O_555,N_28150,N_29118);
nand UO_556 (O_556,N_29395,N_25061);
nand UO_557 (O_557,N_27330,N_25573);
or UO_558 (O_558,N_28058,N_28141);
xor UO_559 (O_559,N_27559,N_27095);
nor UO_560 (O_560,N_28982,N_29087);
xnor UO_561 (O_561,N_26742,N_26601);
nor UO_562 (O_562,N_27394,N_27727);
nand UO_563 (O_563,N_28318,N_25010);
nor UO_564 (O_564,N_28285,N_26414);
and UO_565 (O_565,N_27731,N_29243);
nor UO_566 (O_566,N_26323,N_28945);
and UO_567 (O_567,N_27948,N_26519);
or UO_568 (O_568,N_25711,N_27932);
and UO_569 (O_569,N_26423,N_29797);
nor UO_570 (O_570,N_29886,N_29841);
and UO_571 (O_571,N_28010,N_29236);
xnor UO_572 (O_572,N_29509,N_26492);
and UO_573 (O_573,N_26734,N_26090);
nor UO_574 (O_574,N_26157,N_28393);
xnor UO_575 (O_575,N_26828,N_28136);
and UO_576 (O_576,N_29365,N_29508);
nand UO_577 (O_577,N_29269,N_27091);
nor UO_578 (O_578,N_28430,N_27406);
nor UO_579 (O_579,N_29681,N_27576);
nand UO_580 (O_580,N_27060,N_26844);
nor UO_581 (O_581,N_29959,N_29230);
and UO_582 (O_582,N_26850,N_29036);
nand UO_583 (O_583,N_28434,N_27008);
nor UO_584 (O_584,N_28896,N_29465);
and UO_585 (O_585,N_29466,N_25579);
nor UO_586 (O_586,N_28666,N_25770);
nand UO_587 (O_587,N_27722,N_26199);
or UO_588 (O_588,N_28488,N_28297);
xnor UO_589 (O_589,N_27170,N_25730);
and UO_590 (O_590,N_28897,N_29176);
or UO_591 (O_591,N_25384,N_26082);
or UO_592 (O_592,N_25747,N_27247);
or UO_593 (O_593,N_25118,N_26425);
nand UO_594 (O_594,N_29272,N_28629);
nand UO_595 (O_595,N_25912,N_29293);
or UO_596 (O_596,N_27662,N_27314);
and UO_597 (O_597,N_26319,N_27605);
and UO_598 (O_598,N_29458,N_29529);
and UO_599 (O_599,N_29638,N_29450);
nor UO_600 (O_600,N_26300,N_25365);
or UO_601 (O_601,N_25627,N_28204);
or UO_602 (O_602,N_26000,N_27596);
nor UO_603 (O_603,N_27950,N_26358);
and UO_604 (O_604,N_29723,N_27389);
xor UO_605 (O_605,N_27282,N_29525);
xor UO_606 (O_606,N_26764,N_25888);
and UO_607 (O_607,N_28964,N_29318);
nand UO_608 (O_608,N_25991,N_29411);
nor UO_609 (O_609,N_28887,N_25476);
or UO_610 (O_610,N_25485,N_29626);
or UO_611 (O_611,N_26196,N_25470);
or UO_612 (O_612,N_28944,N_26874);
or UO_613 (O_613,N_26337,N_28839);
and UO_614 (O_614,N_26254,N_26381);
nand UO_615 (O_615,N_27434,N_26522);
nor UO_616 (O_616,N_25249,N_27070);
nor UO_617 (O_617,N_26678,N_29987);
nand UO_618 (O_618,N_29617,N_28725);
nand UO_619 (O_619,N_28686,N_26950);
nand UO_620 (O_620,N_25198,N_28638);
nand UO_621 (O_621,N_28029,N_28060);
nand UO_622 (O_622,N_25697,N_25433);
and UO_623 (O_623,N_26867,N_25736);
nand UO_624 (O_624,N_25742,N_26525);
and UO_625 (O_625,N_26422,N_28849);
nand UO_626 (O_626,N_25574,N_28682);
nand UO_627 (O_627,N_25842,N_29284);
xor UO_628 (O_628,N_29404,N_27418);
or UO_629 (O_629,N_28188,N_27147);
xnor UO_630 (O_630,N_29818,N_28454);
xor UO_631 (O_631,N_25131,N_29784);
nor UO_632 (O_632,N_27053,N_25203);
nand UO_633 (O_633,N_25919,N_28562);
or UO_634 (O_634,N_29533,N_27808);
nand UO_635 (O_635,N_26400,N_27912);
or UO_636 (O_636,N_25829,N_27094);
xnor UO_637 (O_637,N_26065,N_26109);
nand UO_638 (O_638,N_25789,N_29459);
nor UO_639 (O_639,N_25116,N_26729);
and UO_640 (O_640,N_29715,N_28649);
xnor UO_641 (O_641,N_27349,N_26136);
or UO_642 (O_642,N_29261,N_25892);
and UO_643 (O_643,N_28937,N_27623);
xor UO_644 (O_644,N_28732,N_27714);
nand UO_645 (O_645,N_25885,N_26528);
xnor UO_646 (O_646,N_26557,N_25223);
nor UO_647 (O_647,N_28404,N_29556);
and UO_648 (O_648,N_29982,N_26490);
xnor UO_649 (O_649,N_26221,N_28548);
nand UO_650 (O_650,N_29980,N_27360);
nand UO_651 (O_651,N_28851,N_29836);
nand UO_652 (O_652,N_27540,N_29192);
or UO_653 (O_653,N_25437,N_26705);
xnor UO_654 (O_654,N_28965,N_29700);
nand UO_655 (O_655,N_27849,N_26438);
nand UO_656 (O_656,N_29148,N_25315);
nand UO_657 (O_657,N_29157,N_26580);
or UO_658 (O_658,N_26546,N_26006);
and UO_659 (O_659,N_28462,N_25647);
xor UO_660 (O_660,N_26561,N_25707);
xnor UO_661 (O_661,N_28002,N_27589);
nor UO_662 (O_662,N_26197,N_27642);
nand UO_663 (O_663,N_27000,N_29208);
nand UO_664 (O_664,N_26007,N_25555);
xnor UO_665 (O_665,N_26146,N_28729);
and UO_666 (O_666,N_29544,N_28446);
nor UO_667 (O_667,N_29598,N_29362);
nor UO_668 (O_668,N_27538,N_26128);
or UO_669 (O_669,N_25640,N_28277);
and UO_670 (O_670,N_25663,N_29309);
nor UO_671 (O_671,N_26068,N_28192);
nor UO_672 (O_672,N_27341,N_28413);
nand UO_673 (O_673,N_28016,N_26720);
xor UO_674 (O_674,N_29441,N_29590);
xor UO_675 (O_675,N_28391,N_27689);
nand UO_676 (O_676,N_26101,N_25105);
or UO_677 (O_677,N_25563,N_26238);
nor UO_678 (O_678,N_26552,N_26120);
and UO_679 (O_679,N_26264,N_25236);
or UO_680 (O_680,N_28656,N_27422);
or UO_681 (O_681,N_29597,N_28056);
or UO_682 (O_682,N_26613,N_27029);
nand UO_683 (O_683,N_27861,N_25889);
or UO_684 (O_684,N_26677,N_28882);
and UO_685 (O_685,N_28520,N_25784);
or UO_686 (O_686,N_29578,N_27357);
or UO_687 (O_687,N_27963,N_25270);
or UO_688 (O_688,N_28014,N_25455);
or UO_689 (O_689,N_25109,N_25983);
or UO_690 (O_690,N_27827,N_27888);
or UO_691 (O_691,N_25026,N_26798);
xor UO_692 (O_692,N_27831,N_27129);
xor UO_693 (O_693,N_29251,N_25288);
nor UO_694 (O_694,N_29159,N_27416);
or UO_695 (O_695,N_26403,N_25359);
nor UO_696 (O_696,N_28645,N_28160);
xnor UO_697 (O_697,N_27363,N_26773);
nand UO_698 (O_698,N_28067,N_27625);
or UO_699 (O_699,N_26375,N_26617);
nand UO_700 (O_700,N_28470,N_27795);
and UO_701 (O_701,N_28922,N_27678);
nor UO_702 (O_702,N_28095,N_29788);
nand UO_703 (O_703,N_25233,N_27103);
and UO_704 (O_704,N_27529,N_25609);
nand UO_705 (O_705,N_26214,N_29190);
xor UO_706 (O_706,N_25705,N_28031);
nand UO_707 (O_707,N_29256,N_29072);
xor UO_708 (O_708,N_29528,N_27900);
or UO_709 (O_709,N_29147,N_27687);
and UO_710 (O_710,N_28258,N_28667);
nand UO_711 (O_711,N_26286,N_27265);
and UO_712 (O_712,N_25451,N_25292);
nand UO_713 (O_713,N_26806,N_26639);
nor UO_714 (O_714,N_28804,N_27622);
or UO_715 (O_715,N_27609,N_27968);
xnor UO_716 (O_716,N_28880,N_27674);
xor UO_717 (O_717,N_26464,N_25030);
nor UO_718 (O_718,N_26060,N_27489);
nor UO_719 (O_719,N_26312,N_28854);
nand UO_720 (O_720,N_27410,N_25318);
and UO_721 (O_721,N_29312,N_26499);
or UO_722 (O_722,N_26551,N_25572);
nand UO_723 (O_723,N_28006,N_26098);
nand UO_724 (O_724,N_27160,N_27930);
xnor UO_725 (O_725,N_26452,N_25434);
and UO_726 (O_726,N_28902,N_29979);
xor UO_727 (O_727,N_25138,N_29397);
nand UO_728 (O_728,N_28813,N_25989);
nor UO_729 (O_729,N_28924,N_25699);
nand UO_730 (O_730,N_29653,N_28212);
or UO_731 (O_731,N_28558,N_28597);
and UO_732 (O_732,N_27250,N_26881);
xnor UO_733 (O_733,N_27859,N_25252);
xnor UO_734 (O_734,N_25950,N_25708);
nor UO_735 (O_735,N_27485,N_29926);
nand UO_736 (O_736,N_29892,N_26947);
and UO_737 (O_737,N_26442,N_25355);
nand UO_738 (O_738,N_27952,N_27440);
nand UO_739 (O_739,N_25949,N_29126);
nor UO_740 (O_740,N_25334,N_25147);
nor UO_741 (O_741,N_28755,N_29821);
nor UO_742 (O_742,N_29137,N_25457);
nand UO_743 (O_743,N_27555,N_27899);
xor UO_744 (O_744,N_25760,N_28246);
nor UO_745 (O_745,N_25689,N_28089);
nand UO_746 (O_746,N_25951,N_29799);
xor UO_747 (O_747,N_26706,N_27753);
xor UO_748 (O_748,N_29377,N_27921);
or UO_749 (O_749,N_29564,N_29825);
xor UO_750 (O_750,N_25712,N_27308);
or UO_751 (O_751,N_27483,N_27156);
xnor UO_752 (O_752,N_27051,N_28938);
or UO_753 (O_753,N_25486,N_25024);
nand UO_754 (O_754,N_26507,N_28589);
and UO_755 (O_755,N_25197,N_29485);
nand UO_756 (O_756,N_29657,N_27439);
xnor UO_757 (O_757,N_29651,N_26631);
nand UO_758 (O_758,N_27206,N_25801);
nand UO_759 (O_759,N_25881,N_26132);
nand UO_760 (O_760,N_29594,N_29473);
or UO_761 (O_761,N_25741,N_26486);
and UO_762 (O_762,N_29202,N_28068);
or UO_763 (O_763,N_25540,N_26709);
or UO_764 (O_764,N_26667,N_26992);
xnor UO_765 (O_765,N_26373,N_29019);
and UO_766 (O_766,N_25551,N_26194);
nand UO_767 (O_767,N_25055,N_26768);
xor UO_768 (O_768,N_28077,N_25596);
or UO_769 (O_769,N_29180,N_27816);
and UO_770 (O_770,N_26250,N_27185);
and UO_771 (O_771,N_26668,N_29054);
or UO_772 (O_772,N_26395,N_25575);
and UO_773 (O_773,N_28661,N_29752);
nand UO_774 (O_774,N_25381,N_26431);
or UO_775 (O_775,N_26853,N_26816);
nor UO_776 (O_776,N_29234,N_28981);
and UO_777 (O_777,N_28936,N_26715);
nand UO_778 (O_778,N_29955,N_25153);
or UO_779 (O_779,N_28419,N_26856);
or UO_780 (O_780,N_26103,N_26908);
or UO_781 (O_781,N_28220,N_27920);
nand UO_782 (O_782,N_26368,N_25649);
nor UO_783 (O_783,N_26094,N_28779);
and UO_784 (O_784,N_27292,N_29588);
or UO_785 (O_785,N_25658,N_29608);
nand UO_786 (O_786,N_27116,N_28125);
or UO_787 (O_787,N_28082,N_27338);
xor UO_788 (O_788,N_28426,N_27280);
xnor UO_789 (O_789,N_29512,N_29677);
and UO_790 (O_790,N_28398,N_29053);
nand UO_791 (O_791,N_26268,N_26201);
nor UO_792 (O_792,N_25925,N_26483);
nor UO_793 (O_793,N_26872,N_29364);
xnor UO_794 (O_794,N_26498,N_27286);
and UO_795 (O_795,N_25710,N_27344);
xnor UO_796 (O_796,N_29151,N_25652);
nor UO_797 (O_797,N_26555,N_28415);
and UO_798 (O_798,N_25195,N_26622);
xnor UO_799 (O_799,N_28027,N_27802);
and UO_800 (O_800,N_28451,N_26648);
nor UO_801 (O_801,N_26026,N_26024);
xnor UO_802 (O_802,N_29352,N_28600);
nor UO_803 (O_803,N_25124,N_25496);
xor UO_804 (O_804,N_25593,N_26547);
nor UO_805 (O_805,N_25674,N_29305);
nor UO_806 (O_806,N_28359,N_25959);
nand UO_807 (O_807,N_27044,N_26688);
or UO_808 (O_808,N_29742,N_27908);
xnor UO_809 (O_809,N_28689,N_27669);
and UO_810 (O_810,N_28827,N_29727);
and UO_811 (O_811,N_26291,N_29968);
nand UO_812 (O_812,N_29579,N_29407);
nor UO_813 (O_813,N_27403,N_26390);
xor UO_814 (O_814,N_29219,N_27987);
nor UO_815 (O_815,N_27640,N_26860);
or UO_816 (O_816,N_27243,N_29782);
xnor UO_817 (O_817,N_28194,N_28490);
xor UO_818 (O_818,N_28918,N_29863);
xor UO_819 (O_819,N_27455,N_28291);
nor UO_820 (O_820,N_26587,N_25980);
nand UO_821 (O_821,N_29523,N_29448);
or UO_822 (O_822,N_28811,N_27780);
nor UO_823 (O_823,N_25413,N_25656);
xnor UO_824 (O_824,N_27591,N_25623);
nand UO_825 (O_825,N_28330,N_28678);
nand UO_826 (O_826,N_25774,N_25836);
xnor UO_827 (O_827,N_29810,N_29089);
nor UO_828 (O_828,N_29091,N_29487);
nor UO_829 (O_829,N_29879,N_28812);
nand UO_830 (O_830,N_28593,N_28580);
and UO_831 (O_831,N_27719,N_28366);
nand UO_832 (O_832,N_27628,N_27077);
or UO_833 (O_833,N_26450,N_27212);
nor UO_834 (O_834,N_29606,N_25792);
xor UO_835 (O_835,N_28207,N_26303);
nor UO_836 (O_836,N_26051,N_26032);
nand UO_837 (O_837,N_25272,N_29831);
or UO_838 (O_838,N_28245,N_29052);
nand UO_839 (O_839,N_28433,N_25722);
nand UO_840 (O_840,N_26503,N_29361);
nor UO_841 (O_841,N_26099,N_29573);
or UO_842 (O_842,N_28655,N_26270);
nor UO_843 (O_843,N_26124,N_29435);
nand UO_844 (O_844,N_26584,N_29659);
or UO_845 (O_845,N_28577,N_28833);
or UO_846 (O_846,N_28886,N_26363);
nand UO_847 (O_847,N_27438,N_25999);
xor UO_848 (O_848,N_29539,N_27737);
nand UO_849 (O_849,N_29223,N_26100);
nand UO_850 (O_850,N_28906,N_29333);
and UO_851 (O_851,N_28978,N_25379);
xor UO_852 (O_852,N_25008,N_29443);
or UO_853 (O_853,N_25192,N_26399);
xnor UO_854 (O_854,N_25033,N_26028);
and UO_855 (O_855,N_29888,N_27978);
nand UO_856 (O_856,N_27819,N_25860);
nand UO_857 (O_857,N_29930,N_26252);
xnor UO_858 (O_858,N_28720,N_25727);
xnor UO_859 (O_859,N_26809,N_26686);
or UO_860 (O_860,N_27164,N_28983);
xnor UO_861 (O_861,N_28843,N_26793);
nand UO_862 (O_862,N_29792,N_25466);
xor UO_863 (O_863,N_28307,N_29009);
nand UO_864 (O_864,N_29325,N_26888);
and UO_865 (O_865,N_29773,N_29314);
and UO_866 (O_866,N_27319,N_28155);
and UO_867 (O_867,N_29433,N_27806);
nand UO_868 (O_868,N_25521,N_26116);
nand UO_869 (O_869,N_27778,N_28624);
nor UO_870 (O_870,N_27155,N_26249);
nor UO_871 (O_871,N_25160,N_28806);
nor UO_872 (O_872,N_27087,N_27285);
nand UO_873 (O_873,N_25846,N_25941);
nand UO_874 (O_874,N_29670,N_26142);
nor UO_875 (O_875,N_25143,N_25803);
nor UO_876 (O_876,N_27931,N_27150);
xnor UO_877 (O_877,N_26276,N_28376);
and UO_878 (O_878,N_25388,N_28100);
xnor UO_879 (O_879,N_25084,N_27980);
nand UO_880 (O_880,N_28180,N_27643);
and UO_881 (O_881,N_28387,N_25400);
xor UO_882 (O_882,N_28602,N_27926);
nand UO_883 (O_883,N_25254,N_25536);
nand UO_884 (O_884,N_25797,N_27627);
nor UO_885 (O_885,N_25088,N_27812);
nor UO_886 (O_886,N_26901,N_27757);
nand UO_887 (O_887,N_27365,N_25527);
and UO_888 (O_888,N_26787,N_28229);
nand UO_889 (O_889,N_28247,N_27995);
and UO_890 (O_890,N_28857,N_27871);
nor UO_891 (O_891,N_26347,N_26466);
nand UO_892 (O_892,N_28545,N_26318);
nor UO_893 (O_893,N_27502,N_28865);
nor UO_894 (O_894,N_28528,N_29973);
nor UO_895 (O_895,N_25023,N_25182);
and UO_896 (O_896,N_28504,N_28876);
nor UO_897 (O_897,N_25587,N_29561);
nor UO_898 (O_898,N_28890,N_28105);
xnor UO_899 (O_899,N_28115,N_28024);
nor UO_900 (O_900,N_26638,N_26455);
and UO_901 (O_901,N_25036,N_28565);
nand UO_902 (O_902,N_29209,N_28932);
and UO_903 (O_903,N_27303,N_29383);
xor UO_904 (O_904,N_26280,N_25284);
and UO_905 (O_905,N_29672,N_26419);
nor UO_906 (O_906,N_28099,N_25517);
nand UO_907 (O_907,N_28131,N_26177);
xnor UO_908 (O_908,N_27385,N_26121);
nor UO_909 (O_909,N_29701,N_28605);
nand UO_910 (O_910,N_25978,N_28302);
and UO_911 (O_911,N_26027,N_29338);
xor UO_912 (O_912,N_28046,N_25338);
and UO_913 (O_913,N_27466,N_25462);
and UO_914 (O_914,N_25113,N_28535);
xor UO_915 (O_915,N_29826,N_29145);
or UO_916 (O_916,N_29769,N_25861);
nor UO_917 (O_917,N_29360,N_25590);
nor UO_918 (O_918,N_26849,N_27774);
and UO_919 (O_919,N_29461,N_27828);
and UO_920 (O_920,N_25261,N_29929);
nand UO_921 (O_921,N_25974,N_25600);
nor UO_922 (O_922,N_29245,N_29641);
or UO_923 (O_923,N_26756,N_25903);
and UO_924 (O_924,N_29393,N_27683);
xor UO_925 (O_925,N_28525,N_29741);
or UO_926 (O_926,N_26078,N_29096);
xnor UO_927 (O_927,N_25043,N_26751);
and UO_928 (O_928,N_26484,N_29472);
or UO_929 (O_929,N_25887,N_27537);
or UO_930 (O_930,N_28427,N_25883);
or UO_931 (O_931,N_27456,N_28749);
xor UO_932 (O_932,N_29035,N_25256);
and UO_933 (O_933,N_25655,N_26080);
nor UO_934 (O_934,N_29071,N_29279);
and UO_935 (O_935,N_29287,N_29794);
or UO_936 (O_936,N_25049,N_25275);
xnor UO_937 (O_937,N_26494,N_28819);
and UO_938 (O_938,N_25446,N_27446);
nand UO_939 (O_939,N_27208,N_27173);
or UO_940 (O_940,N_29805,N_27738);
and UO_941 (O_941,N_29895,N_26604);
nor UO_942 (O_942,N_25363,N_25063);
or UO_943 (O_943,N_27823,N_26619);
nand UO_944 (O_944,N_28961,N_28841);
xnor UO_945 (O_945,N_26003,N_26892);
nand UO_946 (O_946,N_25838,N_29690);
or UO_947 (O_947,N_28213,N_29281);
nor UO_948 (O_948,N_29369,N_28825);
xor UO_949 (O_949,N_28267,N_25370);
and UO_950 (O_950,N_28641,N_29290);
and UO_951 (O_951,N_27788,N_26919);
nand UO_952 (O_952,N_26531,N_27696);
nand UO_953 (O_953,N_27742,N_29436);
nor UO_954 (O_954,N_28622,N_26478);
nor UO_955 (O_955,N_25339,N_26477);
and UO_956 (O_956,N_26935,N_27531);
and UO_957 (O_957,N_27761,N_28483);
nor UO_958 (O_958,N_28966,N_28073);
nor UO_959 (O_959,N_25548,N_28523);
and UO_960 (O_960,N_27769,N_29541);
nor UO_961 (O_961,N_27409,N_25059);
xor UO_962 (O_962,N_25577,N_25987);
and UO_963 (O_963,N_27328,N_25715);
nor UO_964 (O_964,N_28390,N_25580);
xnor UO_965 (O_965,N_29766,N_27739);
or UO_966 (O_966,N_28790,N_28592);
nand UO_967 (O_967,N_28526,N_28133);
or UO_968 (O_968,N_27105,N_25994);
nand UO_969 (O_969,N_28650,N_28063);
and UO_970 (O_970,N_28331,N_26467);
and UO_971 (O_971,N_26957,N_25076);
or UO_972 (O_972,N_26654,N_25628);
nand UO_973 (O_973,N_29077,N_25698);
and UO_974 (O_974,N_29379,N_26424);
and UO_975 (O_975,N_25335,N_25546);
xor UO_976 (O_976,N_27573,N_25781);
or UO_977 (O_977,N_26269,N_29213);
and UO_978 (O_978,N_26808,N_29476);
nor UO_979 (O_979,N_25653,N_28339);
and UO_980 (O_980,N_29815,N_29874);
nor UO_981 (O_981,N_28685,N_27224);
and UO_982 (O_982,N_29553,N_29066);
or UO_983 (O_983,N_25778,N_27729);
or UO_984 (O_984,N_29058,N_25564);
nor UO_985 (O_985,N_29045,N_26569);
nor UO_986 (O_986,N_28677,N_28660);
xor UO_987 (O_987,N_25104,N_27543);
nand UO_988 (O_988,N_29765,N_25694);
xnor UO_989 (O_989,N_29927,N_26308);
xnor UO_990 (O_990,N_25283,N_29437);
or UO_991 (O_991,N_26412,N_26894);
nand UO_992 (O_992,N_28940,N_28271);
nand UO_993 (O_993,N_29543,N_28400);
nor UO_994 (O_994,N_25166,N_27949);
xor UO_995 (O_995,N_29648,N_27219);
nor UO_996 (O_996,N_27852,N_25242);
and UO_997 (O_997,N_27350,N_25251);
and UO_998 (O_998,N_29028,N_25503);
or UO_999 (O_999,N_25794,N_29135);
and UO_1000 (O_1000,N_27043,N_26949);
nand UO_1001 (O_1001,N_29342,N_25612);
and UO_1002 (O_1002,N_25812,N_29538);
xnor UO_1003 (O_1003,N_26190,N_29398);
xor UO_1004 (O_1004,N_27695,N_29633);
nand UO_1005 (O_1005,N_25924,N_26885);
or UO_1006 (O_1006,N_28313,N_26160);
nand UO_1007 (O_1007,N_25265,N_28693);
and UO_1008 (O_1008,N_26050,N_27550);
nor UO_1009 (O_1009,N_25582,N_27826);
nor UO_1010 (O_1010,N_26750,N_29063);
nor UO_1011 (O_1011,N_25756,N_27712);
or UO_1012 (O_1012,N_27503,N_28569);
nand UO_1013 (O_1013,N_25586,N_25641);
and UO_1014 (O_1014,N_28898,N_26192);
and UO_1015 (O_1015,N_27004,N_25056);
or UO_1016 (O_1016,N_29611,N_27911);
xnor UO_1017 (O_1017,N_27762,N_28644);
or UO_1018 (O_1018,N_26148,N_28489);
xnor UO_1019 (O_1019,N_28552,N_25229);
xor UO_1020 (O_1020,N_29711,N_29370);
nand UO_1021 (O_1021,N_28225,N_27048);
xnor UO_1022 (O_1022,N_28273,N_27614);
nor UO_1023 (O_1023,N_25844,N_27887);
nand UO_1024 (O_1024,N_28298,N_29946);
nor UO_1025 (O_1025,N_27322,N_28726);
nand UO_1026 (O_1026,N_28517,N_29643);
xnor UO_1027 (O_1027,N_25269,N_28370);
and UO_1028 (O_1028,N_25004,N_25969);
xor UO_1029 (O_1029,N_28323,N_28695);
and UO_1030 (O_1030,N_27539,N_25562);
or UO_1031 (O_1031,N_25504,N_29503);
and UO_1032 (O_1032,N_25524,N_28687);
or UO_1033 (O_1033,N_27447,N_28858);
xnor UO_1034 (O_1034,N_26436,N_26794);
xnor UO_1035 (O_1035,N_25210,N_28912);
and UO_1036 (O_1036,N_28479,N_27019);
and UO_1037 (O_1037,N_28072,N_25120);
xor UO_1038 (O_1038,N_28383,N_25650);
or UO_1039 (O_1039,N_25547,N_28440);
or UO_1040 (O_1040,N_28712,N_27084);
and UO_1041 (O_1041,N_27629,N_29520);
or UO_1042 (O_1042,N_28112,N_26704);
nand UO_1043 (O_1043,N_26104,N_27231);
nor UO_1044 (O_1044,N_28013,N_25765);
or UO_1045 (O_1045,N_25394,N_25863);
nand UO_1046 (O_1046,N_28926,N_28165);
or UO_1047 (O_1047,N_25998,N_28394);
or UO_1048 (O_1048,N_25397,N_29074);
xor UO_1049 (O_1049,N_29928,N_25535);
and UO_1050 (O_1050,N_29848,N_27153);
and UO_1051 (O_1051,N_26765,N_28049);
and UO_1052 (O_1052,N_29827,N_27088);
and UO_1053 (O_1053,N_25069,N_29111);
and UO_1054 (O_1054,N_27976,N_29756);
nand UO_1055 (O_1055,N_27509,N_29706);
nand UO_1056 (O_1056,N_25473,N_26417);
or UO_1057 (O_1057,N_27560,N_27526);
or UO_1058 (O_1058,N_28096,N_26293);
or UO_1059 (O_1059,N_29664,N_29574);
and UO_1060 (O_1060,N_28481,N_28933);
or UO_1061 (O_1061,N_28146,N_25161);
or UO_1062 (O_1062,N_25399,N_26999);
and UO_1063 (O_1063,N_26225,N_29094);
and UO_1064 (O_1064,N_29144,N_29417);
nor UO_1065 (O_1065,N_26255,N_29138);
nor UO_1066 (O_1066,N_27524,N_29589);
nor UO_1067 (O_1067,N_29212,N_25324);
or UO_1068 (O_1068,N_29345,N_25149);
and UO_1069 (O_1069,N_26956,N_29871);
xnor UO_1070 (O_1070,N_26980,N_28365);
nand UO_1071 (O_1071,N_26112,N_25452);
or UO_1072 (O_1072,N_26491,N_25075);
xor UO_1073 (O_1073,N_29646,N_28351);
and UO_1074 (O_1074,N_29978,N_29840);
xor UO_1075 (O_1075,N_29614,N_25441);
xor UO_1076 (O_1076,N_29408,N_26481);
nor UO_1077 (O_1077,N_26752,N_28036);
or UO_1078 (O_1078,N_28021,N_28243);
or UO_1079 (O_1079,N_28151,N_25480);
and UO_1080 (O_1080,N_28861,N_26813);
and UO_1081 (O_1081,N_28015,N_26863);
and UO_1082 (O_1082,N_28238,N_27126);
xnor UO_1083 (O_1083,N_26969,N_25390);
xor UO_1084 (O_1084,N_26778,N_27354);
nor UO_1085 (O_1085,N_28913,N_25078);
and UO_1086 (O_1086,N_28290,N_25314);
and UO_1087 (O_1087,N_27553,N_25891);
and UO_1088 (O_1088,N_27267,N_25102);
and UO_1089 (O_1089,N_26559,N_28268);
or UO_1090 (O_1090,N_26884,N_28700);
or UO_1091 (O_1091,N_27171,N_25905);
or UO_1092 (O_1092,N_28190,N_27401);
xnor UO_1093 (O_1093,N_29693,N_25376);
or UO_1094 (O_1094,N_26062,N_25243);
xor UO_1095 (O_1095,N_29178,N_27775);
or UO_1096 (O_1096,N_25635,N_27096);
nand UO_1097 (O_1097,N_29908,N_26019);
xor UO_1098 (O_1098,N_25933,N_25568);
nor UO_1099 (O_1099,N_26865,N_25772);
nand UO_1100 (O_1100,N_27033,N_25835);
and UO_1101 (O_1101,N_29228,N_27235);
nor UO_1102 (O_1102,N_28142,N_29497);
or UO_1103 (O_1103,N_27879,N_28997);
nor UO_1104 (O_1104,N_26566,N_26360);
and UO_1105 (O_1105,N_29596,N_29970);
nand UO_1106 (O_1106,N_29961,N_29322);
xnor UO_1107 (O_1107,N_25092,N_27424);
xor UO_1108 (O_1108,N_25533,N_28282);
nor UO_1109 (O_1109,N_29274,N_28870);
and UO_1110 (O_1110,N_25806,N_28098);
nor UO_1111 (O_1111,N_27395,N_25764);
xor UO_1112 (O_1112,N_25898,N_28191);
nor UO_1113 (O_1113,N_28482,N_26610);
xor UO_1114 (O_1114,N_27124,N_27992);
nor UO_1115 (O_1115,N_26680,N_28822);
xor UO_1116 (O_1116,N_29983,N_26476);
xnor UO_1117 (O_1117,N_26108,N_25753);
nand UO_1118 (O_1118,N_25997,N_25279);
and UO_1119 (O_1119,N_25982,N_27238);
xor UO_1120 (O_1120,N_26346,N_29551);
and UO_1121 (O_1121,N_26523,N_29319);
nor UO_1122 (O_1122,N_26616,N_25357);
nand UO_1123 (O_1123,N_28329,N_27903);
and UO_1124 (O_1124,N_29462,N_28294);
xor UO_1125 (O_1125,N_27460,N_25440);
nand UO_1126 (O_1126,N_29527,N_29095);
xor UO_1127 (O_1127,N_25505,N_28988);
or UO_1128 (O_1128,N_27304,N_27316);
and UO_1129 (O_1129,N_27074,N_25717);
nor UO_1130 (O_1130,N_29724,N_28118);
or UO_1131 (O_1131,N_25266,N_26096);
nor UO_1132 (O_1132,N_26926,N_27461);
and UO_1133 (O_1133,N_25245,N_26975);
nor UO_1134 (O_1134,N_28513,N_28739);
and UO_1135 (O_1135,N_29852,N_28699);
nand UO_1136 (O_1136,N_26342,N_25321);
nand UO_1137 (O_1137,N_26887,N_27977);
and UO_1138 (O_1138,N_26126,N_27880);
and UO_1139 (O_1139,N_29205,N_25728);
nor UO_1140 (O_1140,N_27754,N_27951);
and UO_1141 (O_1141,N_29680,N_26846);
nand UO_1142 (O_1142,N_26278,N_27242);
nand UO_1143 (O_1143,N_29777,N_26457);
and UO_1144 (O_1144,N_27787,N_26659);
nor UO_1145 (O_1145,N_26361,N_26821);
nor UO_1146 (O_1146,N_25896,N_26458);
and UO_1147 (O_1147,N_27260,N_28679);
nand UO_1148 (O_1148,N_27997,N_27488);
or UO_1149 (O_1149,N_25303,N_27123);
xnor UO_1150 (O_1150,N_29231,N_28704);
nor UO_1151 (O_1151,N_25167,N_29278);
nor UO_1152 (O_1152,N_28360,N_25918);
xnor UO_1153 (O_1153,N_26107,N_27062);
xor UO_1154 (O_1154,N_28090,N_29432);
xor UO_1155 (O_1155,N_25954,N_26010);
nand UO_1156 (O_1156,N_29196,N_28547);
and UO_1157 (O_1157,N_25817,N_27134);
nor UO_1158 (O_1158,N_25077,N_27176);
and UO_1159 (O_1159,N_29785,N_25468);
xor UO_1160 (O_1160,N_26448,N_28800);
and UO_1161 (O_1161,N_29932,N_27400);
xnor UO_1162 (O_1162,N_27655,N_26986);
and UO_1163 (O_1163,N_25731,N_27225);
and UO_1164 (O_1164,N_28816,N_27184);
nor UO_1165 (O_1165,N_25567,N_26151);
nand UO_1166 (O_1166,N_26952,N_29750);
nand UO_1167 (O_1167,N_25148,N_27946);
xor UO_1168 (O_1168,N_25444,N_27037);
or UO_1169 (O_1169,N_28684,N_29846);
nand UO_1170 (O_1170,N_28495,N_27407);
and UO_1171 (O_1171,N_28671,N_26282);
or UO_1172 (O_1172,N_28715,N_27841);
nor UO_1173 (O_1173,N_29625,N_28740);
xor UO_1174 (O_1174,N_25141,N_28708);
xnor UO_1175 (O_1175,N_29170,N_25716);
nand UO_1176 (O_1176,N_27960,N_27188);
xnor UO_1177 (O_1177,N_26075,N_27016);
xor UO_1178 (O_1178,N_27568,N_28035);
nor UO_1179 (O_1179,N_28227,N_26805);
nand UO_1180 (O_1180,N_25512,N_27990);
nor UO_1181 (O_1181,N_26297,N_25021);
or UO_1182 (O_1182,N_25435,N_25648);
or UO_1183 (O_1183,N_26296,N_25520);
or UO_1184 (O_1184,N_28874,N_25606);
xnor UO_1185 (O_1185,N_28492,N_26696);
and UO_1186 (O_1186,N_29781,N_25289);
xnor UO_1187 (O_1187,N_28571,N_29046);
and UO_1188 (O_1188,N_26534,N_28973);
xor UO_1189 (O_1189,N_28643,N_25136);
and UO_1190 (O_1190,N_28134,N_29990);
nand UO_1191 (O_1191,N_26016,N_29215);
or UO_1192 (O_1192,N_25420,N_28698);
nand UO_1193 (O_1193,N_27702,N_26598);
nand UO_1194 (O_1194,N_27381,N_29751);
nor UO_1195 (O_1195,N_27404,N_28486);
nor UO_1196 (O_1196,N_28292,N_26161);
and UO_1197 (O_1197,N_25127,N_28020);
nor UO_1198 (O_1198,N_26322,N_27672);
or UO_1199 (O_1199,N_27244,N_29200);
nor UO_1200 (O_1200,N_29083,N_26227);
nand UO_1201 (O_1201,N_28236,N_25970);
xor UO_1202 (O_1202,N_29854,N_27487);
xnor UO_1203 (O_1203,N_29221,N_27552);
nand UO_1204 (O_1204,N_26864,N_28697);
or UO_1205 (O_1205,N_25581,N_28986);
and UO_1206 (O_1206,N_26726,N_26586);
xnor UO_1207 (O_1207,N_25867,N_28321);
nor UO_1208 (O_1208,N_25874,N_28652);
nor UO_1209 (O_1209,N_26506,N_27371);
xor UO_1210 (O_1210,N_26804,N_25108);
xor UO_1211 (O_1211,N_28879,N_28798);
xor UO_1212 (O_1212,N_25180,N_28639);
nand UO_1213 (O_1213,N_25139,N_27984);
xnor UO_1214 (O_1214,N_28363,N_28296);
or UO_1215 (O_1215,N_27616,N_26879);
xor UO_1216 (O_1216,N_25439,N_25132);
nor UO_1217 (O_1217,N_26655,N_25675);
or UO_1218 (O_1218,N_28885,N_29007);
nor UO_1219 (O_1219,N_26626,N_25354);
or UO_1220 (O_1220,N_28970,N_27102);
xor UO_1221 (O_1221,N_27940,N_27897);
nand UO_1222 (O_1222,N_25714,N_29175);
nand UO_1223 (O_1223,N_26851,N_27528);
nand UO_1224 (O_1224,N_27493,N_25777);
and UO_1225 (O_1225,N_28539,N_29482);
or UO_1226 (O_1226,N_26576,N_27142);
nand UO_1227 (O_1227,N_27393,N_26460);
nor UO_1228 (O_1228,N_25804,N_27909);
xnor UO_1229 (O_1229,N_27269,N_26671);
xor UO_1230 (O_1230,N_26870,N_27734);
xnor UO_1231 (O_1231,N_29152,N_28914);
xor UO_1232 (O_1232,N_27776,N_29399);
and UO_1233 (O_1233,N_27673,N_25323);
and UO_1234 (O_1234,N_25248,N_27279);
nand UO_1235 (O_1235,N_29881,N_27876);
nor UO_1236 (O_1236,N_29803,N_27259);
nor UO_1237 (O_1237,N_26345,N_29081);
and UO_1238 (O_1238,N_28171,N_29388);
or UO_1239 (O_1239,N_28037,N_28868);
and UO_1240 (O_1240,N_29684,N_29743);
xnor UO_1241 (O_1241,N_26762,N_26315);
and UO_1242 (O_1242,N_26169,N_26603);
xnor UO_1243 (O_1243,N_26195,N_29297);
nor UO_1244 (O_1244,N_28546,N_26565);
or UO_1245 (O_1245,N_29390,N_25224);
xor UO_1246 (O_1246,N_28957,N_25947);
or UO_1247 (O_1247,N_29812,N_27039);
or UO_1248 (O_1248,N_25025,N_26536);
nand UO_1249 (O_1249,N_25779,N_28803);
or UO_1250 (O_1250,N_26755,N_28611);
nand UO_1251 (O_1251,N_28388,N_28573);
or UO_1252 (O_1252,N_26722,N_28409);
and UO_1253 (O_1253,N_27917,N_29226);
nand UO_1254 (O_1254,N_26047,N_27824);
nand UO_1255 (O_1255,N_25458,N_26407);
or UO_1256 (O_1256,N_25622,N_25333);
and UO_1257 (O_1257,N_28316,N_29282);
and UO_1258 (O_1258,N_29985,N_25201);
nand UO_1259 (O_1259,N_25152,N_26383);
nand UO_1260 (O_1260,N_29003,N_28694);
and UO_1261 (O_1261,N_29210,N_25511);
or UO_1262 (O_1262,N_27593,N_29513);
or UO_1263 (O_1263,N_28226,N_25479);
xor UO_1264 (O_1264,N_26167,N_25326);
or UO_1265 (O_1265,N_28786,N_29130);
and UO_1266 (O_1266,N_29889,N_25140);
nor UO_1267 (O_1267,N_28472,N_26899);
xnor UO_1268 (O_1268,N_29688,N_28108);
and UO_1269 (O_1269,N_25278,N_29537);
xor UO_1270 (O_1270,N_26002,N_26074);
xnor UO_1271 (O_1271,N_25367,N_28783);
nand UO_1272 (O_1272,N_29622,N_29778);
or UO_1273 (O_1273,N_25617,N_27099);
or UO_1274 (O_1274,N_25830,N_28744);
nor UO_1275 (O_1275,N_25135,N_27198);
or UO_1276 (O_1276,N_29505,N_29249);
nand UO_1277 (O_1277,N_28205,N_26134);
nor UO_1278 (O_1278,N_25343,N_28881);
and UO_1279 (O_1279,N_29759,N_26133);
and UO_1280 (O_1280,N_25079,N_27376);
and UO_1281 (O_1281,N_29506,N_25469);
nand UO_1282 (O_1282,N_29254,N_29736);
or UO_1283 (O_1283,N_27511,N_25651);
xnor UO_1284 (O_1284,N_26042,N_28931);
nand UO_1285 (O_1285,N_27118,N_26833);
xor UO_1286 (O_1286,N_28836,N_28996);
xnor UO_1287 (O_1287,N_29833,N_28728);
nand UO_1288 (O_1288,N_28673,N_25282);
or UO_1289 (O_1289,N_28139,N_25541);
or UO_1290 (O_1290,N_26384,N_28306);
nor UO_1291 (O_1291,N_29909,N_26852);
and UO_1292 (O_1292,N_26535,N_25632);
nor UO_1293 (O_1293,N_26607,N_26232);
or UO_1294 (O_1294,N_27895,N_26997);
or UO_1295 (O_1295,N_25401,N_29475);
or UO_1296 (O_1296,N_29934,N_29001);
or UO_1297 (O_1297,N_26508,N_28378);
or UO_1298 (O_1298,N_27794,N_26662);
and UO_1299 (O_1299,N_26740,N_25855);
nand UO_1300 (O_1300,N_26683,N_29729);
and UO_1301 (O_1301,N_25209,N_29469);
nand UO_1302 (O_1302,N_29532,N_28477);
xor UO_1303 (O_1303,N_27209,N_29577);
and UO_1304 (O_1304,N_27713,N_26602);
xor UO_1305 (O_1305,N_27229,N_27942);
and UO_1306 (O_1306,N_25027,N_29217);
nand UO_1307 (O_1307,N_29744,N_26699);
or UO_1308 (O_1308,N_26313,N_28075);
nand UO_1309 (O_1309,N_27391,N_26044);
or UO_1310 (O_1310,N_26810,N_29406);
xor UO_1311 (O_1311,N_25597,N_29593);
or UO_1312 (O_1312,N_26447,N_29005);
nand UO_1313 (O_1313,N_25904,N_26953);
or UO_1314 (O_1314,N_27692,N_27249);
nor UO_1315 (O_1315,N_26265,N_28169);
or UO_1316 (O_1316,N_29040,N_26451);
nor UO_1317 (O_1317,N_27612,N_27475);
nand UO_1318 (O_1318,N_29498,N_25518);
and UO_1319 (O_1319,N_25706,N_27022);
and UO_1320 (O_1320,N_26110,N_26635);
and UO_1321 (O_1321,N_29814,N_26504);
nor UO_1322 (O_1322,N_29327,N_29088);
xnor UO_1323 (O_1323,N_29583,N_27872);
nor UO_1324 (O_1324,N_25615,N_29763);
or UO_1325 (O_1325,N_25208,N_28007);
nor UO_1326 (O_1326,N_25238,N_28086);
nor UO_1327 (O_1327,N_28891,N_26676);
xor UO_1328 (O_1328,N_28405,N_27520);
xor UO_1329 (O_1329,N_27832,N_28242);
or UO_1330 (O_1330,N_26502,N_26568);
xor UO_1331 (O_1331,N_26761,N_27380);
xor UO_1332 (O_1332,N_25328,N_27054);
xnor UO_1333 (O_1333,N_25448,N_28081);
nor UO_1334 (O_1334,N_27991,N_25810);
or UO_1335 (O_1335,N_27706,N_25305);
nand UO_1336 (O_1336,N_25364,N_27157);
nor UO_1337 (O_1337,N_29671,N_27026);
nor UO_1338 (O_1338,N_28999,N_29276);
and UO_1339 (O_1339,N_26961,N_28066);
nor UO_1340 (O_1340,N_25877,N_26147);
or UO_1341 (O_1341,N_29146,N_26636);
xnor UO_1342 (O_1342,N_28867,N_25191);
or UO_1343 (O_1343,N_27362,N_26237);
nand UO_1344 (O_1344,N_29396,N_28239);
xor UO_1345 (O_1345,N_28093,N_25526);
nand UO_1346 (O_1346,N_29061,N_26600);
xnor UO_1347 (O_1347,N_27055,N_25523);
nand UO_1348 (O_1348,N_25454,N_27057);
nor UO_1349 (O_1349,N_27556,N_27793);
xor UO_1350 (O_1350,N_28752,N_27450);
or UO_1351 (O_1351,N_26023,N_29262);
nor UO_1352 (O_1352,N_29504,N_27618);
nor UO_1353 (O_1353,N_28259,N_25531);
nor UO_1354 (O_1354,N_29988,N_27720);
or UO_1355 (O_1355,N_28345,N_27251);
xor UO_1356 (O_1356,N_26093,N_27745);
or UO_1357 (O_1357,N_28230,N_25721);
nand UO_1358 (O_1358,N_29963,N_29642);
xor UO_1359 (O_1359,N_28174,N_25729);
nand UO_1360 (O_1360,N_26305,N_27178);
nor UO_1361 (O_1361,N_27667,N_26955);
nor UO_1362 (O_1362,N_29779,N_27049);
nand UO_1363 (O_1363,N_29495,N_26310);
or UO_1364 (O_1364,N_29093,N_25858);
nand UO_1365 (O_1365,N_29565,N_27010);
and UO_1366 (O_1366,N_27311,N_26394);
and UO_1367 (O_1367,N_29868,N_25811);
or UO_1368 (O_1368,N_26218,N_27317);
and UO_1369 (O_1369,N_25062,N_25412);
nand UO_1370 (O_1370,N_25042,N_26371);
nor UO_1371 (O_1371,N_29572,N_27838);
and UO_1372 (O_1372,N_28401,N_29905);
nor UO_1373 (O_1373,N_25257,N_28324);
nand UO_1374 (O_1374,N_28842,N_27902);
xnor UO_1375 (O_1375,N_29172,N_27708);
and UO_1376 (O_1376,N_27877,N_29907);
and UO_1377 (O_1377,N_29496,N_28057);
nand UO_1378 (O_1378,N_29375,N_25322);
nand UO_1379 (O_1379,N_27335,N_25474);
nand UO_1380 (O_1380,N_27691,N_27855);
nand UO_1381 (O_1381,N_29885,N_26224);
or UO_1382 (O_1382,N_28900,N_28640);
nand UO_1383 (O_1383,N_28664,N_25695);
nor UO_1384 (O_1384,N_28738,N_28439);
nor UO_1385 (O_1385,N_26976,N_27505);
and UO_1386 (O_1386,N_29460,N_25594);
nor UO_1387 (O_1387,N_29735,N_25193);
or UO_1388 (O_1388,N_25690,N_28823);
nor UO_1389 (O_1389,N_29038,N_26350);
xnor UO_1390 (O_1390,N_27325,N_25205);
or UO_1391 (O_1391,N_29265,N_25015);
xnor UO_1392 (O_1392,N_29995,N_27073);
nor UO_1393 (O_1393,N_27299,N_29775);
and UO_1394 (O_1394,N_25815,N_28162);
xnor UO_1395 (O_1395,N_28923,N_25250);
nand UO_1396 (O_1396,N_29357,N_29923);
nand UO_1397 (O_1397,N_29343,N_27913);
and UO_1398 (O_1398,N_28967,N_28828);
xor UO_1399 (O_1399,N_29141,N_29547);
xnor UO_1400 (O_1400,N_26340,N_29890);
or UO_1401 (O_1401,N_28061,N_25028);
and UO_1402 (O_1402,N_25290,N_26202);
nor UO_1403 (O_1403,N_28711,N_27239);
nand UO_1404 (O_1404,N_27481,N_29292);
and UO_1405 (O_1405,N_28864,N_29409);
nand UO_1406 (O_1406,N_28497,N_25007);
nand UO_1407 (O_1407,N_28598,N_29295);
nand UO_1408 (O_1408,N_26207,N_27954);
or UO_1409 (O_1409,N_26627,N_25327);
or UO_1410 (O_1410,N_27069,N_26168);
and UO_1411 (O_1411,N_29181,N_27652);
nor UO_1412 (O_1412,N_26234,N_27276);
xor UO_1413 (O_1413,N_25453,N_26575);
xor UO_1414 (O_1414,N_26634,N_26480);
xnor UO_1415 (O_1415,N_28566,N_26279);
nand UO_1416 (O_1416,N_29400,N_25183);
nand UO_1417 (O_1417,N_26022,N_25754);
nor UO_1418 (O_1418,N_28572,N_26309);
nor UO_1419 (O_1419,N_27768,N_28838);
nor UO_1420 (O_1420,N_27836,N_27444);
or UO_1421 (O_1421,N_27465,N_28468);
and UO_1422 (O_1422,N_25408,N_29602);
and UO_1423 (O_1423,N_26206,N_28853);
nor UO_1424 (O_1424,N_29627,N_25679);
and UO_1425 (O_1425,N_29591,N_25155);
xor UO_1426 (O_1426,N_26749,N_28346);
and UO_1427 (O_1427,N_29106,N_27651);
xor UO_1428 (O_1428,N_29772,N_29582);
xor UO_1429 (O_1429,N_28943,N_28403);
and UO_1430 (O_1430,N_25181,N_25604);
nor UO_1431 (O_1431,N_29603,N_26430);
nand UO_1432 (O_1432,N_27927,N_25620);
and UO_1433 (O_1433,N_29023,N_26548);
nor UO_1434 (O_1434,N_28326,N_25845);
or UO_1435 (O_1435,N_28224,N_28352);
and UO_1436 (O_1436,N_25659,N_25507);
nor UO_1437 (O_1437,N_25134,N_29199);
and UO_1438 (O_1438,N_29056,N_26785);
nor UO_1439 (O_1439,N_26695,N_25294);
nand UO_1440 (O_1440,N_28280,N_28173);
xor UO_1441 (O_1441,N_27232,N_28208);
nand UO_1442 (O_1442,N_29244,N_25206);
xnor UO_1443 (O_1443,N_25296,N_26283);
nand UO_1444 (O_1444,N_27397,N_29502);
or UO_1445 (O_1445,N_29546,N_28647);
nor UO_1446 (O_1446,N_26473,N_25020);
nand UO_1447 (O_1447,N_25624,N_29203);
nor UO_1448 (O_1448,N_26835,N_28757);
nor UO_1449 (O_1449,N_28591,N_29037);
or UO_1450 (O_1450,N_27975,N_26272);
nand UO_1451 (O_1451,N_26854,N_27061);
or UO_1452 (O_1452,N_27236,N_28818);
and UO_1453 (O_1453,N_26057,N_29384);
nor UO_1454 (O_1454,N_28829,N_28536);
or UO_1455 (O_1455,N_27607,N_25404);
xor UO_1456 (O_1456,N_25267,N_29359);
nor UO_1457 (O_1457,N_27462,N_27323);
or UO_1458 (O_1458,N_27180,N_25189);
and UO_1459 (O_1459,N_26385,N_27352);
nand UO_1460 (O_1460,N_27248,N_27121);
nor UO_1461 (O_1461,N_25216,N_25832);
and UO_1462 (O_1462,N_28531,N_29720);
and UO_1463 (O_1463,N_26784,N_29446);
nor UO_1464 (O_1464,N_28311,N_25445);
xor UO_1465 (O_1465,N_28627,N_26795);
xor UO_1466 (O_1466,N_25175,N_27790);
xor UO_1467 (O_1467,N_25037,N_26946);
nand UO_1468 (O_1468,N_26714,N_26832);
xnor UO_1469 (O_1469,N_25843,N_27289);
nor UO_1470 (O_1470,N_27425,N_26725);
nor UO_1471 (O_1471,N_29719,N_28512);
and UO_1472 (O_1472,N_25228,N_28343);
nand UO_1473 (O_1473,N_27943,N_27704);
or UO_1474 (O_1474,N_29424,N_26461);
and UO_1475 (O_1475,N_26866,N_27650);
nand UO_1476 (O_1476,N_25501,N_27825);
and UO_1477 (O_1477,N_27431,N_26369);
nand UO_1478 (O_1478,N_29207,N_28908);
xnor UO_1479 (O_1479,N_29947,N_29143);
or UO_1480 (O_1480,N_26691,N_27429);
nand UO_1481 (O_1481,N_28855,N_26039);
nand UO_1482 (O_1482,N_29952,N_29490);
nand UO_1483 (O_1483,N_28148,N_25499);
nor UO_1484 (O_1484,N_26014,N_29286);
nor UO_1485 (O_1485,N_28272,N_29620);
or UO_1486 (O_1486,N_29733,N_29801);
nand UO_1487 (O_1487,N_25465,N_26083);
nor UO_1488 (O_1488,N_27590,N_25934);
nand UO_1489 (O_1489,N_25164,N_26995);
nor UO_1490 (O_1490,N_25852,N_29085);
xnor UO_1491 (O_1491,N_26965,N_27256);
nor UO_1492 (O_1492,N_29661,N_26053);
xnor UO_1493 (O_1493,N_25064,N_26672);
or UO_1494 (O_1494,N_29195,N_26605);
or UO_1495 (O_1495,N_29501,N_27586);
xnor UO_1496 (O_1496,N_27585,N_29470);
nor UO_1497 (O_1497,N_26760,N_25163);
xnor UO_1498 (O_1498,N_25187,N_26782);
nand UO_1499 (O_1499,N_29787,N_29326);
and UO_1500 (O_1500,N_29557,N_29493);
and UO_1501 (O_1501,N_25330,N_25515);
nand UO_1502 (O_1502,N_27699,N_27564);
and UO_1503 (O_1503,N_28406,N_28542);
nand UO_1504 (O_1504,N_27167,N_26018);
nand UO_1505 (O_1505,N_27781,N_26213);
nor UO_1506 (O_1506,N_27182,N_26690);
nand UO_1507 (O_1507,N_26185,N_26289);
nor UO_1508 (O_1508,N_28603,N_25087);
xor UO_1509 (O_1509,N_26594,N_26843);
xnor UO_1510 (O_1510,N_25549,N_26284);
nand UO_1511 (O_1511,N_26645,N_25639);
nor UO_1512 (O_1512,N_28769,N_25720);
and UO_1513 (O_1513,N_29174,N_25022);
and UO_1514 (O_1514,N_26514,N_29878);
xor UO_1515 (O_1515,N_25150,N_29956);
and UO_1516 (O_1516,N_29548,N_29456);
nand UO_1517 (O_1517,N_28357,N_29193);
nand UO_1518 (O_1518,N_29882,N_25385);
and UO_1519 (O_1519,N_25129,N_27989);
nand UO_1520 (O_1520,N_25837,N_25178);
xor UO_1521 (O_1521,N_29511,N_25227);
and UO_1522 (O_1522,N_25827,N_26072);
and UO_1523 (O_1523,N_29517,N_28862);
and UO_1524 (O_1524,N_26932,N_27884);
nor UO_1525 (O_1525,N_29220,N_27346);
or UO_1526 (O_1526,N_26998,N_29707);
nor UO_1527 (O_1527,N_28607,N_26437);
xor UO_1528 (O_1528,N_29084,N_25856);
nand UO_1529 (O_1529,N_25299,N_26689);
and UO_1530 (O_1530,N_28417,N_28304);
nand UO_1531 (O_1531,N_26102,N_25630);
and UO_1532 (O_1532,N_29233,N_26529);
nor UO_1533 (O_1533,N_25188,N_26262);
nand UO_1534 (O_1534,N_26560,N_25767);
nor UO_1535 (O_1535,N_29649,N_27766);
nor UO_1536 (O_1536,N_29103,N_29171);
xnor UO_1537 (O_1537,N_29605,N_27013);
and UO_1538 (O_1538,N_29894,N_27601);
or UO_1539 (O_1539,N_27597,N_27647);
nand UO_1540 (O_1540,N_27114,N_28567);
nand UO_1541 (O_1541,N_26166,N_28206);
and UO_1542 (O_1542,N_28336,N_27075);
or UO_1543 (O_1543,N_29026,N_25293);
xnor UO_1544 (O_1544,N_26625,N_28333);
xor UO_1545 (O_1545,N_26515,N_27221);
xor UO_1546 (O_1546,N_29761,N_28892);
xnor UO_1547 (O_1547,N_28279,N_27530);
or UO_1548 (O_1548,N_29802,N_28441);
and UO_1549 (O_1549,N_28674,N_29857);
nand UO_1550 (O_1550,N_27620,N_28555);
nor UO_1551 (O_1551,N_29452,N_26409);
nand UO_1552 (O_1552,N_25285,N_28255);
and UO_1553 (O_1553,N_28968,N_28425);
or UO_1554 (O_1554,N_27254,N_27993);
xnor UO_1555 (O_1555,N_27638,N_29098);
nor UO_1556 (O_1556,N_27007,N_29716);
nor UO_1557 (O_1557,N_25392,N_29150);
nand UO_1558 (O_1558,N_25065,N_28305);
nor UO_1559 (O_1559,N_29639,N_28722);
and UO_1560 (O_1560,N_26316,N_29348);
and UO_1561 (O_1561,N_26468,N_25834);
nor UO_1562 (O_1562,N_28642,N_26859);
nor UO_1563 (O_1563,N_26339,N_28808);
or UO_1564 (O_1564,N_26797,N_27602);
and UO_1565 (O_1565,N_28920,N_25145);
nor UO_1566 (O_1566,N_27492,N_26184);
nor UO_1567 (O_1567,N_27106,N_28524);
nand UO_1568 (O_1568,N_28493,N_28584);
xor UO_1569 (O_1569,N_28166,N_26257);
and UO_1570 (O_1570,N_28532,N_29275);
nand UO_1571 (O_1571,N_25341,N_28619);
nor UO_1572 (O_1572,N_25456,N_29514);
nand UO_1573 (O_1573,N_28802,N_28303);
or UO_1574 (O_1574,N_27868,N_29129);
nor UO_1575 (O_1575,N_28019,N_25619);
and UO_1576 (O_1576,N_28210,N_27347);
or UO_1577 (O_1577,N_27805,N_29065);
or UO_1578 (O_1578,N_27312,N_26243);
and UO_1579 (O_1579,N_28514,N_28340);
nand UO_1580 (O_1580,N_29800,N_26086);
nand UO_1581 (O_1581,N_25968,N_26747);
and UO_1582 (O_1582,N_27854,N_26415);
or UO_1583 (O_1583,N_25431,N_28576);
xnor UO_1584 (O_1584,N_28568,N_28494);
xnor UO_1585 (O_1585,N_27850,N_28653);
or UO_1586 (O_1586,N_29906,N_29444);
or UO_1587 (O_1587,N_29225,N_25775);
xnor UO_1588 (O_1588,N_28467,N_28681);
or UO_1589 (O_1589,N_28283,N_25569);
xnor UO_1590 (O_1590,N_28990,N_27009);
nand UO_1591 (O_1591,N_26439,N_26579);
or UO_1592 (O_1592,N_26563,N_28186);
xnor UO_1593 (O_1593,N_26247,N_25126);
nor UO_1594 (O_1594,N_26117,N_28104);
nor UO_1595 (O_1595,N_27834,N_25814);
nand UO_1596 (O_1596,N_27624,N_25688);
nand UO_1597 (O_1597,N_26489,N_25190);
nor UO_1598 (O_1598,N_26694,N_28189);
and UO_1599 (O_1599,N_27470,N_29922);
nand UO_1600 (O_1600,N_25311,N_27964);
xnor UO_1601 (O_1601,N_29754,N_25738);
nand UO_1602 (O_1602,N_29936,N_29378);
nand UO_1603 (O_1603,N_28608,N_27278);
xnor UO_1604 (O_1604,N_28452,N_26521);
nand UO_1605 (O_1605,N_28153,N_26153);
or UO_1606 (O_1606,N_25733,N_29726);
nor UO_1607 (O_1607,N_29806,N_27383);
nor UO_1608 (O_1608,N_27986,N_28768);
nor UO_1609 (O_1609,N_26046,N_28506);
nor UO_1610 (O_1610,N_29903,N_28179);
and UO_1611 (O_1611,N_25463,N_28939);
and UO_1612 (O_1612,N_25975,N_27796);
xor UO_1613 (O_1613,N_26210,N_29218);
or UO_1614 (O_1614,N_26223,N_26138);
nor UO_1615 (O_1615,N_25304,N_27507);
xor UO_1616 (O_1616,N_28221,N_27907);
xor UO_1617 (O_1617,N_26474,N_27293);
xor UO_1618 (O_1618,N_29555,N_29428);
and UO_1619 (O_1619,N_26684,N_25554);
nor UO_1620 (O_1620,N_27300,N_28581);
xor UO_1621 (O_1621,N_28662,N_26349);
nand UO_1622 (O_1622,N_29722,N_29820);
xnor UO_1623 (O_1623,N_26352,N_27811);
nor UO_1624 (O_1624,N_29079,N_28519);
xor UO_1625 (O_1625,N_26803,N_26990);
or UO_1626 (O_1626,N_27545,N_26008);
nand UO_1627 (O_1627,N_25018,N_28765);
xnor UO_1628 (O_1628,N_26180,N_26421);
nor UO_1629 (O_1629,N_28985,N_28848);
or UO_1630 (O_1630,N_25159,N_28110);
xor UO_1631 (O_1631,N_27878,N_27379);
nand UO_1632 (O_1632,N_29385,N_26735);
or UO_1633 (O_1633,N_28557,N_25873);
nand UO_1634 (O_1634,N_29689,N_26517);
or UO_1635 (O_1635,N_29354,N_27040);
and UO_1636 (O_1636,N_28537,N_29967);
or UO_1637 (O_1637,N_29049,N_28149);
nor UO_1638 (O_1638,N_25613,N_26871);
xnor UO_1639 (O_1639,N_28200,N_29016);
and UO_1640 (O_1640,N_28008,N_26692);
or UO_1641 (O_1641,N_26591,N_28659);
nor UO_1642 (O_1642,N_29969,N_28754);
xor UO_1643 (O_1643,N_25758,N_29162);
nor UO_1644 (O_1644,N_29862,N_25093);
nor UO_1645 (O_1645,N_27929,N_26245);
nand UO_1646 (O_1646,N_26058,N_26652);
nor UO_1647 (O_1647,N_26287,N_29600);
nand UO_1648 (O_1648,N_26012,N_28503);
xor UO_1649 (O_1649,N_29042,N_29489);
nor UO_1650 (O_1650,N_29366,N_27580);
nand UO_1651 (O_1651,N_25386,N_26666);
xnor UO_1652 (O_1652,N_26446,N_26858);
nand UO_1653 (O_1653,N_28044,N_29984);
and UO_1654 (O_1654,N_28972,N_29933);
or UO_1655 (O_1655,N_28379,N_28941);
nand UO_1656 (O_1656,N_28508,N_29168);
and UO_1657 (O_1657,N_29524,N_25186);
xor UO_1658 (O_1658,N_27557,N_25383);
nand UO_1659 (O_1659,N_25271,N_27452);
nor UO_1660 (O_1660,N_28791,N_27313);
and UO_1661 (O_1661,N_25967,N_25558);
nor UO_1662 (O_1662,N_27905,N_26398);
or UO_1663 (O_1663,N_29108,N_27996);
and UO_1664 (O_1664,N_29419,N_28766);
or UO_1665 (O_1665,N_27046,N_26845);
and UO_1666 (O_1666,N_26404,N_26925);
nand UO_1667 (O_1667,N_26475,N_26789);
nand UO_1668 (O_1668,N_27241,N_25687);
nand UO_1669 (O_1669,N_29866,N_27015);
xnor UO_1670 (O_1670,N_28301,N_26263);
and UO_1671 (O_1671,N_27390,N_29478);
nor UO_1672 (O_1672,N_29698,N_28815);
xnor UO_1673 (O_1673,N_27355,N_25280);
nand UO_1674 (O_1674,N_28665,N_29060);
nand UO_1675 (O_1675,N_26344,N_25074);
nor UO_1676 (O_1676,N_28534,N_28719);
xor UO_1677 (O_1677,N_25492,N_29687);
and UO_1678 (O_1678,N_25418,N_25718);
nor UO_1679 (O_1679,N_27807,N_29334);
or UO_1680 (O_1680,N_27848,N_28814);
nand UO_1681 (O_1681,N_27028,N_26354);
xnor UO_1682 (O_1682,N_29358,N_28349);
nor UO_1683 (O_1683,N_26628,N_26719);
or UO_1684 (O_1684,N_28087,N_29704);
nor UO_1685 (O_1685,N_26219,N_27549);
nand UO_1686 (O_1686,N_27705,N_25038);
and UO_1687 (O_1687,N_25351,N_25194);
xor UO_1688 (O_1688,N_27220,N_27703);
and UO_1689 (O_1689,N_28774,N_26137);
xnor UO_1690 (O_1690,N_26868,N_27518);
nor UO_1691 (O_1691,N_28078,N_27175);
nor UO_1692 (O_1692,N_27504,N_26165);
and UO_1693 (O_1693,N_27752,N_27851);
or UO_1694 (O_1694,N_29771,N_27789);
nand UO_1695 (O_1695,N_27327,N_29746);
xor UO_1696 (O_1696,N_28921,N_28845);
nor UO_1697 (O_1697,N_27668,N_25158);
nand UO_1698 (O_1698,N_28579,N_27230);
nor UO_1699 (O_1699,N_26432,N_27459);
xnor UO_1700 (O_1700,N_25300,N_28631);
nand UO_1701 (O_1701,N_27399,N_27093);
or UO_1702 (O_1702,N_26883,N_26488);
and UO_1703 (O_1703,N_25402,N_26239);
nor UO_1704 (O_1704,N_29392,N_27649);
xor UO_1705 (O_1705,N_28824,N_25277);
and UO_1706 (O_1706,N_27398,N_29615);
xnor UO_1707 (O_1707,N_28950,N_25545);
nor UO_1708 (O_1708,N_27321,N_28033);
xor UO_1709 (O_1709,N_25773,N_26088);
nand UO_1710 (O_1710,N_28614,N_29851);
nand UO_1711 (O_1711,N_27421,N_28055);
nand UO_1712 (O_1712,N_27003,N_26162);
and UO_1713 (O_1713,N_27203,N_26940);
or UO_1714 (O_1714,N_27656,N_28491);
or UO_1715 (O_1715,N_25425,N_26556);
or UO_1716 (O_1716,N_25522,N_28325);
nor UO_1717 (O_1717,N_26606,N_27130);
nor UO_1718 (O_1718,N_26948,N_29073);
nor UO_1719 (O_1719,N_27283,N_26855);
or UO_1720 (O_1720,N_28915,N_26539);
or UO_1721 (O_1721,N_29014,N_27351);
and UO_1722 (O_1722,N_28269,N_26962);
nand UO_1723 (O_1723,N_28805,N_28487);
nand UO_1724 (O_1724,N_29447,N_26877);
or UO_1725 (O_1725,N_28389,N_29308);
or UO_1726 (O_1726,N_28877,N_26801);
or UO_1727 (O_1727,N_29488,N_25743);
nand UO_1728 (O_1728,N_27047,N_28770);
or UO_1729 (O_1729,N_25739,N_29250);
nor UO_1730 (O_1730,N_26277,N_26064);
xor UO_1731 (O_1731,N_25481,N_26359);
nand UO_1732 (O_1732,N_26370,N_29718);
and UO_1733 (O_1733,N_25631,N_28250);
nand UO_1734 (O_1734,N_28257,N_26372);
nand UO_1735 (O_1735,N_29748,N_28414);
and UO_1736 (O_1736,N_27291,N_25701);
xor UO_1737 (O_1737,N_27858,N_28284);
or UO_1738 (O_1738,N_29728,N_29795);
or UO_1739 (O_1739,N_28646,N_25085);
nand UO_1740 (O_1740,N_29177,N_26246);
nor UO_1741 (O_1741,N_28727,N_27436);
xnor UO_1742 (O_1742,N_27773,N_29373);
or UO_1743 (O_1743,N_26902,N_25588);
xor UO_1744 (O_1744,N_29997,N_28787);
nand UO_1745 (O_1745,N_29403,N_29430);
and UO_1746 (O_1746,N_29076,N_26440);
xor UO_1747 (O_1747,N_26577,N_26972);
nand UO_1748 (O_1748,N_27915,N_29958);
and UO_1749 (O_1749,N_28368,N_29062);
nor UO_1750 (O_1750,N_26171,N_28683);
or UO_1751 (O_1751,N_25095,N_29610);
nor UO_1752 (O_1752,N_27944,N_26416);
or UO_1753 (O_1753,N_25831,N_29948);
xor UO_1754 (O_1754,N_26524,N_29115);
nor UO_1755 (O_1755,N_29242,N_25693);
and UO_1756 (O_1756,N_28496,N_26589);
nor UO_1757 (O_1757,N_26954,N_29296);
xor UO_1758 (O_1758,N_26317,N_29197);
or UO_1759 (O_1759,N_25993,N_29119);
and UO_1760 (O_1760,N_27038,N_28032);
nand UO_1761 (O_1761,N_25965,N_27034);
nor UO_1762 (O_1762,N_26253,N_29998);
and UO_1763 (O_1763,N_27630,N_27730);
xnor UO_1764 (O_1764,N_27925,N_27881);
xnor UO_1765 (O_1765,N_28474,N_26004);
or UO_1766 (O_1766,N_25467,N_25766);
and UO_1767 (O_1767,N_29263,N_25409);
nand UO_1768 (O_1768,N_27131,N_25427);
xor UO_1769 (O_1769,N_26630,N_25337);
xor UO_1770 (O_1770,N_29310,N_25417);
and UO_1771 (O_1771,N_29267,N_26164);
xor UO_1772 (O_1772,N_29337,N_26693);
xor UO_1773 (O_1773,N_27906,N_28570);
and UO_1774 (O_1774,N_25584,N_29055);
and UO_1775 (O_1775,N_27451,N_29972);
xnor UO_1776 (O_1776,N_27122,N_29127);
nor UO_1777 (O_1777,N_29740,N_26135);
xnor UO_1778 (O_1778,N_25173,N_25809);
and UO_1779 (O_1779,N_28969,N_27541);
and UO_1780 (O_1780,N_29012,N_28935);
nand UO_1781 (O_1781,N_28951,N_26274);
or UO_1782 (O_1782,N_28776,N_27307);
xor UO_1783 (O_1783,N_25110,N_28030);
nand UO_1784 (O_1784,N_29668,N_25491);
or UO_1785 (O_1785,N_26928,N_27523);
or UO_1786 (O_1786,N_28658,N_29304);
xnor UO_1787 (O_1787,N_26393,N_29421);
or UO_1788 (O_1788,N_29847,N_28785);
and UO_1789 (O_1789,N_29645,N_27196);
nand UO_1790 (O_1790,N_28083,N_26880);
or UO_1791 (O_1791,N_29758,N_25897);
or UO_1792 (O_1792,N_25894,N_28223);
and UO_1793 (O_1793,N_25137,N_27956);
nor UO_1794 (O_1794,N_26401,N_27471);
nor UO_1795 (O_1795,N_27080,N_26386);
nand UO_1796 (O_1796,N_27658,N_29302);
nor UO_1797 (O_1797,N_27166,N_28550);
nor UO_1798 (O_1798,N_28381,N_29307);
nor UO_1799 (O_1799,N_28062,N_26621);
xor UO_1800 (O_1800,N_29120,N_28767);
xnor UO_1801 (O_1801,N_28040,N_27736);
nand UO_1802 (O_1802,N_28270,N_29994);
or UO_1803 (O_1803,N_29935,N_25826);
and UO_1804 (O_1804,N_29034,N_29427);
nand UO_1805 (O_1805,N_29975,N_27272);
and UO_1806 (O_1806,N_29020,N_25225);
xnor UO_1807 (O_1807,N_28919,N_27508);
nor UO_1808 (O_1808,N_28459,N_27741);
nand UO_1809 (O_1809,N_28680,N_25909);
or UO_1810 (O_1810,N_25559,N_29652);
or UO_1811 (O_1811,N_25165,N_29344);
xor UO_1812 (O_1812,N_29423,N_28676);
nand UO_1813 (O_1813,N_25686,N_26796);
nor UO_1814 (O_1814,N_29039,N_28428);
nand UO_1815 (O_1815,N_27437,N_26331);
or UO_1816 (O_1816,N_26244,N_25156);
nand UO_1817 (O_1817,N_25347,N_25374);
nor UO_1818 (O_1818,N_27716,N_28670);
xor UO_1819 (O_1819,N_26966,N_27227);
xnor UO_1820 (O_1820,N_27588,N_25799);
xnor UO_1821 (O_1821,N_26143,N_25301);
or UO_1822 (O_1822,N_26970,N_25112);
and UO_1823 (O_1823,N_25393,N_27621);
nand UO_1824 (O_1824,N_25142,N_29471);
nor UO_1825 (O_1825,N_28026,N_29949);
and UO_1826 (O_1826,N_26991,N_26203);
xor UO_1827 (O_1827,N_26145,N_29315);
nor UO_1828 (O_1828,N_29568,N_25921);
nor UO_1829 (O_1829,N_25068,N_25923);
nand UO_1830 (O_1830,N_29662,N_28442);
and UO_1831 (O_1831,N_27426,N_29767);
and UO_1832 (O_1832,N_29117,N_25207);
or UO_1833 (O_1833,N_26211,N_29346);
xnor UO_1834 (O_1834,N_26267,N_29165);
nand UO_1835 (O_1835,N_26581,N_28111);
or UO_1836 (O_1836,N_27097,N_27517);
nand UO_1837 (O_1837,N_28380,N_28910);
and UO_1838 (O_1838,N_27567,N_25570);
and UO_1839 (O_1839,N_25050,N_29694);
xnor UO_1840 (O_1840,N_25372,N_26410);
nand UO_1841 (O_1841,N_28312,N_28232);
nor UO_1842 (O_1842,N_28775,N_26230);
and UO_1843 (O_1843,N_26408,N_25442);
xnor UO_1844 (O_1844,N_28480,N_28773);
and UO_1845 (O_1845,N_26994,N_28320);
and UO_1846 (O_1846,N_26271,N_29353);
and UO_1847 (O_1847,N_29057,N_29160);
or UO_1848 (O_1848,N_27939,N_25960);
nor UO_1849 (O_1849,N_26520,N_25910);
nor UO_1850 (O_1850,N_26727,N_26435);
or UO_1851 (O_1851,N_29875,N_28502);
and UO_1852 (O_1852,N_29101,N_26512);
nand UO_1853 (O_1853,N_27810,N_26982);
and UO_1854 (O_1854,N_26822,N_27500);
xnor UO_1855 (O_1855,N_29685,N_27052);
and UO_1856 (O_1856,N_27945,N_29237);
or UO_1857 (O_1857,N_26717,N_27584);
nor UO_1858 (O_1858,N_27767,N_28888);
nand UO_1859 (O_1859,N_27110,N_28109);
nand UO_1860 (O_1860,N_29549,N_26905);
xnor UO_1861 (O_1861,N_26081,N_28561);
and UO_1862 (O_1862,N_25039,N_27090);
and UO_1863 (O_1863,N_26191,N_25917);
and UO_1864 (O_1864,N_26837,N_28011);
and UO_1865 (O_1865,N_29090,N_28735);
and UO_1866 (O_1866,N_25971,N_25566);
nor UO_1867 (O_1867,N_28782,N_26097);
and UO_1868 (O_1868,N_27065,N_29798);
nor UO_1869 (O_1869,N_27717,N_29048);
xnor UO_1870 (O_1870,N_26382,N_25920);
nor UO_1871 (O_1871,N_25185,N_26842);
or UO_1872 (O_1872,N_29991,N_29229);
nand UO_1873 (O_1873,N_27162,N_26362);
and UO_1874 (O_1874,N_26445,N_29189);
nor UO_1875 (O_1875,N_28461,N_25133);
nor UO_1876 (O_1876,N_29413,N_29031);
and UO_1877 (O_1877,N_27867,N_28385);
nand UO_1878 (O_1878,N_27045,N_26215);
and UO_1879 (O_1879,N_25725,N_29032);
xor UO_1880 (O_1880,N_27829,N_27755);
xnor UO_1881 (O_1881,N_26511,N_28300);
nand UO_1882 (O_1882,N_25769,N_26898);
nand UO_1883 (O_1883,N_28170,N_27217);
and UO_1884 (O_1884,N_25634,N_27336);
nor UO_1885 (O_1885,N_27281,N_27494);
and UO_1886 (O_1886,N_29149,N_25344);
nand UO_1887 (O_1887,N_25986,N_28723);
and UO_1888 (O_1888,N_27295,N_26054);
xor UO_1889 (O_1889,N_29516,N_26723);
xor UO_1890 (O_1890,N_29655,N_26355);
or UO_1891 (O_1891,N_28436,N_28837);
nand UO_1892 (O_1892,N_25638,N_28585);
or UO_1893 (O_1893,N_25672,N_25011);
and UO_1894 (O_1894,N_27498,N_28181);
nor UO_1895 (O_1895,N_26364,N_27059);
nor UO_1896 (O_1896,N_28702,N_26934);
nor UO_1897 (O_1897,N_27369,N_29817);
nand UO_1898 (O_1898,N_25660,N_29368);
nor UO_1899 (O_1899,N_28669,N_25497);
xnor UO_1900 (O_1900,N_25915,N_27957);
nand UO_1901 (O_1901,N_28079,N_26766);
nand UO_1902 (O_1902,N_26895,N_27515);
nor UO_1903 (O_1903,N_26281,N_29112);
nand UO_1904 (O_1904,N_25081,N_26441);
nor UO_1905 (O_1905,N_26670,N_29696);
and UO_1906 (O_1906,N_27749,N_28157);
nor UO_1907 (O_1907,N_29350,N_27113);
or UO_1908 (O_1908,N_29099,N_28369);
and UO_1909 (O_1909,N_25489,N_26186);
xor UO_1910 (O_1910,N_26325,N_26380);
xnor UO_1911 (O_1911,N_28384,N_26037);
nand UO_1912 (O_1912,N_27733,N_25561);
nor UO_1913 (O_1913,N_27554,N_29270);
and UO_1914 (O_1914,N_25851,N_25072);
and UO_1915 (O_1915,N_27916,N_28909);
xnor UO_1916 (O_1916,N_27866,N_27420);
xnor UO_1917 (O_1917,N_27201,N_26127);
and UO_1918 (O_1918,N_27758,N_28742);
nor UO_1919 (O_1919,N_28392,N_28691);
and UO_1920 (O_1920,N_28234,N_28114);
xor UO_1921 (O_1921,N_29464,N_25940);
nor UO_1922 (O_1922,N_27972,N_28126);
nor UO_1923 (O_1923,N_25001,N_26673);
nand UO_1924 (O_1924,N_29010,N_28510);
or UO_1925 (O_1925,N_29169,N_27744);
xor UO_1926 (O_1926,N_25530,N_29838);
nor UO_1927 (O_1927,N_25340,N_25680);
nor UO_1928 (O_1928,N_28763,N_25740);
or UO_1929 (O_1929,N_29986,N_29331);
or UO_1930 (O_1930,N_28154,N_27138);
or UO_1931 (O_1931,N_25066,N_27718);
nor UO_1932 (O_1932,N_29843,N_25325);
xor UO_1933 (O_1933,N_28347,N_26513);
or UO_1934 (O_1934,N_26711,N_27035);
and UO_1935 (O_1935,N_28734,N_27898);
nand UO_1936 (O_1936,N_26981,N_29822);
nand UO_1937 (O_1937,N_26084,N_27690);
or UO_1938 (O_1938,N_27375,N_29113);
xnor UO_1939 (O_1939,N_28564,N_26259);
and UO_1940 (O_1940,N_26228,N_28821);
and UO_1941 (O_1941,N_27358,N_26791);
nand UO_1942 (O_1942,N_26216,N_25459);
and UO_1943 (O_1943,N_28672,N_29732);
and UO_1944 (O_1944,N_28793,N_28460);
or UO_1945 (O_1945,N_25067,N_29122);
and UO_1946 (O_1946,N_25607,N_26663);
xnor UO_1947 (O_1947,N_28810,N_26049);
nand UO_1948 (O_1948,N_25214,N_25603);
and UO_1949 (O_1949,N_29491,N_27194);
nor UO_1950 (O_1950,N_25168,N_27453);
and UO_1951 (O_1951,N_25047,N_29796);
nand UO_1952 (O_1952,N_28064,N_25702);
nor UO_1953 (O_1953,N_25543,N_26343);
xnor UO_1954 (O_1954,N_25352,N_29850);
and UO_1955 (O_1955,N_26674,N_27764);
or UO_1956 (O_1956,N_28737,N_29484);
nand UO_1957 (O_1957,N_26077,N_26927);
nand UO_1958 (O_1958,N_26487,N_26298);
nand UO_1959 (O_1959,N_26933,N_27961);
xor UO_1960 (O_1960,N_26649,N_26220);
xor UO_1961 (O_1961,N_28135,N_27615);
nand UO_1962 (O_1962,N_28059,N_27025);
nor UO_1963 (O_1963,N_27904,N_26459);
xor UO_1964 (O_1964,N_28582,N_29842);
or UO_1965 (O_1965,N_26665,N_25542);
nor UO_1966 (O_1966,N_25429,N_27408);
and UO_1967 (O_1967,N_29510,N_29644);
xnor UO_1968 (O_1968,N_25071,N_29481);
or UO_1969 (O_1969,N_29813,N_27723);
or UO_1970 (O_1970,N_29451,N_28852);
xnor UO_1971 (O_1971,N_25963,N_26141);
nand UO_1972 (O_1972,N_26176,N_26951);
and UO_1973 (O_1973,N_26036,N_29474);
and UO_1974 (O_1974,N_27726,N_25944);
and UO_1975 (O_1975,N_27893,N_25629);
nor UO_1976 (O_1976,N_25783,N_29463);
nor UO_1977 (O_1977,N_25316,N_25461);
nand UO_1978 (O_1978,N_29017,N_29861);
nor UO_1979 (O_1979,N_27918,N_28097);
nor UO_1980 (O_1980,N_28375,N_28432);
nand UO_1981 (O_1981,N_28835,N_25348);
nor UO_1982 (O_1982,N_28410,N_25298);
nor UO_1983 (O_1983,N_27076,N_27670);
and UO_1984 (O_1984,N_27865,N_26198);
nand UO_1985 (O_1985,N_29303,N_29710);
and UO_1986 (O_1986,N_29635,N_26609);
and UO_1987 (O_1987,N_25853,N_25964);
xnor UO_1988 (O_1988,N_27890,N_26656);
or UO_1989 (O_1989,N_25162,N_25389);
or UO_1990 (O_1990,N_29977,N_29919);
nand UO_1991 (O_1991,N_25864,N_27463);
or UO_1992 (O_1992,N_29900,N_26608);
xor UO_1993 (O_1993,N_25807,N_26599);
xnor UO_1994 (O_1994,N_28278,N_28894);
xor UO_1995 (O_1995,N_27154,N_25375);
and UO_1996 (O_1996,N_29755,N_27565);
or UO_1997 (O_1997,N_26973,N_27857);
or UO_1998 (O_1998,N_26658,N_29440);
nand UO_1999 (O_1999,N_29264,N_25665);
nor UO_2000 (O_2000,N_28696,N_25244);
nor UO_2001 (O_2001,N_29454,N_25212);
nand UO_2002 (O_2002,N_29540,N_26497);
or UO_2003 (O_2003,N_29563,N_25014);
and UO_2004 (O_2004,N_28750,N_25128);
and UO_2005 (O_2005,N_29951,N_25054);
nand UO_2006 (O_2006,N_29844,N_29601);
xor UO_2007 (O_2007,N_28731,N_29709);
and UO_2008 (O_2008,N_26163,N_29306);
nand UO_2009 (O_2009,N_27571,N_28018);
or UO_2010 (O_2010,N_26644,N_27981);
nand UO_2011 (O_2011,N_29865,N_26139);
xnor UO_2012 (O_2012,N_27356,N_29837);
and UO_2013 (O_2013,N_28287,N_26226);
nor UO_2014 (O_2014,N_28116,N_25262);
nand UO_2015 (O_2015,N_27305,N_29288);
and UO_2016 (O_2016,N_27449,N_25576);
xor UO_2017 (O_2017,N_28954,N_27482);
nand UO_2018 (O_2018,N_29674,N_26071);
nor UO_2019 (O_2019,N_26533,N_25621);
nand UO_2020 (O_2020,N_26781,N_26241);
nor UO_2021 (O_2021,N_29161,N_25199);
nor UO_2022 (O_2022,N_26043,N_27158);
nand UO_2023 (O_2023,N_25748,N_27415);
nand UO_2024 (O_2024,N_25495,N_26923);
nand UO_2025 (O_2025,N_28421,N_27843);
and UO_2026 (O_2026,N_28651,N_28991);
and UO_2027 (O_2027,N_29380,N_27012);
or UO_2028 (O_2028,N_29576,N_28617);
and UO_2029 (O_2029,N_28553,N_28457);
nor UO_2030 (O_2030,N_28216,N_25016);
nor UO_2031 (O_2031,N_25751,N_25902);
xnor UO_2032 (O_2032,N_27941,N_29248);
nor UO_2033 (O_2033,N_29616,N_29043);
nor UO_2034 (O_2034,N_28856,N_27469);
nor UO_2035 (O_2035,N_27183,N_26891);
nor UO_2036 (O_2036,N_28648,N_29323);
nor UO_2037 (O_2037,N_27297,N_27697);
nand UO_2038 (O_2038,N_25291,N_28402);
nor UO_2039 (O_2039,N_27966,N_25935);
or UO_2040 (O_2040,N_27863,N_28762);
xor UO_2041 (O_2041,N_28714,N_28172);
nor UO_2042 (O_2042,N_27747,N_28332);
xnor UO_2043 (O_2043,N_26454,N_26664);
nand UO_2044 (O_2044,N_27869,N_25510);
nor UO_2045 (O_2045,N_26646,N_27611);
nand UO_2046 (O_2046,N_29442,N_25958);
nor UO_2047 (O_2047,N_27973,N_27771);
nand UO_2048 (O_2048,N_29790,N_27388);
xnor UO_2049 (O_2049,N_26205,N_25768);
or UO_2050 (O_2050,N_27329,N_27411);
nor UO_2051 (O_2051,N_28799,N_25669);
xor UO_2052 (O_2052,N_28507,N_28632);
or UO_2053 (O_2053,N_25146,N_28144);
and UO_2054 (O_2054,N_26988,N_26537);
and UO_2055 (O_2055,N_26396,N_25796);
xor UO_2056 (O_2056,N_25281,N_27513);
xor UO_2057 (O_2057,N_25482,N_26936);
and UO_2058 (O_2058,N_26882,N_26958);
and UO_2059 (O_2059,N_29654,N_25336);
xnor UO_2060 (O_2060,N_29227,N_25086);
nor UO_2061 (O_2061,N_25313,N_29041);
or UO_2062 (O_2062,N_25115,N_25857);
xnor UO_2063 (O_2063,N_27815,N_26056);
xor UO_2064 (O_2064,N_26356,N_26067);
xnor UO_2065 (O_2065,N_25319,N_25977);
or UO_2066 (O_2066,N_27632,N_25787);
nand UO_2067 (O_2067,N_29291,N_25154);
and UO_2068 (O_2068,N_25117,N_28167);
or UO_2069 (O_2069,N_27412,N_28471);
nor UO_2070 (O_2070,N_26518,N_28709);
xnor UO_2071 (O_2071,N_27264,N_25045);
nor UO_2072 (O_2072,N_26079,N_27190);
nand UO_2073 (O_2073,N_27193,N_28751);
or UO_2074 (O_2074,N_27082,N_27081);
nand UO_2075 (O_2075,N_25260,N_28443);
nand UO_2076 (O_2076,N_26757,N_26131);
or UO_2077 (O_2077,N_28903,N_25353);
and UO_2078 (O_2078,N_28088,N_26063);
xor UO_2079 (O_2079,N_29663,N_27253);
nand UO_2080 (O_2080,N_28124,N_25833);
nor UO_2081 (O_2081,N_26174,N_26496);
xor UO_2082 (O_2082,N_27128,N_26527);
xnor UO_2083 (O_2083,N_25447,N_26152);
or UO_2084 (O_2084,N_28071,N_29477);
nor UO_2085 (O_2085,N_27189,N_29336);
or UO_2086 (O_2086,N_26984,N_29521);
nor UO_2087 (O_2087,N_29753,N_27579);
xnor UO_2088 (O_2088,N_25529,N_27284);
nand UO_2089 (O_2089,N_28960,N_25003);
nor UO_2090 (O_2090,N_25312,N_29912);
or UO_2091 (O_2091,N_29259,N_25785);
nand UO_2092 (O_2092,N_27835,N_25031);
xor UO_2093 (O_2093,N_26306,N_28012);
nand UO_2094 (O_2094,N_28201,N_28759);
nor UO_2095 (O_2095,N_28955,N_29235);
or UO_2096 (O_2096,N_25371,N_29102);
nand UO_2097 (O_2097,N_28023,N_28140);
and UO_2098 (O_2098,N_27883,N_29976);
nand UO_2099 (O_2099,N_28299,N_26426);
nand UO_2100 (O_2100,N_25464,N_26553);
xor UO_2101 (O_2101,N_29624,N_26875);
xnor UO_2102 (O_2102,N_26839,N_29943);
and UO_2103 (O_2103,N_29695,N_28203);
nor UO_2104 (O_2104,N_27833,N_27005);
and UO_2105 (O_2105,N_26085,N_25032);
xnor UO_2106 (O_2106,N_26275,N_29289);
and UO_2107 (O_2107,N_25752,N_25878);
nor UO_2108 (O_2108,N_26979,N_28222);
or UO_2109 (O_2109,N_25040,N_27636);
nor UO_2110 (O_2110,N_27337,N_26572);
and UO_2111 (O_2111,N_25932,N_26324);
nand UO_2112 (O_2112,N_29068,N_29992);
xnor UO_2113 (O_2113,N_26501,N_26411);
or UO_2114 (O_2114,N_29186,N_28807);
nand UO_2115 (O_2115,N_28540,N_26376);
xor UO_2116 (O_2116,N_28408,N_28335);
xnor UO_2117 (O_2117,N_26329,N_29535);
or UO_2118 (O_2118,N_25589,N_25550);
or UO_2119 (O_2119,N_28476,N_25802);
nand UO_2120 (O_2120,N_27969,N_26943);
nand UO_2121 (O_2121,N_29125,N_28253);
nor UO_2122 (O_2122,N_27634,N_25945);
nor UO_2123 (O_2123,N_28475,N_25119);
nor UO_2124 (O_2124,N_29911,N_25378);
nand UO_2125 (O_2125,N_26724,N_26187);
nand UO_2126 (O_2126,N_26661,N_29356);
xnor UO_2127 (O_2127,N_26703,N_25952);
and UO_2128 (O_2128,N_26929,N_27512);
and UO_2129 (O_2129,N_28254,N_28050);
nor UO_2130 (O_2130,N_27958,N_25308);
nand UO_2131 (O_2131,N_26921,N_28628);
nand UO_2132 (O_2132,N_27821,N_29745);
nor UO_2133 (O_2133,N_29656,N_26295);
or UO_2134 (O_2134,N_27521,N_29136);
or UO_2135 (O_2135,N_28028,N_28947);
and UO_2136 (O_2136,N_26336,N_28795);
or UO_2137 (O_2137,N_25602,N_29807);
xor UO_2138 (O_2138,N_26155,N_27092);
or UO_2139 (O_2139,N_27798,N_26469);
or UO_2140 (O_2140,N_26978,N_27688);
nand UO_2141 (O_2141,N_29518,N_28533);
nand UO_2142 (O_2142,N_29013,N_27800);
nor UO_2143 (O_2143,N_26493,N_27715);
xor UO_2144 (O_2144,N_27546,N_28065);
or UO_2145 (O_2145,N_29612,N_29301);
xor UO_2146 (O_2146,N_29401,N_25907);
nor UO_2147 (O_2147,N_25358,N_25368);
nor UO_2148 (O_2148,N_29211,N_26041);
or UO_2149 (O_2149,N_26495,N_26453);
nand UO_2150 (O_2150,N_25407,N_27215);
or UO_2151 (O_2151,N_28143,N_26301);
and UO_2152 (O_2152,N_27574,N_25821);
or UO_2153 (O_2153,N_25317,N_28753);
or UO_2154 (O_2154,N_25094,N_27271);
and UO_2155 (O_2155,N_26912,N_28760);
and UO_2156 (O_2156,N_29507,N_27468);
nor UO_2157 (O_2157,N_29355,N_26583);
and UO_2158 (O_2158,N_29901,N_25012);
nand UO_2159 (O_2159,N_25070,N_29587);
nor UO_2160 (O_2160,N_25657,N_25713);
and UO_2161 (O_2161,N_25749,N_27382);
xnor UO_2162 (O_2162,N_26170,N_28554);
nand UO_2163 (O_2163,N_27063,N_29823);
or UO_2164 (O_2164,N_27414,N_29558);
or UO_2165 (O_2165,N_27143,N_25416);
nor UO_2166 (O_2166,N_25179,N_27663);
or UO_2167 (O_2167,N_29739,N_28198);
xor UO_2168 (O_2168,N_27608,N_25556);
or UO_2169 (O_2169,N_27202,N_26009);
nor UO_2170 (O_2170,N_29232,N_26505);
nand UO_2171 (O_2171,N_25073,N_25882);
nand UO_2172 (O_2172,N_27818,N_28182);
nand UO_2173 (O_2173,N_27681,N_25419);
and UO_2174 (O_2174,N_28998,N_25091);
or UO_2175 (O_2175,N_27724,N_27641);
nor UO_2176 (O_2176,N_25098,N_25976);
nand UO_2177 (O_2177,N_28989,N_27364);
nand UO_2178 (O_2178,N_28196,N_26173);
xnor UO_2179 (O_2179,N_29867,N_29859);
nand UO_2180 (O_2180,N_29273,N_26285);
or UO_2181 (O_2181,N_29575,N_29702);
xor UO_2182 (O_2182,N_25895,N_27572);
and UO_2183 (O_2183,N_29027,N_29372);
and UO_2184 (O_2184,N_25380,N_27191);
xor UO_2185 (O_2185,N_28974,N_25678);
or UO_2186 (O_2186,N_28445,N_29789);
xnor UO_2187 (O_2187,N_25422,N_27801);
xnor UO_2188 (O_2188,N_25211,N_29619);
nand UO_2189 (O_2189,N_28396,N_28948);
nand UO_2190 (O_2190,N_25106,N_28780);
nor UO_2191 (O_2191,N_27372,N_27839);
nor UO_2192 (O_2192,N_28251,N_29104);
and UO_2193 (O_2193,N_29339,N_29238);
xor UO_2194 (O_2194,N_26792,N_29570);
nor UO_2195 (O_2195,N_26156,N_29500);
and UO_2196 (O_2196,N_28070,N_28883);
or UO_2197 (O_2197,N_27205,N_25276);
nand UO_2198 (O_2198,N_26017,N_28596);
or UO_2199 (O_2199,N_29993,N_28559);
or UO_2200 (O_2200,N_29021,N_29829);
or UO_2201 (O_2201,N_25349,N_29809);
xnor UO_2202 (O_2202,N_25172,N_26095);
xor UO_2203 (O_2203,N_27448,N_26826);
or UO_2204 (O_2204,N_25953,N_29075);
or UO_2205 (O_2205,N_29757,N_26708);
nor UO_2206 (O_2206,N_25226,N_26700);
or UO_2207 (O_2207,N_29853,N_25625);
nor UO_2208 (O_2208,N_28372,N_29595);
nor UO_2209 (O_2209,N_28626,N_25171);
and UO_2210 (O_2210,N_27197,N_27262);
nand UO_2211 (O_2211,N_29483,N_28113);
xor UO_2212 (O_2212,N_28995,N_26710);
or UO_2213 (O_2213,N_29808,N_29585);
xnor UO_2214 (O_2214,N_25560,N_29439);
or UO_2215 (O_2215,N_28437,N_27953);
and UO_2216 (O_2216,N_26918,N_29623);
or UO_2217 (O_2217,N_27606,N_25992);
or UO_2218 (O_2218,N_29015,N_25819);
nor UO_2219 (O_2219,N_27784,N_29971);
nor UO_2220 (O_2220,N_25493,N_26034);
or UO_2221 (O_2221,N_29184,N_26338);
or UO_2222 (O_2222,N_25840,N_26302);
nand UO_2223 (O_2223,N_27428,N_28463);
and UO_2224 (O_2224,N_25681,N_28041);
and UO_2225 (O_2225,N_27914,N_28138);
nand UO_2226 (O_2226,N_29560,N_27595);
nor UO_2227 (O_2227,N_27213,N_29786);
and UO_2228 (O_2228,N_27021,N_29965);
xnor UO_2229 (O_2229,N_29191,N_26570);
nor UO_2230 (O_2230,N_29260,N_28846);
and UO_2231 (O_2231,N_26472,N_26470);
nor UO_2232 (O_2232,N_29070,N_29599);
or UO_2233 (O_2233,N_25096,N_29142);
and UO_2234 (O_2234,N_26261,N_26573);
nand UO_2235 (O_2235,N_25009,N_28663);
nor UO_2236 (O_2236,N_29774,N_25460);
and UO_2237 (O_2237,N_25746,N_27127);
or UO_2238 (O_2238,N_26193,N_26273);
nand UO_2239 (O_2239,N_25103,N_29697);
or UO_2240 (O_2240,N_28556,N_25111);
nand UO_2241 (O_2241,N_25438,N_28707);
or UO_2242 (O_2242,N_26831,N_28764);
xnor UO_2243 (O_2243,N_28448,N_26585);
and UO_2244 (O_2244,N_28416,N_26510);
or UO_2245 (O_2245,N_26748,N_26236);
nand UO_2246 (O_2246,N_27635,N_28522);
nor UO_2247 (O_2247,N_25822,N_26055);
and UO_2248 (O_2248,N_26045,N_26326);
nand UO_2249 (O_2249,N_27599,N_28039);
and UO_2250 (O_2250,N_27495,N_26029);
and UO_2251 (O_2251,N_28382,N_29675);
xor UO_2252 (O_2252,N_28455,N_25204);
and UO_2253 (O_2253,N_29884,N_28478);
nor UO_2254 (O_2254,N_29154,N_29630);
xor UO_2255 (O_2255,N_26294,N_27679);
or UO_2256 (O_2256,N_28074,N_25626);
and UO_2257 (O_2257,N_27922,N_28197);
or UO_2258 (O_2258,N_27675,N_25605);
and UO_2259 (O_2259,N_28447,N_28635);
nand UO_2260 (O_2260,N_27384,N_25666);
nand UO_2261 (O_2261,N_29132,N_25633);
xnor UO_2262 (O_2262,N_28288,N_28293);
nor UO_2263 (O_2263,N_25704,N_29891);
nor UO_2264 (O_2264,N_28942,N_26070);
xnor UO_2265 (O_2265,N_27653,N_26248);
or UO_2266 (O_2266,N_28456,N_25213);
nor UO_2267 (O_2267,N_28233,N_28145);
xnor UO_2268 (O_2268,N_26959,N_28473);
nor UO_2269 (O_2269,N_29363,N_29201);
xnor UO_2270 (O_2270,N_27163,N_26989);
and UO_2271 (O_2271,N_27671,N_27222);
and UO_2272 (O_2272,N_28710,N_27392);
or UO_2273 (O_2273,N_25525,N_27144);
nor UO_2274 (O_2274,N_25676,N_25196);
xor UO_2275 (O_2275,N_25995,N_26471);
and UO_2276 (O_2276,N_28962,N_29329);
nand UO_2277 (O_2277,N_27499,N_27419);
nor UO_2278 (O_2278,N_25696,N_27603);
nand UO_2279 (O_2279,N_28356,N_29156);
or UO_2280 (O_2280,N_28703,N_25000);
nor UO_2281 (O_2281,N_26545,N_26848);
or UO_2282 (O_2282,N_25757,N_25414);
xnor UO_2283 (O_2283,N_25513,N_29897);
xor UO_2284 (O_2284,N_28772,N_27938);
xor UO_2285 (O_2285,N_28777,N_28675);
and UO_2286 (O_2286,N_26767,N_29410);
nor UO_2287 (O_2287,N_25880,N_26679);
xnor UO_2288 (O_2288,N_26732,N_25871);
xnor UO_2289 (O_2289,N_27442,N_28889);
nand UO_2290 (O_2290,N_28281,N_26836);
nor UO_2291 (O_2291,N_25677,N_26834);
or UO_2292 (O_2292,N_28244,N_26647);
xor UO_2293 (O_2293,N_26769,N_25483);
or UO_2294 (O_2294,N_26651,N_28850);
and UO_2295 (O_2295,N_27842,N_29550);
nand UO_2296 (O_2296,N_29166,N_27152);
or UO_2297 (O_2297,N_28511,N_26754);
xnor UO_2298 (O_2298,N_29255,N_28407);
nand UO_2299 (O_2299,N_28202,N_25805);
and UO_2300 (O_2300,N_25177,N_26389);
xor UO_2301 (O_2301,N_27050,N_26038);
nor UO_2302 (O_2302,N_28758,N_26596);
nor UO_2303 (O_2303,N_28214,N_26707);
nor UO_2304 (O_2304,N_26567,N_26367);
or UO_2305 (O_2305,N_28034,N_26048);
or UO_2306 (O_2306,N_27086,N_27011);
nand UO_2307 (O_2307,N_28373,N_25636);
and UO_2308 (O_2308,N_27998,N_27665);
nand UO_2309 (O_2309,N_26129,N_25870);
xnor UO_2310 (O_2310,N_28163,N_29791);
nand UO_2311 (O_2311,N_27870,N_28928);
xnor UO_2312 (O_2312,N_26251,N_28328);
or UO_2313 (O_2313,N_27558,N_28916);
or UO_2314 (O_2314,N_25901,N_25114);
xor UO_2315 (O_2315,N_25823,N_25519);
nor UO_2316 (O_2316,N_25426,N_29050);
and UO_2317 (O_2317,N_28310,N_25591);
and UO_2318 (O_2318,N_25988,N_26869);
xor UO_2319 (O_2319,N_25592,N_28899);
nand UO_2320 (O_2320,N_27159,N_26687);
nor UO_2321 (O_2321,N_28733,N_25670);
xor UO_2322 (O_2322,N_26463,N_26824);
nor UO_2323 (O_2323,N_27919,N_27343);
or UO_2324 (O_2324,N_27562,N_28832);
nand UO_2325 (O_2325,N_25866,N_27115);
or UO_2326 (O_2326,N_27274,N_26830);
and UO_2327 (O_2327,N_26873,N_26434);
nor UO_2328 (O_2328,N_27684,N_29412);
and UO_2329 (O_2329,N_26730,N_25490);
xor UO_2330 (O_2330,N_28741,N_28612);
and UO_2331 (O_2331,N_27275,N_29438);
nor UO_2332 (O_2332,N_26595,N_25528);
nor UO_2333 (O_2333,N_29131,N_26753);
xor UO_2334 (O_2334,N_27847,N_29673);
nor UO_2335 (O_2335,N_27270,N_25387);
nor UO_2336 (O_2336,N_28527,N_28901);
xnor UO_2337 (O_2337,N_29628,N_29320);
xnor UO_2338 (O_2338,N_26900,N_25373);
and UO_2339 (O_2339,N_29768,N_27860);
or UO_2340 (O_2340,N_27763,N_27132);
nand UO_2341 (O_2341,N_27396,N_29351);
xor UO_2342 (O_2342,N_28953,N_25046);
nor UO_2343 (O_2343,N_27979,N_28117);
nor UO_2344 (O_2344,N_28866,N_28449);
and UO_2345 (O_2345,N_28736,N_28979);
and UO_2346 (O_2346,N_25219,N_29425);
xnor UO_2347 (O_2347,N_26914,N_27467);
or UO_2348 (O_2348,N_26260,N_29915);
and UO_2349 (O_2349,N_26653,N_27067);
or UO_2350 (O_2350,N_25538,N_26612);
or UO_2351 (O_2351,N_27803,N_26066);
nor UO_2352 (O_2352,N_29869,N_28831);
nor UO_2353 (O_2353,N_25692,N_25611);
and UO_2354 (O_2354,N_25818,N_25423);
nor UO_2355 (O_2355,N_28315,N_26332);
or UO_2356 (O_2356,N_27999,N_28123);
xor UO_2357 (O_2357,N_27151,N_27648);
or UO_2358 (O_2358,N_29321,N_26420);
or UO_2359 (O_2359,N_26743,N_27534);
nor UO_2360 (O_2360,N_29194,N_28984);
or UO_2361 (O_2361,N_27141,N_26744);
nand UO_2362 (O_2362,N_28054,N_27519);
and UO_2363 (O_2363,N_29105,N_29445);
xnor UO_2364 (O_2364,N_28784,N_28610);
nand UO_2365 (O_2365,N_28980,N_27889);
nor UO_2366 (O_2366,N_25956,N_27266);
nand UO_2367 (O_2367,N_25926,N_28228);
nor UO_2368 (O_2368,N_29607,N_29666);
or UO_2369 (O_2369,N_27296,N_27104);
and UO_2370 (O_2370,N_27484,N_27101);
xnor UO_2371 (O_2371,N_27613,N_28429);
and UO_2372 (O_2372,N_27583,N_28595);
or UO_2373 (O_2373,N_27089,N_26886);
and UO_2374 (O_2374,N_28354,N_27728);
or UO_2375 (O_2375,N_26597,N_29632);
nand UO_2376 (O_2376,N_26465,N_28761);
and UO_2377 (O_2377,N_25514,N_28549);
nor UO_2378 (O_2378,N_29239,N_29004);
nor UO_2379 (O_2379,N_27427,N_27445);
xor UO_2380 (O_2380,N_29328,N_27245);
or UO_2381 (O_2381,N_28217,N_25886);
or UO_2382 (O_2382,N_29945,N_27148);
xnor UO_2383 (O_2383,N_27413,N_27617);
or UO_2384 (O_2384,N_25029,N_27306);
and UO_2385 (O_2385,N_26212,N_28265);
or UO_2386 (O_2386,N_26154,N_26823);
xor UO_2387 (O_2387,N_29914,N_27959);
or UO_2388 (O_2388,N_26538,N_25121);
nor UO_2389 (O_2389,N_28830,N_28465);
or UO_2390 (O_2390,N_29530,N_27604);
nor UO_2391 (O_2391,N_27367,N_27873);
nand UO_2392 (O_2392,N_28164,N_25759);
or UO_2393 (O_2393,N_28337,N_28604);
xor UO_2394 (O_2394,N_25745,N_25302);
xor UO_2395 (O_2395,N_29941,N_29340);
and UO_2396 (O_2396,N_29415,N_27032);
xnor UO_2397 (O_2397,N_29534,N_29311);
xnor UO_2398 (O_2398,N_29374,N_26069);
nand UO_2399 (O_2399,N_27476,N_26040);
and UO_2400 (O_2400,N_25295,N_27547);
xor UO_2401 (O_2401,N_29887,N_28187);
or UO_2402 (O_2402,N_28231,N_29938);
nor UO_2403 (O_2403,N_26001,N_25793);
nand UO_2404 (O_2404,N_28132,N_28623);
xnor UO_2405 (O_2405,N_26554,N_26348);
xnor UO_2406 (O_2406,N_26377,N_27694);
xor UO_2407 (O_2407,N_26543,N_27721);
or UO_2408 (O_2408,N_26402,N_29367);
or UO_2409 (O_2409,N_25859,N_27386);
or UO_2410 (O_2410,N_28038,N_26775);
and UO_2411 (O_2411,N_28724,N_26235);
nand UO_2412 (O_2412,N_28185,N_28159);
nor UO_2413 (O_2413,N_26812,N_28069);
xnor UO_2414 (O_2414,N_27177,N_26915);
nand UO_2415 (O_2415,N_28485,N_29816);
nor UO_2416 (O_2416,N_27477,N_29182);
nor UO_2417 (O_2417,N_29870,N_28353);
xor UO_2418 (O_2418,N_29631,N_29059);
and UO_2419 (O_2419,N_29133,N_28274);
nor UO_2420 (O_2420,N_27661,N_26122);
or UO_2421 (O_2421,N_29002,N_25449);
nor UO_2422 (O_2422,N_27246,N_27136);
or UO_2423 (O_2423,N_28103,N_29222);
nor UO_2424 (O_2424,N_25661,N_26820);
xor UO_2425 (O_2425,N_26985,N_27117);
nor UO_2426 (O_2426,N_28237,N_29542);
nand UO_2427 (O_2427,N_28563,N_27837);
and UO_2428 (O_2428,N_26682,N_26924);
nand UO_2429 (O_2429,N_26939,N_28521);
nor UO_2430 (O_2430,N_27610,N_28176);
and UO_2431 (O_2431,N_29240,N_27947);
xor UO_2432 (O_2432,N_27822,N_26712);
xnor UO_2433 (O_2433,N_25218,N_25800);
and UO_2434 (O_2434,N_29783,N_27535);
xnor UO_2435 (O_2435,N_27882,N_29989);
or UO_2436 (O_2436,N_29855,N_27760);
or UO_2437 (O_2437,N_28538,N_29480);
and UO_2438 (O_2438,N_28469,N_28241);
or UO_2439 (O_2439,N_25035,N_25539);
xnor UO_2440 (O_2440,N_29246,N_29613);
nor UO_2441 (O_2441,N_29486,N_29731);
nor UO_2442 (O_2442,N_28076,N_29258);
xnor UO_2443 (O_2443,N_28917,N_26119);
xnor UO_2444 (O_2444,N_28688,N_28797);
xnor UO_2445 (O_2445,N_26123,N_29669);
and UO_2446 (O_2446,N_25083,N_29479);
nor UO_2447 (O_2447,N_26005,N_29330);
and UO_2448 (O_2448,N_25005,N_26413);
and UO_2449 (O_2449,N_29316,N_28344);
nand UO_2450 (O_2450,N_25048,N_27258);
and UO_2451 (O_2451,N_25411,N_25398);
and UO_2452 (O_2452,N_28609,N_27320);
nor UO_2453 (O_2453,N_25890,N_26857);
or UO_2454 (O_2454,N_28048,N_27041);
nand UO_2455 (O_2455,N_27853,N_25184);
xor UO_2456 (O_2456,N_26379,N_25578);
nor UO_2457 (O_2457,N_27965,N_25174);
or UO_2458 (O_2458,N_29420,N_25391);
nand UO_2459 (O_2459,N_29864,N_26013);
or UO_2460 (O_2460,N_25258,N_28971);
nor UO_2461 (O_2461,N_29880,N_27165);
or UO_2462 (O_2462,N_28129,N_25824);
and UO_2463 (O_2463,N_27582,N_26971);
nand UO_2464 (O_2464,N_28119,N_26172);
and UO_2465 (O_2465,N_26564,N_27432);
nand UO_2466 (O_2466,N_28747,N_28412);
or UO_2467 (O_2467,N_27598,N_27682);
and UO_2468 (O_2468,N_25911,N_26641);
xnor UO_2469 (O_2469,N_25222,N_25430);
or UO_2470 (O_2470,N_26229,N_26130);
nand UO_2471 (O_2471,N_26209,N_25737);
nor UO_2472 (O_2472,N_28122,N_28424);
nand UO_2473 (O_2473,N_29214,N_26911);
nand UO_2474 (O_2474,N_27886,N_28934);
and UO_2475 (O_2475,N_26188,N_27072);
or UO_2476 (O_2476,N_28423,N_27974);
nand UO_2477 (O_2477,N_29621,N_26829);
nand UO_2478 (O_2478,N_26736,N_29429);
nor UO_2479 (O_2479,N_27204,N_27186);
nand UO_2480 (O_2480,N_27536,N_26031);
xnor UO_2481 (O_2481,N_26571,N_29402);
nand UO_2482 (O_2482,N_27441,N_26304);
nand UO_2483 (O_2483,N_25616,N_25813);
nand UO_2484 (O_2484,N_28601,N_26758);
nor UO_2485 (O_2485,N_28518,N_29394);
xnor UO_2486 (O_2486,N_25494,N_26222);
and UO_2487 (O_2487,N_26741,N_29519);
and UO_2488 (O_2488,N_29294,N_25599);
nand UO_2489 (O_2489,N_29691,N_27187);
xor UO_2490 (O_2490,N_27353,N_26825);
or UO_2491 (O_2491,N_28264,N_29562);
or UO_2492 (O_2492,N_27334,N_25268);
xor UO_2493 (O_2493,N_27569,N_26615);
nor UO_2494 (O_2494,N_25099,N_26011);
and UO_2495 (O_2495,N_27845,N_26105);
xnor UO_2496 (O_2496,N_26183,N_25130);
or UO_2497 (O_2497,N_26840,N_26479);
or UO_2498 (O_2498,N_25051,N_29153);
nor UO_2499 (O_2499,N_27575,N_25990);
nand UO_2500 (O_2500,N_29385,N_28790);
or UO_2501 (O_2501,N_27228,N_25629);
and UO_2502 (O_2502,N_26747,N_25441);
nor UO_2503 (O_2503,N_27060,N_25837);
nor UO_2504 (O_2504,N_28020,N_29230);
xnor UO_2505 (O_2505,N_28718,N_28653);
or UO_2506 (O_2506,N_28967,N_29891);
nor UO_2507 (O_2507,N_28424,N_28441);
nor UO_2508 (O_2508,N_26702,N_26963);
nor UO_2509 (O_2509,N_25556,N_28321);
and UO_2510 (O_2510,N_29717,N_28343);
or UO_2511 (O_2511,N_27026,N_26017);
or UO_2512 (O_2512,N_28546,N_25046);
xnor UO_2513 (O_2513,N_25399,N_26313);
nand UO_2514 (O_2514,N_27637,N_27427);
or UO_2515 (O_2515,N_26076,N_29022);
or UO_2516 (O_2516,N_28390,N_28420);
nor UO_2517 (O_2517,N_25875,N_29420);
or UO_2518 (O_2518,N_25988,N_26346);
nor UO_2519 (O_2519,N_28205,N_26621);
nand UO_2520 (O_2520,N_26068,N_28118);
xnor UO_2521 (O_2521,N_25825,N_26349);
nor UO_2522 (O_2522,N_28732,N_26350);
nor UO_2523 (O_2523,N_26901,N_25671);
xor UO_2524 (O_2524,N_26129,N_29790);
nor UO_2525 (O_2525,N_29157,N_27864);
nor UO_2526 (O_2526,N_29492,N_26358);
nor UO_2527 (O_2527,N_29453,N_26063);
and UO_2528 (O_2528,N_26169,N_26182);
or UO_2529 (O_2529,N_29280,N_26240);
xnor UO_2530 (O_2530,N_27249,N_28394);
nor UO_2531 (O_2531,N_29935,N_27866);
nand UO_2532 (O_2532,N_28341,N_27369);
xor UO_2533 (O_2533,N_26591,N_29432);
or UO_2534 (O_2534,N_29608,N_29667);
nor UO_2535 (O_2535,N_26097,N_26931);
nor UO_2536 (O_2536,N_28726,N_25166);
nand UO_2537 (O_2537,N_29318,N_26252);
nand UO_2538 (O_2538,N_28751,N_25436);
nor UO_2539 (O_2539,N_28155,N_27801);
and UO_2540 (O_2540,N_25466,N_27603);
xor UO_2541 (O_2541,N_27616,N_28540);
nor UO_2542 (O_2542,N_26648,N_29475);
or UO_2543 (O_2543,N_28559,N_29921);
or UO_2544 (O_2544,N_29406,N_26442);
nor UO_2545 (O_2545,N_27851,N_29083);
nand UO_2546 (O_2546,N_29871,N_26156);
and UO_2547 (O_2547,N_26903,N_26784);
xor UO_2548 (O_2548,N_27183,N_29488);
or UO_2549 (O_2549,N_28586,N_25638);
and UO_2550 (O_2550,N_27440,N_28711);
nor UO_2551 (O_2551,N_27111,N_29837);
nand UO_2552 (O_2552,N_26071,N_25478);
xnor UO_2553 (O_2553,N_28871,N_26503);
nor UO_2554 (O_2554,N_26600,N_25291);
and UO_2555 (O_2555,N_27593,N_25912);
or UO_2556 (O_2556,N_29033,N_28473);
xnor UO_2557 (O_2557,N_28150,N_25553);
nor UO_2558 (O_2558,N_27045,N_26446);
nor UO_2559 (O_2559,N_25945,N_25748);
xnor UO_2560 (O_2560,N_26893,N_25777);
nand UO_2561 (O_2561,N_29389,N_25076);
and UO_2562 (O_2562,N_26676,N_29755);
nand UO_2563 (O_2563,N_26279,N_25676);
and UO_2564 (O_2564,N_25116,N_25363);
or UO_2565 (O_2565,N_26816,N_27621);
or UO_2566 (O_2566,N_26781,N_28047);
nor UO_2567 (O_2567,N_25221,N_25450);
xnor UO_2568 (O_2568,N_28188,N_29146);
xnor UO_2569 (O_2569,N_26637,N_28644);
nor UO_2570 (O_2570,N_26803,N_28746);
xor UO_2571 (O_2571,N_25409,N_28140);
nor UO_2572 (O_2572,N_28238,N_28680);
and UO_2573 (O_2573,N_28985,N_28572);
xor UO_2574 (O_2574,N_25714,N_27698);
or UO_2575 (O_2575,N_29725,N_29924);
and UO_2576 (O_2576,N_26758,N_27274);
xor UO_2577 (O_2577,N_29808,N_28415);
or UO_2578 (O_2578,N_28647,N_26882);
or UO_2579 (O_2579,N_25020,N_25494);
or UO_2580 (O_2580,N_27990,N_26787);
xor UO_2581 (O_2581,N_25223,N_28139);
xnor UO_2582 (O_2582,N_27708,N_26578);
nor UO_2583 (O_2583,N_25084,N_27661);
xnor UO_2584 (O_2584,N_29906,N_29466);
nor UO_2585 (O_2585,N_25600,N_26240);
nand UO_2586 (O_2586,N_29595,N_29979);
nand UO_2587 (O_2587,N_28676,N_29228);
xor UO_2588 (O_2588,N_29873,N_25771);
nor UO_2589 (O_2589,N_28885,N_25272);
nor UO_2590 (O_2590,N_25462,N_26489);
nand UO_2591 (O_2591,N_29865,N_25190);
nand UO_2592 (O_2592,N_29739,N_27883);
xnor UO_2593 (O_2593,N_25290,N_27199);
nand UO_2594 (O_2594,N_28986,N_28462);
or UO_2595 (O_2595,N_25103,N_28015);
or UO_2596 (O_2596,N_25761,N_25128);
nand UO_2597 (O_2597,N_29559,N_28387);
nor UO_2598 (O_2598,N_25369,N_29218);
or UO_2599 (O_2599,N_27152,N_25348);
nand UO_2600 (O_2600,N_29443,N_26144);
nor UO_2601 (O_2601,N_27331,N_27136);
nor UO_2602 (O_2602,N_29775,N_29356);
and UO_2603 (O_2603,N_25781,N_25921);
xnor UO_2604 (O_2604,N_28123,N_26945);
nand UO_2605 (O_2605,N_27833,N_27691);
nand UO_2606 (O_2606,N_28279,N_26008);
xor UO_2607 (O_2607,N_25884,N_27125);
xnor UO_2608 (O_2608,N_26824,N_25566);
xor UO_2609 (O_2609,N_26682,N_28978);
and UO_2610 (O_2610,N_26477,N_28487);
xnor UO_2611 (O_2611,N_28329,N_28932);
nand UO_2612 (O_2612,N_26199,N_27834);
xor UO_2613 (O_2613,N_26728,N_25058);
and UO_2614 (O_2614,N_25639,N_25626);
xor UO_2615 (O_2615,N_26930,N_29752);
nand UO_2616 (O_2616,N_27322,N_25008);
and UO_2617 (O_2617,N_29046,N_29762);
and UO_2618 (O_2618,N_25903,N_28444);
or UO_2619 (O_2619,N_29498,N_25731);
nand UO_2620 (O_2620,N_26829,N_29403);
xnor UO_2621 (O_2621,N_26628,N_27446);
or UO_2622 (O_2622,N_25722,N_29103);
nor UO_2623 (O_2623,N_29383,N_25547);
xnor UO_2624 (O_2624,N_29550,N_29632);
nand UO_2625 (O_2625,N_26456,N_25031);
or UO_2626 (O_2626,N_29023,N_25634);
nor UO_2627 (O_2627,N_27159,N_28038);
or UO_2628 (O_2628,N_27959,N_28171);
nor UO_2629 (O_2629,N_26011,N_25392);
xor UO_2630 (O_2630,N_28720,N_29103);
nor UO_2631 (O_2631,N_25907,N_29355);
or UO_2632 (O_2632,N_27211,N_25032);
or UO_2633 (O_2633,N_27269,N_29299);
or UO_2634 (O_2634,N_29717,N_26505);
or UO_2635 (O_2635,N_25800,N_25851);
nand UO_2636 (O_2636,N_29710,N_29807);
and UO_2637 (O_2637,N_25368,N_26220);
xnor UO_2638 (O_2638,N_25017,N_29817);
nand UO_2639 (O_2639,N_25055,N_28512);
nand UO_2640 (O_2640,N_26924,N_26099);
xnor UO_2641 (O_2641,N_26747,N_28989);
and UO_2642 (O_2642,N_28849,N_27678);
nand UO_2643 (O_2643,N_28663,N_26781);
nor UO_2644 (O_2644,N_28069,N_26510);
nor UO_2645 (O_2645,N_27874,N_29001);
xnor UO_2646 (O_2646,N_26259,N_26646);
nor UO_2647 (O_2647,N_28938,N_29860);
xor UO_2648 (O_2648,N_25634,N_29551);
and UO_2649 (O_2649,N_28771,N_29252);
or UO_2650 (O_2650,N_28464,N_25842);
xnor UO_2651 (O_2651,N_28108,N_29488);
nor UO_2652 (O_2652,N_27597,N_26205);
nand UO_2653 (O_2653,N_28308,N_29775);
xor UO_2654 (O_2654,N_28751,N_26544);
nor UO_2655 (O_2655,N_25549,N_27521);
xnor UO_2656 (O_2656,N_25121,N_26301);
or UO_2657 (O_2657,N_25212,N_25334);
xnor UO_2658 (O_2658,N_28492,N_28427);
xnor UO_2659 (O_2659,N_27918,N_28272);
and UO_2660 (O_2660,N_29165,N_25492);
and UO_2661 (O_2661,N_25759,N_28979);
nand UO_2662 (O_2662,N_29402,N_27598);
nor UO_2663 (O_2663,N_26012,N_28468);
nor UO_2664 (O_2664,N_26846,N_26050);
nand UO_2665 (O_2665,N_27520,N_28346);
xnor UO_2666 (O_2666,N_29304,N_28919);
and UO_2667 (O_2667,N_25230,N_26224);
or UO_2668 (O_2668,N_29184,N_28092);
nand UO_2669 (O_2669,N_25245,N_27422);
nor UO_2670 (O_2670,N_28081,N_29446);
xor UO_2671 (O_2671,N_26776,N_29797);
or UO_2672 (O_2672,N_25671,N_25323);
nand UO_2673 (O_2673,N_29064,N_29678);
and UO_2674 (O_2674,N_25229,N_29778);
and UO_2675 (O_2675,N_29959,N_28338);
nand UO_2676 (O_2676,N_28686,N_29470);
or UO_2677 (O_2677,N_26532,N_25969);
xnor UO_2678 (O_2678,N_27706,N_25279);
or UO_2679 (O_2679,N_28034,N_26356);
or UO_2680 (O_2680,N_25105,N_26031);
nand UO_2681 (O_2681,N_25825,N_27039);
and UO_2682 (O_2682,N_27044,N_26414);
xor UO_2683 (O_2683,N_29236,N_26484);
nor UO_2684 (O_2684,N_28740,N_29472);
or UO_2685 (O_2685,N_28099,N_26829);
nand UO_2686 (O_2686,N_29559,N_26322);
xnor UO_2687 (O_2687,N_27578,N_28560);
xor UO_2688 (O_2688,N_27078,N_28648);
nor UO_2689 (O_2689,N_25771,N_28531);
nand UO_2690 (O_2690,N_25442,N_26225);
nand UO_2691 (O_2691,N_26650,N_27190);
nor UO_2692 (O_2692,N_29616,N_29447);
or UO_2693 (O_2693,N_27242,N_29335);
xor UO_2694 (O_2694,N_25611,N_28197);
and UO_2695 (O_2695,N_29957,N_25856);
xor UO_2696 (O_2696,N_28996,N_29369);
and UO_2697 (O_2697,N_26062,N_29831);
and UO_2698 (O_2698,N_28896,N_29682);
and UO_2699 (O_2699,N_25806,N_26337);
nor UO_2700 (O_2700,N_28969,N_28990);
and UO_2701 (O_2701,N_28570,N_27386);
nor UO_2702 (O_2702,N_28677,N_29584);
xor UO_2703 (O_2703,N_27030,N_28812);
nor UO_2704 (O_2704,N_29344,N_25701);
xnor UO_2705 (O_2705,N_28847,N_27470);
nor UO_2706 (O_2706,N_26692,N_28784);
xor UO_2707 (O_2707,N_26769,N_28139);
and UO_2708 (O_2708,N_26393,N_29907);
nor UO_2709 (O_2709,N_29514,N_26726);
nor UO_2710 (O_2710,N_28939,N_26225);
and UO_2711 (O_2711,N_28507,N_25954);
nand UO_2712 (O_2712,N_29425,N_27209);
xnor UO_2713 (O_2713,N_29118,N_26438);
nand UO_2714 (O_2714,N_28596,N_27288);
or UO_2715 (O_2715,N_27191,N_28303);
or UO_2716 (O_2716,N_29661,N_28400);
and UO_2717 (O_2717,N_27325,N_29396);
or UO_2718 (O_2718,N_29226,N_27230);
or UO_2719 (O_2719,N_26626,N_29073);
or UO_2720 (O_2720,N_25277,N_26302);
or UO_2721 (O_2721,N_27088,N_28762);
nor UO_2722 (O_2722,N_26725,N_29565);
or UO_2723 (O_2723,N_26617,N_28786);
and UO_2724 (O_2724,N_25524,N_29959);
nand UO_2725 (O_2725,N_25681,N_29174);
nor UO_2726 (O_2726,N_27791,N_27749);
or UO_2727 (O_2727,N_29754,N_26250);
nor UO_2728 (O_2728,N_26367,N_27107);
nand UO_2729 (O_2729,N_27057,N_26436);
or UO_2730 (O_2730,N_28845,N_27910);
and UO_2731 (O_2731,N_25107,N_29093);
nand UO_2732 (O_2732,N_26380,N_27110);
nand UO_2733 (O_2733,N_27589,N_28921);
nor UO_2734 (O_2734,N_29884,N_26369);
xnor UO_2735 (O_2735,N_27017,N_25962);
and UO_2736 (O_2736,N_28211,N_27710);
xor UO_2737 (O_2737,N_27863,N_25067);
xor UO_2738 (O_2738,N_26015,N_26814);
xnor UO_2739 (O_2739,N_29876,N_28896);
nor UO_2740 (O_2740,N_28118,N_29325);
nand UO_2741 (O_2741,N_25404,N_27449);
or UO_2742 (O_2742,N_28517,N_29587);
and UO_2743 (O_2743,N_25048,N_29522);
nor UO_2744 (O_2744,N_28216,N_29887);
nand UO_2745 (O_2745,N_26782,N_26486);
or UO_2746 (O_2746,N_27121,N_27644);
or UO_2747 (O_2747,N_27438,N_28903);
nor UO_2748 (O_2748,N_27319,N_25976);
xnor UO_2749 (O_2749,N_26385,N_28350);
nor UO_2750 (O_2750,N_25803,N_27517);
xor UO_2751 (O_2751,N_28138,N_27757);
nand UO_2752 (O_2752,N_29405,N_27120);
and UO_2753 (O_2753,N_25789,N_28743);
or UO_2754 (O_2754,N_26582,N_26118);
and UO_2755 (O_2755,N_26101,N_25833);
and UO_2756 (O_2756,N_29461,N_26841);
nor UO_2757 (O_2757,N_28922,N_25144);
xnor UO_2758 (O_2758,N_29719,N_25591);
xnor UO_2759 (O_2759,N_27535,N_29919);
or UO_2760 (O_2760,N_27763,N_28633);
or UO_2761 (O_2761,N_29364,N_25407);
nor UO_2762 (O_2762,N_27727,N_29179);
and UO_2763 (O_2763,N_29578,N_29929);
xnor UO_2764 (O_2764,N_26386,N_26056);
nand UO_2765 (O_2765,N_27600,N_28391);
xnor UO_2766 (O_2766,N_25541,N_27335);
xnor UO_2767 (O_2767,N_29304,N_28414);
or UO_2768 (O_2768,N_26438,N_26081);
nand UO_2769 (O_2769,N_26374,N_26851);
nand UO_2770 (O_2770,N_28897,N_29403);
and UO_2771 (O_2771,N_27337,N_25475);
nand UO_2772 (O_2772,N_27245,N_29298);
nor UO_2773 (O_2773,N_28873,N_25782);
nand UO_2774 (O_2774,N_26282,N_29400);
nor UO_2775 (O_2775,N_28905,N_27663);
nand UO_2776 (O_2776,N_25439,N_29323);
nand UO_2777 (O_2777,N_27614,N_26075);
or UO_2778 (O_2778,N_27320,N_29005);
xnor UO_2779 (O_2779,N_26208,N_27811);
and UO_2780 (O_2780,N_25578,N_28540);
nor UO_2781 (O_2781,N_27881,N_27317);
xor UO_2782 (O_2782,N_28641,N_26929);
xnor UO_2783 (O_2783,N_25079,N_29249);
or UO_2784 (O_2784,N_25358,N_27336);
xor UO_2785 (O_2785,N_25716,N_27878);
xor UO_2786 (O_2786,N_29121,N_29290);
nor UO_2787 (O_2787,N_29427,N_28479);
xnor UO_2788 (O_2788,N_28299,N_28240);
xor UO_2789 (O_2789,N_29589,N_28815);
nor UO_2790 (O_2790,N_27866,N_29438);
nand UO_2791 (O_2791,N_28790,N_29750);
nor UO_2792 (O_2792,N_29794,N_28124);
xnor UO_2793 (O_2793,N_25598,N_27059);
or UO_2794 (O_2794,N_25216,N_28782);
and UO_2795 (O_2795,N_29880,N_26652);
or UO_2796 (O_2796,N_27055,N_29600);
or UO_2797 (O_2797,N_29135,N_28459);
and UO_2798 (O_2798,N_29258,N_29155);
nor UO_2799 (O_2799,N_27009,N_27612);
nor UO_2800 (O_2800,N_25299,N_26123);
or UO_2801 (O_2801,N_28382,N_28750);
nand UO_2802 (O_2802,N_29530,N_27990);
and UO_2803 (O_2803,N_26579,N_29142);
and UO_2804 (O_2804,N_25634,N_26175);
xor UO_2805 (O_2805,N_29979,N_27265);
nor UO_2806 (O_2806,N_26452,N_27525);
xor UO_2807 (O_2807,N_26922,N_25789);
xnor UO_2808 (O_2808,N_29766,N_26849);
or UO_2809 (O_2809,N_29571,N_26864);
and UO_2810 (O_2810,N_25225,N_25090);
nor UO_2811 (O_2811,N_25262,N_28539);
or UO_2812 (O_2812,N_27684,N_28388);
or UO_2813 (O_2813,N_28860,N_29347);
or UO_2814 (O_2814,N_25756,N_26291);
or UO_2815 (O_2815,N_28068,N_26247);
and UO_2816 (O_2816,N_27588,N_27237);
and UO_2817 (O_2817,N_28748,N_29449);
xor UO_2818 (O_2818,N_27179,N_29397);
or UO_2819 (O_2819,N_26543,N_29057);
nor UO_2820 (O_2820,N_25192,N_26904);
nor UO_2821 (O_2821,N_25600,N_25241);
or UO_2822 (O_2822,N_27828,N_27795);
nor UO_2823 (O_2823,N_28760,N_26314);
xnor UO_2824 (O_2824,N_27025,N_29211);
nor UO_2825 (O_2825,N_29271,N_28911);
xor UO_2826 (O_2826,N_28042,N_26164);
or UO_2827 (O_2827,N_27901,N_28535);
xnor UO_2828 (O_2828,N_29382,N_29727);
nand UO_2829 (O_2829,N_27104,N_29660);
or UO_2830 (O_2830,N_25972,N_29015);
xnor UO_2831 (O_2831,N_29710,N_26519);
xnor UO_2832 (O_2832,N_29620,N_26996);
nand UO_2833 (O_2833,N_29694,N_28371);
and UO_2834 (O_2834,N_29526,N_25585);
or UO_2835 (O_2835,N_25121,N_26430);
nand UO_2836 (O_2836,N_26962,N_26708);
nand UO_2837 (O_2837,N_28454,N_26233);
and UO_2838 (O_2838,N_27953,N_27832);
nand UO_2839 (O_2839,N_28967,N_28597);
xnor UO_2840 (O_2840,N_29092,N_26616);
and UO_2841 (O_2841,N_25603,N_29627);
or UO_2842 (O_2842,N_26242,N_28950);
nand UO_2843 (O_2843,N_27437,N_25096);
nand UO_2844 (O_2844,N_29336,N_25857);
xnor UO_2845 (O_2845,N_28392,N_28550);
or UO_2846 (O_2846,N_28678,N_28279);
nand UO_2847 (O_2847,N_28238,N_29484);
and UO_2848 (O_2848,N_28014,N_25056);
nor UO_2849 (O_2849,N_25895,N_27184);
or UO_2850 (O_2850,N_28696,N_28048);
and UO_2851 (O_2851,N_26073,N_27474);
xnor UO_2852 (O_2852,N_26101,N_27710);
or UO_2853 (O_2853,N_25282,N_27909);
nand UO_2854 (O_2854,N_27545,N_25307);
xnor UO_2855 (O_2855,N_26188,N_26562);
nor UO_2856 (O_2856,N_26092,N_29584);
xnor UO_2857 (O_2857,N_27859,N_26927);
nor UO_2858 (O_2858,N_26140,N_27600);
xnor UO_2859 (O_2859,N_26089,N_29743);
or UO_2860 (O_2860,N_26996,N_26351);
and UO_2861 (O_2861,N_25898,N_26403);
nand UO_2862 (O_2862,N_26545,N_28235);
nor UO_2863 (O_2863,N_28673,N_26254);
and UO_2864 (O_2864,N_27724,N_25582);
nand UO_2865 (O_2865,N_29986,N_25634);
and UO_2866 (O_2866,N_26328,N_25430);
xnor UO_2867 (O_2867,N_25030,N_29006);
nor UO_2868 (O_2868,N_27913,N_28749);
nand UO_2869 (O_2869,N_25673,N_25622);
or UO_2870 (O_2870,N_26761,N_25857);
nand UO_2871 (O_2871,N_27873,N_27342);
nor UO_2872 (O_2872,N_28547,N_29877);
or UO_2873 (O_2873,N_26903,N_26914);
or UO_2874 (O_2874,N_26253,N_25793);
xor UO_2875 (O_2875,N_29680,N_28337);
nand UO_2876 (O_2876,N_26376,N_25998);
xor UO_2877 (O_2877,N_28122,N_28603);
nand UO_2878 (O_2878,N_26186,N_28749);
nor UO_2879 (O_2879,N_29200,N_27293);
and UO_2880 (O_2880,N_26739,N_25227);
xor UO_2881 (O_2881,N_25243,N_26064);
nor UO_2882 (O_2882,N_29633,N_28518);
nand UO_2883 (O_2883,N_25621,N_27666);
xnor UO_2884 (O_2884,N_26805,N_25546);
or UO_2885 (O_2885,N_26024,N_29943);
and UO_2886 (O_2886,N_29864,N_28071);
or UO_2887 (O_2887,N_27444,N_25149);
nand UO_2888 (O_2888,N_27288,N_26420);
nand UO_2889 (O_2889,N_26264,N_28725);
or UO_2890 (O_2890,N_25220,N_29435);
or UO_2891 (O_2891,N_27026,N_28830);
or UO_2892 (O_2892,N_28698,N_25304);
or UO_2893 (O_2893,N_29564,N_29151);
nor UO_2894 (O_2894,N_28937,N_29461);
nand UO_2895 (O_2895,N_25385,N_26897);
nor UO_2896 (O_2896,N_27493,N_29305);
xor UO_2897 (O_2897,N_25755,N_28571);
nand UO_2898 (O_2898,N_27407,N_28178);
and UO_2899 (O_2899,N_29870,N_25412);
xor UO_2900 (O_2900,N_27244,N_27803);
xnor UO_2901 (O_2901,N_29431,N_28018);
nor UO_2902 (O_2902,N_27613,N_29190);
nor UO_2903 (O_2903,N_27063,N_25082);
and UO_2904 (O_2904,N_28669,N_27903);
and UO_2905 (O_2905,N_27396,N_29843);
nor UO_2906 (O_2906,N_29561,N_28189);
and UO_2907 (O_2907,N_25153,N_25572);
and UO_2908 (O_2908,N_27126,N_28381);
and UO_2909 (O_2909,N_27879,N_25918);
or UO_2910 (O_2910,N_29976,N_29056);
nand UO_2911 (O_2911,N_28895,N_25582);
nand UO_2912 (O_2912,N_29145,N_25197);
or UO_2913 (O_2913,N_26159,N_25825);
nor UO_2914 (O_2914,N_26296,N_26492);
and UO_2915 (O_2915,N_26331,N_28032);
nor UO_2916 (O_2916,N_26760,N_25775);
nand UO_2917 (O_2917,N_25881,N_25158);
or UO_2918 (O_2918,N_27325,N_29392);
or UO_2919 (O_2919,N_28440,N_27160);
nand UO_2920 (O_2920,N_29322,N_25636);
nand UO_2921 (O_2921,N_29744,N_25134);
nand UO_2922 (O_2922,N_27853,N_25220);
or UO_2923 (O_2923,N_29805,N_27544);
xnor UO_2924 (O_2924,N_26941,N_28437);
xor UO_2925 (O_2925,N_25881,N_26310);
xnor UO_2926 (O_2926,N_28454,N_28308);
or UO_2927 (O_2927,N_25210,N_25750);
xor UO_2928 (O_2928,N_25397,N_28380);
and UO_2929 (O_2929,N_27437,N_28052);
xor UO_2930 (O_2930,N_26652,N_26001);
or UO_2931 (O_2931,N_29366,N_27079);
nand UO_2932 (O_2932,N_28670,N_27185);
and UO_2933 (O_2933,N_29188,N_28992);
xnor UO_2934 (O_2934,N_29535,N_29825);
or UO_2935 (O_2935,N_27012,N_25251);
and UO_2936 (O_2936,N_29187,N_25263);
and UO_2937 (O_2937,N_29209,N_27892);
xnor UO_2938 (O_2938,N_25393,N_27638);
xnor UO_2939 (O_2939,N_27323,N_25746);
nand UO_2940 (O_2940,N_25312,N_27505);
or UO_2941 (O_2941,N_27042,N_25756);
or UO_2942 (O_2942,N_25472,N_29009);
xnor UO_2943 (O_2943,N_28390,N_28492);
or UO_2944 (O_2944,N_29533,N_25834);
nand UO_2945 (O_2945,N_27682,N_29112);
and UO_2946 (O_2946,N_25751,N_29867);
nand UO_2947 (O_2947,N_27334,N_29668);
xor UO_2948 (O_2948,N_28549,N_26778);
nor UO_2949 (O_2949,N_26038,N_28448);
nor UO_2950 (O_2950,N_27167,N_25134);
or UO_2951 (O_2951,N_25085,N_25459);
xor UO_2952 (O_2952,N_28728,N_27654);
and UO_2953 (O_2953,N_29245,N_28307);
and UO_2954 (O_2954,N_28518,N_28831);
nand UO_2955 (O_2955,N_25402,N_26415);
xor UO_2956 (O_2956,N_28413,N_26058);
and UO_2957 (O_2957,N_28286,N_26344);
xor UO_2958 (O_2958,N_28296,N_29446);
and UO_2959 (O_2959,N_25631,N_26470);
xor UO_2960 (O_2960,N_28950,N_29611);
and UO_2961 (O_2961,N_28502,N_25433);
or UO_2962 (O_2962,N_25112,N_27608);
or UO_2963 (O_2963,N_29368,N_25396);
and UO_2964 (O_2964,N_29571,N_29023);
nand UO_2965 (O_2965,N_27784,N_27501);
or UO_2966 (O_2966,N_26940,N_26675);
and UO_2967 (O_2967,N_27276,N_28621);
and UO_2968 (O_2968,N_27231,N_28637);
nand UO_2969 (O_2969,N_27296,N_28971);
nand UO_2970 (O_2970,N_28655,N_25160);
or UO_2971 (O_2971,N_29757,N_28903);
nor UO_2972 (O_2972,N_28056,N_27485);
xnor UO_2973 (O_2973,N_27016,N_28112);
or UO_2974 (O_2974,N_29946,N_25569);
nand UO_2975 (O_2975,N_29002,N_29024);
or UO_2976 (O_2976,N_25584,N_26562);
or UO_2977 (O_2977,N_29239,N_27138);
nor UO_2978 (O_2978,N_29415,N_26672);
xnor UO_2979 (O_2979,N_28336,N_25888);
nor UO_2980 (O_2980,N_25883,N_25060);
xor UO_2981 (O_2981,N_29262,N_29003);
nor UO_2982 (O_2982,N_25993,N_29645);
xnor UO_2983 (O_2983,N_28644,N_28167);
nand UO_2984 (O_2984,N_26458,N_25399);
or UO_2985 (O_2985,N_29745,N_28654);
nand UO_2986 (O_2986,N_25618,N_28799);
or UO_2987 (O_2987,N_25768,N_27430);
xor UO_2988 (O_2988,N_27082,N_26184);
nor UO_2989 (O_2989,N_27975,N_26816);
or UO_2990 (O_2990,N_27646,N_26424);
nor UO_2991 (O_2991,N_28623,N_26625);
and UO_2992 (O_2992,N_29193,N_29291);
nand UO_2993 (O_2993,N_25546,N_28048);
xnor UO_2994 (O_2994,N_26566,N_26591);
and UO_2995 (O_2995,N_28982,N_25065);
xnor UO_2996 (O_2996,N_25308,N_29516);
xnor UO_2997 (O_2997,N_26329,N_27320);
nand UO_2998 (O_2998,N_26588,N_29201);
or UO_2999 (O_2999,N_25373,N_29775);
xnor UO_3000 (O_3000,N_27026,N_25339);
xor UO_3001 (O_3001,N_29467,N_26509);
or UO_3002 (O_3002,N_28197,N_26642);
or UO_3003 (O_3003,N_25124,N_25662);
and UO_3004 (O_3004,N_28043,N_29602);
nand UO_3005 (O_3005,N_27743,N_26210);
and UO_3006 (O_3006,N_27785,N_25605);
nand UO_3007 (O_3007,N_25189,N_29721);
nand UO_3008 (O_3008,N_29860,N_27761);
xnor UO_3009 (O_3009,N_29937,N_27253);
xnor UO_3010 (O_3010,N_25252,N_25199);
and UO_3011 (O_3011,N_28534,N_26543);
xnor UO_3012 (O_3012,N_27676,N_28490);
or UO_3013 (O_3013,N_28233,N_25183);
xnor UO_3014 (O_3014,N_28843,N_29307);
and UO_3015 (O_3015,N_28214,N_29938);
or UO_3016 (O_3016,N_25991,N_28676);
or UO_3017 (O_3017,N_28114,N_28780);
or UO_3018 (O_3018,N_26776,N_27155);
xor UO_3019 (O_3019,N_28350,N_27364);
nor UO_3020 (O_3020,N_26253,N_28732);
xnor UO_3021 (O_3021,N_29983,N_28569);
and UO_3022 (O_3022,N_27853,N_25961);
nor UO_3023 (O_3023,N_25497,N_25581);
nand UO_3024 (O_3024,N_25240,N_28815);
nand UO_3025 (O_3025,N_27975,N_26890);
xor UO_3026 (O_3026,N_29742,N_28497);
xnor UO_3027 (O_3027,N_26032,N_25277);
xor UO_3028 (O_3028,N_29274,N_25865);
and UO_3029 (O_3029,N_29537,N_28753);
and UO_3030 (O_3030,N_25460,N_28898);
nand UO_3031 (O_3031,N_28064,N_27504);
xnor UO_3032 (O_3032,N_26134,N_27274);
nor UO_3033 (O_3033,N_26438,N_28298);
or UO_3034 (O_3034,N_25433,N_26929);
or UO_3035 (O_3035,N_25720,N_29948);
and UO_3036 (O_3036,N_26023,N_28668);
and UO_3037 (O_3037,N_27612,N_28221);
nor UO_3038 (O_3038,N_29670,N_27549);
or UO_3039 (O_3039,N_28042,N_29343);
xnor UO_3040 (O_3040,N_26115,N_27891);
and UO_3041 (O_3041,N_29097,N_25683);
and UO_3042 (O_3042,N_29717,N_25606);
nand UO_3043 (O_3043,N_27577,N_28790);
nor UO_3044 (O_3044,N_26056,N_27432);
xor UO_3045 (O_3045,N_27610,N_27854);
nor UO_3046 (O_3046,N_29260,N_29291);
and UO_3047 (O_3047,N_27871,N_27855);
nor UO_3048 (O_3048,N_29978,N_25054);
nor UO_3049 (O_3049,N_27328,N_25643);
xnor UO_3050 (O_3050,N_25437,N_29231);
or UO_3051 (O_3051,N_29127,N_26539);
nor UO_3052 (O_3052,N_27606,N_29578);
and UO_3053 (O_3053,N_27179,N_27838);
nor UO_3054 (O_3054,N_28879,N_28208);
nor UO_3055 (O_3055,N_29924,N_27444);
xor UO_3056 (O_3056,N_27901,N_25014);
nor UO_3057 (O_3057,N_25867,N_28594);
nand UO_3058 (O_3058,N_27179,N_27976);
nand UO_3059 (O_3059,N_25663,N_26255);
or UO_3060 (O_3060,N_29816,N_27467);
and UO_3061 (O_3061,N_29010,N_27864);
or UO_3062 (O_3062,N_26959,N_25427);
nand UO_3063 (O_3063,N_26275,N_29479);
nor UO_3064 (O_3064,N_27304,N_25222);
or UO_3065 (O_3065,N_25690,N_27286);
or UO_3066 (O_3066,N_27320,N_25328);
nand UO_3067 (O_3067,N_27616,N_29964);
xor UO_3068 (O_3068,N_29536,N_25532);
nand UO_3069 (O_3069,N_26514,N_29328);
nand UO_3070 (O_3070,N_29767,N_25247);
xnor UO_3071 (O_3071,N_28259,N_27466);
nand UO_3072 (O_3072,N_28999,N_29033);
or UO_3073 (O_3073,N_27998,N_25867);
nor UO_3074 (O_3074,N_27303,N_29903);
nor UO_3075 (O_3075,N_28454,N_29750);
xor UO_3076 (O_3076,N_29907,N_25223);
or UO_3077 (O_3077,N_26147,N_26273);
xor UO_3078 (O_3078,N_26603,N_26321);
or UO_3079 (O_3079,N_28099,N_25227);
xnor UO_3080 (O_3080,N_25562,N_28680);
xnor UO_3081 (O_3081,N_29921,N_28641);
xor UO_3082 (O_3082,N_25617,N_27068);
nand UO_3083 (O_3083,N_28097,N_25807);
or UO_3084 (O_3084,N_27214,N_26840);
nor UO_3085 (O_3085,N_28363,N_26317);
and UO_3086 (O_3086,N_25592,N_25910);
and UO_3087 (O_3087,N_28535,N_29572);
or UO_3088 (O_3088,N_26128,N_28852);
or UO_3089 (O_3089,N_26782,N_25462);
nor UO_3090 (O_3090,N_25657,N_26209);
or UO_3091 (O_3091,N_27033,N_29869);
nor UO_3092 (O_3092,N_28185,N_28431);
and UO_3093 (O_3093,N_26543,N_25608);
or UO_3094 (O_3094,N_25270,N_27558);
nand UO_3095 (O_3095,N_25660,N_26555);
nand UO_3096 (O_3096,N_29978,N_26853);
or UO_3097 (O_3097,N_29264,N_29963);
and UO_3098 (O_3098,N_25515,N_25223);
nand UO_3099 (O_3099,N_27899,N_25175);
xnor UO_3100 (O_3100,N_26657,N_25747);
nand UO_3101 (O_3101,N_27094,N_26896);
xor UO_3102 (O_3102,N_25550,N_29504);
or UO_3103 (O_3103,N_29343,N_25371);
or UO_3104 (O_3104,N_28453,N_28115);
nand UO_3105 (O_3105,N_27348,N_27099);
nor UO_3106 (O_3106,N_28656,N_26455);
nand UO_3107 (O_3107,N_28993,N_28228);
xnor UO_3108 (O_3108,N_25714,N_26679);
nor UO_3109 (O_3109,N_26232,N_26903);
or UO_3110 (O_3110,N_28381,N_28063);
and UO_3111 (O_3111,N_27488,N_25107);
nor UO_3112 (O_3112,N_25676,N_25550);
or UO_3113 (O_3113,N_28635,N_25316);
xor UO_3114 (O_3114,N_26674,N_26901);
nand UO_3115 (O_3115,N_25986,N_28138);
nand UO_3116 (O_3116,N_28484,N_25336);
and UO_3117 (O_3117,N_28745,N_27595);
nand UO_3118 (O_3118,N_29590,N_27872);
or UO_3119 (O_3119,N_27149,N_25984);
and UO_3120 (O_3120,N_27468,N_27932);
nor UO_3121 (O_3121,N_28675,N_29403);
nand UO_3122 (O_3122,N_29750,N_27695);
nand UO_3123 (O_3123,N_29344,N_27867);
xor UO_3124 (O_3124,N_27478,N_28011);
or UO_3125 (O_3125,N_27437,N_25760);
or UO_3126 (O_3126,N_26042,N_28533);
nand UO_3127 (O_3127,N_27512,N_25180);
xnor UO_3128 (O_3128,N_28102,N_26771);
and UO_3129 (O_3129,N_29159,N_28498);
and UO_3130 (O_3130,N_28004,N_29675);
xor UO_3131 (O_3131,N_29890,N_26961);
and UO_3132 (O_3132,N_28374,N_25388);
nor UO_3133 (O_3133,N_29779,N_27226);
nand UO_3134 (O_3134,N_28414,N_26646);
or UO_3135 (O_3135,N_26816,N_28359);
or UO_3136 (O_3136,N_26728,N_27214);
and UO_3137 (O_3137,N_27372,N_29172);
nor UO_3138 (O_3138,N_26156,N_26159);
xnor UO_3139 (O_3139,N_26223,N_27470);
or UO_3140 (O_3140,N_27557,N_29609);
or UO_3141 (O_3141,N_28327,N_26278);
xor UO_3142 (O_3142,N_29259,N_25350);
xnor UO_3143 (O_3143,N_26821,N_25549);
xor UO_3144 (O_3144,N_26227,N_27584);
nand UO_3145 (O_3145,N_28408,N_27136);
nand UO_3146 (O_3146,N_26164,N_28115);
xnor UO_3147 (O_3147,N_29093,N_27860);
and UO_3148 (O_3148,N_26631,N_25382);
nand UO_3149 (O_3149,N_28267,N_28055);
nand UO_3150 (O_3150,N_25411,N_29957);
xor UO_3151 (O_3151,N_26666,N_29063);
or UO_3152 (O_3152,N_28022,N_27555);
nand UO_3153 (O_3153,N_29857,N_27030);
or UO_3154 (O_3154,N_29322,N_26405);
nand UO_3155 (O_3155,N_27613,N_26127);
and UO_3156 (O_3156,N_29936,N_28450);
and UO_3157 (O_3157,N_25699,N_28321);
nor UO_3158 (O_3158,N_26490,N_25557);
or UO_3159 (O_3159,N_27030,N_25766);
nand UO_3160 (O_3160,N_25184,N_27201);
or UO_3161 (O_3161,N_27450,N_27977);
nand UO_3162 (O_3162,N_26103,N_28079);
or UO_3163 (O_3163,N_29837,N_29576);
nor UO_3164 (O_3164,N_28583,N_27528);
and UO_3165 (O_3165,N_25854,N_29108);
or UO_3166 (O_3166,N_26118,N_27678);
xor UO_3167 (O_3167,N_27878,N_25560);
nor UO_3168 (O_3168,N_28038,N_28981);
or UO_3169 (O_3169,N_25342,N_26327);
xor UO_3170 (O_3170,N_27249,N_27416);
xnor UO_3171 (O_3171,N_29756,N_28604);
xor UO_3172 (O_3172,N_28561,N_27525);
xor UO_3173 (O_3173,N_25074,N_25458);
nand UO_3174 (O_3174,N_27508,N_28037);
nor UO_3175 (O_3175,N_27549,N_27565);
nand UO_3176 (O_3176,N_28177,N_27275);
nand UO_3177 (O_3177,N_26237,N_28820);
and UO_3178 (O_3178,N_29403,N_28611);
and UO_3179 (O_3179,N_25500,N_27056);
nand UO_3180 (O_3180,N_26578,N_28750);
and UO_3181 (O_3181,N_25421,N_28990);
nand UO_3182 (O_3182,N_26798,N_29441);
nand UO_3183 (O_3183,N_27067,N_26229);
and UO_3184 (O_3184,N_26203,N_29699);
and UO_3185 (O_3185,N_29192,N_26065);
nor UO_3186 (O_3186,N_29172,N_27132);
nor UO_3187 (O_3187,N_29101,N_25747);
xor UO_3188 (O_3188,N_29060,N_26537);
and UO_3189 (O_3189,N_25900,N_27433);
xnor UO_3190 (O_3190,N_25723,N_28685);
and UO_3191 (O_3191,N_28213,N_26379);
xnor UO_3192 (O_3192,N_28235,N_25459);
nand UO_3193 (O_3193,N_27229,N_29274);
or UO_3194 (O_3194,N_29172,N_28335);
nor UO_3195 (O_3195,N_25767,N_28409);
xor UO_3196 (O_3196,N_29052,N_27250);
and UO_3197 (O_3197,N_28076,N_26853);
and UO_3198 (O_3198,N_26565,N_25476);
or UO_3199 (O_3199,N_29325,N_27853);
xnor UO_3200 (O_3200,N_29960,N_27508);
or UO_3201 (O_3201,N_26800,N_28320);
nand UO_3202 (O_3202,N_27005,N_27081);
nand UO_3203 (O_3203,N_29230,N_26322);
nor UO_3204 (O_3204,N_27485,N_27693);
nor UO_3205 (O_3205,N_28409,N_27887);
or UO_3206 (O_3206,N_27873,N_26000);
nand UO_3207 (O_3207,N_28223,N_26194);
and UO_3208 (O_3208,N_28362,N_27778);
or UO_3209 (O_3209,N_29904,N_25167);
nand UO_3210 (O_3210,N_28437,N_27727);
nand UO_3211 (O_3211,N_27243,N_29419);
xor UO_3212 (O_3212,N_26449,N_26864);
xor UO_3213 (O_3213,N_25014,N_25151);
nor UO_3214 (O_3214,N_27812,N_25844);
or UO_3215 (O_3215,N_29747,N_28430);
xnor UO_3216 (O_3216,N_27662,N_28495);
or UO_3217 (O_3217,N_25537,N_28868);
nand UO_3218 (O_3218,N_27016,N_25209);
or UO_3219 (O_3219,N_27780,N_29553);
nand UO_3220 (O_3220,N_25957,N_25937);
xor UO_3221 (O_3221,N_25155,N_26050);
nand UO_3222 (O_3222,N_25668,N_29335);
nor UO_3223 (O_3223,N_25419,N_29986);
nor UO_3224 (O_3224,N_27653,N_27794);
nor UO_3225 (O_3225,N_28127,N_25886);
nor UO_3226 (O_3226,N_29500,N_25695);
and UO_3227 (O_3227,N_29956,N_27744);
or UO_3228 (O_3228,N_29030,N_27694);
nor UO_3229 (O_3229,N_27312,N_27272);
or UO_3230 (O_3230,N_29142,N_25251);
xor UO_3231 (O_3231,N_25063,N_28206);
nand UO_3232 (O_3232,N_29609,N_28702);
or UO_3233 (O_3233,N_28196,N_26896);
or UO_3234 (O_3234,N_29725,N_27451);
or UO_3235 (O_3235,N_28102,N_27908);
or UO_3236 (O_3236,N_28619,N_25862);
nand UO_3237 (O_3237,N_25148,N_25711);
xor UO_3238 (O_3238,N_26852,N_29191);
or UO_3239 (O_3239,N_27277,N_26540);
and UO_3240 (O_3240,N_28820,N_28733);
xor UO_3241 (O_3241,N_27992,N_28442);
or UO_3242 (O_3242,N_28616,N_29599);
xnor UO_3243 (O_3243,N_26796,N_26119);
xor UO_3244 (O_3244,N_25380,N_27103);
nor UO_3245 (O_3245,N_27817,N_28400);
or UO_3246 (O_3246,N_27325,N_29032);
nor UO_3247 (O_3247,N_26709,N_27205);
and UO_3248 (O_3248,N_28244,N_28457);
and UO_3249 (O_3249,N_25610,N_26060);
nor UO_3250 (O_3250,N_28912,N_25321);
and UO_3251 (O_3251,N_27004,N_29320);
and UO_3252 (O_3252,N_29664,N_25439);
or UO_3253 (O_3253,N_29986,N_29698);
xor UO_3254 (O_3254,N_28200,N_28714);
xor UO_3255 (O_3255,N_28390,N_26378);
nor UO_3256 (O_3256,N_28746,N_29229);
and UO_3257 (O_3257,N_25658,N_26528);
or UO_3258 (O_3258,N_27265,N_28989);
or UO_3259 (O_3259,N_27512,N_25708);
xnor UO_3260 (O_3260,N_26802,N_28172);
xnor UO_3261 (O_3261,N_29210,N_25161);
or UO_3262 (O_3262,N_28507,N_27549);
xor UO_3263 (O_3263,N_26919,N_27730);
and UO_3264 (O_3264,N_27443,N_25225);
nand UO_3265 (O_3265,N_26516,N_25227);
and UO_3266 (O_3266,N_29105,N_27895);
or UO_3267 (O_3267,N_28518,N_26031);
nand UO_3268 (O_3268,N_26308,N_27352);
nand UO_3269 (O_3269,N_27384,N_25380);
or UO_3270 (O_3270,N_28844,N_29794);
and UO_3271 (O_3271,N_27467,N_28082);
or UO_3272 (O_3272,N_27263,N_29470);
nor UO_3273 (O_3273,N_25843,N_29215);
nand UO_3274 (O_3274,N_28725,N_25821);
or UO_3275 (O_3275,N_27590,N_25392);
or UO_3276 (O_3276,N_28658,N_27382);
nand UO_3277 (O_3277,N_29391,N_28220);
nor UO_3278 (O_3278,N_28694,N_27671);
nand UO_3279 (O_3279,N_29906,N_25168);
nor UO_3280 (O_3280,N_28634,N_26911);
nor UO_3281 (O_3281,N_27048,N_27421);
or UO_3282 (O_3282,N_26565,N_25796);
and UO_3283 (O_3283,N_28716,N_29591);
and UO_3284 (O_3284,N_26393,N_26446);
or UO_3285 (O_3285,N_29430,N_26555);
xor UO_3286 (O_3286,N_29870,N_28100);
and UO_3287 (O_3287,N_29641,N_26835);
nor UO_3288 (O_3288,N_26843,N_25408);
xor UO_3289 (O_3289,N_27055,N_29318);
or UO_3290 (O_3290,N_29958,N_25736);
nor UO_3291 (O_3291,N_28133,N_25790);
and UO_3292 (O_3292,N_26268,N_27717);
xor UO_3293 (O_3293,N_28752,N_27335);
or UO_3294 (O_3294,N_28669,N_26885);
and UO_3295 (O_3295,N_26895,N_29832);
and UO_3296 (O_3296,N_26066,N_29659);
and UO_3297 (O_3297,N_26251,N_25211);
nand UO_3298 (O_3298,N_29925,N_25399);
and UO_3299 (O_3299,N_28305,N_27631);
nand UO_3300 (O_3300,N_29915,N_28245);
nand UO_3301 (O_3301,N_26180,N_29173);
or UO_3302 (O_3302,N_26919,N_27434);
and UO_3303 (O_3303,N_28804,N_27160);
nor UO_3304 (O_3304,N_27869,N_25652);
nand UO_3305 (O_3305,N_27860,N_26367);
nor UO_3306 (O_3306,N_27275,N_26084);
or UO_3307 (O_3307,N_28036,N_28321);
nand UO_3308 (O_3308,N_28673,N_29813);
xnor UO_3309 (O_3309,N_27813,N_25436);
nor UO_3310 (O_3310,N_26103,N_26264);
and UO_3311 (O_3311,N_28959,N_25884);
or UO_3312 (O_3312,N_29405,N_27160);
xor UO_3313 (O_3313,N_25656,N_25542);
nand UO_3314 (O_3314,N_27113,N_28974);
nor UO_3315 (O_3315,N_29032,N_26020);
and UO_3316 (O_3316,N_28200,N_27362);
and UO_3317 (O_3317,N_29935,N_26438);
and UO_3318 (O_3318,N_28226,N_26751);
nor UO_3319 (O_3319,N_25732,N_25587);
nand UO_3320 (O_3320,N_29520,N_26550);
xor UO_3321 (O_3321,N_27099,N_28812);
and UO_3322 (O_3322,N_26369,N_28323);
xnor UO_3323 (O_3323,N_29628,N_29313);
or UO_3324 (O_3324,N_28017,N_27980);
or UO_3325 (O_3325,N_28591,N_28276);
xor UO_3326 (O_3326,N_29994,N_28792);
xnor UO_3327 (O_3327,N_26508,N_26553);
nand UO_3328 (O_3328,N_26266,N_29196);
or UO_3329 (O_3329,N_28421,N_26643);
xor UO_3330 (O_3330,N_26203,N_26837);
xnor UO_3331 (O_3331,N_28263,N_27004);
nand UO_3332 (O_3332,N_27575,N_29660);
nor UO_3333 (O_3333,N_28378,N_28157);
or UO_3334 (O_3334,N_29636,N_26787);
xor UO_3335 (O_3335,N_25320,N_27303);
nand UO_3336 (O_3336,N_28312,N_26708);
xor UO_3337 (O_3337,N_29868,N_28292);
nor UO_3338 (O_3338,N_29105,N_27767);
nand UO_3339 (O_3339,N_28397,N_25912);
nand UO_3340 (O_3340,N_29548,N_26849);
xor UO_3341 (O_3341,N_29077,N_26156);
nand UO_3342 (O_3342,N_25287,N_29374);
nor UO_3343 (O_3343,N_29167,N_26475);
and UO_3344 (O_3344,N_26325,N_29974);
and UO_3345 (O_3345,N_26089,N_29028);
xor UO_3346 (O_3346,N_28517,N_25517);
nand UO_3347 (O_3347,N_28949,N_26176);
nor UO_3348 (O_3348,N_29487,N_26100);
xor UO_3349 (O_3349,N_25673,N_26197);
and UO_3350 (O_3350,N_29317,N_29565);
and UO_3351 (O_3351,N_25235,N_29905);
or UO_3352 (O_3352,N_26814,N_29066);
and UO_3353 (O_3353,N_28966,N_29165);
and UO_3354 (O_3354,N_29435,N_29542);
and UO_3355 (O_3355,N_29514,N_27743);
nor UO_3356 (O_3356,N_28730,N_28549);
or UO_3357 (O_3357,N_27066,N_26238);
or UO_3358 (O_3358,N_27234,N_28826);
nand UO_3359 (O_3359,N_25824,N_26316);
nor UO_3360 (O_3360,N_26028,N_26563);
nand UO_3361 (O_3361,N_25746,N_29278);
or UO_3362 (O_3362,N_25738,N_29470);
nand UO_3363 (O_3363,N_29304,N_29068);
or UO_3364 (O_3364,N_25462,N_26445);
xor UO_3365 (O_3365,N_29567,N_27298);
nor UO_3366 (O_3366,N_26204,N_25776);
xnor UO_3367 (O_3367,N_27181,N_25660);
and UO_3368 (O_3368,N_28724,N_25643);
and UO_3369 (O_3369,N_26653,N_25845);
nor UO_3370 (O_3370,N_29127,N_28624);
nand UO_3371 (O_3371,N_28436,N_26171);
nand UO_3372 (O_3372,N_28753,N_25165);
nor UO_3373 (O_3373,N_28351,N_25000);
or UO_3374 (O_3374,N_25274,N_26476);
or UO_3375 (O_3375,N_27665,N_26948);
nand UO_3376 (O_3376,N_28799,N_29029);
nand UO_3377 (O_3377,N_27243,N_25791);
and UO_3378 (O_3378,N_26475,N_27402);
or UO_3379 (O_3379,N_26690,N_29298);
and UO_3380 (O_3380,N_28922,N_25236);
nand UO_3381 (O_3381,N_29094,N_29195);
xnor UO_3382 (O_3382,N_25856,N_25401);
and UO_3383 (O_3383,N_25990,N_26385);
nor UO_3384 (O_3384,N_28885,N_25027);
or UO_3385 (O_3385,N_29306,N_26715);
nand UO_3386 (O_3386,N_25754,N_29857);
or UO_3387 (O_3387,N_28030,N_27959);
and UO_3388 (O_3388,N_27447,N_26261);
nand UO_3389 (O_3389,N_28775,N_25762);
and UO_3390 (O_3390,N_26638,N_27948);
nor UO_3391 (O_3391,N_25383,N_28667);
and UO_3392 (O_3392,N_29107,N_25876);
or UO_3393 (O_3393,N_29570,N_28961);
nor UO_3394 (O_3394,N_28086,N_28109);
nand UO_3395 (O_3395,N_29643,N_27265);
xnor UO_3396 (O_3396,N_26482,N_28475);
nor UO_3397 (O_3397,N_28750,N_25289);
and UO_3398 (O_3398,N_28036,N_26221);
or UO_3399 (O_3399,N_27912,N_27657);
and UO_3400 (O_3400,N_27029,N_27558);
xnor UO_3401 (O_3401,N_25925,N_25795);
nand UO_3402 (O_3402,N_25240,N_25909);
or UO_3403 (O_3403,N_28389,N_27710);
or UO_3404 (O_3404,N_27645,N_26242);
nor UO_3405 (O_3405,N_28365,N_25692);
nand UO_3406 (O_3406,N_26782,N_27496);
xor UO_3407 (O_3407,N_28067,N_29225);
or UO_3408 (O_3408,N_28282,N_29607);
xor UO_3409 (O_3409,N_27354,N_28321);
nor UO_3410 (O_3410,N_25197,N_25734);
nor UO_3411 (O_3411,N_26079,N_26898);
nor UO_3412 (O_3412,N_29252,N_29261);
and UO_3413 (O_3413,N_28307,N_26002);
nand UO_3414 (O_3414,N_29665,N_25361);
nand UO_3415 (O_3415,N_26923,N_27986);
or UO_3416 (O_3416,N_28820,N_28544);
nor UO_3417 (O_3417,N_25860,N_28006);
and UO_3418 (O_3418,N_26080,N_29053);
and UO_3419 (O_3419,N_29073,N_26039);
nand UO_3420 (O_3420,N_29298,N_25675);
or UO_3421 (O_3421,N_26635,N_26751);
and UO_3422 (O_3422,N_27332,N_26829);
or UO_3423 (O_3423,N_29922,N_26706);
nand UO_3424 (O_3424,N_26563,N_28200);
xnor UO_3425 (O_3425,N_26093,N_28657);
nor UO_3426 (O_3426,N_27822,N_29364);
nor UO_3427 (O_3427,N_26660,N_28674);
nand UO_3428 (O_3428,N_28739,N_26015);
xnor UO_3429 (O_3429,N_26276,N_28122);
nor UO_3430 (O_3430,N_26202,N_28465);
nand UO_3431 (O_3431,N_29433,N_29441);
xnor UO_3432 (O_3432,N_26314,N_28827);
or UO_3433 (O_3433,N_28512,N_26010);
and UO_3434 (O_3434,N_27117,N_25475);
or UO_3435 (O_3435,N_27304,N_27581);
and UO_3436 (O_3436,N_27134,N_26922);
and UO_3437 (O_3437,N_29590,N_25485);
or UO_3438 (O_3438,N_27698,N_26859);
nor UO_3439 (O_3439,N_29906,N_29350);
xor UO_3440 (O_3440,N_26462,N_28378);
nor UO_3441 (O_3441,N_25078,N_29986);
nand UO_3442 (O_3442,N_29788,N_29913);
or UO_3443 (O_3443,N_29957,N_27951);
nor UO_3444 (O_3444,N_28908,N_26827);
or UO_3445 (O_3445,N_26275,N_25695);
nor UO_3446 (O_3446,N_25611,N_27039);
nor UO_3447 (O_3447,N_29842,N_25469);
nor UO_3448 (O_3448,N_26023,N_26671);
xnor UO_3449 (O_3449,N_26957,N_28406);
and UO_3450 (O_3450,N_28278,N_29554);
xnor UO_3451 (O_3451,N_29980,N_26252);
or UO_3452 (O_3452,N_29525,N_27415);
nor UO_3453 (O_3453,N_26656,N_29168);
and UO_3454 (O_3454,N_28082,N_28772);
and UO_3455 (O_3455,N_26958,N_25744);
nor UO_3456 (O_3456,N_28696,N_26905);
or UO_3457 (O_3457,N_27693,N_26463);
xnor UO_3458 (O_3458,N_26898,N_25267);
nor UO_3459 (O_3459,N_28731,N_29324);
nand UO_3460 (O_3460,N_29157,N_29566);
or UO_3461 (O_3461,N_28814,N_27794);
nand UO_3462 (O_3462,N_28968,N_25416);
or UO_3463 (O_3463,N_25131,N_27781);
nand UO_3464 (O_3464,N_28713,N_27027);
and UO_3465 (O_3465,N_29803,N_26986);
nand UO_3466 (O_3466,N_28204,N_26529);
or UO_3467 (O_3467,N_28982,N_26200);
or UO_3468 (O_3468,N_26362,N_28590);
xnor UO_3469 (O_3469,N_28209,N_28680);
nor UO_3470 (O_3470,N_26377,N_25350);
nor UO_3471 (O_3471,N_28886,N_25115);
or UO_3472 (O_3472,N_29223,N_26777);
and UO_3473 (O_3473,N_29128,N_26460);
and UO_3474 (O_3474,N_26418,N_26511);
and UO_3475 (O_3475,N_29095,N_25848);
or UO_3476 (O_3476,N_25405,N_27334);
nor UO_3477 (O_3477,N_28912,N_27436);
and UO_3478 (O_3478,N_26564,N_29604);
and UO_3479 (O_3479,N_27665,N_25392);
or UO_3480 (O_3480,N_27857,N_28305);
xnor UO_3481 (O_3481,N_25791,N_26629);
and UO_3482 (O_3482,N_26965,N_28401);
nor UO_3483 (O_3483,N_25945,N_25826);
or UO_3484 (O_3484,N_27297,N_29970);
xnor UO_3485 (O_3485,N_28249,N_26882);
nand UO_3486 (O_3486,N_27463,N_28549);
and UO_3487 (O_3487,N_28095,N_29448);
or UO_3488 (O_3488,N_29474,N_27437);
nand UO_3489 (O_3489,N_28179,N_27036);
nor UO_3490 (O_3490,N_29085,N_27121);
nor UO_3491 (O_3491,N_26938,N_29823);
and UO_3492 (O_3492,N_26477,N_29952);
nor UO_3493 (O_3493,N_27047,N_28964);
nor UO_3494 (O_3494,N_26914,N_27317);
or UO_3495 (O_3495,N_29369,N_28648);
nand UO_3496 (O_3496,N_27026,N_26359);
or UO_3497 (O_3497,N_29332,N_27751);
nor UO_3498 (O_3498,N_27666,N_27383);
and UO_3499 (O_3499,N_26829,N_28237);
endmodule