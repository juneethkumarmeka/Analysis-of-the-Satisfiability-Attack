module basic_1500_15000_2000_20_levels_5xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
xor U0 (N_0,In_102,In_1246);
or U1 (N_1,In_266,In_616);
and U2 (N_2,In_1218,In_1138);
nand U3 (N_3,In_762,In_823);
nand U4 (N_4,In_1332,In_600);
and U5 (N_5,In_827,In_481);
and U6 (N_6,In_105,In_1245);
and U7 (N_7,In_617,In_1328);
nand U8 (N_8,In_1206,In_1354);
nand U9 (N_9,In_455,In_1152);
and U10 (N_10,In_807,In_963);
xnor U11 (N_11,In_190,In_619);
and U12 (N_12,In_690,In_528);
nor U13 (N_13,In_1068,In_903);
nor U14 (N_14,In_755,In_35);
nand U15 (N_15,In_192,In_1244);
nor U16 (N_16,In_951,In_529);
and U17 (N_17,In_911,In_220);
and U18 (N_18,In_391,In_1471);
nand U19 (N_19,In_921,In_1454);
or U20 (N_20,In_221,In_649);
or U21 (N_21,In_277,In_1326);
and U22 (N_22,In_939,In_1358);
nor U23 (N_23,In_889,In_1385);
nor U24 (N_24,In_1440,In_1472);
or U25 (N_25,In_1459,In_106);
nand U26 (N_26,In_203,In_381);
or U27 (N_27,In_31,In_1367);
nor U28 (N_28,In_1172,In_1382);
nor U29 (N_29,In_744,In_21);
or U30 (N_30,In_95,In_885);
or U31 (N_31,In_270,In_626);
nor U32 (N_32,In_522,In_1429);
nor U33 (N_33,In_1297,In_441);
and U34 (N_34,In_1123,In_1029);
or U35 (N_35,In_1431,In_1415);
and U36 (N_36,In_235,In_394);
and U37 (N_37,In_197,In_593);
and U38 (N_38,In_1341,In_1254);
or U39 (N_39,In_677,In_533);
nand U40 (N_40,In_1443,In_151);
or U41 (N_41,In_1181,In_965);
and U42 (N_42,In_90,In_931);
nor U43 (N_43,In_970,In_1339);
nand U44 (N_44,In_797,In_377);
xnor U45 (N_45,In_412,In_1421);
nand U46 (N_46,In_19,In_1122);
nor U47 (N_47,In_1176,In_309);
or U48 (N_48,In_680,In_3);
xor U49 (N_49,In_919,In_1002);
xnor U50 (N_50,In_263,In_325);
and U51 (N_51,In_557,In_176);
or U52 (N_52,In_1369,In_443);
and U53 (N_53,In_374,In_682);
nand U54 (N_54,In_365,In_85);
nor U55 (N_55,In_205,In_702);
nor U56 (N_56,In_851,In_1248);
or U57 (N_57,In_524,In_743);
xnor U58 (N_58,In_125,In_375);
and U59 (N_59,In_1252,In_163);
or U60 (N_60,In_713,In_242);
and U61 (N_61,In_378,In_438);
nand U62 (N_62,In_218,In_1311);
nor U63 (N_63,In_1357,In_1491);
nand U64 (N_64,In_346,In_62);
nor U65 (N_65,In_1222,In_298);
or U66 (N_66,In_1427,In_1072);
xnor U67 (N_67,In_1204,In_356);
nand U68 (N_68,In_737,In_578);
nand U69 (N_69,In_767,In_818);
or U70 (N_70,In_511,In_282);
or U71 (N_71,In_369,In_1110);
nand U72 (N_72,In_1209,In_1470);
nand U73 (N_73,In_445,In_69);
nor U74 (N_74,In_312,In_1322);
nand U75 (N_75,In_780,In_1462);
and U76 (N_76,In_265,In_367);
and U77 (N_77,In_305,In_1196);
nor U78 (N_78,In_1379,In_1488);
or U79 (N_79,In_43,In_761);
or U80 (N_80,In_981,In_29);
and U81 (N_81,In_654,In_1126);
or U82 (N_82,In_845,In_139);
or U83 (N_83,In_1094,In_161);
nor U84 (N_84,In_523,In_512);
and U85 (N_85,In_558,In_450);
or U86 (N_86,In_491,In_787);
and U87 (N_87,In_354,In_1154);
or U88 (N_88,In_422,In_666);
or U89 (N_89,In_1098,In_754);
nor U90 (N_90,In_1109,In_1085);
and U91 (N_91,In_728,In_130);
nor U92 (N_92,In_1120,In_448);
nor U93 (N_93,In_841,In_1046);
nor U94 (N_94,In_1225,In_793);
nor U95 (N_95,In_212,In_1145);
and U96 (N_96,In_335,In_295);
nor U97 (N_97,In_293,In_543);
nand U98 (N_98,In_829,In_1489);
nand U99 (N_99,In_627,In_509);
nand U100 (N_100,In_1399,In_1477);
nand U101 (N_101,In_1082,In_238);
and U102 (N_102,In_147,In_722);
xnor U103 (N_103,In_1381,In_819);
or U104 (N_104,In_1307,In_414);
or U105 (N_105,In_494,In_956);
or U106 (N_106,In_1131,In_925);
and U107 (N_107,In_261,In_1093);
nor U108 (N_108,In_1166,In_1057);
and U109 (N_109,In_531,In_1139);
nand U110 (N_110,In_1346,In_526);
nand U111 (N_111,In_968,In_673);
nand U112 (N_112,In_742,In_363);
nor U113 (N_113,In_824,In_16);
or U114 (N_114,In_456,In_368);
nor U115 (N_115,In_1352,In_1115);
and U116 (N_116,In_255,In_1273);
nor U117 (N_117,In_294,In_167);
nor U118 (N_118,In_904,In_639);
nand U119 (N_119,In_186,In_870);
and U120 (N_120,In_124,In_561);
or U121 (N_121,In_988,In_338);
nor U122 (N_122,In_237,In_606);
nor U123 (N_123,In_1320,In_983);
nor U124 (N_124,In_916,In_707);
nand U125 (N_125,In_1490,In_60);
nor U126 (N_126,In_1242,In_143);
or U127 (N_127,In_1272,In_894);
or U128 (N_128,In_960,In_901);
nor U129 (N_129,In_1410,In_663);
xor U130 (N_130,In_646,In_103);
nor U131 (N_131,In_185,In_1069);
nand U132 (N_132,In_97,In_588);
nand U133 (N_133,In_556,In_679);
nand U134 (N_134,In_1052,In_1264);
nor U135 (N_135,In_1387,In_301);
nand U136 (N_136,In_315,In_1373);
or U137 (N_137,In_1496,In_625);
and U138 (N_138,In_248,In_1301);
and U139 (N_139,In_539,In_624);
or U140 (N_140,In_936,In_891);
nor U141 (N_141,In_1392,In_1370);
nand U142 (N_142,In_1480,In_678);
or U143 (N_143,In_120,In_1420);
nor U144 (N_144,In_1251,In_250);
nand U145 (N_145,In_1193,In_168);
nand U146 (N_146,In_995,In_207);
or U147 (N_147,In_183,In_1147);
or U148 (N_148,In_1366,In_935);
or U149 (N_149,In_188,In_1444);
nand U150 (N_150,In_38,In_739);
nor U151 (N_151,In_590,In_882);
and U152 (N_152,In_407,In_244);
nor U153 (N_153,In_1185,In_57);
nand U154 (N_154,In_1405,In_1050);
and U155 (N_155,In_842,In_174);
or U156 (N_156,In_1450,In_213);
and U157 (N_157,In_286,In_803);
nor U158 (N_158,In_436,In_217);
xor U159 (N_159,In_1282,In_1389);
and U160 (N_160,In_1079,In_1200);
nand U161 (N_161,In_403,In_432);
or U162 (N_162,In_339,In_599);
and U163 (N_163,In_740,In_608);
and U164 (N_164,In_1287,In_78);
nor U165 (N_165,In_859,In_1487);
xor U166 (N_166,In_34,In_1195);
nand U167 (N_167,In_108,In_961);
xnor U168 (N_168,In_1034,In_421);
and U169 (N_169,In_1021,In_5);
nand U170 (N_170,In_607,In_877);
and U171 (N_171,In_347,In_300);
nand U172 (N_172,In_763,In_598);
nor U173 (N_173,In_764,In_75);
and U174 (N_174,In_1237,In_1055);
nand U175 (N_175,In_1375,In_1157);
nand U176 (N_176,In_1359,In_1304);
nor U177 (N_177,In_292,In_1080);
and U178 (N_178,In_209,In_1127);
and U179 (N_179,In_836,In_835);
and U180 (N_180,In_1062,In_1128);
nand U181 (N_181,In_1058,In_199);
nor U182 (N_182,In_1309,In_1087);
nor U183 (N_183,In_955,In_538);
and U184 (N_184,In_10,In_1411);
or U185 (N_185,In_1347,In_579);
nor U186 (N_186,In_1108,In_1016);
nand U187 (N_187,In_1001,In_264);
and U188 (N_188,In_439,In_714);
and U189 (N_189,In_1011,In_506);
nor U190 (N_190,In_359,In_283);
xnor U191 (N_191,In_136,In_789);
and U192 (N_192,In_938,In_906);
or U193 (N_193,In_26,In_149);
nand U194 (N_194,In_989,In_37);
nor U195 (N_195,In_1111,In_1153);
or U196 (N_196,In_50,In_311);
and U197 (N_197,In_631,In_554);
nor U198 (N_198,In_817,In_379);
nor U199 (N_199,In_513,In_1344);
nand U200 (N_200,In_618,In_344);
or U201 (N_201,In_676,In_279);
or U202 (N_202,In_1289,In_1164);
and U203 (N_203,In_245,In_1025);
nor U204 (N_204,In_826,In_451);
or U205 (N_205,In_734,In_1099);
or U206 (N_206,In_1476,In_974);
and U207 (N_207,In_1168,In_405);
and U208 (N_208,In_1310,In_380);
nand U209 (N_209,In_285,In_474);
xnor U210 (N_210,In_975,In_310);
nor U211 (N_211,In_1231,In_1299);
nand U212 (N_212,In_1239,In_861);
nor U213 (N_213,In_322,In_642);
nand U214 (N_214,In_1250,In_1019);
xor U215 (N_215,In_1407,In_427);
or U216 (N_216,In_1140,In_794);
xnor U217 (N_217,In_792,In_1194);
or U218 (N_218,In_729,In_419);
nand U219 (N_219,In_905,In_475);
and U220 (N_220,In_100,In_700);
nand U221 (N_221,In_1014,In_1107);
nor U222 (N_222,In_45,In_162);
and U223 (N_223,In_1278,In_636);
or U224 (N_224,In_1372,In_635);
nor U225 (N_225,In_1092,In_483);
nand U226 (N_226,In_1292,In_630);
or U227 (N_227,In_316,In_349);
and U228 (N_228,In_1060,In_1066);
nor U229 (N_229,In_92,In_1283);
nand U230 (N_230,In_896,In_434);
nor U231 (N_231,In_1319,In_423);
nand U232 (N_232,In_401,In_71);
nand U233 (N_233,In_887,In_1054);
xnor U234 (N_234,In_6,In_495);
or U235 (N_235,In_18,In_1217);
and U236 (N_236,In_542,In_850);
nand U237 (N_237,In_1170,In_1497);
or U238 (N_238,In_417,In_775);
or U239 (N_239,In_1028,In_949);
or U240 (N_240,In_831,In_121);
nor U241 (N_241,In_1018,In_1048);
nor U242 (N_242,In_1324,In_144);
xor U243 (N_243,In_520,In_478);
or U244 (N_244,In_675,In_820);
and U245 (N_245,In_269,In_1269);
nand U246 (N_246,In_1355,In_604);
and U247 (N_247,In_281,In_937);
and U248 (N_248,In_719,In_1404);
and U249 (N_249,In_1081,In_692);
nand U250 (N_250,In_1067,In_546);
or U251 (N_251,In_798,In_908);
and U252 (N_252,In_28,In_537);
and U253 (N_253,In_321,In_156);
nand U254 (N_254,In_759,In_1412);
nor U255 (N_255,In_150,In_133);
or U256 (N_256,In_1143,In_442);
or U257 (N_257,In_716,In_204);
nand U258 (N_258,In_671,In_648);
nand U259 (N_259,In_726,In_997);
nor U260 (N_260,In_1312,In_1163);
or U261 (N_261,In_643,In_788);
nand U262 (N_262,In_385,In_544);
and U263 (N_263,In_247,In_1306);
nand U264 (N_264,In_944,In_1013);
nor U265 (N_265,In_1277,In_146);
nand U266 (N_266,In_1174,In_1484);
and U267 (N_267,In_530,In_917);
or U268 (N_268,In_1268,In_484);
nand U269 (N_269,In_516,In_540);
or U270 (N_270,In_1158,In_148);
xnor U271 (N_271,In_771,In_1467);
nor U272 (N_272,In_1474,In_1056);
nor U273 (N_273,In_249,In_1229);
or U274 (N_274,In_206,In_1286);
and U275 (N_275,In_79,In_527);
nand U276 (N_276,In_652,In_596);
nor U277 (N_277,In_1033,In_736);
and U278 (N_278,In_73,In_230);
nor U279 (N_279,In_198,In_465);
and U280 (N_280,In_1485,In_228);
xnor U281 (N_281,In_1343,In_1228);
nand U282 (N_282,In_592,In_697);
nor U283 (N_283,In_765,In_1119);
or U284 (N_284,In_262,In_155);
nor U285 (N_285,In_259,In_813);
nand U286 (N_286,In_1220,In_909);
or U287 (N_287,In_1134,In_660);
nor U288 (N_288,In_1409,In_776);
nor U289 (N_289,In_801,In_65);
nor U290 (N_290,In_480,In_1468);
or U291 (N_291,In_1430,In_66);
nor U292 (N_292,In_1378,In_131);
nor U293 (N_293,In_1116,In_950);
and U294 (N_294,In_517,In_211);
nand U295 (N_295,In_810,In_994);
or U296 (N_296,In_881,In_802);
nand U297 (N_297,In_668,In_1465);
nor U298 (N_298,In_1223,In_572);
nand U299 (N_299,In_1362,In_233);
nand U300 (N_300,In_387,In_865);
nand U301 (N_301,In_202,In_685);
or U302 (N_302,In_1267,In_138);
and U303 (N_303,In_748,In_1070);
nor U304 (N_304,In_1064,In_1447);
and U305 (N_305,In_398,In_973);
nand U306 (N_306,In_651,In_548);
and U307 (N_307,In_1183,In_932);
xnor U308 (N_308,In_1148,In_429);
nand U309 (N_309,In_957,In_98);
xor U310 (N_310,In_996,In_560);
and U311 (N_311,In_805,In_562);
xnor U312 (N_312,In_396,In_1149);
and U313 (N_313,In_1142,In_1247);
nor U314 (N_314,In_966,In_382);
and U315 (N_315,In_760,In_738);
nand U316 (N_316,In_603,In_1401);
and U317 (N_317,In_1363,In_366);
and U318 (N_318,In_234,In_469);
nand U319 (N_319,In_622,In_757);
nor U320 (N_320,In_1102,In_782);
nand U321 (N_321,In_900,In_123);
nand U322 (N_322,In_458,In_1380);
and U323 (N_323,In_32,In_1049);
and U324 (N_324,In_834,In_637);
and U325 (N_325,In_11,In_1043);
and U326 (N_326,In_825,In_541);
xnor U327 (N_327,In_425,In_1161);
nand U328 (N_328,In_376,In_89);
nor U329 (N_329,In_532,In_597);
and U330 (N_330,In_515,In_30);
and U331 (N_331,In_437,In_371);
or U332 (N_332,In_110,In_501);
nor U333 (N_333,In_866,In_927);
or U334 (N_334,In_240,In_534);
or U335 (N_335,In_1232,In_1088);
xnor U336 (N_336,In_1325,In_504);
or U337 (N_337,In_647,In_1159);
nand U338 (N_338,In_402,In_140);
nand U339 (N_339,In_1479,In_1336);
nand U340 (N_340,In_1483,In_661);
xnor U341 (N_341,In_634,In_843);
nor U342 (N_342,In_777,In_778);
nor U343 (N_343,In_1408,In_308);
xor U344 (N_344,In_122,In_1000);
xnor U345 (N_345,In_662,In_2);
nand U346 (N_346,In_1213,In_674);
or U347 (N_347,In_327,In_84);
or U348 (N_348,In_610,In_855);
or U349 (N_349,In_223,In_849);
or U350 (N_350,In_628,In_934);
nand U351 (N_351,In_940,In_681);
xnor U352 (N_352,In_926,In_733);
xnor U353 (N_353,In_113,In_486);
nor U354 (N_354,In_201,In_1432);
nand U355 (N_355,In_1114,In_1135);
nor U356 (N_356,In_397,In_1449);
and U357 (N_357,In_361,In_1270);
and U358 (N_358,In_1300,In_1235);
xnor U359 (N_359,In_51,In_452);
and U360 (N_360,In_1302,In_306);
nand U361 (N_361,In_1027,In_137);
xor U362 (N_362,In_1020,In_1285);
xnor U363 (N_363,In_64,In_1463);
nor U364 (N_364,In_165,In_1191);
nand U365 (N_365,In_94,In_977);
nand U366 (N_366,In_992,In_1323);
and U367 (N_367,In_153,In_547);
nor U368 (N_368,In_1199,In_470);
nand U369 (N_369,In_118,In_930);
nor U370 (N_370,In_418,In_166);
or U371 (N_371,In_1426,In_1210);
nand U372 (N_372,In_336,In_1065);
or U373 (N_373,In_468,In_1275);
nand U374 (N_374,In_880,In_948);
xnor U375 (N_375,In_864,In_567);
nor U376 (N_376,In_1318,In_128);
and U377 (N_377,In_979,In_847);
nand U378 (N_378,In_169,In_224);
xnor U379 (N_379,In_758,In_4);
nand U380 (N_380,In_1475,In_1439);
nand U381 (N_381,In_959,In_779);
xor U382 (N_382,In_1495,In_1331);
or U383 (N_383,In_698,In_246);
and U384 (N_384,In_46,In_857);
nor U385 (N_385,In_521,In_1418);
and U386 (N_386,In_1469,In_1010);
and U387 (N_387,In_252,In_1457);
nor U388 (N_388,In_1041,In_899);
nand U389 (N_389,In_1263,In_222);
nor U390 (N_390,In_1243,In_821);
nor U391 (N_391,In_587,In_268);
nor U392 (N_392,In_329,In_157);
nand U393 (N_393,In_725,In_431);
and U394 (N_394,In_187,In_574);
nand U395 (N_395,In_447,In_1321);
nand U396 (N_396,In_783,In_969);
nor U397 (N_397,In_1342,In_1039);
or U398 (N_398,In_806,In_735);
and U399 (N_399,In_72,In_967);
or U400 (N_400,In_1208,In_164);
and U401 (N_401,In_753,In_337);
xnor U402 (N_402,In_1132,In_1315);
or U403 (N_403,In_119,In_1478);
nand U404 (N_404,In_1221,In_351);
nand U405 (N_405,In_1190,In_471);
nand U406 (N_406,In_145,In_229);
nor U407 (N_407,In_493,In_297);
and U408 (N_408,In_946,In_127);
or U409 (N_409,In_179,In_1047);
nand U410 (N_410,In_769,In_695);
xnor U411 (N_411,In_1156,In_1042);
nand U412 (N_412,In_1051,In_355);
and U413 (N_413,In_884,In_920);
or U414 (N_414,In_77,In_1075);
nand U415 (N_415,In_796,In_406);
or U416 (N_416,In_61,In_575);
xor U417 (N_417,In_1155,In_47);
nor U418 (N_418,In_809,In_952);
or U419 (N_419,In_345,In_879);
and U420 (N_420,In_1086,In_814);
nand U421 (N_421,In_485,In_576);
nor U422 (N_422,In_1274,In_559);
nor U423 (N_423,In_1071,In_444);
and U424 (N_424,In_341,In_1423);
nand U425 (N_425,In_462,In_709);
nor U426 (N_426,In_586,In_160);
or U427 (N_427,In_696,In_86);
and U428 (N_428,In_291,In_1189);
and U429 (N_429,In_68,In_773);
nor U430 (N_430,In_833,In_1394);
nand U431 (N_431,In_918,In_1162);
and U432 (N_432,In_180,In_258);
nand U433 (N_433,In_1305,In_732);
and U434 (N_434,In_1337,In_116);
and U435 (N_435,In_941,In_569);
nand U436 (N_436,In_388,In_563);
nor U437 (N_437,In_227,In_1233);
nand U438 (N_438,In_41,In_1446);
xnor U439 (N_439,In_473,In_1433);
nor U440 (N_440,In_840,In_1303);
nor U441 (N_441,In_1197,In_585);
or U442 (N_442,In_514,In_1376);
nand U443 (N_443,In_1097,In_1351);
and U444 (N_444,In_871,In_1249);
nand U445 (N_445,In_1493,In_890);
and U446 (N_446,In_1089,In_1340);
or U447 (N_447,In_1073,In_27);
nand U448 (N_448,In_1173,In_307);
nand U449 (N_449,In_632,In_741);
or U450 (N_450,In_54,In_1117);
nand U451 (N_451,In_1452,In_1255);
xor U452 (N_452,In_1486,In_621);
or U453 (N_453,In_104,In_1413);
or U454 (N_454,In_768,In_340);
nor U455 (N_455,In_1038,In_644);
or U456 (N_456,In_785,In_1040);
nor U457 (N_457,In_1461,In_1211);
xor U458 (N_458,In_1160,In_770);
nand U459 (N_459,In_980,In_594);
nor U460 (N_460,In_1276,In_1017);
nor U461 (N_461,In_1428,In_290);
nor U462 (N_462,In_1226,In_200);
and U463 (N_463,In_457,In_177);
or U464 (N_464,In_348,In_984);
and U465 (N_465,In_278,In_1494);
nand U466 (N_466,In_314,In_689);
or U467 (N_467,In_853,In_232);
nand U468 (N_468,In_1256,In_749);
or U469 (N_469,In_1112,In_1146);
nand U470 (N_470,In_1003,In_1374);
nor U471 (N_471,In_1422,In_114);
nor U472 (N_472,In_76,In_1290);
nor U473 (N_473,In_1205,In_87);
nand U474 (N_474,In_1473,In_208);
nor U475 (N_475,In_525,In_962);
or U476 (N_476,In_1403,In_815);
xnor U477 (N_477,In_352,In_446);
or U478 (N_478,In_795,In_56);
and U479 (N_479,In_99,In_583);
nor U480 (N_480,In_1383,In_489);
nor U481 (N_481,In_1313,In_440);
nand U482 (N_482,In_717,In_657);
nor U483 (N_483,In_658,In_490);
and U484 (N_484,In_1314,In_1150);
xnor U485 (N_485,In_605,In_170);
or U486 (N_486,In_129,In_1214);
nand U487 (N_487,In_112,In_874);
nor U488 (N_488,In_1498,In_786);
nor U489 (N_489,In_1182,In_318);
nor U490 (N_490,In_459,In_1133);
or U491 (N_491,In_830,In_404);
or U492 (N_492,In_1258,In_1386);
xor U493 (N_493,In_22,In_1201);
xnor U494 (N_494,In_498,In_1044);
and U495 (N_495,In_577,In_132);
or U496 (N_496,In_159,In_1371);
nor U497 (N_497,In_1434,In_878);
or U498 (N_498,In_1350,In_1104);
or U499 (N_499,In_433,In_426);
nor U500 (N_500,In_858,In_1437);
nand U501 (N_501,In_655,In_832);
and U502 (N_502,In_756,In_415);
and U503 (N_503,In_111,In_1045);
nor U504 (N_504,In_1438,In_1406);
or U505 (N_505,In_500,In_1187);
and U506 (N_506,In_91,In_115);
nor U507 (N_507,In_313,In_1400);
nand U508 (N_508,In_611,In_924);
or U509 (N_509,In_1460,In_1333);
xor U510 (N_510,In_747,In_175);
or U511 (N_511,In_1393,In_373);
nand U512 (N_512,In_463,In_774);
nor U513 (N_513,In_1230,In_914);
nor U514 (N_514,In_273,In_1348);
or U515 (N_515,In_1455,In_48);
nand U516 (N_516,In_645,In_623);
xor U517 (N_517,In_1171,In_1091);
nand U518 (N_518,In_52,In_1425);
xor U519 (N_519,In_1448,In_1262);
xnor U520 (N_520,In_691,In_1424);
xnor U521 (N_521,In_875,In_1053);
and U522 (N_522,In_411,In_392);
nor U523 (N_523,In_1360,In_1240);
nor U524 (N_524,In_615,In_410);
nand U525 (N_525,In_466,In_499);
nor U526 (N_526,In_191,In_1026);
and U527 (N_527,In_892,In_568);
nor U528 (N_528,In_1353,In_852);
or U529 (N_529,In_1391,In_822);
nand U530 (N_530,In_828,In_1482);
nand U531 (N_531,In_63,In_1456);
xnor U532 (N_532,In_693,In_573);
and U533 (N_533,In_923,In_1203);
nand U534 (N_534,In_602,In_362);
and U535 (N_535,In_1464,In_1224);
nor U536 (N_536,In_1090,In_1365);
and U537 (N_537,In_343,In_194);
and U538 (N_538,In_260,In_497);
or U539 (N_539,In_296,In_505);
or U540 (N_540,In_910,In_667);
xor U541 (N_541,In_196,In_1451);
and U542 (N_542,In_724,In_1345);
or U543 (N_543,In_1202,In_808);
and U544 (N_544,In_620,In_1436);
and U545 (N_545,In_650,In_1012);
and U546 (N_546,In_971,In_550);
and U547 (N_547,In_182,In_751);
or U548 (N_548,In_342,In_88);
and U549 (N_549,In_36,In_323);
nand U550 (N_550,In_55,In_134);
or U551 (N_551,In_686,In_1151);
nor U552 (N_552,In_353,In_1212);
and U553 (N_553,In_326,In_536);
or U554 (N_554,In_328,In_750);
nor U555 (N_555,In_876,In_929);
or U556 (N_556,In_320,In_1004);
and U557 (N_557,In_154,In_848);
nand U558 (N_558,In_1442,In_584);
or U559 (N_559,In_704,In_791);
or U560 (N_560,In_552,In_898);
or U561 (N_561,In_1398,In_1063);
nor U562 (N_562,In_510,In_784);
and U563 (N_563,In_897,In_181);
and U564 (N_564,In_1481,In_612);
nand U565 (N_565,In_332,In_854);
nand U566 (N_566,In_1192,In_210);
nor U567 (N_567,In_1207,In_1396);
nor U568 (N_568,In_449,In_1106);
nand U569 (N_569,In_289,In_1124);
or U570 (N_570,In_42,In_254);
or U571 (N_571,In_1,In_812);
nand U572 (N_572,In_659,In_1024);
or U573 (N_573,In_1308,In_488);
and U574 (N_574,In_869,In_991);
nand U575 (N_575,In_985,In_1022);
or U576 (N_576,In_752,In_1130);
or U577 (N_577,In_1435,In_928);
xnor U578 (N_578,In_1035,In_1280);
nor U579 (N_579,In_1334,In_1327);
and U580 (N_580,In_93,In_1167);
nand U581 (N_581,In_49,In_236);
nand U582 (N_582,In_684,In_288);
nand U583 (N_583,In_333,In_372);
xnor U584 (N_584,In_731,In_1007);
and U585 (N_585,In_708,In_1083);
or U586 (N_586,In_1458,In_1178);
nor U587 (N_587,In_409,In_1384);
or U588 (N_588,In_1180,In_8);
and U589 (N_589,In_712,In_720);
and U590 (N_590,In_14,In_317);
or U591 (N_591,In_964,In_82);
xnor U592 (N_592,In_141,In_1335);
nor U593 (N_593,In_553,In_389);
and U594 (N_594,In_1284,In_253);
xnor U595 (N_595,In_976,In_867);
or U596 (N_596,In_564,In_101);
or U597 (N_597,In_1219,In_503);
or U598 (N_598,In_274,In_888);
nor U599 (N_599,In_256,In_730);
or U600 (N_600,In_267,In_9);
nor U601 (N_601,In_545,In_287);
or U602 (N_602,In_251,In_954);
nand U603 (N_603,In_225,In_1402);
nand U604 (N_604,In_1129,In_15);
nor U605 (N_605,In_74,In_799);
nand U606 (N_606,In_641,In_1416);
nand U607 (N_607,In_1074,In_629);
and U608 (N_608,In_257,In_1492);
nor U609 (N_609,In_816,In_216);
nor U610 (N_610,In_1241,In_360);
nor U611 (N_611,In_863,In_280);
and U612 (N_612,In_58,In_868);
or U613 (N_613,In_370,In_601);
nor U614 (N_614,In_496,In_1023);
and U615 (N_615,In_383,In_1077);
xor U616 (N_616,In_838,In_464);
xor U617 (N_617,In_476,In_711);
and U618 (N_618,In_913,In_721);
or U619 (N_619,In_13,In_633);
and U620 (N_620,In_856,In_319);
nor U621 (N_621,In_1377,In_1257);
nand U622 (N_622,In_1036,In_430);
or U623 (N_623,In_1296,In_986);
nor U624 (N_624,In_1281,In_1136);
nor U625 (N_625,In_1030,In_135);
or U626 (N_626,In_59,In_416);
nor U627 (N_627,In_1293,In_1103);
or U628 (N_628,In_570,In_1165);
or U629 (N_629,In_1101,In_715);
and U630 (N_630,In_912,In_482);
nor U631 (N_631,In_1390,In_1188);
nand U632 (N_632,In_1329,In_862);
or U633 (N_633,In_1395,In_1261);
nand U634 (N_634,In_670,In_358);
nand U635 (N_635,In_1445,In_171);
and U636 (N_636,In_978,In_1414);
nand U637 (N_637,In_334,In_1100);
or U638 (N_638,In_549,In_1009);
nand U639 (N_639,In_1234,In_1364);
xnor U640 (N_640,In_454,In_844);
and U641 (N_641,In_428,In_271);
nor U642 (N_642,In_555,In_1137);
nand U643 (N_643,In_1084,In_1141);
and U644 (N_644,In_565,In_173);
and U645 (N_645,In_656,In_126);
nor U646 (N_646,In_420,In_640);
xnor U647 (N_647,In_1031,In_998);
nor U648 (N_648,In_987,In_551);
and U649 (N_649,In_1015,In_435);
and U650 (N_650,In_942,In_811);
or U651 (N_651,In_395,In_1216);
and U652 (N_652,In_1061,In_20);
or U653 (N_653,In_453,In_189);
and U654 (N_654,In_331,In_492);
nand U655 (N_655,In_982,In_653);
nand U656 (N_656,In_589,In_142);
or U657 (N_657,In_609,In_1259);
nand U658 (N_658,In_688,In_1125);
xor U659 (N_659,In_800,In_1453);
and U660 (N_660,In_508,In_947);
nand U661 (N_661,In_25,In_1330);
and U662 (N_662,In_81,In_893);
or U663 (N_663,In_804,In_1419);
nand U664 (N_664,In_665,In_1499);
nor U665 (N_665,In_638,In_53);
nand U666 (N_666,In_364,In_1279);
nand U667 (N_667,In_1295,In_614);
or U668 (N_668,In_846,In_860);
nor U669 (N_669,In_324,In_276);
and U670 (N_670,In_883,In_595);
or U671 (N_671,In_502,In_24);
or U672 (N_672,In_945,In_1466);
and U673 (N_673,In_518,In_284);
and U674 (N_674,In_1417,In_193);
nand U675 (N_675,In_1266,In_1397);
nor U676 (N_676,In_718,In_1076);
nor U677 (N_677,In_687,In_1184);
nor U678 (N_678,In_272,In_1175);
xnor U679 (N_679,In_1169,In_96);
nand U680 (N_680,In_999,In_781);
and U681 (N_681,In_1227,In_195);
xnor U682 (N_682,In_461,In_460);
or U683 (N_683,In_304,In_571);
nor U684 (N_684,In_184,In_1059);
and U685 (N_685,In_535,In_672);
xnor U686 (N_686,In_1095,In_40);
nand U687 (N_687,In_699,In_107);
nor U688 (N_688,In_39,In_472);
or U689 (N_689,In_1260,In_1349);
nor U690 (N_690,In_933,In_1338);
nand U691 (N_691,In_746,In_581);
nor U692 (N_692,In_710,In_766);
or U693 (N_693,In_993,In_67);
nor U694 (N_694,In_487,In_582);
and U695 (N_695,In_23,In_1005);
nand U696 (N_696,In_243,In_705);
or U697 (N_697,In_790,In_1215);
nand U698 (N_698,In_384,In_1265);
or U699 (N_699,In_178,In_386);
and U700 (N_700,In_1078,In_580);
nand U701 (N_701,In_839,In_424);
nand U702 (N_702,In_239,In_837);
or U703 (N_703,In_886,In_727);
xnor U704 (N_704,In_330,In_109);
nor U705 (N_705,In_0,In_479);
nand U706 (N_706,In_703,In_1032);
or U707 (N_707,In_613,In_12);
nor U708 (N_708,In_70,In_477);
or U709 (N_709,In_275,In_1006);
nand U710 (N_710,In_302,In_507);
nand U711 (N_711,In_390,In_172);
nand U712 (N_712,In_1271,In_915);
or U713 (N_713,In_7,In_1356);
xnor U714 (N_714,In_902,In_44);
or U715 (N_715,In_214,In_241);
xnor U716 (N_716,In_357,In_299);
or U717 (N_717,In_80,In_226);
nand U718 (N_718,In_1298,In_1177);
nor U719 (N_719,In_1238,In_1294);
nand U720 (N_720,In_943,In_33);
nor U721 (N_721,In_772,In_1096);
and U722 (N_722,In_873,In_400);
and U723 (N_723,In_1198,In_872);
or U724 (N_724,In_1317,In_1186);
or U725 (N_725,In_1253,In_303);
nand U726 (N_726,In_83,In_158);
and U727 (N_727,In_215,In_152);
xor U728 (N_728,In_591,In_745);
xor U729 (N_729,In_1361,In_408);
or U730 (N_730,In_1008,In_669);
and U731 (N_731,In_350,In_953);
or U732 (N_732,In_701,In_1113);
xor U733 (N_733,In_1388,In_683);
and U734 (N_734,In_219,In_231);
nand U735 (N_735,In_1291,In_467);
or U736 (N_736,In_706,In_1441);
nor U737 (N_737,In_990,In_566);
xnor U738 (N_738,In_1368,In_1037);
or U739 (N_739,In_1105,In_393);
xnor U740 (N_740,In_922,In_907);
and U741 (N_741,In_1118,In_17);
nand U742 (N_742,In_399,In_117);
nand U743 (N_743,In_694,In_1316);
nand U744 (N_744,In_1288,In_958);
or U745 (N_745,In_895,In_1121);
or U746 (N_746,In_664,In_1236);
nor U747 (N_747,In_723,In_413);
nor U748 (N_748,In_519,In_1144);
or U749 (N_749,In_972,In_1179);
nor U750 (N_750,N_426,N_670);
and U751 (N_751,N_330,N_290);
nand U752 (N_752,N_421,N_232);
nor U753 (N_753,N_239,N_193);
and U754 (N_754,N_257,N_500);
or U755 (N_755,N_139,N_334);
or U756 (N_756,N_361,N_648);
nor U757 (N_757,N_737,N_225);
nand U758 (N_758,N_517,N_64);
or U759 (N_759,N_480,N_604);
and U760 (N_760,N_574,N_52);
or U761 (N_761,N_98,N_716);
and U762 (N_762,N_730,N_204);
or U763 (N_763,N_159,N_739);
nand U764 (N_764,N_355,N_601);
nor U765 (N_765,N_173,N_196);
xor U766 (N_766,N_405,N_635);
nor U767 (N_767,N_178,N_710);
nand U768 (N_768,N_510,N_580);
and U769 (N_769,N_206,N_721);
nand U770 (N_770,N_133,N_434);
and U771 (N_771,N_276,N_566);
and U772 (N_772,N_532,N_261);
nand U773 (N_773,N_283,N_85);
xnor U774 (N_774,N_651,N_265);
or U775 (N_775,N_288,N_570);
or U776 (N_776,N_121,N_630);
nor U777 (N_777,N_294,N_57);
xor U778 (N_778,N_735,N_218);
xor U779 (N_779,N_62,N_609);
or U780 (N_780,N_299,N_612);
or U781 (N_781,N_297,N_199);
nand U782 (N_782,N_7,N_594);
and U783 (N_783,N_715,N_528);
and U784 (N_784,N_745,N_310);
and U785 (N_785,N_89,N_189);
nor U786 (N_786,N_47,N_95);
nor U787 (N_787,N_148,N_45);
xor U788 (N_788,N_460,N_124);
xor U789 (N_789,N_593,N_567);
nand U790 (N_790,N_430,N_511);
and U791 (N_791,N_63,N_669);
xor U792 (N_792,N_701,N_97);
nor U793 (N_793,N_37,N_616);
nand U794 (N_794,N_38,N_625);
nor U795 (N_795,N_87,N_191);
xnor U796 (N_796,N_524,N_584);
nor U797 (N_797,N_126,N_269);
and U798 (N_798,N_514,N_111);
nand U799 (N_799,N_321,N_492);
nand U800 (N_800,N_342,N_679);
nand U801 (N_801,N_181,N_53);
xor U802 (N_802,N_263,N_585);
nor U803 (N_803,N_676,N_262);
nand U804 (N_804,N_72,N_114);
nand U805 (N_805,N_92,N_33);
or U806 (N_806,N_315,N_116);
nor U807 (N_807,N_543,N_314);
nor U808 (N_808,N_392,N_234);
or U809 (N_809,N_203,N_546);
and U810 (N_810,N_1,N_741);
nor U811 (N_811,N_266,N_352);
and U812 (N_812,N_446,N_661);
nand U813 (N_813,N_591,N_354);
or U814 (N_814,N_496,N_388);
or U815 (N_815,N_638,N_120);
xnor U816 (N_816,N_311,N_190);
xor U817 (N_817,N_439,N_305);
nand U818 (N_818,N_639,N_699);
nand U819 (N_819,N_744,N_526);
or U820 (N_820,N_200,N_668);
nor U821 (N_821,N_647,N_12);
or U822 (N_822,N_449,N_665);
xor U823 (N_823,N_40,N_530);
and U824 (N_824,N_689,N_558);
or U825 (N_825,N_579,N_633);
or U826 (N_826,N_478,N_158);
nand U827 (N_827,N_373,N_337);
nand U828 (N_828,N_219,N_141);
and U829 (N_829,N_484,N_435);
xnor U830 (N_830,N_274,N_350);
and U831 (N_831,N_589,N_748);
nand U832 (N_832,N_508,N_652);
xnor U833 (N_833,N_101,N_734);
nor U834 (N_834,N_367,N_43);
and U835 (N_835,N_226,N_340);
nand U836 (N_836,N_258,N_403);
or U837 (N_837,N_260,N_731);
or U838 (N_838,N_27,N_73);
nor U839 (N_839,N_51,N_212);
or U840 (N_840,N_105,N_614);
and U841 (N_841,N_497,N_55);
nand U842 (N_842,N_18,N_666);
nor U843 (N_843,N_685,N_658);
nand U844 (N_844,N_391,N_390);
nand U845 (N_845,N_680,N_109);
or U846 (N_846,N_255,N_413);
and U847 (N_847,N_143,N_254);
and U848 (N_848,N_417,N_119);
xnor U849 (N_849,N_194,N_175);
nand U850 (N_850,N_91,N_19);
nand U851 (N_851,N_100,N_729);
nor U852 (N_852,N_207,N_36);
and U853 (N_853,N_621,N_402);
or U854 (N_854,N_166,N_533);
and U855 (N_855,N_375,N_78);
xor U856 (N_856,N_397,N_182);
and U857 (N_857,N_581,N_582);
or U858 (N_858,N_736,N_586);
xor U859 (N_859,N_523,N_184);
and U860 (N_860,N_235,N_214);
nor U861 (N_861,N_695,N_171);
nand U862 (N_862,N_383,N_90);
and U863 (N_863,N_479,N_606);
or U864 (N_864,N_2,N_146);
and U865 (N_865,N_197,N_664);
or U866 (N_866,N_487,N_195);
and U867 (N_867,N_698,N_285);
or U868 (N_868,N_592,N_519);
nand U869 (N_869,N_0,N_169);
or U870 (N_870,N_549,N_600);
xnor U871 (N_871,N_252,N_180);
and U872 (N_872,N_281,N_505);
nor U873 (N_873,N_371,N_231);
and U874 (N_874,N_291,N_327);
and U875 (N_875,N_167,N_369);
and U876 (N_876,N_335,N_248);
and U877 (N_877,N_747,N_718);
or U878 (N_878,N_351,N_83);
nor U879 (N_879,N_565,N_39);
or U880 (N_880,N_289,N_712);
nand U881 (N_881,N_551,N_316);
and U882 (N_882,N_536,N_153);
or U883 (N_883,N_11,N_14);
and U884 (N_884,N_401,N_270);
nand U885 (N_885,N_389,N_576);
or U886 (N_886,N_690,N_432);
nor U887 (N_887,N_564,N_448);
or U888 (N_888,N_458,N_722);
nor U889 (N_889,N_209,N_429);
and U890 (N_890,N_339,N_470);
or U891 (N_891,N_293,N_74);
and U892 (N_892,N_451,N_475);
nand U893 (N_893,N_694,N_509);
or U894 (N_894,N_221,N_140);
nor U895 (N_895,N_468,N_151);
and U896 (N_896,N_675,N_704);
nor U897 (N_897,N_702,N_697);
or U898 (N_898,N_58,N_28);
or U899 (N_899,N_346,N_10);
xor U900 (N_900,N_548,N_372);
or U901 (N_901,N_75,N_147);
nor U902 (N_902,N_466,N_740);
nor U903 (N_903,N_251,N_185);
nand U904 (N_904,N_296,N_208);
nand U905 (N_905,N_317,N_393);
nor U906 (N_906,N_682,N_366);
nor U907 (N_907,N_220,N_309);
nor U908 (N_908,N_476,N_501);
nand U909 (N_909,N_172,N_483);
or U910 (N_910,N_65,N_368);
nand U911 (N_911,N_336,N_253);
nor U912 (N_912,N_202,N_643);
nor U913 (N_913,N_272,N_99);
xor U914 (N_914,N_404,N_469);
nor U915 (N_915,N_556,N_452);
or U916 (N_916,N_130,N_619);
nand U917 (N_917,N_198,N_80);
and U918 (N_918,N_241,N_280);
nor U919 (N_919,N_110,N_507);
nand U920 (N_920,N_686,N_132);
and U921 (N_921,N_138,N_3);
or U922 (N_922,N_81,N_325);
and U923 (N_923,N_59,N_525);
and U924 (N_924,N_539,N_410);
nand U925 (N_925,N_168,N_738);
and U926 (N_926,N_152,N_513);
and U927 (N_927,N_673,N_442);
nand U928 (N_928,N_450,N_406);
nand U929 (N_929,N_424,N_343);
and U930 (N_930,N_603,N_544);
and U931 (N_931,N_16,N_136);
nand U932 (N_932,N_622,N_211);
and U933 (N_933,N_17,N_632);
xor U934 (N_934,N_654,N_646);
nor U935 (N_935,N_590,N_268);
or U936 (N_936,N_54,N_433);
nand U937 (N_937,N_481,N_323);
nand U938 (N_938,N_245,N_610);
and U939 (N_939,N_22,N_333);
and U940 (N_940,N_127,N_418);
nand U941 (N_941,N_502,N_719);
nor U942 (N_942,N_620,N_550);
and U943 (N_943,N_286,N_284);
or U944 (N_944,N_408,N_428);
nor U945 (N_945,N_400,N_331);
nor U946 (N_946,N_308,N_29);
nor U947 (N_947,N_527,N_84);
nand U948 (N_948,N_642,N_504);
nor U949 (N_949,N_34,N_471);
xor U950 (N_950,N_31,N_279);
nand U951 (N_951,N_444,N_568);
or U952 (N_952,N_250,N_332);
nor U953 (N_953,N_687,N_44);
xnor U954 (N_954,N_298,N_596);
or U955 (N_955,N_644,N_660);
nor U956 (N_956,N_681,N_453);
and U957 (N_957,N_683,N_246);
nor U958 (N_958,N_443,N_287);
or U959 (N_959,N_77,N_615);
xnor U960 (N_960,N_608,N_282);
or U961 (N_961,N_46,N_613);
xnor U962 (N_962,N_559,N_709);
and U963 (N_963,N_467,N_490);
nor U964 (N_964,N_457,N_278);
nor U965 (N_965,N_678,N_599);
or U966 (N_966,N_617,N_123);
and U967 (N_967,N_376,N_650);
nand U968 (N_968,N_577,N_228);
and U969 (N_969,N_672,N_176);
and U970 (N_970,N_300,N_463);
xnor U971 (N_971,N_521,N_149);
or U972 (N_972,N_267,N_144);
or U973 (N_973,N_223,N_349);
nor U974 (N_974,N_156,N_649);
nor U975 (N_975,N_96,N_9);
nand U976 (N_976,N_531,N_318);
or U977 (N_977,N_381,N_137);
nand U978 (N_978,N_529,N_94);
nand U979 (N_979,N_32,N_708);
nor U980 (N_980,N_386,N_436);
nor U981 (N_981,N_724,N_150);
nor U982 (N_982,N_216,N_135);
nand U983 (N_983,N_322,N_636);
and U984 (N_984,N_423,N_707);
and U985 (N_985,N_345,N_24);
or U986 (N_986,N_498,N_705);
nand U987 (N_987,N_555,N_416);
nor U988 (N_988,N_359,N_117);
or U989 (N_989,N_237,N_233);
or U990 (N_990,N_86,N_360);
nor U991 (N_991,N_569,N_485);
or U992 (N_992,N_247,N_552);
xnor U993 (N_993,N_387,N_720);
nand U994 (N_994,N_573,N_611);
or U995 (N_995,N_303,N_542);
xnor U996 (N_996,N_499,N_422);
and U997 (N_997,N_562,N_142);
nand U998 (N_998,N_411,N_727);
nand U999 (N_999,N_347,N_183);
and U1000 (N_1000,N_465,N_627);
or U1001 (N_1001,N_348,N_362);
and U1002 (N_1002,N_662,N_482);
or U1003 (N_1003,N_71,N_48);
xor U1004 (N_1004,N_363,N_61);
nand U1005 (N_1005,N_742,N_656);
nor U1006 (N_1006,N_455,N_50);
nand U1007 (N_1007,N_595,N_688);
and U1008 (N_1008,N_629,N_503);
xnor U1009 (N_1009,N_93,N_412);
or U1010 (N_1010,N_201,N_431);
xor U1011 (N_1011,N_437,N_186);
nand U1012 (N_1012,N_82,N_165);
nor U1013 (N_1013,N_634,N_560);
nor U1014 (N_1014,N_653,N_456);
nand U1015 (N_1015,N_491,N_399);
nand U1016 (N_1016,N_671,N_227);
or U1017 (N_1017,N_8,N_242);
nor U1018 (N_1018,N_728,N_15);
and U1019 (N_1019,N_474,N_42);
and U1020 (N_1020,N_711,N_364);
or U1021 (N_1021,N_192,N_13);
nor U1022 (N_1022,N_541,N_554);
and U1023 (N_1023,N_398,N_547);
nor U1024 (N_1024,N_161,N_215);
or U1025 (N_1025,N_88,N_696);
or U1026 (N_1026,N_409,N_69);
and U1027 (N_1027,N_425,N_494);
nand U1028 (N_1028,N_396,N_229);
or U1029 (N_1029,N_329,N_67);
and U1030 (N_1030,N_217,N_462);
nand U1031 (N_1031,N_370,N_575);
nor U1032 (N_1032,N_657,N_518);
xnor U1033 (N_1033,N_495,N_717);
nor U1034 (N_1034,N_598,N_545);
nand U1035 (N_1035,N_420,N_306);
and U1036 (N_1036,N_684,N_438);
and U1037 (N_1037,N_512,N_113);
or U1038 (N_1038,N_112,N_441);
nand U1039 (N_1039,N_240,N_749);
nand U1040 (N_1040,N_243,N_20);
and U1041 (N_1041,N_553,N_49);
nand U1042 (N_1042,N_743,N_353);
nor U1043 (N_1043,N_273,N_746);
nand U1044 (N_1044,N_578,N_691);
or U1045 (N_1045,N_56,N_640);
or U1046 (N_1046,N_128,N_377);
and U1047 (N_1047,N_641,N_256);
or U1048 (N_1048,N_703,N_160);
nor U1049 (N_1049,N_374,N_328);
and U1050 (N_1050,N_713,N_108);
nand U1051 (N_1051,N_125,N_414);
nor U1052 (N_1052,N_179,N_407);
nor U1053 (N_1053,N_131,N_464);
or U1054 (N_1054,N_302,N_25);
nor U1055 (N_1055,N_395,N_597);
and U1056 (N_1056,N_106,N_385);
nand U1057 (N_1057,N_725,N_520);
and U1058 (N_1058,N_259,N_6);
nor U1059 (N_1059,N_70,N_26);
or U1060 (N_1060,N_4,N_170);
and U1061 (N_1061,N_312,N_493);
nand U1062 (N_1062,N_540,N_394);
nor U1063 (N_1063,N_213,N_236);
and U1064 (N_1064,N_714,N_21);
nand U1065 (N_1065,N_304,N_655);
nand U1066 (N_1066,N_104,N_628);
and U1067 (N_1067,N_378,N_733);
and U1068 (N_1068,N_459,N_571);
and U1069 (N_1069,N_489,N_174);
and U1070 (N_1070,N_522,N_382);
nor U1071 (N_1071,N_326,N_275);
nand U1072 (N_1072,N_30,N_103);
nor U1073 (N_1073,N_427,N_588);
nor U1074 (N_1074,N_230,N_277);
and U1075 (N_1075,N_177,N_440);
xnor U1076 (N_1076,N_380,N_320);
and U1077 (N_1077,N_488,N_118);
xnor U1078 (N_1078,N_605,N_626);
or U1079 (N_1079,N_473,N_631);
nand U1080 (N_1080,N_292,N_66);
nand U1081 (N_1081,N_618,N_623);
nor U1082 (N_1082,N_472,N_5);
nor U1083 (N_1083,N_538,N_637);
or U1084 (N_1084,N_723,N_115);
or U1085 (N_1085,N_358,N_344);
xor U1086 (N_1086,N_607,N_301);
or U1087 (N_1087,N_692,N_319);
or U1088 (N_1088,N_107,N_244);
or U1089 (N_1089,N_324,N_122);
or U1090 (N_1090,N_356,N_357);
nor U1091 (N_1091,N_341,N_659);
nor U1092 (N_1092,N_129,N_561);
or U1093 (N_1093,N_145,N_205);
nor U1094 (N_1094,N_379,N_693);
and U1095 (N_1095,N_155,N_60);
or U1096 (N_1096,N_516,N_102);
nor U1097 (N_1097,N_587,N_506);
nand U1098 (N_1098,N_79,N_164);
xor U1099 (N_1099,N_645,N_187);
or U1100 (N_1100,N_445,N_583);
or U1101 (N_1101,N_726,N_537);
and U1102 (N_1102,N_534,N_535);
and U1103 (N_1103,N_134,N_76);
or U1104 (N_1104,N_624,N_677);
nand U1105 (N_1105,N_188,N_447);
and U1106 (N_1106,N_157,N_461);
or U1107 (N_1107,N_674,N_23);
xor U1108 (N_1108,N_384,N_515);
or U1109 (N_1109,N_35,N_264);
nor U1110 (N_1110,N_572,N_307);
or U1111 (N_1111,N_313,N_454);
nor U1112 (N_1112,N_338,N_162);
or U1113 (N_1113,N_667,N_271);
nor U1114 (N_1114,N_238,N_224);
or U1115 (N_1115,N_706,N_415);
or U1116 (N_1116,N_602,N_68);
nor U1117 (N_1117,N_41,N_563);
or U1118 (N_1118,N_557,N_365);
or U1119 (N_1119,N_700,N_163);
and U1120 (N_1120,N_210,N_222);
and U1121 (N_1121,N_732,N_154);
xor U1122 (N_1122,N_663,N_486);
or U1123 (N_1123,N_477,N_419);
and U1124 (N_1124,N_249,N_295);
nor U1125 (N_1125,N_417,N_19);
nand U1126 (N_1126,N_28,N_181);
or U1127 (N_1127,N_688,N_427);
xor U1128 (N_1128,N_511,N_404);
nor U1129 (N_1129,N_724,N_707);
xor U1130 (N_1130,N_347,N_5);
nor U1131 (N_1131,N_153,N_444);
and U1132 (N_1132,N_36,N_324);
nand U1133 (N_1133,N_705,N_64);
nor U1134 (N_1134,N_136,N_407);
and U1135 (N_1135,N_512,N_709);
or U1136 (N_1136,N_152,N_213);
and U1137 (N_1137,N_642,N_207);
nor U1138 (N_1138,N_597,N_468);
xor U1139 (N_1139,N_454,N_93);
nor U1140 (N_1140,N_674,N_606);
nand U1141 (N_1141,N_334,N_348);
nor U1142 (N_1142,N_580,N_22);
nor U1143 (N_1143,N_721,N_452);
or U1144 (N_1144,N_336,N_627);
xnor U1145 (N_1145,N_22,N_248);
nand U1146 (N_1146,N_630,N_101);
or U1147 (N_1147,N_535,N_342);
or U1148 (N_1148,N_24,N_388);
xor U1149 (N_1149,N_570,N_488);
and U1150 (N_1150,N_316,N_35);
xnor U1151 (N_1151,N_571,N_305);
or U1152 (N_1152,N_137,N_431);
nand U1153 (N_1153,N_716,N_108);
or U1154 (N_1154,N_606,N_632);
nor U1155 (N_1155,N_491,N_384);
and U1156 (N_1156,N_34,N_157);
nand U1157 (N_1157,N_632,N_194);
and U1158 (N_1158,N_392,N_374);
or U1159 (N_1159,N_228,N_400);
and U1160 (N_1160,N_717,N_626);
nand U1161 (N_1161,N_120,N_62);
or U1162 (N_1162,N_77,N_132);
or U1163 (N_1163,N_419,N_46);
and U1164 (N_1164,N_534,N_664);
or U1165 (N_1165,N_749,N_428);
and U1166 (N_1166,N_492,N_156);
and U1167 (N_1167,N_129,N_435);
xor U1168 (N_1168,N_744,N_124);
nand U1169 (N_1169,N_27,N_608);
nand U1170 (N_1170,N_105,N_486);
nand U1171 (N_1171,N_626,N_265);
or U1172 (N_1172,N_416,N_512);
nand U1173 (N_1173,N_478,N_571);
nand U1174 (N_1174,N_133,N_542);
nor U1175 (N_1175,N_410,N_236);
nand U1176 (N_1176,N_642,N_33);
nand U1177 (N_1177,N_720,N_548);
or U1178 (N_1178,N_113,N_246);
and U1179 (N_1179,N_449,N_640);
xnor U1180 (N_1180,N_508,N_4);
and U1181 (N_1181,N_79,N_262);
or U1182 (N_1182,N_380,N_504);
or U1183 (N_1183,N_643,N_109);
and U1184 (N_1184,N_92,N_538);
nand U1185 (N_1185,N_592,N_354);
nand U1186 (N_1186,N_121,N_1);
nor U1187 (N_1187,N_148,N_609);
or U1188 (N_1188,N_606,N_557);
nor U1189 (N_1189,N_204,N_320);
or U1190 (N_1190,N_507,N_257);
and U1191 (N_1191,N_263,N_232);
xor U1192 (N_1192,N_645,N_128);
or U1193 (N_1193,N_291,N_42);
and U1194 (N_1194,N_538,N_84);
and U1195 (N_1195,N_505,N_665);
nor U1196 (N_1196,N_703,N_613);
and U1197 (N_1197,N_682,N_488);
nor U1198 (N_1198,N_34,N_710);
and U1199 (N_1199,N_489,N_180);
or U1200 (N_1200,N_667,N_130);
nand U1201 (N_1201,N_684,N_377);
xnor U1202 (N_1202,N_346,N_80);
nand U1203 (N_1203,N_471,N_49);
nor U1204 (N_1204,N_644,N_383);
nor U1205 (N_1205,N_51,N_355);
and U1206 (N_1206,N_337,N_712);
nor U1207 (N_1207,N_452,N_182);
nor U1208 (N_1208,N_82,N_138);
nor U1209 (N_1209,N_25,N_389);
and U1210 (N_1210,N_5,N_223);
nand U1211 (N_1211,N_121,N_641);
or U1212 (N_1212,N_664,N_626);
xnor U1213 (N_1213,N_561,N_280);
or U1214 (N_1214,N_198,N_152);
xnor U1215 (N_1215,N_405,N_446);
or U1216 (N_1216,N_330,N_641);
nor U1217 (N_1217,N_139,N_212);
or U1218 (N_1218,N_222,N_534);
and U1219 (N_1219,N_128,N_385);
or U1220 (N_1220,N_729,N_476);
nor U1221 (N_1221,N_260,N_686);
nor U1222 (N_1222,N_595,N_219);
or U1223 (N_1223,N_151,N_82);
xnor U1224 (N_1224,N_659,N_595);
nand U1225 (N_1225,N_39,N_542);
nand U1226 (N_1226,N_310,N_300);
nand U1227 (N_1227,N_136,N_302);
xnor U1228 (N_1228,N_700,N_546);
and U1229 (N_1229,N_343,N_415);
nand U1230 (N_1230,N_64,N_112);
or U1231 (N_1231,N_490,N_23);
or U1232 (N_1232,N_435,N_194);
nand U1233 (N_1233,N_541,N_24);
nand U1234 (N_1234,N_711,N_601);
nor U1235 (N_1235,N_317,N_74);
and U1236 (N_1236,N_386,N_211);
or U1237 (N_1237,N_320,N_208);
and U1238 (N_1238,N_405,N_155);
and U1239 (N_1239,N_61,N_317);
nand U1240 (N_1240,N_558,N_478);
nor U1241 (N_1241,N_591,N_121);
nor U1242 (N_1242,N_372,N_497);
or U1243 (N_1243,N_270,N_50);
xor U1244 (N_1244,N_8,N_525);
nor U1245 (N_1245,N_408,N_271);
xor U1246 (N_1246,N_315,N_590);
nor U1247 (N_1247,N_80,N_414);
nand U1248 (N_1248,N_641,N_488);
nor U1249 (N_1249,N_709,N_549);
and U1250 (N_1250,N_532,N_700);
xor U1251 (N_1251,N_369,N_570);
nor U1252 (N_1252,N_89,N_153);
and U1253 (N_1253,N_696,N_263);
nand U1254 (N_1254,N_88,N_55);
nand U1255 (N_1255,N_223,N_505);
and U1256 (N_1256,N_688,N_728);
or U1257 (N_1257,N_228,N_667);
or U1258 (N_1258,N_630,N_300);
xnor U1259 (N_1259,N_735,N_724);
and U1260 (N_1260,N_593,N_317);
nand U1261 (N_1261,N_743,N_718);
or U1262 (N_1262,N_314,N_682);
or U1263 (N_1263,N_494,N_141);
and U1264 (N_1264,N_124,N_502);
nand U1265 (N_1265,N_638,N_717);
and U1266 (N_1266,N_404,N_327);
and U1267 (N_1267,N_121,N_609);
nand U1268 (N_1268,N_149,N_279);
and U1269 (N_1269,N_97,N_243);
nor U1270 (N_1270,N_572,N_12);
nand U1271 (N_1271,N_671,N_267);
or U1272 (N_1272,N_416,N_695);
xor U1273 (N_1273,N_533,N_321);
nand U1274 (N_1274,N_477,N_596);
xnor U1275 (N_1275,N_624,N_399);
or U1276 (N_1276,N_257,N_282);
and U1277 (N_1277,N_0,N_166);
or U1278 (N_1278,N_724,N_593);
nor U1279 (N_1279,N_319,N_68);
nor U1280 (N_1280,N_502,N_310);
xor U1281 (N_1281,N_432,N_156);
nand U1282 (N_1282,N_62,N_19);
and U1283 (N_1283,N_64,N_634);
or U1284 (N_1284,N_217,N_356);
or U1285 (N_1285,N_36,N_171);
or U1286 (N_1286,N_631,N_441);
or U1287 (N_1287,N_410,N_419);
nor U1288 (N_1288,N_289,N_288);
nor U1289 (N_1289,N_97,N_40);
or U1290 (N_1290,N_120,N_174);
nor U1291 (N_1291,N_741,N_140);
or U1292 (N_1292,N_385,N_173);
or U1293 (N_1293,N_684,N_66);
and U1294 (N_1294,N_126,N_656);
or U1295 (N_1295,N_48,N_611);
nand U1296 (N_1296,N_676,N_251);
nor U1297 (N_1297,N_631,N_229);
or U1298 (N_1298,N_498,N_362);
or U1299 (N_1299,N_178,N_303);
or U1300 (N_1300,N_445,N_685);
nand U1301 (N_1301,N_198,N_445);
and U1302 (N_1302,N_2,N_697);
nand U1303 (N_1303,N_62,N_410);
and U1304 (N_1304,N_77,N_264);
and U1305 (N_1305,N_360,N_20);
nor U1306 (N_1306,N_63,N_297);
xor U1307 (N_1307,N_389,N_376);
nand U1308 (N_1308,N_332,N_381);
xor U1309 (N_1309,N_204,N_327);
nand U1310 (N_1310,N_31,N_122);
xnor U1311 (N_1311,N_111,N_58);
and U1312 (N_1312,N_168,N_201);
or U1313 (N_1313,N_322,N_544);
and U1314 (N_1314,N_152,N_510);
or U1315 (N_1315,N_111,N_241);
and U1316 (N_1316,N_441,N_251);
xnor U1317 (N_1317,N_78,N_203);
and U1318 (N_1318,N_154,N_195);
nor U1319 (N_1319,N_571,N_450);
nor U1320 (N_1320,N_488,N_695);
nand U1321 (N_1321,N_489,N_27);
nor U1322 (N_1322,N_273,N_293);
and U1323 (N_1323,N_426,N_330);
or U1324 (N_1324,N_321,N_104);
nor U1325 (N_1325,N_600,N_648);
or U1326 (N_1326,N_346,N_185);
or U1327 (N_1327,N_358,N_149);
nand U1328 (N_1328,N_700,N_371);
nor U1329 (N_1329,N_66,N_517);
or U1330 (N_1330,N_718,N_371);
or U1331 (N_1331,N_576,N_57);
or U1332 (N_1332,N_407,N_564);
nand U1333 (N_1333,N_10,N_181);
and U1334 (N_1334,N_187,N_447);
nand U1335 (N_1335,N_136,N_94);
or U1336 (N_1336,N_394,N_591);
xnor U1337 (N_1337,N_669,N_370);
or U1338 (N_1338,N_335,N_169);
nand U1339 (N_1339,N_606,N_93);
and U1340 (N_1340,N_180,N_361);
or U1341 (N_1341,N_692,N_406);
nor U1342 (N_1342,N_386,N_108);
nor U1343 (N_1343,N_120,N_147);
and U1344 (N_1344,N_258,N_256);
nor U1345 (N_1345,N_466,N_663);
nor U1346 (N_1346,N_43,N_673);
nor U1347 (N_1347,N_82,N_501);
nand U1348 (N_1348,N_503,N_301);
nor U1349 (N_1349,N_573,N_46);
nand U1350 (N_1350,N_82,N_360);
nand U1351 (N_1351,N_120,N_86);
and U1352 (N_1352,N_182,N_185);
nand U1353 (N_1353,N_521,N_121);
nor U1354 (N_1354,N_485,N_383);
nor U1355 (N_1355,N_701,N_40);
and U1356 (N_1356,N_132,N_414);
or U1357 (N_1357,N_560,N_359);
nand U1358 (N_1358,N_619,N_639);
xnor U1359 (N_1359,N_451,N_505);
or U1360 (N_1360,N_576,N_448);
nor U1361 (N_1361,N_458,N_617);
and U1362 (N_1362,N_220,N_161);
or U1363 (N_1363,N_648,N_398);
nand U1364 (N_1364,N_48,N_248);
or U1365 (N_1365,N_455,N_694);
or U1366 (N_1366,N_467,N_621);
nor U1367 (N_1367,N_53,N_476);
and U1368 (N_1368,N_379,N_67);
and U1369 (N_1369,N_488,N_397);
xor U1370 (N_1370,N_205,N_479);
or U1371 (N_1371,N_0,N_362);
and U1372 (N_1372,N_160,N_70);
nand U1373 (N_1373,N_213,N_323);
nor U1374 (N_1374,N_341,N_557);
and U1375 (N_1375,N_515,N_621);
nor U1376 (N_1376,N_91,N_581);
or U1377 (N_1377,N_739,N_591);
or U1378 (N_1378,N_379,N_465);
or U1379 (N_1379,N_422,N_145);
and U1380 (N_1380,N_551,N_244);
and U1381 (N_1381,N_93,N_402);
or U1382 (N_1382,N_634,N_100);
nor U1383 (N_1383,N_77,N_442);
and U1384 (N_1384,N_120,N_598);
xor U1385 (N_1385,N_16,N_584);
nand U1386 (N_1386,N_645,N_313);
nor U1387 (N_1387,N_296,N_599);
or U1388 (N_1388,N_648,N_603);
nor U1389 (N_1389,N_127,N_130);
and U1390 (N_1390,N_604,N_612);
nor U1391 (N_1391,N_12,N_359);
and U1392 (N_1392,N_441,N_700);
nor U1393 (N_1393,N_294,N_446);
and U1394 (N_1394,N_742,N_175);
and U1395 (N_1395,N_455,N_681);
and U1396 (N_1396,N_537,N_356);
and U1397 (N_1397,N_365,N_371);
or U1398 (N_1398,N_269,N_118);
or U1399 (N_1399,N_141,N_696);
or U1400 (N_1400,N_124,N_88);
nor U1401 (N_1401,N_515,N_666);
nand U1402 (N_1402,N_165,N_678);
xnor U1403 (N_1403,N_118,N_437);
nor U1404 (N_1404,N_242,N_311);
xor U1405 (N_1405,N_272,N_285);
and U1406 (N_1406,N_201,N_573);
nor U1407 (N_1407,N_19,N_66);
nand U1408 (N_1408,N_496,N_102);
nand U1409 (N_1409,N_668,N_211);
xor U1410 (N_1410,N_165,N_101);
and U1411 (N_1411,N_746,N_509);
xor U1412 (N_1412,N_0,N_260);
or U1413 (N_1413,N_150,N_372);
nor U1414 (N_1414,N_351,N_28);
or U1415 (N_1415,N_593,N_236);
or U1416 (N_1416,N_16,N_50);
xor U1417 (N_1417,N_248,N_164);
nand U1418 (N_1418,N_116,N_405);
nor U1419 (N_1419,N_482,N_442);
nand U1420 (N_1420,N_649,N_255);
xnor U1421 (N_1421,N_678,N_381);
nor U1422 (N_1422,N_386,N_742);
and U1423 (N_1423,N_293,N_75);
nand U1424 (N_1424,N_415,N_659);
xor U1425 (N_1425,N_426,N_733);
or U1426 (N_1426,N_505,N_30);
and U1427 (N_1427,N_60,N_393);
xnor U1428 (N_1428,N_413,N_143);
or U1429 (N_1429,N_191,N_97);
nor U1430 (N_1430,N_635,N_172);
nand U1431 (N_1431,N_451,N_124);
nand U1432 (N_1432,N_616,N_540);
and U1433 (N_1433,N_182,N_85);
and U1434 (N_1434,N_87,N_330);
nand U1435 (N_1435,N_360,N_129);
xnor U1436 (N_1436,N_545,N_417);
or U1437 (N_1437,N_581,N_208);
and U1438 (N_1438,N_573,N_187);
and U1439 (N_1439,N_509,N_570);
and U1440 (N_1440,N_630,N_594);
nand U1441 (N_1441,N_72,N_298);
or U1442 (N_1442,N_290,N_102);
and U1443 (N_1443,N_671,N_202);
or U1444 (N_1444,N_531,N_221);
nor U1445 (N_1445,N_266,N_125);
nor U1446 (N_1446,N_93,N_642);
and U1447 (N_1447,N_267,N_226);
nand U1448 (N_1448,N_600,N_262);
nand U1449 (N_1449,N_401,N_1);
nand U1450 (N_1450,N_341,N_58);
nor U1451 (N_1451,N_562,N_570);
or U1452 (N_1452,N_116,N_9);
nor U1453 (N_1453,N_73,N_548);
xor U1454 (N_1454,N_164,N_323);
nor U1455 (N_1455,N_310,N_508);
nand U1456 (N_1456,N_260,N_592);
xor U1457 (N_1457,N_381,N_487);
xnor U1458 (N_1458,N_583,N_633);
xor U1459 (N_1459,N_378,N_434);
or U1460 (N_1460,N_123,N_602);
nand U1461 (N_1461,N_234,N_304);
nand U1462 (N_1462,N_262,N_340);
xor U1463 (N_1463,N_437,N_708);
nor U1464 (N_1464,N_744,N_458);
nor U1465 (N_1465,N_264,N_83);
nand U1466 (N_1466,N_4,N_308);
and U1467 (N_1467,N_438,N_152);
nand U1468 (N_1468,N_455,N_704);
and U1469 (N_1469,N_626,N_150);
and U1470 (N_1470,N_213,N_530);
or U1471 (N_1471,N_87,N_83);
or U1472 (N_1472,N_223,N_554);
nand U1473 (N_1473,N_672,N_281);
nor U1474 (N_1474,N_201,N_178);
nor U1475 (N_1475,N_65,N_672);
and U1476 (N_1476,N_421,N_93);
xor U1477 (N_1477,N_8,N_99);
nand U1478 (N_1478,N_490,N_152);
nand U1479 (N_1479,N_10,N_142);
and U1480 (N_1480,N_381,N_618);
nand U1481 (N_1481,N_208,N_436);
nor U1482 (N_1482,N_530,N_116);
nand U1483 (N_1483,N_558,N_189);
or U1484 (N_1484,N_291,N_323);
nand U1485 (N_1485,N_454,N_160);
nand U1486 (N_1486,N_592,N_89);
or U1487 (N_1487,N_180,N_618);
nand U1488 (N_1488,N_84,N_573);
nand U1489 (N_1489,N_492,N_124);
and U1490 (N_1490,N_173,N_610);
and U1491 (N_1491,N_705,N_408);
nand U1492 (N_1492,N_575,N_116);
nor U1493 (N_1493,N_460,N_75);
nand U1494 (N_1494,N_470,N_162);
and U1495 (N_1495,N_95,N_173);
or U1496 (N_1496,N_559,N_257);
nand U1497 (N_1497,N_192,N_519);
or U1498 (N_1498,N_435,N_642);
nand U1499 (N_1499,N_397,N_585);
nor U1500 (N_1500,N_1476,N_1395);
nand U1501 (N_1501,N_785,N_1268);
or U1502 (N_1502,N_762,N_1046);
or U1503 (N_1503,N_1221,N_1052);
and U1504 (N_1504,N_956,N_860);
and U1505 (N_1505,N_1400,N_1024);
nor U1506 (N_1506,N_1014,N_993);
nand U1507 (N_1507,N_1007,N_784);
and U1508 (N_1508,N_989,N_1102);
and U1509 (N_1509,N_1488,N_1027);
nor U1510 (N_1510,N_824,N_960);
xor U1511 (N_1511,N_1183,N_1434);
nor U1512 (N_1512,N_1460,N_1124);
and U1513 (N_1513,N_872,N_1015);
or U1514 (N_1514,N_958,N_1265);
and U1515 (N_1515,N_1304,N_1185);
or U1516 (N_1516,N_861,N_812);
nor U1517 (N_1517,N_1163,N_1390);
nand U1518 (N_1518,N_927,N_1469);
nor U1519 (N_1519,N_1241,N_1199);
nand U1520 (N_1520,N_985,N_1252);
nor U1521 (N_1521,N_754,N_1438);
nand U1522 (N_1522,N_909,N_1250);
nor U1523 (N_1523,N_1166,N_818);
or U1524 (N_1524,N_1466,N_929);
and U1525 (N_1525,N_1378,N_799);
and U1526 (N_1526,N_1055,N_976);
or U1527 (N_1527,N_1332,N_1448);
and U1528 (N_1528,N_780,N_966);
and U1529 (N_1529,N_1149,N_1232);
nor U1530 (N_1530,N_923,N_1405);
and U1531 (N_1531,N_1051,N_1272);
nor U1532 (N_1532,N_1396,N_1392);
or U1533 (N_1533,N_1213,N_804);
and U1534 (N_1534,N_1454,N_839);
and U1535 (N_1535,N_1230,N_850);
or U1536 (N_1536,N_1133,N_919);
or U1537 (N_1537,N_1417,N_1098);
xor U1538 (N_1538,N_880,N_1349);
and U1539 (N_1539,N_992,N_1299);
nor U1540 (N_1540,N_1427,N_891);
or U1541 (N_1541,N_1408,N_1115);
nor U1542 (N_1542,N_1394,N_1292);
nor U1543 (N_1543,N_1309,N_1442);
or U1544 (N_1544,N_805,N_1415);
nand U1545 (N_1545,N_937,N_939);
or U1546 (N_1546,N_1354,N_819);
nor U1547 (N_1547,N_1347,N_1082);
and U1548 (N_1548,N_1182,N_997);
nand U1549 (N_1549,N_874,N_761);
nand U1550 (N_1550,N_853,N_1203);
or U1551 (N_1551,N_836,N_1079);
or U1552 (N_1552,N_757,N_1487);
or U1553 (N_1553,N_1470,N_1491);
nor U1554 (N_1554,N_1087,N_1177);
nor U1555 (N_1555,N_1356,N_772);
or U1556 (N_1556,N_1063,N_1481);
or U1557 (N_1557,N_1219,N_935);
nand U1558 (N_1558,N_1225,N_962);
nor U1559 (N_1559,N_1353,N_1075);
or U1560 (N_1560,N_1017,N_803);
or U1561 (N_1561,N_1071,N_1237);
and U1562 (N_1562,N_791,N_1464);
and U1563 (N_1563,N_1239,N_1031);
nand U1564 (N_1564,N_917,N_986);
and U1565 (N_1565,N_933,N_924);
nor U1566 (N_1566,N_1385,N_938);
nand U1567 (N_1567,N_1473,N_1441);
nor U1568 (N_1568,N_1229,N_1382);
nor U1569 (N_1569,N_848,N_934);
nand U1570 (N_1570,N_1452,N_1251);
nor U1571 (N_1571,N_1422,N_1076);
and U1572 (N_1572,N_994,N_981);
nand U1573 (N_1573,N_867,N_1145);
nand U1574 (N_1574,N_967,N_904);
and U1575 (N_1575,N_1139,N_1041);
or U1576 (N_1576,N_920,N_1281);
and U1577 (N_1577,N_1215,N_1016);
and U1578 (N_1578,N_1044,N_1106);
and U1579 (N_1579,N_1423,N_1092);
nand U1580 (N_1580,N_1424,N_1123);
nand U1581 (N_1581,N_1257,N_1413);
or U1582 (N_1582,N_779,N_1165);
or U1583 (N_1583,N_863,N_1223);
and U1584 (N_1584,N_1181,N_877);
nor U1585 (N_1585,N_1338,N_817);
or U1586 (N_1586,N_1249,N_978);
nor U1587 (N_1587,N_903,N_1457);
nand U1588 (N_1588,N_1231,N_807);
nand U1589 (N_1589,N_1303,N_832);
or U1590 (N_1590,N_946,N_1243);
nand U1591 (N_1591,N_1032,N_795);
or U1592 (N_1592,N_782,N_1267);
nor U1593 (N_1593,N_844,N_996);
nor U1594 (N_1594,N_889,N_1381);
and U1595 (N_1595,N_755,N_1290);
or U1596 (N_1596,N_1371,N_1254);
or U1597 (N_1597,N_1446,N_1320);
xnor U1598 (N_1598,N_1253,N_887);
and U1599 (N_1599,N_1148,N_1263);
and U1600 (N_1600,N_1029,N_1323);
nand U1601 (N_1601,N_1198,N_1398);
nor U1602 (N_1602,N_1285,N_1426);
or U1603 (N_1603,N_1286,N_1449);
nor U1604 (N_1604,N_1121,N_856);
or U1605 (N_1605,N_1489,N_1137);
nand U1606 (N_1606,N_1386,N_1404);
nand U1607 (N_1607,N_1120,N_1058);
nor U1608 (N_1608,N_1194,N_1069);
xnor U1609 (N_1609,N_1066,N_1499);
and U1610 (N_1610,N_1479,N_1348);
or U1611 (N_1611,N_1244,N_928);
nand U1612 (N_1612,N_1428,N_1492);
xnor U1613 (N_1613,N_1370,N_1319);
or U1614 (N_1614,N_1196,N_810);
nor U1615 (N_1615,N_1172,N_1278);
or U1616 (N_1616,N_852,N_1377);
and U1617 (N_1617,N_1284,N_1274);
or U1618 (N_1618,N_1147,N_1212);
nor U1619 (N_1619,N_1184,N_1006);
nor U1620 (N_1620,N_949,N_1154);
nand U1621 (N_1621,N_1220,N_1195);
or U1622 (N_1622,N_1068,N_1022);
nor U1623 (N_1623,N_1380,N_1111);
or U1624 (N_1624,N_787,N_1401);
nor U1625 (N_1625,N_1372,N_1202);
nor U1626 (N_1626,N_921,N_881);
or U1627 (N_1627,N_814,N_1037);
and U1628 (N_1628,N_838,N_1351);
or U1629 (N_1629,N_1078,N_1062);
xnor U1630 (N_1630,N_1206,N_1170);
nand U1631 (N_1631,N_1297,N_1316);
or U1632 (N_1632,N_1205,N_947);
or U1633 (N_1633,N_875,N_940);
nor U1634 (N_1634,N_1156,N_1298);
nand U1635 (N_1635,N_847,N_783);
and U1636 (N_1636,N_1064,N_1486);
nand U1637 (N_1637,N_901,N_876);
nor U1638 (N_1638,N_1150,N_965);
nor U1639 (N_1639,N_769,N_1368);
nor U1640 (N_1640,N_879,N_1142);
or U1641 (N_1641,N_1009,N_882);
or U1642 (N_1642,N_1146,N_1339);
xor U1643 (N_1643,N_963,N_1050);
and U1644 (N_1644,N_1093,N_1141);
or U1645 (N_1645,N_1095,N_890);
and U1646 (N_1646,N_1236,N_1126);
and U1647 (N_1647,N_1471,N_1101);
nand U1648 (N_1648,N_760,N_1313);
nor U1649 (N_1649,N_945,N_1116);
nor U1650 (N_1650,N_764,N_931);
nor U1651 (N_1651,N_1393,N_1033);
nand U1652 (N_1652,N_991,N_767);
nor U1653 (N_1653,N_1402,N_1472);
nand U1654 (N_1654,N_1389,N_1451);
nor U1655 (N_1655,N_1119,N_1228);
nor U1656 (N_1656,N_833,N_977);
nand U1657 (N_1657,N_1025,N_987);
nor U1658 (N_1658,N_944,N_1409);
or U1659 (N_1659,N_1461,N_790);
and U1660 (N_1660,N_906,N_1334);
or U1661 (N_1661,N_1161,N_815);
nand U1662 (N_1662,N_1085,N_813);
nor U1663 (N_1663,N_883,N_980);
nor U1664 (N_1664,N_859,N_857);
xnor U1665 (N_1665,N_1099,N_1279);
nor U1666 (N_1666,N_1346,N_1056);
nor U1667 (N_1667,N_1342,N_913);
or U1668 (N_1668,N_825,N_1399);
nand U1669 (N_1669,N_884,N_802);
xnor U1670 (N_1670,N_763,N_1406);
and U1671 (N_1671,N_1084,N_1217);
nand U1672 (N_1672,N_1057,N_1131);
nand U1673 (N_1673,N_1384,N_816);
and U1674 (N_1674,N_1480,N_1010);
nand U1675 (N_1675,N_952,N_789);
nand U1676 (N_1676,N_1034,N_866);
nand U1677 (N_1677,N_1122,N_1197);
xnor U1678 (N_1678,N_1222,N_936);
or U1679 (N_1679,N_1047,N_1109);
nor U1680 (N_1680,N_752,N_900);
nand U1681 (N_1681,N_1162,N_1157);
nand U1682 (N_1682,N_1042,N_1416);
and U1683 (N_1683,N_855,N_1336);
and U1684 (N_1684,N_908,N_1361);
or U1685 (N_1685,N_1352,N_1322);
and U1686 (N_1686,N_1374,N_1048);
nand U1687 (N_1687,N_1360,N_1186);
nand U1688 (N_1688,N_1295,N_775);
or U1689 (N_1689,N_1397,N_1248);
and U1690 (N_1690,N_1328,N_1053);
nor U1691 (N_1691,N_1337,N_1288);
nor U1692 (N_1692,N_1435,N_1040);
or U1693 (N_1693,N_998,N_1373);
xor U1694 (N_1694,N_1324,N_1483);
nand U1695 (N_1695,N_1301,N_751);
and U1696 (N_1696,N_854,N_766);
nor U1697 (N_1697,N_1412,N_1496);
or U1698 (N_1698,N_905,N_1482);
nor U1699 (N_1699,N_862,N_864);
nand U1700 (N_1700,N_1114,N_1218);
nand U1701 (N_1701,N_1314,N_786);
or U1702 (N_1702,N_1282,N_873);
and U1703 (N_1703,N_1321,N_1362);
nor U1704 (N_1704,N_1180,N_1103);
nor U1705 (N_1705,N_1160,N_1383);
or U1706 (N_1706,N_897,N_1028);
or U1707 (N_1707,N_1012,N_1478);
or U1708 (N_1708,N_1468,N_840);
nor U1709 (N_1709,N_1127,N_1045);
nand U1710 (N_1710,N_1238,N_1072);
or U1711 (N_1711,N_801,N_914);
nand U1712 (N_1712,N_1011,N_955);
or U1713 (N_1713,N_1453,N_1269);
or U1714 (N_1714,N_796,N_1311);
and U1715 (N_1715,N_1358,N_831);
xnor U1716 (N_1716,N_1317,N_1411);
nor U1717 (N_1717,N_1467,N_1107);
and U1718 (N_1718,N_843,N_1113);
nor U1719 (N_1719,N_776,N_830);
or U1720 (N_1720,N_1443,N_1246);
nor U1721 (N_1721,N_1344,N_778);
and U1722 (N_1722,N_1117,N_1108);
or U1723 (N_1723,N_1333,N_926);
nand U1724 (N_1724,N_969,N_1159);
nand U1725 (N_1725,N_1445,N_888);
nor U1726 (N_1726,N_1305,N_1002);
nand U1727 (N_1727,N_1070,N_1280);
or U1728 (N_1728,N_1135,N_1129);
nand U1729 (N_1729,N_1379,N_979);
nor U1730 (N_1730,N_1327,N_1429);
and U1731 (N_1731,N_1433,N_1245);
or U1732 (N_1732,N_1271,N_1289);
nor U1733 (N_1733,N_842,N_1077);
and U1734 (N_1734,N_1112,N_1188);
and U1735 (N_1735,N_1214,N_1456);
nor U1736 (N_1736,N_851,N_1110);
nor U1737 (N_1737,N_1226,N_916);
nor U1738 (N_1738,N_918,N_1008);
nand U1739 (N_1739,N_1410,N_1357);
xor U1740 (N_1740,N_1340,N_1151);
nor U1741 (N_1741,N_971,N_1414);
or U1742 (N_1742,N_828,N_1256);
and U1743 (N_1743,N_878,N_1430);
nor U1744 (N_1744,N_1059,N_1345);
and U1745 (N_1745,N_1296,N_1233);
and U1746 (N_1746,N_1359,N_1211);
and U1747 (N_1747,N_788,N_858);
or U1748 (N_1748,N_1136,N_915);
nor U1749 (N_1749,N_1266,N_1407);
nand U1750 (N_1750,N_1096,N_988);
and U1751 (N_1751,N_972,N_777);
nand U1752 (N_1752,N_1094,N_1018);
and U1753 (N_1753,N_1049,N_1100);
and U1754 (N_1754,N_1283,N_765);
xnor U1755 (N_1755,N_845,N_1363);
nor U1756 (N_1756,N_1128,N_894);
nor U1757 (N_1757,N_1235,N_750);
and U1758 (N_1758,N_1440,N_1169);
nor U1759 (N_1759,N_1138,N_1432);
and U1760 (N_1760,N_1447,N_1287);
nand U1761 (N_1761,N_942,N_1485);
nand U1762 (N_1762,N_1270,N_1125);
nand U1763 (N_1763,N_1302,N_1097);
or U1764 (N_1764,N_1291,N_1164);
nor U1765 (N_1765,N_792,N_1403);
nor U1766 (N_1766,N_954,N_1001);
or U1767 (N_1767,N_1036,N_1021);
and U1768 (N_1768,N_964,N_984);
nand U1769 (N_1769,N_1167,N_1081);
or U1770 (N_1770,N_1105,N_1247);
nand U1771 (N_1771,N_822,N_975);
or U1772 (N_1772,N_1493,N_1365);
nor U1773 (N_1773,N_898,N_841);
nand U1774 (N_1774,N_1325,N_1090);
or U1775 (N_1775,N_1035,N_794);
xnor U1776 (N_1776,N_1061,N_1255);
nand U1777 (N_1777,N_768,N_871);
and U1778 (N_1778,N_1437,N_1003);
xor U1779 (N_1779,N_1350,N_773);
nor U1780 (N_1780,N_865,N_990);
and U1781 (N_1781,N_1300,N_1065);
nor U1782 (N_1782,N_1306,N_800);
or U1783 (N_1783,N_911,N_1312);
and U1784 (N_1784,N_892,N_1355);
or U1785 (N_1785,N_1477,N_793);
or U1786 (N_1786,N_1495,N_770);
nand U1787 (N_1787,N_1143,N_1369);
or U1788 (N_1788,N_1039,N_753);
and U1789 (N_1789,N_771,N_869);
and U1790 (N_1790,N_1174,N_899);
or U1791 (N_1791,N_1375,N_756);
and U1792 (N_1792,N_959,N_1260);
or U1793 (N_1793,N_837,N_1227);
and U1794 (N_1794,N_1019,N_1294);
xor U1795 (N_1795,N_781,N_1153);
and U1796 (N_1796,N_820,N_982);
nand U1797 (N_1797,N_1155,N_1026);
and U1798 (N_1798,N_1086,N_902);
and U1799 (N_1799,N_1341,N_1074);
xor U1800 (N_1800,N_953,N_907);
nor U1801 (N_1801,N_1458,N_1210);
or U1802 (N_1802,N_983,N_1091);
nand U1803 (N_1803,N_1152,N_1073);
nor U1804 (N_1804,N_1130,N_941);
nand U1805 (N_1805,N_948,N_1420);
nand U1806 (N_1806,N_826,N_834);
nand U1807 (N_1807,N_973,N_974);
and U1808 (N_1808,N_1030,N_1261);
xnor U1809 (N_1809,N_1475,N_1388);
xor U1810 (N_1810,N_1308,N_1176);
or U1811 (N_1811,N_1104,N_895);
and U1812 (N_1812,N_1330,N_1000);
or U1813 (N_1813,N_1175,N_1439);
nand U1814 (N_1814,N_1455,N_1273);
nand U1815 (N_1815,N_932,N_1436);
or U1816 (N_1816,N_1173,N_1418);
or U1817 (N_1817,N_1387,N_995);
and U1818 (N_1818,N_1240,N_1140);
or U1819 (N_1819,N_1179,N_1208);
nor U1820 (N_1820,N_1277,N_1171);
xnor U1821 (N_1821,N_759,N_870);
nor U1822 (N_1822,N_930,N_1310);
nand U1823 (N_1823,N_1275,N_922);
nor U1824 (N_1824,N_1315,N_829);
and U1825 (N_1825,N_811,N_1067);
or U1826 (N_1826,N_1262,N_910);
nor U1827 (N_1827,N_970,N_1224);
or U1828 (N_1828,N_1005,N_1462);
and U1829 (N_1829,N_1118,N_1158);
nor U1830 (N_1830,N_1080,N_1004);
and U1831 (N_1831,N_1259,N_1193);
nand U1832 (N_1832,N_1421,N_1307);
or U1833 (N_1833,N_1463,N_1060);
and U1834 (N_1834,N_1258,N_1023);
nand U1835 (N_1835,N_1490,N_1331);
nor U1836 (N_1836,N_1088,N_849);
and U1837 (N_1837,N_999,N_806);
or U1838 (N_1838,N_951,N_1234);
or U1839 (N_1839,N_912,N_885);
or U1840 (N_1840,N_1465,N_797);
and U1841 (N_1841,N_1054,N_758);
or U1842 (N_1842,N_1089,N_1391);
or U1843 (N_1843,N_1200,N_950);
and U1844 (N_1844,N_1144,N_1459);
nor U1845 (N_1845,N_896,N_1450);
or U1846 (N_1846,N_1020,N_1326);
nor U1847 (N_1847,N_823,N_968);
nor U1848 (N_1848,N_1376,N_925);
nand U1849 (N_1849,N_1329,N_809);
or U1850 (N_1850,N_1364,N_1335);
or U1851 (N_1851,N_1192,N_1083);
nor U1852 (N_1852,N_774,N_1431);
nand U1853 (N_1853,N_1264,N_1201);
nand U1854 (N_1854,N_1216,N_846);
nor U1855 (N_1855,N_886,N_1276);
and U1856 (N_1856,N_1187,N_1038);
or U1857 (N_1857,N_893,N_1366);
and U1858 (N_1858,N_1190,N_1343);
nor U1859 (N_1859,N_1043,N_1191);
or U1860 (N_1860,N_1484,N_1207);
nand U1861 (N_1861,N_1497,N_835);
nand U1862 (N_1862,N_1189,N_821);
and U1863 (N_1863,N_1178,N_1419);
nor U1864 (N_1864,N_1494,N_1132);
nor U1865 (N_1865,N_1204,N_1474);
or U1866 (N_1866,N_1293,N_1318);
nor U1867 (N_1867,N_1242,N_808);
nand U1868 (N_1868,N_943,N_1013);
xnor U1869 (N_1869,N_1209,N_1498);
nand U1870 (N_1870,N_798,N_961);
nand U1871 (N_1871,N_868,N_1425);
nor U1872 (N_1872,N_1168,N_827);
xnor U1873 (N_1873,N_1367,N_1444);
nand U1874 (N_1874,N_957,N_1134);
or U1875 (N_1875,N_1158,N_849);
nor U1876 (N_1876,N_1022,N_940);
and U1877 (N_1877,N_791,N_1399);
nand U1878 (N_1878,N_883,N_1331);
nor U1879 (N_1879,N_1317,N_771);
or U1880 (N_1880,N_896,N_1446);
nand U1881 (N_1881,N_1346,N_775);
or U1882 (N_1882,N_1060,N_1054);
nor U1883 (N_1883,N_1001,N_1487);
nor U1884 (N_1884,N_1092,N_1216);
nor U1885 (N_1885,N_803,N_817);
xnor U1886 (N_1886,N_1352,N_887);
nor U1887 (N_1887,N_1168,N_987);
xor U1888 (N_1888,N_860,N_1345);
xor U1889 (N_1889,N_859,N_1318);
nor U1890 (N_1890,N_773,N_826);
and U1891 (N_1891,N_779,N_820);
xnor U1892 (N_1892,N_1009,N_894);
or U1893 (N_1893,N_1204,N_1002);
or U1894 (N_1894,N_1426,N_1023);
or U1895 (N_1895,N_757,N_826);
nor U1896 (N_1896,N_1292,N_1467);
and U1897 (N_1897,N_1126,N_1028);
or U1898 (N_1898,N_945,N_923);
xnor U1899 (N_1899,N_1043,N_1068);
or U1900 (N_1900,N_1338,N_911);
and U1901 (N_1901,N_1048,N_1261);
nand U1902 (N_1902,N_1434,N_1150);
and U1903 (N_1903,N_1248,N_1247);
nand U1904 (N_1904,N_887,N_846);
or U1905 (N_1905,N_1136,N_1489);
or U1906 (N_1906,N_950,N_883);
nor U1907 (N_1907,N_1460,N_1050);
or U1908 (N_1908,N_847,N_1432);
or U1909 (N_1909,N_1177,N_900);
nor U1910 (N_1910,N_1115,N_1055);
nand U1911 (N_1911,N_807,N_910);
nand U1912 (N_1912,N_1072,N_1282);
nand U1913 (N_1913,N_1246,N_1047);
nand U1914 (N_1914,N_978,N_1096);
nor U1915 (N_1915,N_856,N_1403);
nand U1916 (N_1916,N_1456,N_1121);
or U1917 (N_1917,N_1299,N_771);
nor U1918 (N_1918,N_895,N_970);
or U1919 (N_1919,N_1093,N_1360);
and U1920 (N_1920,N_1391,N_800);
or U1921 (N_1921,N_1291,N_1375);
or U1922 (N_1922,N_797,N_1146);
nand U1923 (N_1923,N_816,N_1048);
nor U1924 (N_1924,N_1412,N_1165);
or U1925 (N_1925,N_1101,N_866);
or U1926 (N_1926,N_902,N_1370);
nor U1927 (N_1927,N_1475,N_1037);
nand U1928 (N_1928,N_1137,N_927);
or U1929 (N_1929,N_1021,N_937);
nand U1930 (N_1930,N_994,N_1141);
xor U1931 (N_1931,N_1366,N_1199);
nand U1932 (N_1932,N_1089,N_1116);
or U1933 (N_1933,N_1271,N_995);
or U1934 (N_1934,N_849,N_1352);
xnor U1935 (N_1935,N_770,N_791);
xor U1936 (N_1936,N_1450,N_918);
nand U1937 (N_1937,N_1331,N_782);
nor U1938 (N_1938,N_1259,N_1278);
nand U1939 (N_1939,N_1182,N_1311);
or U1940 (N_1940,N_801,N_1247);
or U1941 (N_1941,N_1088,N_1008);
or U1942 (N_1942,N_1208,N_1032);
nand U1943 (N_1943,N_1027,N_1106);
nand U1944 (N_1944,N_1140,N_840);
or U1945 (N_1945,N_1035,N_1450);
and U1946 (N_1946,N_1261,N_1110);
nor U1947 (N_1947,N_1328,N_1316);
and U1948 (N_1948,N_853,N_941);
nor U1949 (N_1949,N_837,N_1369);
or U1950 (N_1950,N_915,N_1049);
nand U1951 (N_1951,N_1014,N_1470);
or U1952 (N_1952,N_1183,N_843);
or U1953 (N_1953,N_778,N_1072);
nand U1954 (N_1954,N_1220,N_846);
nor U1955 (N_1955,N_785,N_860);
nor U1956 (N_1956,N_1011,N_1293);
nand U1957 (N_1957,N_1396,N_963);
nand U1958 (N_1958,N_790,N_1211);
or U1959 (N_1959,N_957,N_1251);
nor U1960 (N_1960,N_1183,N_1483);
or U1961 (N_1961,N_1011,N_1054);
nor U1962 (N_1962,N_893,N_1214);
nor U1963 (N_1963,N_902,N_963);
and U1964 (N_1964,N_1221,N_1479);
xnor U1965 (N_1965,N_1067,N_1206);
or U1966 (N_1966,N_857,N_1167);
and U1967 (N_1967,N_1278,N_786);
nand U1968 (N_1968,N_785,N_798);
or U1969 (N_1969,N_887,N_928);
and U1970 (N_1970,N_1216,N_1109);
nand U1971 (N_1971,N_1451,N_1488);
or U1972 (N_1972,N_1008,N_776);
or U1973 (N_1973,N_1213,N_796);
xor U1974 (N_1974,N_1278,N_818);
and U1975 (N_1975,N_1432,N_940);
and U1976 (N_1976,N_782,N_974);
or U1977 (N_1977,N_1264,N_1328);
and U1978 (N_1978,N_785,N_1138);
xor U1979 (N_1979,N_1270,N_888);
nand U1980 (N_1980,N_1033,N_1291);
nor U1981 (N_1981,N_1314,N_1492);
or U1982 (N_1982,N_861,N_952);
nand U1983 (N_1983,N_971,N_1227);
xnor U1984 (N_1984,N_980,N_846);
and U1985 (N_1985,N_1048,N_1044);
xnor U1986 (N_1986,N_780,N_1017);
xnor U1987 (N_1987,N_1415,N_800);
nor U1988 (N_1988,N_1253,N_1461);
xor U1989 (N_1989,N_1387,N_850);
and U1990 (N_1990,N_884,N_909);
and U1991 (N_1991,N_911,N_1224);
or U1992 (N_1992,N_754,N_1459);
nor U1993 (N_1993,N_1172,N_1081);
nand U1994 (N_1994,N_1179,N_804);
nand U1995 (N_1995,N_916,N_1239);
and U1996 (N_1996,N_1243,N_1488);
nand U1997 (N_1997,N_1395,N_1188);
or U1998 (N_1998,N_1423,N_1123);
and U1999 (N_1999,N_1095,N_1446);
nor U2000 (N_2000,N_987,N_1479);
or U2001 (N_2001,N_1097,N_895);
nand U2002 (N_2002,N_969,N_1241);
nor U2003 (N_2003,N_1306,N_1201);
or U2004 (N_2004,N_761,N_943);
and U2005 (N_2005,N_910,N_1400);
nand U2006 (N_2006,N_1144,N_799);
and U2007 (N_2007,N_1435,N_879);
nor U2008 (N_2008,N_812,N_1431);
and U2009 (N_2009,N_1368,N_1337);
nand U2010 (N_2010,N_1455,N_859);
or U2011 (N_2011,N_1268,N_952);
or U2012 (N_2012,N_973,N_785);
nor U2013 (N_2013,N_765,N_1417);
or U2014 (N_2014,N_898,N_1224);
and U2015 (N_2015,N_1253,N_768);
xor U2016 (N_2016,N_1085,N_809);
or U2017 (N_2017,N_1309,N_900);
xor U2018 (N_2018,N_992,N_1134);
nand U2019 (N_2019,N_1382,N_1492);
and U2020 (N_2020,N_1047,N_1057);
nand U2021 (N_2021,N_1196,N_1346);
and U2022 (N_2022,N_1382,N_938);
and U2023 (N_2023,N_799,N_1450);
and U2024 (N_2024,N_764,N_1498);
and U2025 (N_2025,N_1281,N_1417);
nor U2026 (N_2026,N_879,N_1299);
nand U2027 (N_2027,N_1271,N_826);
xor U2028 (N_2028,N_1061,N_1405);
or U2029 (N_2029,N_1162,N_924);
or U2030 (N_2030,N_894,N_964);
xnor U2031 (N_2031,N_835,N_898);
or U2032 (N_2032,N_945,N_1345);
or U2033 (N_2033,N_824,N_940);
nor U2034 (N_2034,N_1338,N_1192);
xnor U2035 (N_2035,N_1366,N_934);
and U2036 (N_2036,N_1453,N_1152);
nand U2037 (N_2037,N_1320,N_1486);
nand U2038 (N_2038,N_1097,N_1429);
or U2039 (N_2039,N_1194,N_1452);
xor U2040 (N_2040,N_1203,N_1244);
nand U2041 (N_2041,N_933,N_805);
nor U2042 (N_2042,N_876,N_763);
nand U2043 (N_2043,N_1110,N_1432);
nand U2044 (N_2044,N_1439,N_894);
nor U2045 (N_2045,N_955,N_897);
and U2046 (N_2046,N_1258,N_921);
nand U2047 (N_2047,N_835,N_1049);
nor U2048 (N_2048,N_777,N_823);
nand U2049 (N_2049,N_1041,N_1430);
nand U2050 (N_2050,N_1494,N_1423);
nor U2051 (N_2051,N_1092,N_906);
nand U2052 (N_2052,N_1467,N_950);
xor U2053 (N_2053,N_1067,N_818);
or U2054 (N_2054,N_1094,N_1109);
and U2055 (N_2055,N_1465,N_981);
and U2056 (N_2056,N_1318,N_1004);
nor U2057 (N_2057,N_1086,N_1173);
xor U2058 (N_2058,N_1006,N_878);
nand U2059 (N_2059,N_1284,N_1086);
or U2060 (N_2060,N_983,N_1428);
nand U2061 (N_2061,N_823,N_931);
nor U2062 (N_2062,N_846,N_1043);
and U2063 (N_2063,N_1482,N_1241);
nor U2064 (N_2064,N_1265,N_1249);
nor U2065 (N_2065,N_848,N_1352);
or U2066 (N_2066,N_1497,N_993);
or U2067 (N_2067,N_1225,N_952);
nand U2068 (N_2068,N_1335,N_1404);
nand U2069 (N_2069,N_1071,N_1334);
and U2070 (N_2070,N_1394,N_970);
or U2071 (N_2071,N_1022,N_1263);
nor U2072 (N_2072,N_814,N_990);
and U2073 (N_2073,N_1462,N_1224);
and U2074 (N_2074,N_1155,N_1477);
or U2075 (N_2075,N_1101,N_1303);
and U2076 (N_2076,N_1386,N_1400);
nor U2077 (N_2077,N_790,N_880);
and U2078 (N_2078,N_773,N_1444);
nor U2079 (N_2079,N_929,N_1059);
nor U2080 (N_2080,N_1098,N_1306);
nand U2081 (N_2081,N_1195,N_1475);
and U2082 (N_2082,N_1035,N_826);
and U2083 (N_2083,N_778,N_1408);
xnor U2084 (N_2084,N_1096,N_1201);
nand U2085 (N_2085,N_773,N_1122);
nor U2086 (N_2086,N_912,N_1131);
xor U2087 (N_2087,N_775,N_824);
nor U2088 (N_2088,N_1465,N_1169);
nor U2089 (N_2089,N_1294,N_977);
nand U2090 (N_2090,N_1288,N_1134);
nand U2091 (N_2091,N_970,N_1341);
and U2092 (N_2092,N_1305,N_1302);
and U2093 (N_2093,N_1493,N_1337);
nand U2094 (N_2094,N_1440,N_773);
nor U2095 (N_2095,N_1107,N_1019);
and U2096 (N_2096,N_875,N_930);
or U2097 (N_2097,N_1155,N_1405);
nand U2098 (N_2098,N_1012,N_1364);
or U2099 (N_2099,N_1276,N_884);
or U2100 (N_2100,N_1028,N_1294);
and U2101 (N_2101,N_1196,N_999);
nor U2102 (N_2102,N_1405,N_1136);
or U2103 (N_2103,N_1171,N_783);
xnor U2104 (N_2104,N_1402,N_1211);
nand U2105 (N_2105,N_1244,N_1322);
and U2106 (N_2106,N_1478,N_893);
nor U2107 (N_2107,N_1033,N_1188);
or U2108 (N_2108,N_1246,N_769);
or U2109 (N_2109,N_986,N_1003);
nand U2110 (N_2110,N_875,N_791);
nor U2111 (N_2111,N_1204,N_828);
xor U2112 (N_2112,N_1441,N_1238);
nand U2113 (N_2113,N_874,N_1443);
or U2114 (N_2114,N_929,N_1242);
nor U2115 (N_2115,N_802,N_1043);
and U2116 (N_2116,N_1026,N_1438);
nor U2117 (N_2117,N_1128,N_1354);
nand U2118 (N_2118,N_1456,N_1486);
or U2119 (N_2119,N_1489,N_1111);
xor U2120 (N_2120,N_1079,N_1302);
or U2121 (N_2121,N_879,N_779);
nand U2122 (N_2122,N_884,N_1132);
and U2123 (N_2123,N_1109,N_1474);
or U2124 (N_2124,N_852,N_911);
or U2125 (N_2125,N_797,N_1367);
and U2126 (N_2126,N_1485,N_1389);
and U2127 (N_2127,N_770,N_1471);
nand U2128 (N_2128,N_1422,N_921);
or U2129 (N_2129,N_849,N_1429);
and U2130 (N_2130,N_1247,N_1222);
nand U2131 (N_2131,N_988,N_1485);
xnor U2132 (N_2132,N_920,N_1380);
nor U2133 (N_2133,N_1381,N_1287);
nand U2134 (N_2134,N_1407,N_1222);
or U2135 (N_2135,N_1323,N_824);
xor U2136 (N_2136,N_1093,N_1353);
and U2137 (N_2137,N_1210,N_1151);
and U2138 (N_2138,N_1152,N_1169);
nand U2139 (N_2139,N_1337,N_1013);
or U2140 (N_2140,N_804,N_1096);
xnor U2141 (N_2141,N_1183,N_1085);
nand U2142 (N_2142,N_1413,N_1161);
or U2143 (N_2143,N_753,N_1422);
or U2144 (N_2144,N_1445,N_1349);
nand U2145 (N_2145,N_1292,N_1315);
xor U2146 (N_2146,N_1308,N_1137);
nand U2147 (N_2147,N_1080,N_778);
xor U2148 (N_2148,N_1474,N_1382);
nor U2149 (N_2149,N_1497,N_1365);
nor U2150 (N_2150,N_1082,N_912);
nor U2151 (N_2151,N_888,N_782);
and U2152 (N_2152,N_1120,N_1170);
xor U2153 (N_2153,N_1407,N_847);
nand U2154 (N_2154,N_866,N_1118);
nand U2155 (N_2155,N_1486,N_886);
nand U2156 (N_2156,N_1043,N_1021);
nand U2157 (N_2157,N_1004,N_900);
nand U2158 (N_2158,N_863,N_1327);
or U2159 (N_2159,N_1332,N_1247);
nand U2160 (N_2160,N_1185,N_1441);
nor U2161 (N_2161,N_795,N_1317);
nand U2162 (N_2162,N_1018,N_778);
and U2163 (N_2163,N_1485,N_920);
and U2164 (N_2164,N_1077,N_1042);
and U2165 (N_2165,N_826,N_983);
xor U2166 (N_2166,N_1353,N_1244);
nand U2167 (N_2167,N_1460,N_813);
or U2168 (N_2168,N_1043,N_1454);
nor U2169 (N_2169,N_863,N_1145);
nand U2170 (N_2170,N_1384,N_1432);
nor U2171 (N_2171,N_955,N_766);
nand U2172 (N_2172,N_1009,N_1026);
or U2173 (N_2173,N_803,N_809);
nor U2174 (N_2174,N_1311,N_1415);
or U2175 (N_2175,N_1332,N_1345);
xor U2176 (N_2176,N_1193,N_1284);
or U2177 (N_2177,N_1232,N_1418);
nor U2178 (N_2178,N_1025,N_1118);
and U2179 (N_2179,N_823,N_1333);
nor U2180 (N_2180,N_1135,N_1189);
or U2181 (N_2181,N_1194,N_1170);
and U2182 (N_2182,N_1452,N_945);
or U2183 (N_2183,N_1344,N_1276);
and U2184 (N_2184,N_857,N_1080);
nor U2185 (N_2185,N_831,N_1127);
nand U2186 (N_2186,N_1264,N_1097);
nand U2187 (N_2187,N_1193,N_1139);
or U2188 (N_2188,N_1466,N_891);
nand U2189 (N_2189,N_1401,N_1109);
or U2190 (N_2190,N_890,N_884);
nand U2191 (N_2191,N_1065,N_1256);
nand U2192 (N_2192,N_1486,N_769);
nor U2193 (N_2193,N_1444,N_1158);
nor U2194 (N_2194,N_996,N_1106);
nor U2195 (N_2195,N_1300,N_1369);
xnor U2196 (N_2196,N_1089,N_1058);
and U2197 (N_2197,N_1218,N_752);
nor U2198 (N_2198,N_1238,N_1135);
and U2199 (N_2199,N_1234,N_1210);
nand U2200 (N_2200,N_842,N_776);
nand U2201 (N_2201,N_1286,N_1443);
or U2202 (N_2202,N_1215,N_782);
xnor U2203 (N_2203,N_1488,N_1468);
nor U2204 (N_2204,N_1107,N_1062);
or U2205 (N_2205,N_1025,N_988);
nand U2206 (N_2206,N_1209,N_1346);
nor U2207 (N_2207,N_1283,N_1389);
or U2208 (N_2208,N_1030,N_888);
or U2209 (N_2209,N_1312,N_949);
nor U2210 (N_2210,N_1372,N_766);
nand U2211 (N_2211,N_1388,N_930);
xnor U2212 (N_2212,N_1033,N_807);
and U2213 (N_2213,N_1394,N_868);
nor U2214 (N_2214,N_1324,N_893);
nand U2215 (N_2215,N_1020,N_939);
nand U2216 (N_2216,N_1146,N_1429);
nor U2217 (N_2217,N_1478,N_1248);
xor U2218 (N_2218,N_1129,N_1286);
and U2219 (N_2219,N_1002,N_1159);
or U2220 (N_2220,N_1169,N_1407);
nor U2221 (N_2221,N_1027,N_1129);
or U2222 (N_2222,N_1433,N_1244);
or U2223 (N_2223,N_1253,N_1489);
nand U2224 (N_2224,N_876,N_1435);
xnor U2225 (N_2225,N_755,N_1395);
or U2226 (N_2226,N_1270,N_1327);
or U2227 (N_2227,N_1288,N_1479);
nand U2228 (N_2228,N_1076,N_1487);
nor U2229 (N_2229,N_990,N_886);
nand U2230 (N_2230,N_1046,N_792);
and U2231 (N_2231,N_1223,N_1288);
xor U2232 (N_2232,N_1341,N_1292);
nor U2233 (N_2233,N_923,N_1286);
nor U2234 (N_2234,N_1332,N_1310);
or U2235 (N_2235,N_1477,N_1364);
and U2236 (N_2236,N_1411,N_1089);
nor U2237 (N_2237,N_953,N_916);
and U2238 (N_2238,N_907,N_945);
or U2239 (N_2239,N_1497,N_1477);
or U2240 (N_2240,N_944,N_1443);
or U2241 (N_2241,N_971,N_904);
nor U2242 (N_2242,N_1195,N_751);
nand U2243 (N_2243,N_1455,N_1476);
and U2244 (N_2244,N_1105,N_793);
nand U2245 (N_2245,N_1478,N_753);
nand U2246 (N_2246,N_963,N_1230);
or U2247 (N_2247,N_1099,N_795);
or U2248 (N_2248,N_1160,N_954);
or U2249 (N_2249,N_892,N_816);
and U2250 (N_2250,N_1955,N_2022);
nand U2251 (N_2251,N_1660,N_1783);
nor U2252 (N_2252,N_1735,N_1877);
and U2253 (N_2253,N_1593,N_2003);
nor U2254 (N_2254,N_1915,N_1539);
nor U2255 (N_2255,N_1981,N_1625);
nand U2256 (N_2256,N_1702,N_1950);
or U2257 (N_2257,N_2121,N_2074);
and U2258 (N_2258,N_1816,N_1703);
and U2259 (N_2259,N_1532,N_1841);
and U2260 (N_2260,N_2115,N_2164);
nand U2261 (N_2261,N_2112,N_2055);
nor U2262 (N_2262,N_2075,N_2067);
nand U2263 (N_2263,N_2197,N_1884);
nor U2264 (N_2264,N_1600,N_1644);
nor U2265 (N_2265,N_1529,N_1568);
nand U2266 (N_2266,N_1585,N_2206);
or U2267 (N_2267,N_2072,N_1807);
or U2268 (N_2268,N_2047,N_1962);
nor U2269 (N_2269,N_2013,N_1558);
or U2270 (N_2270,N_2183,N_2227);
or U2271 (N_2271,N_2059,N_1795);
or U2272 (N_2272,N_1716,N_1998);
nor U2273 (N_2273,N_1595,N_2123);
nand U2274 (N_2274,N_1867,N_1746);
or U2275 (N_2275,N_1919,N_1829);
xor U2276 (N_2276,N_2160,N_1898);
and U2277 (N_2277,N_1632,N_2133);
nor U2278 (N_2278,N_1990,N_1775);
or U2279 (N_2279,N_1963,N_2130);
and U2280 (N_2280,N_1940,N_1588);
nor U2281 (N_2281,N_1861,N_1742);
xor U2282 (N_2282,N_1538,N_1824);
or U2283 (N_2283,N_1774,N_1821);
nand U2284 (N_2284,N_1996,N_1729);
nor U2285 (N_2285,N_2126,N_2065);
or U2286 (N_2286,N_2118,N_1573);
nor U2287 (N_2287,N_1779,N_2032);
nand U2288 (N_2288,N_1823,N_1960);
or U2289 (N_2289,N_1605,N_2114);
nand U2290 (N_2290,N_1606,N_2180);
and U2291 (N_2291,N_2066,N_1806);
and U2292 (N_2292,N_1750,N_1731);
nand U2293 (N_2293,N_1518,N_2189);
and U2294 (N_2294,N_1516,N_2037);
and U2295 (N_2295,N_1914,N_2246);
nor U2296 (N_2296,N_2007,N_2150);
nand U2297 (N_2297,N_2175,N_1843);
nor U2298 (N_2298,N_1946,N_1726);
nor U2299 (N_2299,N_1834,N_2058);
nor U2300 (N_2300,N_1511,N_2000);
or U2301 (N_2301,N_2182,N_1679);
and U2302 (N_2302,N_1601,N_1769);
nor U2303 (N_2303,N_1790,N_2129);
nand U2304 (N_2304,N_2196,N_1965);
xnor U2305 (N_2305,N_1688,N_2177);
nand U2306 (N_2306,N_1840,N_1700);
nor U2307 (N_2307,N_1924,N_2042);
nand U2308 (N_2308,N_2033,N_1740);
or U2309 (N_2309,N_1942,N_1904);
or U2310 (N_2310,N_1530,N_1671);
and U2311 (N_2311,N_2139,N_1853);
or U2312 (N_2312,N_2140,N_1669);
nor U2313 (N_2313,N_1611,N_1762);
and U2314 (N_2314,N_1552,N_1693);
nand U2315 (N_2315,N_1627,N_2245);
xor U2316 (N_2316,N_1613,N_2169);
and U2317 (N_2317,N_1901,N_2117);
or U2318 (N_2318,N_2024,N_1794);
or U2319 (N_2319,N_2184,N_1744);
or U2320 (N_2320,N_2199,N_2011);
nor U2321 (N_2321,N_1564,N_1948);
or U2322 (N_2322,N_2030,N_1674);
nor U2323 (N_2323,N_1888,N_1586);
nand U2324 (N_2324,N_1665,N_1859);
and U2325 (N_2325,N_1912,N_2028);
nand U2326 (N_2326,N_1567,N_1999);
and U2327 (N_2327,N_1819,N_2219);
nand U2328 (N_2328,N_2190,N_1645);
nand U2329 (N_2329,N_2050,N_2009);
and U2330 (N_2330,N_1850,N_1690);
and U2331 (N_2331,N_2104,N_2076);
or U2332 (N_2332,N_2052,N_1730);
nand U2333 (N_2333,N_2044,N_2156);
nor U2334 (N_2334,N_1534,N_1609);
or U2335 (N_2335,N_1577,N_1933);
or U2336 (N_2336,N_1725,N_2127);
and U2337 (N_2337,N_1865,N_2023);
or U2338 (N_2338,N_2069,N_1533);
and U2339 (N_2339,N_2012,N_1637);
nand U2340 (N_2340,N_2103,N_1974);
and U2341 (N_2341,N_2064,N_1624);
nor U2342 (N_2342,N_1891,N_1868);
xnor U2343 (N_2343,N_2077,N_1984);
nor U2344 (N_2344,N_1696,N_1808);
and U2345 (N_2345,N_1668,N_2082);
or U2346 (N_2346,N_1612,N_1559);
or U2347 (N_2347,N_2017,N_1755);
and U2348 (N_2348,N_1957,N_2101);
xnor U2349 (N_2349,N_2040,N_2053);
xor U2350 (N_2350,N_2031,N_1785);
or U2351 (N_2351,N_1581,N_1563);
nor U2352 (N_2352,N_2242,N_1846);
nor U2353 (N_2353,N_1712,N_2014);
nor U2354 (N_2354,N_2231,N_1952);
and U2355 (N_2355,N_1592,N_1943);
nor U2356 (N_2356,N_1681,N_1907);
and U2357 (N_2357,N_2135,N_1886);
nor U2358 (N_2358,N_1995,N_1972);
and U2359 (N_2359,N_1780,N_2084);
or U2360 (N_2360,N_1699,N_1708);
nand U2361 (N_2361,N_2217,N_1911);
and U2362 (N_2362,N_1504,N_1903);
or U2363 (N_2363,N_1797,N_1992);
xor U2364 (N_2364,N_1749,N_2096);
nor U2365 (N_2365,N_1626,N_1872);
and U2366 (N_2366,N_1923,N_1607);
nor U2367 (N_2367,N_1721,N_1893);
xor U2368 (N_2368,N_1747,N_1964);
nor U2369 (N_2369,N_1856,N_2211);
and U2370 (N_2370,N_2005,N_2157);
and U2371 (N_2371,N_2098,N_1851);
and U2372 (N_2372,N_1500,N_1618);
or U2373 (N_2373,N_1845,N_1709);
and U2374 (N_2374,N_1805,N_1959);
nand U2375 (N_2375,N_1881,N_2167);
or U2376 (N_2376,N_1522,N_1766);
nand U2377 (N_2377,N_1895,N_1835);
nor U2378 (N_2378,N_1936,N_2116);
or U2379 (N_2379,N_1727,N_1953);
and U2380 (N_2380,N_1608,N_1773);
nor U2381 (N_2381,N_2068,N_2155);
or U2382 (N_2382,N_1728,N_1997);
or U2383 (N_2383,N_1734,N_1935);
nor U2384 (N_2384,N_1815,N_1880);
nand U2385 (N_2385,N_1741,N_1509);
or U2386 (N_2386,N_1582,N_1908);
and U2387 (N_2387,N_2201,N_1528);
xnor U2388 (N_2388,N_1890,N_1630);
or U2389 (N_2389,N_1926,N_1689);
or U2390 (N_2390,N_1883,N_1958);
nand U2391 (N_2391,N_2240,N_1508);
xnor U2392 (N_2392,N_2236,N_2146);
or U2393 (N_2393,N_2132,N_1673);
nor U2394 (N_2394,N_2095,N_1574);
or U2395 (N_2395,N_1858,N_1598);
nor U2396 (N_2396,N_2202,N_1547);
nor U2397 (N_2397,N_2234,N_1772);
and U2398 (N_2398,N_1930,N_1869);
or U2399 (N_2399,N_1803,N_1782);
or U2400 (N_2400,N_2247,N_1855);
xnor U2401 (N_2401,N_1575,N_2224);
nor U2402 (N_2402,N_1555,N_1658);
or U2403 (N_2403,N_2086,N_1583);
nand U2404 (N_2404,N_2147,N_1651);
nor U2405 (N_2405,N_1542,N_1887);
nand U2406 (N_2406,N_1871,N_1659);
and U2407 (N_2407,N_2036,N_1704);
and U2408 (N_2408,N_2089,N_2239);
xnor U2409 (N_2409,N_2181,N_1980);
and U2410 (N_2410,N_1506,N_1737);
and U2411 (N_2411,N_2046,N_1666);
nand U2412 (N_2412,N_1971,N_1767);
xnor U2413 (N_2413,N_2008,N_1531);
nor U2414 (N_2414,N_1937,N_2016);
and U2415 (N_2415,N_1722,N_1710);
and U2416 (N_2416,N_1839,N_1672);
and U2417 (N_2417,N_1594,N_2020);
nand U2418 (N_2418,N_2237,N_1988);
xor U2419 (N_2419,N_1879,N_1813);
and U2420 (N_2420,N_2062,N_1793);
xor U2421 (N_2421,N_1944,N_2045);
or U2422 (N_2422,N_2185,N_1641);
or U2423 (N_2423,N_2105,N_1550);
and U2424 (N_2424,N_1643,N_2142);
and U2425 (N_2425,N_2195,N_1844);
and U2426 (N_2426,N_2018,N_1922);
nand U2427 (N_2427,N_2244,N_1620);
nor U2428 (N_2428,N_1553,N_1633);
xnor U2429 (N_2429,N_2214,N_2145);
nor U2430 (N_2430,N_1597,N_1849);
nand U2431 (N_2431,N_1572,N_1697);
or U2432 (N_2432,N_1521,N_2080);
xnor U2433 (N_2433,N_1765,N_1913);
nand U2434 (N_2434,N_2148,N_2079);
or U2435 (N_2435,N_1897,N_1546);
and U2436 (N_2436,N_1791,N_1610);
or U2437 (N_2437,N_2194,N_2138);
or U2438 (N_2438,N_1866,N_1975);
nand U2439 (N_2439,N_1870,N_1571);
or U2440 (N_2440,N_2026,N_2153);
nor U2441 (N_2441,N_1758,N_1677);
nor U2442 (N_2442,N_2204,N_1655);
nor U2443 (N_2443,N_2019,N_1968);
nor U2444 (N_2444,N_1544,N_1678);
nor U2445 (N_2445,N_1818,N_2097);
or U2446 (N_2446,N_1809,N_1885);
nand U2447 (N_2447,N_2122,N_2203);
nor U2448 (N_2448,N_2039,N_1757);
or U2449 (N_2449,N_1847,N_2109);
xor U2450 (N_2450,N_2187,N_1661);
or U2451 (N_2451,N_1642,N_1691);
nand U2452 (N_2452,N_2091,N_2001);
nor U2453 (N_2453,N_1842,N_1776);
or U2454 (N_2454,N_1502,N_1587);
nand U2455 (N_2455,N_1501,N_1622);
nand U2456 (N_2456,N_1848,N_1812);
nand U2457 (N_2457,N_1723,N_2171);
xor U2458 (N_2458,N_1978,N_1536);
or U2459 (N_2459,N_2048,N_2083);
or U2460 (N_2460,N_1650,N_2060);
xor U2461 (N_2461,N_1902,N_1987);
and U2462 (N_2462,N_2090,N_1820);
nor U2463 (N_2463,N_2220,N_2221);
nor U2464 (N_2464,N_1640,N_1896);
or U2465 (N_2465,N_2006,N_1694);
and U2466 (N_2466,N_1949,N_1802);
nor U2467 (N_2467,N_1753,N_1695);
and U2468 (N_2468,N_2162,N_2152);
nor U2469 (N_2469,N_1543,N_1771);
or U2470 (N_2470,N_1526,N_2212);
nand U2471 (N_2471,N_1875,N_1917);
nor U2472 (N_2472,N_1811,N_1604);
or U2473 (N_2473,N_1628,N_1591);
nand U2474 (N_2474,N_2073,N_1910);
and U2475 (N_2475,N_1584,N_1636);
xnor U2476 (N_2476,N_1649,N_2179);
xor U2477 (N_2477,N_1863,N_1894);
and U2478 (N_2478,N_1786,N_2092);
nor U2479 (N_2479,N_1751,N_1961);
and U2480 (N_2480,N_1639,N_1525);
and U2481 (N_2481,N_2210,N_2191);
or U2482 (N_2482,N_1970,N_1985);
or U2483 (N_2483,N_2102,N_1510);
xnor U2484 (N_2484,N_1579,N_2056);
and U2485 (N_2485,N_1635,N_1733);
nand U2486 (N_2486,N_2004,N_1732);
nand U2487 (N_2487,N_2172,N_1991);
nand U2488 (N_2488,N_1882,N_2034);
or U2489 (N_2489,N_2233,N_1993);
or U2490 (N_2490,N_1994,N_1570);
nor U2491 (N_2491,N_1599,N_2107);
nor U2492 (N_2492,N_1580,N_1557);
nor U2493 (N_2493,N_2228,N_1687);
nand U2494 (N_2494,N_1535,N_1692);
and U2495 (N_2495,N_1878,N_1675);
nand U2496 (N_2496,N_2208,N_1556);
or U2497 (N_2497,N_1864,N_2110);
or U2498 (N_2498,N_1837,N_1724);
and U2499 (N_2499,N_1826,N_1739);
nor U2500 (N_2500,N_1921,N_2061);
or U2501 (N_2501,N_1513,N_2041);
nand U2502 (N_2502,N_2168,N_1938);
and U2503 (N_2503,N_2188,N_2015);
and U2504 (N_2504,N_1801,N_2161);
or U2505 (N_2505,N_2232,N_1939);
or U2506 (N_2506,N_1973,N_1663);
nor U2507 (N_2507,N_1947,N_2166);
nand U2508 (N_2508,N_1596,N_1934);
or U2509 (N_2509,N_1832,N_2002);
nand U2510 (N_2510,N_1646,N_1514);
xor U2511 (N_2511,N_1623,N_1562);
or U2512 (N_2512,N_2106,N_2049);
nand U2513 (N_2513,N_1761,N_1752);
and U2514 (N_2514,N_1720,N_1931);
and U2515 (N_2515,N_1541,N_1977);
nand U2516 (N_2516,N_1754,N_1551);
xor U2517 (N_2517,N_1527,N_1860);
and U2518 (N_2518,N_1928,N_1828);
nand U2519 (N_2519,N_2081,N_2051);
or U2520 (N_2520,N_1590,N_1667);
and U2521 (N_2521,N_1784,N_1540);
xnor U2522 (N_2522,N_1670,N_1825);
nor U2523 (N_2523,N_2099,N_2057);
nor U2524 (N_2524,N_2213,N_2093);
nand U2525 (N_2525,N_2222,N_2021);
or U2526 (N_2526,N_1715,N_2154);
or U2527 (N_2527,N_1778,N_1874);
xnor U2528 (N_2528,N_1830,N_1787);
nor U2529 (N_2529,N_1956,N_1760);
and U2530 (N_2530,N_1634,N_1519);
nand U2531 (N_2531,N_2223,N_1686);
or U2532 (N_2532,N_1792,N_1713);
nor U2533 (N_2533,N_2087,N_2136);
nand U2534 (N_2534,N_1954,N_1905);
and U2535 (N_2535,N_1906,N_2113);
and U2536 (N_2536,N_1983,N_2027);
nand U2537 (N_2537,N_1916,N_2070);
or U2538 (N_2538,N_1810,N_2111);
xnor U2539 (N_2539,N_1814,N_1892);
nor U2540 (N_2540,N_1569,N_1682);
and U2541 (N_2541,N_1537,N_2125);
and U2542 (N_2542,N_2149,N_1621);
and U2543 (N_2543,N_1831,N_2128);
nor U2544 (N_2544,N_1900,N_1602);
nand U2545 (N_2545,N_2235,N_1838);
or U2546 (N_2546,N_1698,N_1523);
and U2547 (N_2547,N_2207,N_1929);
or U2548 (N_2548,N_2200,N_2205);
xor U2549 (N_2549,N_2151,N_2144);
nor U2550 (N_2550,N_1515,N_2241);
or U2551 (N_2551,N_1909,N_1549);
nor U2552 (N_2552,N_1756,N_1748);
xnor U2553 (N_2553,N_2193,N_2094);
and U2554 (N_2554,N_1664,N_1576);
nand U2555 (N_2555,N_1631,N_1578);
nand U2556 (N_2556,N_2120,N_2225);
or U2557 (N_2557,N_2063,N_1927);
nand U2558 (N_2558,N_2124,N_1736);
xnor U2559 (N_2559,N_1873,N_1662);
xnor U2560 (N_2560,N_1979,N_1683);
and U2561 (N_2561,N_1654,N_1548);
nor U2562 (N_2562,N_1619,N_1711);
and U2563 (N_2563,N_1804,N_1560);
and U2564 (N_2564,N_1701,N_1706);
nand U2565 (N_2565,N_1788,N_2108);
and U2566 (N_2566,N_2134,N_1966);
nand U2567 (N_2567,N_1989,N_2038);
and U2568 (N_2568,N_1918,N_2248);
and U2569 (N_2569,N_1889,N_1616);
xor U2570 (N_2570,N_1617,N_1524);
nand U2571 (N_2571,N_1833,N_1759);
nand U2572 (N_2572,N_1554,N_1862);
xnor U2573 (N_2573,N_2165,N_1512);
or U2574 (N_2574,N_2029,N_2226);
or U2575 (N_2575,N_1507,N_2143);
nor U2576 (N_2576,N_1717,N_1676);
or U2577 (N_2577,N_1781,N_1561);
and U2578 (N_2578,N_2218,N_2230);
or U2579 (N_2579,N_2215,N_1614);
or U2580 (N_2580,N_2229,N_1777);
nor U2581 (N_2581,N_1876,N_2163);
nor U2582 (N_2582,N_1857,N_2209);
nand U2583 (N_2583,N_1789,N_1517);
nor U2584 (N_2584,N_2043,N_1738);
xor U2585 (N_2585,N_2192,N_1680);
nor U2586 (N_2586,N_1718,N_1763);
nand U2587 (N_2587,N_1503,N_2137);
and U2588 (N_2588,N_2158,N_1836);
nor U2589 (N_2589,N_2054,N_2010);
nand U2590 (N_2590,N_1505,N_1705);
and U2591 (N_2591,N_1899,N_2178);
nand U2592 (N_2592,N_1986,N_1817);
nor U2593 (N_2593,N_1638,N_1764);
or U2594 (N_2594,N_2119,N_1796);
and U2595 (N_2595,N_1920,N_1565);
xor U2596 (N_2596,N_1982,N_1657);
nand U2597 (N_2597,N_2071,N_1656);
and U2598 (N_2598,N_2170,N_1932);
or U2599 (N_2599,N_1545,N_2198);
nand U2600 (N_2600,N_1925,N_2173);
nand U2601 (N_2601,N_2249,N_2174);
nand U2602 (N_2602,N_1743,N_1648);
nor U2603 (N_2603,N_1647,N_1566);
or U2604 (N_2604,N_2176,N_1629);
xor U2605 (N_2605,N_1827,N_1714);
and U2606 (N_2606,N_2186,N_1520);
or U2607 (N_2607,N_1603,N_2243);
or U2608 (N_2608,N_1799,N_2141);
or U2609 (N_2609,N_1745,N_2100);
and U2610 (N_2610,N_2035,N_2085);
or U2611 (N_2611,N_1652,N_1800);
or U2612 (N_2612,N_2131,N_1976);
or U2613 (N_2613,N_1589,N_1941);
nor U2614 (N_2614,N_1852,N_2216);
nor U2615 (N_2615,N_1770,N_2025);
nand U2616 (N_2616,N_1615,N_1967);
or U2617 (N_2617,N_1685,N_1798);
nor U2618 (N_2618,N_1684,N_2078);
and U2619 (N_2619,N_1854,N_2238);
and U2620 (N_2620,N_1822,N_1969);
nor U2621 (N_2621,N_1707,N_1653);
nand U2622 (N_2622,N_1768,N_2159);
nor U2623 (N_2623,N_2088,N_1945);
nor U2624 (N_2624,N_1951,N_1719);
nand U2625 (N_2625,N_2137,N_1847);
nand U2626 (N_2626,N_1867,N_1620);
nor U2627 (N_2627,N_1555,N_1525);
nor U2628 (N_2628,N_2088,N_1500);
and U2629 (N_2629,N_1846,N_1796);
and U2630 (N_2630,N_1801,N_1716);
nor U2631 (N_2631,N_1799,N_1875);
and U2632 (N_2632,N_2081,N_2157);
and U2633 (N_2633,N_1568,N_1674);
nand U2634 (N_2634,N_2044,N_1578);
nand U2635 (N_2635,N_2124,N_2143);
nand U2636 (N_2636,N_2067,N_1654);
or U2637 (N_2637,N_1627,N_1725);
or U2638 (N_2638,N_2022,N_1531);
and U2639 (N_2639,N_1801,N_2215);
and U2640 (N_2640,N_1869,N_2075);
xnor U2641 (N_2641,N_2047,N_1869);
and U2642 (N_2642,N_1538,N_1641);
xnor U2643 (N_2643,N_1628,N_1833);
xnor U2644 (N_2644,N_1562,N_2078);
or U2645 (N_2645,N_2120,N_2128);
and U2646 (N_2646,N_1824,N_1827);
or U2647 (N_2647,N_1875,N_1544);
nand U2648 (N_2648,N_2230,N_1881);
and U2649 (N_2649,N_1712,N_2154);
nor U2650 (N_2650,N_2102,N_1593);
nand U2651 (N_2651,N_1731,N_1954);
and U2652 (N_2652,N_2099,N_1544);
xor U2653 (N_2653,N_2110,N_1787);
or U2654 (N_2654,N_1778,N_2049);
nand U2655 (N_2655,N_1575,N_1706);
and U2656 (N_2656,N_2154,N_2162);
nor U2657 (N_2657,N_2013,N_2179);
nor U2658 (N_2658,N_2136,N_1535);
and U2659 (N_2659,N_1958,N_1967);
and U2660 (N_2660,N_2006,N_2004);
nor U2661 (N_2661,N_1977,N_2119);
and U2662 (N_2662,N_1935,N_1823);
and U2663 (N_2663,N_2115,N_1924);
and U2664 (N_2664,N_1667,N_1869);
or U2665 (N_2665,N_1912,N_1958);
nand U2666 (N_2666,N_1539,N_2092);
and U2667 (N_2667,N_1891,N_1827);
and U2668 (N_2668,N_1568,N_1785);
and U2669 (N_2669,N_2070,N_1935);
nand U2670 (N_2670,N_1851,N_1668);
or U2671 (N_2671,N_2047,N_2017);
xnor U2672 (N_2672,N_1989,N_1714);
xor U2673 (N_2673,N_1788,N_1500);
nor U2674 (N_2674,N_1857,N_1642);
and U2675 (N_2675,N_1936,N_2065);
and U2676 (N_2676,N_2137,N_1741);
or U2677 (N_2677,N_1569,N_2144);
nor U2678 (N_2678,N_1816,N_1717);
and U2679 (N_2679,N_1782,N_2103);
or U2680 (N_2680,N_2144,N_1790);
or U2681 (N_2681,N_2104,N_1613);
and U2682 (N_2682,N_2235,N_2181);
and U2683 (N_2683,N_2170,N_2245);
xor U2684 (N_2684,N_2145,N_1646);
and U2685 (N_2685,N_1510,N_1812);
nor U2686 (N_2686,N_1857,N_1529);
nand U2687 (N_2687,N_1841,N_2076);
nand U2688 (N_2688,N_2158,N_2206);
or U2689 (N_2689,N_2064,N_1508);
and U2690 (N_2690,N_1625,N_1822);
or U2691 (N_2691,N_2040,N_2051);
nand U2692 (N_2692,N_1972,N_2204);
nand U2693 (N_2693,N_2078,N_1919);
nor U2694 (N_2694,N_1887,N_1602);
or U2695 (N_2695,N_2124,N_1569);
or U2696 (N_2696,N_1742,N_2233);
or U2697 (N_2697,N_1708,N_2076);
nor U2698 (N_2698,N_1587,N_2184);
nand U2699 (N_2699,N_1793,N_2078);
and U2700 (N_2700,N_1617,N_1895);
nand U2701 (N_2701,N_1775,N_1558);
nand U2702 (N_2702,N_1958,N_1551);
and U2703 (N_2703,N_1662,N_2177);
nand U2704 (N_2704,N_1756,N_1754);
nor U2705 (N_2705,N_1643,N_2150);
and U2706 (N_2706,N_1942,N_1869);
and U2707 (N_2707,N_1634,N_2010);
and U2708 (N_2708,N_1581,N_1951);
or U2709 (N_2709,N_2193,N_1919);
or U2710 (N_2710,N_2084,N_1853);
and U2711 (N_2711,N_1555,N_1824);
nand U2712 (N_2712,N_1852,N_1715);
nor U2713 (N_2713,N_2169,N_2145);
nor U2714 (N_2714,N_1865,N_2208);
and U2715 (N_2715,N_1885,N_2184);
nand U2716 (N_2716,N_1658,N_2018);
and U2717 (N_2717,N_2096,N_1746);
nand U2718 (N_2718,N_1825,N_1559);
nand U2719 (N_2719,N_1767,N_1621);
nor U2720 (N_2720,N_1633,N_2151);
nand U2721 (N_2721,N_2086,N_2089);
and U2722 (N_2722,N_1629,N_1789);
nand U2723 (N_2723,N_1683,N_1851);
or U2724 (N_2724,N_2206,N_1801);
nand U2725 (N_2725,N_1680,N_2235);
nand U2726 (N_2726,N_2056,N_1748);
nand U2727 (N_2727,N_2220,N_1605);
and U2728 (N_2728,N_2210,N_2124);
nor U2729 (N_2729,N_1682,N_1712);
nor U2730 (N_2730,N_1734,N_1806);
and U2731 (N_2731,N_2029,N_1746);
nand U2732 (N_2732,N_1997,N_1573);
or U2733 (N_2733,N_1989,N_2033);
nand U2734 (N_2734,N_1539,N_1625);
or U2735 (N_2735,N_2137,N_1778);
nand U2736 (N_2736,N_1740,N_1634);
or U2737 (N_2737,N_2054,N_2196);
and U2738 (N_2738,N_1680,N_2080);
nor U2739 (N_2739,N_1830,N_1621);
and U2740 (N_2740,N_2217,N_2098);
and U2741 (N_2741,N_2095,N_2197);
nor U2742 (N_2742,N_1750,N_1696);
nor U2743 (N_2743,N_1754,N_2027);
nand U2744 (N_2744,N_2148,N_1989);
nand U2745 (N_2745,N_2072,N_1888);
or U2746 (N_2746,N_1941,N_2201);
or U2747 (N_2747,N_2041,N_2045);
nand U2748 (N_2748,N_1978,N_2184);
xor U2749 (N_2749,N_2185,N_1899);
xor U2750 (N_2750,N_2088,N_2153);
nand U2751 (N_2751,N_1650,N_2230);
nand U2752 (N_2752,N_1785,N_1935);
nand U2753 (N_2753,N_2231,N_1536);
nor U2754 (N_2754,N_1594,N_1622);
or U2755 (N_2755,N_1624,N_1883);
nor U2756 (N_2756,N_1815,N_1621);
xor U2757 (N_2757,N_1553,N_1680);
nand U2758 (N_2758,N_2188,N_2236);
nand U2759 (N_2759,N_2035,N_2099);
or U2760 (N_2760,N_1950,N_2191);
nand U2761 (N_2761,N_1661,N_1929);
or U2762 (N_2762,N_1809,N_1735);
nand U2763 (N_2763,N_1730,N_1893);
nor U2764 (N_2764,N_2232,N_2148);
nor U2765 (N_2765,N_2087,N_1938);
nand U2766 (N_2766,N_1637,N_1866);
nand U2767 (N_2767,N_1804,N_2115);
nand U2768 (N_2768,N_1964,N_1611);
xor U2769 (N_2769,N_1706,N_2036);
nor U2770 (N_2770,N_1844,N_1542);
and U2771 (N_2771,N_1790,N_2025);
xor U2772 (N_2772,N_1742,N_2195);
xnor U2773 (N_2773,N_1564,N_1860);
or U2774 (N_2774,N_1855,N_1869);
and U2775 (N_2775,N_1779,N_2022);
nand U2776 (N_2776,N_1969,N_1600);
and U2777 (N_2777,N_1701,N_1631);
and U2778 (N_2778,N_1828,N_1905);
nand U2779 (N_2779,N_1871,N_1850);
nand U2780 (N_2780,N_2183,N_2077);
or U2781 (N_2781,N_2136,N_2172);
and U2782 (N_2782,N_2011,N_1950);
or U2783 (N_2783,N_1554,N_2097);
and U2784 (N_2784,N_1835,N_2059);
or U2785 (N_2785,N_1504,N_1779);
or U2786 (N_2786,N_1807,N_1611);
and U2787 (N_2787,N_1758,N_2128);
nor U2788 (N_2788,N_1568,N_1657);
nor U2789 (N_2789,N_1841,N_2051);
or U2790 (N_2790,N_1801,N_2085);
nor U2791 (N_2791,N_1504,N_1522);
or U2792 (N_2792,N_1526,N_1656);
and U2793 (N_2793,N_1651,N_1731);
nor U2794 (N_2794,N_2073,N_2175);
xnor U2795 (N_2795,N_1762,N_2002);
and U2796 (N_2796,N_1971,N_2191);
xor U2797 (N_2797,N_1567,N_2220);
and U2798 (N_2798,N_1557,N_2170);
nor U2799 (N_2799,N_2184,N_1607);
and U2800 (N_2800,N_2206,N_1619);
nand U2801 (N_2801,N_2024,N_1729);
nand U2802 (N_2802,N_1659,N_1539);
nand U2803 (N_2803,N_1622,N_1854);
nand U2804 (N_2804,N_1850,N_1802);
or U2805 (N_2805,N_1639,N_1624);
nand U2806 (N_2806,N_1517,N_1998);
nor U2807 (N_2807,N_1936,N_2072);
xor U2808 (N_2808,N_1879,N_1503);
or U2809 (N_2809,N_1799,N_1562);
or U2810 (N_2810,N_2102,N_1932);
xor U2811 (N_2811,N_1889,N_1808);
or U2812 (N_2812,N_1735,N_1697);
and U2813 (N_2813,N_1900,N_1726);
nand U2814 (N_2814,N_1764,N_1759);
nor U2815 (N_2815,N_1697,N_1869);
xnor U2816 (N_2816,N_1684,N_1807);
xor U2817 (N_2817,N_2052,N_1558);
or U2818 (N_2818,N_1767,N_1882);
xnor U2819 (N_2819,N_1913,N_1607);
nand U2820 (N_2820,N_2119,N_1785);
or U2821 (N_2821,N_2039,N_1947);
or U2822 (N_2822,N_1573,N_1706);
nor U2823 (N_2823,N_2177,N_1691);
xnor U2824 (N_2824,N_1907,N_1810);
nand U2825 (N_2825,N_2188,N_1700);
xor U2826 (N_2826,N_2073,N_1603);
and U2827 (N_2827,N_1620,N_1639);
nor U2828 (N_2828,N_1578,N_1935);
nand U2829 (N_2829,N_2051,N_1951);
xor U2830 (N_2830,N_1608,N_2145);
nor U2831 (N_2831,N_2153,N_2016);
nor U2832 (N_2832,N_1913,N_1932);
or U2833 (N_2833,N_1631,N_2010);
xor U2834 (N_2834,N_1557,N_2187);
nand U2835 (N_2835,N_2010,N_2034);
or U2836 (N_2836,N_1926,N_1823);
or U2837 (N_2837,N_1838,N_2133);
or U2838 (N_2838,N_2030,N_1593);
or U2839 (N_2839,N_1821,N_1662);
or U2840 (N_2840,N_2183,N_1558);
xor U2841 (N_2841,N_1956,N_1714);
and U2842 (N_2842,N_2186,N_1940);
nand U2843 (N_2843,N_1974,N_1898);
nor U2844 (N_2844,N_2116,N_1508);
nor U2845 (N_2845,N_1823,N_1951);
or U2846 (N_2846,N_1780,N_2168);
and U2847 (N_2847,N_1982,N_1983);
and U2848 (N_2848,N_1720,N_1956);
or U2849 (N_2849,N_2150,N_1659);
and U2850 (N_2850,N_2177,N_2064);
xor U2851 (N_2851,N_1613,N_1858);
nand U2852 (N_2852,N_1752,N_1725);
nor U2853 (N_2853,N_1943,N_2243);
or U2854 (N_2854,N_2155,N_1500);
and U2855 (N_2855,N_1990,N_1503);
and U2856 (N_2856,N_1539,N_2127);
nor U2857 (N_2857,N_1508,N_1896);
and U2858 (N_2858,N_2162,N_2063);
and U2859 (N_2859,N_1706,N_1829);
nand U2860 (N_2860,N_2173,N_1763);
nand U2861 (N_2861,N_1721,N_1669);
or U2862 (N_2862,N_1903,N_2230);
and U2863 (N_2863,N_1806,N_1838);
or U2864 (N_2864,N_1860,N_1870);
and U2865 (N_2865,N_1751,N_1803);
or U2866 (N_2866,N_1501,N_1693);
nor U2867 (N_2867,N_2117,N_2167);
or U2868 (N_2868,N_1948,N_2246);
xor U2869 (N_2869,N_1533,N_1534);
nor U2870 (N_2870,N_1919,N_1828);
nor U2871 (N_2871,N_1977,N_1548);
nor U2872 (N_2872,N_1567,N_1794);
or U2873 (N_2873,N_2002,N_1989);
xnor U2874 (N_2874,N_1905,N_1595);
and U2875 (N_2875,N_1805,N_2158);
and U2876 (N_2876,N_2191,N_2083);
xnor U2877 (N_2877,N_2217,N_2090);
nor U2878 (N_2878,N_2230,N_2071);
or U2879 (N_2879,N_1782,N_1657);
and U2880 (N_2880,N_2207,N_1691);
and U2881 (N_2881,N_1999,N_2156);
xnor U2882 (N_2882,N_1693,N_2223);
and U2883 (N_2883,N_1568,N_2104);
nand U2884 (N_2884,N_1551,N_1931);
nor U2885 (N_2885,N_1700,N_1890);
nand U2886 (N_2886,N_1546,N_1831);
nor U2887 (N_2887,N_2032,N_1585);
nand U2888 (N_2888,N_2032,N_1543);
or U2889 (N_2889,N_1876,N_2064);
or U2890 (N_2890,N_1749,N_2155);
or U2891 (N_2891,N_2065,N_1848);
and U2892 (N_2892,N_1994,N_1842);
or U2893 (N_2893,N_1952,N_2124);
and U2894 (N_2894,N_2019,N_1707);
and U2895 (N_2895,N_1722,N_2153);
or U2896 (N_2896,N_1935,N_2135);
and U2897 (N_2897,N_1983,N_1964);
and U2898 (N_2898,N_1943,N_2169);
nor U2899 (N_2899,N_1701,N_1601);
nor U2900 (N_2900,N_2226,N_1671);
and U2901 (N_2901,N_1782,N_2213);
and U2902 (N_2902,N_2243,N_1539);
or U2903 (N_2903,N_1976,N_2066);
nor U2904 (N_2904,N_1922,N_1731);
nand U2905 (N_2905,N_1805,N_1730);
or U2906 (N_2906,N_1635,N_2168);
xor U2907 (N_2907,N_1679,N_1878);
nor U2908 (N_2908,N_1921,N_1636);
or U2909 (N_2909,N_2144,N_1884);
nor U2910 (N_2910,N_1653,N_1967);
nor U2911 (N_2911,N_1851,N_2245);
and U2912 (N_2912,N_1700,N_1694);
nor U2913 (N_2913,N_2146,N_2187);
nor U2914 (N_2914,N_1704,N_2077);
and U2915 (N_2915,N_1704,N_1880);
or U2916 (N_2916,N_1716,N_1730);
or U2917 (N_2917,N_1870,N_1724);
nor U2918 (N_2918,N_1517,N_1927);
or U2919 (N_2919,N_1516,N_1951);
and U2920 (N_2920,N_2035,N_1657);
nand U2921 (N_2921,N_1924,N_1597);
and U2922 (N_2922,N_2138,N_1897);
or U2923 (N_2923,N_2001,N_1517);
nor U2924 (N_2924,N_2023,N_1708);
or U2925 (N_2925,N_1533,N_1625);
or U2926 (N_2926,N_2051,N_1759);
nor U2927 (N_2927,N_2194,N_2182);
nand U2928 (N_2928,N_2223,N_2092);
nand U2929 (N_2929,N_1708,N_1574);
or U2930 (N_2930,N_2215,N_1806);
or U2931 (N_2931,N_1875,N_1638);
nor U2932 (N_2932,N_1891,N_1900);
nand U2933 (N_2933,N_1550,N_1791);
nor U2934 (N_2934,N_2201,N_2085);
nor U2935 (N_2935,N_1644,N_1789);
and U2936 (N_2936,N_2185,N_1675);
or U2937 (N_2937,N_1860,N_1936);
and U2938 (N_2938,N_1974,N_2152);
nand U2939 (N_2939,N_1523,N_1606);
nor U2940 (N_2940,N_2011,N_1925);
nand U2941 (N_2941,N_1782,N_1985);
nor U2942 (N_2942,N_1638,N_1960);
xor U2943 (N_2943,N_1621,N_2183);
nand U2944 (N_2944,N_2096,N_1531);
and U2945 (N_2945,N_2123,N_2139);
and U2946 (N_2946,N_1920,N_1580);
nor U2947 (N_2947,N_1522,N_1755);
and U2948 (N_2948,N_2002,N_2179);
nand U2949 (N_2949,N_1755,N_2194);
and U2950 (N_2950,N_2197,N_2135);
and U2951 (N_2951,N_2146,N_1570);
xor U2952 (N_2952,N_2045,N_2099);
nor U2953 (N_2953,N_1953,N_1571);
and U2954 (N_2954,N_1859,N_1677);
and U2955 (N_2955,N_1729,N_1726);
and U2956 (N_2956,N_2144,N_1861);
and U2957 (N_2957,N_1955,N_1757);
nor U2958 (N_2958,N_2086,N_2075);
and U2959 (N_2959,N_1815,N_1642);
or U2960 (N_2960,N_2037,N_1571);
nand U2961 (N_2961,N_1687,N_1839);
and U2962 (N_2962,N_1521,N_1910);
nand U2963 (N_2963,N_1810,N_2097);
nand U2964 (N_2964,N_2028,N_2047);
or U2965 (N_2965,N_1992,N_2212);
and U2966 (N_2966,N_1792,N_1515);
or U2967 (N_2967,N_1713,N_1691);
nor U2968 (N_2968,N_2099,N_1945);
nor U2969 (N_2969,N_1608,N_1503);
or U2970 (N_2970,N_1781,N_2230);
nand U2971 (N_2971,N_1952,N_2200);
nor U2972 (N_2972,N_2000,N_1805);
or U2973 (N_2973,N_1948,N_2173);
nor U2974 (N_2974,N_2152,N_1989);
nand U2975 (N_2975,N_1915,N_1980);
nor U2976 (N_2976,N_1783,N_1839);
and U2977 (N_2977,N_1869,N_2044);
and U2978 (N_2978,N_1605,N_1681);
nor U2979 (N_2979,N_1890,N_2148);
xor U2980 (N_2980,N_1628,N_1580);
or U2981 (N_2981,N_2192,N_1563);
nand U2982 (N_2982,N_1583,N_2158);
or U2983 (N_2983,N_2235,N_2066);
or U2984 (N_2984,N_1679,N_1858);
and U2985 (N_2985,N_1515,N_1588);
and U2986 (N_2986,N_1870,N_2152);
nor U2987 (N_2987,N_2211,N_2227);
nor U2988 (N_2988,N_1667,N_1511);
nor U2989 (N_2989,N_2159,N_2154);
nor U2990 (N_2990,N_1559,N_1683);
and U2991 (N_2991,N_2127,N_2207);
nand U2992 (N_2992,N_1529,N_1739);
nand U2993 (N_2993,N_1860,N_1932);
nand U2994 (N_2994,N_2014,N_2070);
nand U2995 (N_2995,N_2205,N_1535);
nor U2996 (N_2996,N_1937,N_1696);
nor U2997 (N_2997,N_2092,N_1917);
nor U2998 (N_2998,N_1615,N_1773);
nand U2999 (N_2999,N_1920,N_1951);
xnor U3000 (N_3000,N_2562,N_2936);
or U3001 (N_3001,N_2296,N_2655);
xor U3002 (N_3002,N_2552,N_2255);
nand U3003 (N_3003,N_2368,N_2875);
or U3004 (N_3004,N_2627,N_2793);
and U3005 (N_3005,N_2880,N_2436);
or U3006 (N_3006,N_2832,N_2277);
nand U3007 (N_3007,N_2459,N_2488);
xnor U3008 (N_3008,N_2509,N_2857);
and U3009 (N_3009,N_2814,N_2555);
or U3010 (N_3010,N_2365,N_2886);
nand U3011 (N_3011,N_2478,N_2588);
nand U3012 (N_3012,N_2926,N_2749);
nor U3013 (N_3013,N_2645,N_2716);
nand U3014 (N_3014,N_2523,N_2802);
nand U3015 (N_3015,N_2896,N_2809);
xnor U3016 (N_3016,N_2270,N_2499);
xor U3017 (N_3017,N_2288,N_2884);
xnor U3018 (N_3018,N_2556,N_2981);
or U3019 (N_3019,N_2479,N_2739);
nor U3020 (N_3020,N_2625,N_2691);
or U3021 (N_3021,N_2601,N_2890);
or U3022 (N_3022,N_2976,N_2966);
nand U3023 (N_3023,N_2912,N_2514);
nor U3024 (N_3024,N_2983,N_2780);
and U3025 (N_3025,N_2569,N_2399);
and U3026 (N_3026,N_2619,N_2755);
and U3027 (N_3027,N_2495,N_2414);
nor U3028 (N_3028,N_2431,N_2456);
nor U3029 (N_3029,N_2615,N_2674);
nand U3030 (N_3030,N_2901,N_2502);
nor U3031 (N_3031,N_2786,N_2358);
nand U3032 (N_3032,N_2433,N_2761);
nor U3033 (N_3033,N_2341,N_2476);
and U3034 (N_3034,N_2993,N_2961);
or U3035 (N_3035,N_2692,N_2975);
nor U3036 (N_3036,N_2818,N_2529);
and U3037 (N_3037,N_2375,N_2672);
nor U3038 (N_3038,N_2913,N_2520);
or U3039 (N_3039,N_2524,N_2577);
nand U3040 (N_3040,N_2776,N_2256);
nand U3041 (N_3041,N_2335,N_2825);
xor U3042 (N_3042,N_2357,N_2503);
or U3043 (N_3043,N_2799,N_2643);
nor U3044 (N_3044,N_2383,N_2889);
nand U3045 (N_3045,N_2564,N_2883);
and U3046 (N_3046,N_2282,N_2711);
xnor U3047 (N_3047,N_2989,N_2957);
nand U3048 (N_3048,N_2977,N_2455);
nor U3049 (N_3049,N_2589,N_2508);
nand U3050 (N_3050,N_2690,N_2490);
or U3051 (N_3051,N_2254,N_2516);
nor U3052 (N_3052,N_2581,N_2699);
nor U3053 (N_3053,N_2421,N_2602);
or U3054 (N_3054,N_2487,N_2658);
nand U3055 (N_3055,N_2385,N_2806);
nand U3056 (N_3056,N_2424,N_2262);
or U3057 (N_3057,N_2554,N_2994);
nor U3058 (N_3058,N_2572,N_2822);
nand U3059 (N_3059,N_2428,N_2921);
or U3060 (N_3060,N_2693,N_2485);
and U3061 (N_3061,N_2752,N_2475);
nand U3062 (N_3062,N_2534,N_2733);
or U3063 (N_3063,N_2486,N_2967);
nor U3064 (N_3064,N_2550,N_2662);
nand U3065 (N_3065,N_2607,N_2997);
nor U3066 (N_3066,N_2865,N_2449);
nor U3067 (N_3067,N_2530,N_2613);
xor U3068 (N_3068,N_2753,N_2984);
or U3069 (N_3069,N_2960,N_2535);
nor U3070 (N_3070,N_2506,N_2267);
xnor U3071 (N_3071,N_2732,N_2784);
or U3072 (N_3072,N_2268,N_2393);
or U3073 (N_3073,N_2673,N_2945);
nand U3074 (N_3074,N_2548,N_2726);
nor U3075 (N_3075,N_2877,N_2561);
nand U3076 (N_3076,N_2338,N_2911);
or U3077 (N_3077,N_2898,N_2264);
or U3078 (N_3078,N_2764,N_2763);
and U3079 (N_3079,N_2782,N_2578);
nor U3080 (N_3080,N_2582,N_2873);
nor U3081 (N_3081,N_2702,N_2489);
or U3082 (N_3082,N_2316,N_2311);
and U3083 (N_3083,N_2861,N_2930);
nor U3084 (N_3084,N_2986,N_2928);
nor U3085 (N_3085,N_2531,N_2415);
xor U3086 (N_3086,N_2999,N_2418);
nor U3087 (N_3087,N_2622,N_2280);
xnor U3088 (N_3088,N_2309,N_2794);
and U3089 (N_3089,N_2330,N_2988);
nor U3090 (N_3090,N_2656,N_2536);
or U3091 (N_3091,N_2964,N_2423);
and U3092 (N_3092,N_2949,N_2305);
nor U3093 (N_3093,N_2453,N_2891);
nand U3094 (N_3094,N_2532,N_2855);
or U3095 (N_3095,N_2633,N_2778);
nand U3096 (N_3096,N_2797,N_2298);
nand U3097 (N_3097,N_2512,N_2491);
nor U3098 (N_3098,N_2819,N_2319);
nand U3099 (N_3099,N_2969,N_2637);
nor U3100 (N_3100,N_2852,N_2540);
and U3101 (N_3101,N_2329,N_2481);
nor U3102 (N_3102,N_2370,N_2679);
nor U3103 (N_3103,N_2392,N_2354);
and U3104 (N_3104,N_2844,N_2477);
and U3105 (N_3105,N_2683,N_2566);
nor U3106 (N_3106,N_2751,N_2841);
nand U3107 (N_3107,N_2652,N_2834);
nand U3108 (N_3108,N_2703,N_2501);
nor U3109 (N_3109,N_2823,N_2366);
and U3110 (N_3110,N_2545,N_2632);
or U3111 (N_3111,N_2468,N_2629);
and U3112 (N_3112,N_2259,N_2792);
and U3113 (N_3113,N_2680,N_2798);
nor U3114 (N_3114,N_2342,N_2482);
nand U3115 (N_3115,N_2695,N_2253);
nor U3116 (N_3116,N_2642,N_2933);
xnor U3117 (N_3117,N_2351,N_2850);
and U3118 (N_3118,N_2729,N_2777);
or U3119 (N_3119,N_2483,N_2304);
xor U3120 (N_3120,N_2738,N_2575);
nand U3121 (N_3121,N_2872,N_2878);
nand U3122 (N_3122,N_2323,N_2686);
nor U3123 (N_3123,N_2346,N_2942);
nand U3124 (N_3124,N_2671,N_2888);
xnor U3125 (N_3125,N_2598,N_2467);
or U3126 (N_3126,N_2684,N_2522);
nor U3127 (N_3127,N_2462,N_2331);
nand U3128 (N_3128,N_2756,N_2694);
or U3129 (N_3129,N_2263,N_2987);
nor U3130 (N_3130,N_2829,N_2731);
xnor U3131 (N_3131,N_2376,N_2381);
or U3132 (N_3132,N_2845,N_2626);
xnor U3133 (N_3133,N_2868,N_2294);
nor U3134 (N_3134,N_2864,N_2546);
nor U3135 (N_3135,N_2286,N_2922);
or U3136 (N_3136,N_2271,N_2412);
nor U3137 (N_3137,N_2905,N_2608);
or U3138 (N_3138,N_2448,N_2718);
or U3139 (N_3139,N_2741,N_2333);
nor U3140 (N_3140,N_2876,N_2874);
or U3141 (N_3141,N_2526,N_2434);
nor U3142 (N_3142,N_2301,N_2353);
or U3143 (N_3143,N_2585,N_2343);
xnor U3144 (N_3144,N_2590,N_2340);
and U3145 (N_3145,N_2973,N_2881);
or U3146 (N_3146,N_2696,N_2635);
nor U3147 (N_3147,N_2879,N_2668);
nor U3148 (N_3148,N_2885,N_2549);
nand U3149 (N_3149,N_2442,N_2371);
nor U3150 (N_3150,N_2398,N_2283);
or U3151 (N_3151,N_2750,N_2909);
nand U3152 (N_3152,N_2307,N_2728);
nor U3153 (N_3153,N_2599,N_2722);
xor U3154 (N_3154,N_2473,N_2787);
xor U3155 (N_3155,N_2836,N_2712);
nor U3156 (N_3156,N_2273,N_2929);
nor U3157 (N_3157,N_2854,N_2406);
and U3158 (N_3158,N_2427,N_2788);
and U3159 (N_3159,N_2952,N_2510);
nand U3160 (N_3160,N_2355,N_2466);
nor U3161 (N_3161,N_2742,N_2859);
or U3162 (N_3162,N_2367,N_2736);
or U3163 (N_3163,N_2458,N_2943);
or U3164 (N_3164,N_2940,N_2946);
xnor U3165 (N_3165,N_2820,N_2443);
nor U3166 (N_3166,N_2372,N_2916);
nand U3167 (N_3167,N_2297,N_2789);
nand U3168 (N_3168,N_2727,N_2407);
and U3169 (N_3169,N_2700,N_2541);
nand U3170 (N_3170,N_2647,N_2849);
or U3171 (N_3171,N_2698,N_2308);
nor U3172 (N_3172,N_2828,N_2609);
and U3173 (N_3173,N_2397,N_2269);
or U3174 (N_3174,N_2306,N_2646);
nand U3175 (N_3175,N_2639,N_2597);
and U3176 (N_3176,N_2616,N_2528);
nand U3177 (N_3177,N_2663,N_2801);
and U3178 (N_3178,N_2285,N_2903);
or U3179 (N_3179,N_2725,N_2650);
nand U3180 (N_3180,N_2737,N_2363);
and U3181 (N_3181,N_2498,N_2471);
or U3182 (N_3182,N_2402,N_2720);
and U3183 (N_3183,N_2920,N_2278);
nor U3184 (N_3184,N_2866,N_2704);
nor U3185 (N_3185,N_2312,N_2826);
nor U3186 (N_3186,N_2551,N_2317);
or U3187 (N_3187,N_2553,N_2678);
or U3188 (N_3188,N_2580,N_2250);
nand U3189 (N_3189,N_2387,N_2507);
and U3190 (N_3190,N_2290,N_2900);
or U3191 (N_3191,N_2527,N_2303);
xnor U3192 (N_3192,N_2446,N_2604);
nand U3193 (N_3193,N_2992,N_2915);
nor U3194 (N_3194,N_2591,N_2848);
nor U3195 (N_3195,N_2902,N_2813);
or U3196 (N_3196,N_2817,N_2723);
and U3197 (N_3197,N_2324,N_2759);
nor U3198 (N_3198,N_2935,N_2557);
and U3199 (N_3199,N_2361,N_2500);
nor U3200 (N_3200,N_2775,N_2724);
xor U3201 (N_3201,N_2537,N_2416);
or U3202 (N_3202,N_2746,N_2587);
nand U3203 (N_3203,N_2745,N_2917);
nand U3204 (N_3204,N_2380,N_2260);
and U3205 (N_3205,N_2839,N_2411);
nor U3206 (N_3206,N_2689,N_2925);
nand U3207 (N_3207,N_2560,N_2653);
nor U3208 (N_3208,N_2785,N_2707);
nand U3209 (N_3209,N_2605,N_2706);
or U3210 (N_3210,N_2772,N_2377);
and U3211 (N_3211,N_2369,N_2544);
or U3212 (N_3212,N_2413,N_2719);
xnor U3213 (N_3213,N_2594,N_2677);
nor U3214 (N_3214,N_2675,N_2420);
nor U3215 (N_3215,N_2640,N_2621);
or U3216 (N_3216,N_2807,N_2440);
nor U3217 (N_3217,N_2687,N_2291);
or U3218 (N_3218,N_2451,N_2388);
nand U3219 (N_3219,N_2505,N_2571);
and U3220 (N_3220,N_2394,N_2948);
nor U3221 (N_3221,N_2344,N_2757);
nor U3222 (N_3222,N_2904,N_2570);
nor U3223 (N_3223,N_2810,N_2617);
xnor U3224 (N_3224,N_2284,N_2403);
nand U3225 (N_3225,N_2941,N_2827);
or U3226 (N_3226,N_2417,N_2261);
xnor U3227 (N_3227,N_2676,N_2714);
nand U3228 (N_3228,N_2539,N_2595);
nor U3229 (N_3229,N_2337,N_2493);
and U3230 (N_3230,N_2908,N_2389);
nor U3231 (N_3231,N_2321,N_2334);
and U3232 (N_3232,N_2887,N_2944);
and U3233 (N_3233,N_2795,N_2513);
nor U3234 (N_3234,N_2592,N_2390);
and U3235 (N_3235,N_2325,N_2979);
nand U3236 (N_3236,N_2894,N_2644);
nand U3237 (N_3237,N_2910,N_2584);
or U3238 (N_3238,N_2767,N_2740);
nor U3239 (N_3239,N_2950,N_2408);
nand U3240 (N_3240,N_2982,N_2669);
or U3241 (N_3241,N_2766,N_2435);
nor U3242 (N_3242,N_2519,N_2842);
xor U3243 (N_3243,N_2563,N_2295);
or U3244 (N_3244,N_2314,N_2445);
nand U3245 (N_3245,N_2614,N_2636);
nor U3246 (N_3246,N_2892,N_2754);
xor U3247 (N_3247,N_2790,N_2847);
and U3248 (N_3248,N_2744,N_2279);
nand U3249 (N_3249,N_2918,N_2897);
or U3250 (N_3250,N_2391,N_2927);
and U3251 (N_3251,N_2631,N_2893);
xnor U3252 (N_3252,N_2300,N_2715);
nor U3253 (N_3253,N_2618,N_2538);
nand U3254 (N_3254,N_2292,N_2426);
and U3255 (N_3255,N_2914,N_2439);
nor U3256 (N_3256,N_2939,N_2934);
nand U3257 (N_3257,N_2606,N_2452);
xor U3258 (N_3258,N_2543,N_2252);
and U3259 (N_3259,N_2593,N_2313);
nand U3260 (N_3260,N_2734,N_2947);
and U3261 (N_3261,N_2289,N_2705);
nand U3262 (N_3262,N_2400,N_2923);
xnor U3263 (N_3263,N_2821,N_2919);
and U3264 (N_3264,N_2511,N_2359);
xnor U3265 (N_3265,N_2410,N_2469);
nand U3266 (N_3266,N_2525,N_2721);
nor U3267 (N_3267,N_2717,N_2634);
or U3268 (N_3268,N_2474,N_2956);
or U3269 (N_3269,N_2611,N_2480);
or U3270 (N_3270,N_2871,N_2816);
and U3271 (N_3271,N_2762,N_2275);
or U3272 (N_3272,N_2257,N_2951);
xnor U3273 (N_3273,N_2743,N_2974);
nor U3274 (N_3274,N_2460,N_2838);
nand U3275 (N_3275,N_2612,N_2293);
nor U3276 (N_3276,N_2339,N_2573);
nand U3277 (N_3277,N_2781,N_2384);
and U3278 (N_3278,N_2444,N_2515);
nor U3279 (N_3279,N_2968,N_2990);
and U3280 (N_3280,N_2345,N_2962);
nor U3281 (N_3281,N_2463,N_2682);
or U3282 (N_3282,N_2980,N_2830);
and U3283 (N_3283,N_2831,N_2701);
nor U3284 (N_3284,N_2840,N_2533);
nor U3285 (N_3285,N_2559,N_2867);
nor U3286 (N_3286,N_2379,N_2299);
nor U3287 (N_3287,N_2266,N_2657);
nand U3288 (N_3288,N_2382,N_2396);
or U3289 (N_3289,N_2765,N_2998);
nor U3290 (N_3290,N_2791,N_2464);
nor U3291 (N_3291,N_2862,N_2352);
nand U3292 (N_3292,N_2659,N_2709);
or U3293 (N_3293,N_2437,N_2438);
and U3294 (N_3294,N_2496,N_2708);
or U3295 (N_3295,N_2747,N_2362);
xnor U3296 (N_3296,N_2378,N_2758);
or U3297 (N_3297,N_2858,N_2425);
and U3298 (N_3298,N_2666,N_2815);
or U3299 (N_3299,N_2651,N_2472);
or U3300 (N_3300,N_2447,N_2336);
nor U3301 (N_3301,N_2600,N_2805);
and U3302 (N_3302,N_2837,N_2504);
and U3303 (N_3303,N_2863,N_2924);
nand U3304 (N_3304,N_2688,N_2386);
or U3305 (N_3305,N_2395,N_2628);
nand U3306 (N_3306,N_2985,N_2931);
nand U3307 (N_3307,N_2429,N_2735);
nand U3308 (N_3308,N_2995,N_2641);
or U3309 (N_3309,N_2310,N_2665);
nand U3310 (N_3310,N_2853,N_2347);
nand U3311 (N_3311,N_2547,N_2567);
nor U3312 (N_3312,N_2374,N_2409);
nor U3313 (N_3313,N_2586,N_2484);
and U3314 (N_3314,N_2565,N_2610);
and U3315 (N_3315,N_2405,N_2970);
or U3316 (N_3316,N_2661,N_2856);
and U3317 (N_3317,N_2769,N_2860);
and U3318 (N_3318,N_2518,N_2870);
nand U3319 (N_3319,N_2664,N_2667);
nand U3320 (N_3320,N_2251,N_2326);
nand U3321 (N_3321,N_2649,N_2364);
and U3322 (N_3322,N_2517,N_2457);
nand U3323 (N_3323,N_2978,N_2835);
or U3324 (N_3324,N_2470,N_2596);
or U3325 (N_3325,N_2265,N_2783);
and U3326 (N_3326,N_2521,N_2274);
or U3327 (N_3327,N_2302,N_2349);
nor U3328 (N_3328,N_2497,N_2328);
nand U3329 (N_3329,N_2558,N_2869);
and U3330 (N_3330,N_2670,N_2315);
nor U3331 (N_3331,N_2846,N_2938);
and U3332 (N_3332,N_2373,N_2465);
and U3333 (N_3333,N_2630,N_2954);
xor U3334 (N_3334,N_2771,N_2322);
and U3335 (N_3335,N_2603,N_2811);
nand U3336 (N_3336,N_2430,N_2620);
and U3337 (N_3337,N_2906,N_2350);
or U3338 (N_3338,N_2958,N_2287);
nor U3339 (N_3339,N_2895,N_2937);
nand U3340 (N_3340,N_2419,N_2851);
xor U3341 (N_3341,N_2422,N_2360);
and U3342 (N_3342,N_2272,N_2624);
or U3343 (N_3343,N_2576,N_2320);
nand U3344 (N_3344,N_2685,N_2332);
nor U3345 (N_3345,N_2568,N_2730);
and U3346 (N_3346,N_2773,N_2404);
and U3347 (N_3347,N_2774,N_2401);
nor U3348 (N_3348,N_2972,N_2996);
nor U3349 (N_3349,N_2681,N_2779);
and U3350 (N_3350,N_2899,N_2281);
nand U3351 (N_3351,N_2760,N_2971);
xor U3352 (N_3352,N_2450,N_2804);
nand U3353 (N_3353,N_2623,N_2770);
nand U3354 (N_3354,N_2648,N_2824);
or U3355 (N_3355,N_2492,N_2348);
nand U3356 (N_3356,N_2713,N_2638);
nor U3357 (N_3357,N_2991,N_2276);
or U3358 (N_3358,N_2953,N_2454);
xnor U3359 (N_3359,N_2579,N_2882);
or U3360 (N_3360,N_2494,N_2808);
and U3361 (N_3361,N_2318,N_2812);
nor U3362 (N_3362,N_2461,N_2258);
and U3363 (N_3363,N_2654,N_2748);
nor U3364 (N_3364,N_2965,N_2327);
or U3365 (N_3365,N_2542,N_2697);
nor U3366 (N_3366,N_2441,N_2959);
and U3367 (N_3367,N_2768,N_2710);
nor U3368 (N_3368,N_2796,N_2574);
and U3369 (N_3369,N_2432,N_2907);
nor U3370 (N_3370,N_2833,N_2583);
or U3371 (N_3371,N_2800,N_2803);
and U3372 (N_3372,N_2963,N_2356);
nand U3373 (N_3373,N_2660,N_2843);
nand U3374 (N_3374,N_2955,N_2932);
nand U3375 (N_3375,N_2339,N_2827);
or U3376 (N_3376,N_2304,N_2839);
nor U3377 (N_3377,N_2539,N_2259);
or U3378 (N_3378,N_2494,N_2631);
and U3379 (N_3379,N_2284,N_2445);
nand U3380 (N_3380,N_2371,N_2542);
nand U3381 (N_3381,N_2643,N_2716);
nand U3382 (N_3382,N_2939,N_2730);
and U3383 (N_3383,N_2793,N_2615);
and U3384 (N_3384,N_2516,N_2454);
nor U3385 (N_3385,N_2677,N_2609);
nand U3386 (N_3386,N_2352,N_2918);
and U3387 (N_3387,N_2479,N_2748);
and U3388 (N_3388,N_2253,N_2345);
or U3389 (N_3389,N_2438,N_2908);
or U3390 (N_3390,N_2259,N_2614);
or U3391 (N_3391,N_2934,N_2793);
nor U3392 (N_3392,N_2650,N_2489);
nand U3393 (N_3393,N_2563,N_2626);
and U3394 (N_3394,N_2843,N_2852);
nand U3395 (N_3395,N_2333,N_2378);
or U3396 (N_3396,N_2522,N_2979);
nor U3397 (N_3397,N_2618,N_2331);
and U3398 (N_3398,N_2699,N_2451);
nor U3399 (N_3399,N_2492,N_2910);
and U3400 (N_3400,N_2969,N_2946);
and U3401 (N_3401,N_2631,N_2421);
and U3402 (N_3402,N_2513,N_2579);
xor U3403 (N_3403,N_2970,N_2839);
or U3404 (N_3404,N_2916,N_2571);
or U3405 (N_3405,N_2539,N_2677);
nor U3406 (N_3406,N_2437,N_2604);
or U3407 (N_3407,N_2377,N_2326);
nand U3408 (N_3408,N_2344,N_2712);
nand U3409 (N_3409,N_2255,N_2570);
nand U3410 (N_3410,N_2400,N_2634);
nand U3411 (N_3411,N_2706,N_2583);
and U3412 (N_3412,N_2323,N_2540);
or U3413 (N_3413,N_2555,N_2822);
and U3414 (N_3414,N_2970,N_2946);
nand U3415 (N_3415,N_2722,N_2721);
and U3416 (N_3416,N_2932,N_2778);
and U3417 (N_3417,N_2493,N_2366);
nor U3418 (N_3418,N_2555,N_2570);
xor U3419 (N_3419,N_2427,N_2693);
nor U3420 (N_3420,N_2929,N_2353);
nor U3421 (N_3421,N_2967,N_2564);
xor U3422 (N_3422,N_2622,N_2323);
nand U3423 (N_3423,N_2999,N_2684);
xnor U3424 (N_3424,N_2360,N_2464);
and U3425 (N_3425,N_2794,N_2458);
nor U3426 (N_3426,N_2275,N_2695);
nand U3427 (N_3427,N_2892,N_2280);
and U3428 (N_3428,N_2337,N_2949);
nand U3429 (N_3429,N_2582,N_2864);
nand U3430 (N_3430,N_2387,N_2455);
or U3431 (N_3431,N_2563,N_2777);
nand U3432 (N_3432,N_2701,N_2364);
or U3433 (N_3433,N_2728,N_2383);
or U3434 (N_3434,N_2929,N_2698);
and U3435 (N_3435,N_2892,N_2376);
nor U3436 (N_3436,N_2652,N_2697);
or U3437 (N_3437,N_2328,N_2312);
or U3438 (N_3438,N_2732,N_2656);
and U3439 (N_3439,N_2915,N_2256);
nand U3440 (N_3440,N_2993,N_2859);
or U3441 (N_3441,N_2618,N_2286);
nand U3442 (N_3442,N_2830,N_2615);
nor U3443 (N_3443,N_2558,N_2722);
or U3444 (N_3444,N_2715,N_2794);
and U3445 (N_3445,N_2938,N_2851);
xnor U3446 (N_3446,N_2605,N_2839);
and U3447 (N_3447,N_2802,N_2671);
nand U3448 (N_3448,N_2756,N_2948);
or U3449 (N_3449,N_2339,N_2952);
or U3450 (N_3450,N_2780,N_2848);
and U3451 (N_3451,N_2673,N_2295);
and U3452 (N_3452,N_2645,N_2733);
or U3453 (N_3453,N_2932,N_2351);
nor U3454 (N_3454,N_2523,N_2876);
or U3455 (N_3455,N_2885,N_2944);
and U3456 (N_3456,N_2914,N_2940);
nor U3457 (N_3457,N_2726,N_2399);
nand U3458 (N_3458,N_2823,N_2624);
or U3459 (N_3459,N_2407,N_2266);
and U3460 (N_3460,N_2710,N_2706);
nor U3461 (N_3461,N_2740,N_2738);
xnor U3462 (N_3462,N_2748,N_2504);
xor U3463 (N_3463,N_2320,N_2926);
xor U3464 (N_3464,N_2949,N_2894);
nand U3465 (N_3465,N_2733,N_2943);
or U3466 (N_3466,N_2498,N_2890);
or U3467 (N_3467,N_2917,N_2801);
nand U3468 (N_3468,N_2541,N_2714);
or U3469 (N_3469,N_2487,N_2925);
or U3470 (N_3470,N_2650,N_2736);
and U3471 (N_3471,N_2371,N_2687);
nand U3472 (N_3472,N_2550,N_2641);
nor U3473 (N_3473,N_2753,N_2678);
xor U3474 (N_3474,N_2879,N_2462);
or U3475 (N_3475,N_2353,N_2989);
or U3476 (N_3476,N_2338,N_2344);
nand U3477 (N_3477,N_2432,N_2933);
nand U3478 (N_3478,N_2261,N_2626);
and U3479 (N_3479,N_2404,N_2937);
or U3480 (N_3480,N_2662,N_2276);
or U3481 (N_3481,N_2893,N_2360);
or U3482 (N_3482,N_2939,N_2404);
nor U3483 (N_3483,N_2678,N_2386);
xor U3484 (N_3484,N_2517,N_2409);
and U3485 (N_3485,N_2340,N_2519);
xnor U3486 (N_3486,N_2396,N_2916);
nand U3487 (N_3487,N_2649,N_2335);
nand U3488 (N_3488,N_2717,N_2426);
and U3489 (N_3489,N_2724,N_2965);
or U3490 (N_3490,N_2292,N_2817);
nor U3491 (N_3491,N_2307,N_2941);
or U3492 (N_3492,N_2844,N_2362);
or U3493 (N_3493,N_2738,N_2959);
and U3494 (N_3494,N_2407,N_2256);
and U3495 (N_3495,N_2448,N_2584);
or U3496 (N_3496,N_2840,N_2499);
nor U3497 (N_3497,N_2601,N_2809);
and U3498 (N_3498,N_2293,N_2743);
nand U3499 (N_3499,N_2933,N_2824);
nor U3500 (N_3500,N_2672,N_2986);
and U3501 (N_3501,N_2566,N_2312);
xnor U3502 (N_3502,N_2575,N_2879);
or U3503 (N_3503,N_2460,N_2752);
nor U3504 (N_3504,N_2554,N_2409);
or U3505 (N_3505,N_2845,N_2889);
nor U3506 (N_3506,N_2553,N_2495);
nand U3507 (N_3507,N_2376,N_2678);
nand U3508 (N_3508,N_2604,N_2411);
and U3509 (N_3509,N_2348,N_2636);
nand U3510 (N_3510,N_2882,N_2549);
or U3511 (N_3511,N_2410,N_2467);
nand U3512 (N_3512,N_2442,N_2785);
nand U3513 (N_3513,N_2382,N_2778);
xor U3514 (N_3514,N_2904,N_2961);
or U3515 (N_3515,N_2740,N_2692);
and U3516 (N_3516,N_2642,N_2564);
or U3517 (N_3517,N_2388,N_2394);
nand U3518 (N_3518,N_2267,N_2334);
nand U3519 (N_3519,N_2321,N_2317);
or U3520 (N_3520,N_2962,N_2673);
and U3521 (N_3521,N_2797,N_2560);
nor U3522 (N_3522,N_2370,N_2826);
xor U3523 (N_3523,N_2676,N_2732);
nor U3524 (N_3524,N_2364,N_2309);
nor U3525 (N_3525,N_2828,N_2900);
or U3526 (N_3526,N_2934,N_2638);
or U3527 (N_3527,N_2861,N_2821);
or U3528 (N_3528,N_2456,N_2301);
nor U3529 (N_3529,N_2795,N_2881);
nand U3530 (N_3530,N_2661,N_2294);
and U3531 (N_3531,N_2685,N_2908);
and U3532 (N_3532,N_2808,N_2666);
or U3533 (N_3533,N_2355,N_2740);
nor U3534 (N_3534,N_2616,N_2316);
nor U3535 (N_3535,N_2409,N_2280);
and U3536 (N_3536,N_2595,N_2885);
nand U3537 (N_3537,N_2981,N_2320);
nor U3538 (N_3538,N_2298,N_2645);
nor U3539 (N_3539,N_2362,N_2688);
nor U3540 (N_3540,N_2373,N_2878);
nor U3541 (N_3541,N_2912,N_2852);
and U3542 (N_3542,N_2890,N_2336);
nor U3543 (N_3543,N_2595,N_2625);
or U3544 (N_3544,N_2387,N_2702);
nand U3545 (N_3545,N_2377,N_2469);
or U3546 (N_3546,N_2959,N_2708);
and U3547 (N_3547,N_2919,N_2377);
xor U3548 (N_3548,N_2541,N_2362);
nor U3549 (N_3549,N_2727,N_2862);
and U3550 (N_3550,N_2669,N_2663);
nor U3551 (N_3551,N_2577,N_2763);
and U3552 (N_3552,N_2275,N_2303);
nand U3553 (N_3553,N_2608,N_2432);
nor U3554 (N_3554,N_2444,N_2681);
or U3555 (N_3555,N_2304,N_2383);
and U3556 (N_3556,N_2341,N_2888);
xor U3557 (N_3557,N_2943,N_2450);
or U3558 (N_3558,N_2936,N_2741);
or U3559 (N_3559,N_2581,N_2770);
nand U3560 (N_3560,N_2505,N_2360);
and U3561 (N_3561,N_2472,N_2896);
nor U3562 (N_3562,N_2900,N_2686);
or U3563 (N_3563,N_2536,N_2520);
or U3564 (N_3564,N_2775,N_2593);
xor U3565 (N_3565,N_2761,N_2351);
nor U3566 (N_3566,N_2336,N_2814);
nor U3567 (N_3567,N_2637,N_2356);
xor U3568 (N_3568,N_2608,N_2267);
nand U3569 (N_3569,N_2867,N_2511);
or U3570 (N_3570,N_2576,N_2724);
or U3571 (N_3571,N_2751,N_2484);
and U3572 (N_3572,N_2693,N_2372);
or U3573 (N_3573,N_2405,N_2792);
and U3574 (N_3574,N_2741,N_2723);
or U3575 (N_3575,N_2646,N_2872);
nand U3576 (N_3576,N_2732,N_2295);
nor U3577 (N_3577,N_2256,N_2337);
nor U3578 (N_3578,N_2281,N_2636);
and U3579 (N_3579,N_2642,N_2846);
nor U3580 (N_3580,N_2606,N_2803);
xor U3581 (N_3581,N_2656,N_2364);
xor U3582 (N_3582,N_2915,N_2857);
nand U3583 (N_3583,N_2278,N_2867);
nor U3584 (N_3584,N_2970,N_2760);
nand U3585 (N_3585,N_2888,N_2572);
nand U3586 (N_3586,N_2533,N_2690);
nor U3587 (N_3587,N_2619,N_2654);
xnor U3588 (N_3588,N_2731,N_2764);
xnor U3589 (N_3589,N_2890,N_2585);
and U3590 (N_3590,N_2838,N_2727);
or U3591 (N_3591,N_2628,N_2254);
and U3592 (N_3592,N_2728,N_2443);
nand U3593 (N_3593,N_2821,N_2626);
nor U3594 (N_3594,N_2712,N_2319);
nor U3595 (N_3595,N_2254,N_2579);
nand U3596 (N_3596,N_2974,N_2899);
nand U3597 (N_3597,N_2570,N_2834);
nor U3598 (N_3598,N_2515,N_2665);
nand U3599 (N_3599,N_2705,N_2597);
nor U3600 (N_3600,N_2404,N_2876);
nor U3601 (N_3601,N_2664,N_2473);
nor U3602 (N_3602,N_2709,N_2995);
nor U3603 (N_3603,N_2776,N_2305);
or U3604 (N_3604,N_2643,N_2990);
nand U3605 (N_3605,N_2616,N_2758);
xor U3606 (N_3606,N_2788,N_2844);
nor U3607 (N_3607,N_2920,N_2542);
and U3608 (N_3608,N_2572,N_2968);
and U3609 (N_3609,N_2654,N_2983);
or U3610 (N_3610,N_2756,N_2670);
nor U3611 (N_3611,N_2677,N_2852);
nor U3612 (N_3612,N_2810,N_2409);
and U3613 (N_3613,N_2791,N_2436);
xor U3614 (N_3614,N_2492,N_2781);
nand U3615 (N_3615,N_2700,N_2396);
xnor U3616 (N_3616,N_2946,N_2280);
nor U3617 (N_3617,N_2651,N_2703);
or U3618 (N_3618,N_2973,N_2272);
or U3619 (N_3619,N_2528,N_2379);
xor U3620 (N_3620,N_2552,N_2504);
or U3621 (N_3621,N_2488,N_2960);
nand U3622 (N_3622,N_2507,N_2860);
and U3623 (N_3623,N_2355,N_2767);
nor U3624 (N_3624,N_2811,N_2396);
nand U3625 (N_3625,N_2273,N_2338);
nor U3626 (N_3626,N_2483,N_2564);
nand U3627 (N_3627,N_2866,N_2951);
nor U3628 (N_3628,N_2408,N_2852);
and U3629 (N_3629,N_2521,N_2972);
and U3630 (N_3630,N_2397,N_2904);
or U3631 (N_3631,N_2621,N_2499);
or U3632 (N_3632,N_2294,N_2670);
nor U3633 (N_3633,N_2666,N_2488);
xor U3634 (N_3634,N_2931,N_2937);
nor U3635 (N_3635,N_2780,N_2636);
or U3636 (N_3636,N_2402,N_2809);
xor U3637 (N_3637,N_2565,N_2270);
or U3638 (N_3638,N_2266,N_2711);
nand U3639 (N_3639,N_2358,N_2905);
nand U3640 (N_3640,N_2808,N_2388);
xor U3641 (N_3641,N_2934,N_2957);
nand U3642 (N_3642,N_2376,N_2363);
nand U3643 (N_3643,N_2923,N_2372);
nor U3644 (N_3644,N_2443,N_2891);
nand U3645 (N_3645,N_2500,N_2379);
nand U3646 (N_3646,N_2933,N_2351);
and U3647 (N_3647,N_2908,N_2992);
nor U3648 (N_3648,N_2369,N_2626);
or U3649 (N_3649,N_2970,N_2634);
nand U3650 (N_3650,N_2713,N_2549);
nand U3651 (N_3651,N_2921,N_2619);
and U3652 (N_3652,N_2699,N_2962);
or U3653 (N_3653,N_2762,N_2944);
and U3654 (N_3654,N_2575,N_2725);
and U3655 (N_3655,N_2422,N_2339);
nand U3656 (N_3656,N_2958,N_2971);
nor U3657 (N_3657,N_2597,N_2839);
xnor U3658 (N_3658,N_2433,N_2776);
nand U3659 (N_3659,N_2988,N_2773);
nor U3660 (N_3660,N_2973,N_2292);
or U3661 (N_3661,N_2295,N_2250);
nand U3662 (N_3662,N_2429,N_2328);
or U3663 (N_3663,N_2977,N_2605);
nor U3664 (N_3664,N_2969,N_2440);
nand U3665 (N_3665,N_2959,N_2372);
nand U3666 (N_3666,N_2779,N_2598);
xor U3667 (N_3667,N_2841,N_2783);
or U3668 (N_3668,N_2700,N_2438);
xor U3669 (N_3669,N_2959,N_2527);
nor U3670 (N_3670,N_2886,N_2261);
or U3671 (N_3671,N_2725,N_2715);
nor U3672 (N_3672,N_2302,N_2492);
and U3673 (N_3673,N_2993,N_2650);
nand U3674 (N_3674,N_2944,N_2625);
xor U3675 (N_3675,N_2282,N_2858);
and U3676 (N_3676,N_2763,N_2690);
and U3677 (N_3677,N_2764,N_2391);
nand U3678 (N_3678,N_2940,N_2287);
nand U3679 (N_3679,N_2734,N_2730);
nand U3680 (N_3680,N_2918,N_2750);
nor U3681 (N_3681,N_2792,N_2787);
nor U3682 (N_3682,N_2601,N_2785);
or U3683 (N_3683,N_2904,N_2712);
or U3684 (N_3684,N_2552,N_2887);
xnor U3685 (N_3685,N_2438,N_2668);
or U3686 (N_3686,N_2945,N_2744);
xnor U3687 (N_3687,N_2847,N_2401);
nor U3688 (N_3688,N_2411,N_2433);
and U3689 (N_3689,N_2283,N_2381);
and U3690 (N_3690,N_2250,N_2474);
nor U3691 (N_3691,N_2707,N_2861);
nor U3692 (N_3692,N_2580,N_2734);
and U3693 (N_3693,N_2327,N_2493);
nand U3694 (N_3694,N_2599,N_2871);
or U3695 (N_3695,N_2592,N_2938);
and U3696 (N_3696,N_2987,N_2319);
nor U3697 (N_3697,N_2628,N_2371);
and U3698 (N_3698,N_2470,N_2314);
nand U3699 (N_3699,N_2943,N_2547);
and U3700 (N_3700,N_2499,N_2677);
or U3701 (N_3701,N_2979,N_2910);
and U3702 (N_3702,N_2848,N_2940);
nand U3703 (N_3703,N_2861,N_2306);
nand U3704 (N_3704,N_2611,N_2748);
or U3705 (N_3705,N_2532,N_2882);
and U3706 (N_3706,N_2837,N_2744);
or U3707 (N_3707,N_2290,N_2480);
or U3708 (N_3708,N_2936,N_2858);
or U3709 (N_3709,N_2512,N_2887);
or U3710 (N_3710,N_2295,N_2970);
and U3711 (N_3711,N_2367,N_2958);
and U3712 (N_3712,N_2282,N_2260);
or U3713 (N_3713,N_2290,N_2479);
and U3714 (N_3714,N_2397,N_2492);
nand U3715 (N_3715,N_2636,N_2546);
nand U3716 (N_3716,N_2575,N_2859);
xor U3717 (N_3717,N_2408,N_2808);
or U3718 (N_3718,N_2967,N_2645);
or U3719 (N_3719,N_2539,N_2651);
and U3720 (N_3720,N_2856,N_2311);
nand U3721 (N_3721,N_2581,N_2673);
and U3722 (N_3722,N_2735,N_2715);
and U3723 (N_3723,N_2439,N_2698);
nor U3724 (N_3724,N_2844,N_2777);
nor U3725 (N_3725,N_2998,N_2360);
and U3726 (N_3726,N_2574,N_2682);
nand U3727 (N_3727,N_2900,N_2322);
nand U3728 (N_3728,N_2573,N_2901);
or U3729 (N_3729,N_2534,N_2631);
or U3730 (N_3730,N_2533,N_2291);
and U3731 (N_3731,N_2396,N_2570);
nor U3732 (N_3732,N_2714,N_2342);
nor U3733 (N_3733,N_2886,N_2464);
nor U3734 (N_3734,N_2294,N_2362);
nor U3735 (N_3735,N_2603,N_2902);
and U3736 (N_3736,N_2529,N_2966);
and U3737 (N_3737,N_2687,N_2638);
xor U3738 (N_3738,N_2579,N_2864);
or U3739 (N_3739,N_2619,N_2482);
and U3740 (N_3740,N_2545,N_2666);
nand U3741 (N_3741,N_2842,N_2798);
xor U3742 (N_3742,N_2289,N_2835);
or U3743 (N_3743,N_2979,N_2353);
nor U3744 (N_3744,N_2940,N_2901);
xor U3745 (N_3745,N_2674,N_2265);
nand U3746 (N_3746,N_2402,N_2849);
nand U3747 (N_3747,N_2918,N_2317);
and U3748 (N_3748,N_2634,N_2398);
nor U3749 (N_3749,N_2317,N_2690);
xor U3750 (N_3750,N_3101,N_3428);
or U3751 (N_3751,N_3155,N_3073);
or U3752 (N_3752,N_3743,N_3429);
nand U3753 (N_3753,N_3515,N_3041);
and U3754 (N_3754,N_3538,N_3660);
or U3755 (N_3755,N_3489,N_3116);
nand U3756 (N_3756,N_3677,N_3707);
nor U3757 (N_3757,N_3164,N_3220);
or U3758 (N_3758,N_3350,N_3355);
nor U3759 (N_3759,N_3369,N_3390);
or U3760 (N_3760,N_3175,N_3518);
nand U3761 (N_3761,N_3201,N_3718);
nor U3762 (N_3762,N_3023,N_3345);
nor U3763 (N_3763,N_3712,N_3179);
xor U3764 (N_3764,N_3230,N_3208);
and U3765 (N_3765,N_3168,N_3466);
and U3766 (N_3766,N_3348,N_3254);
and U3767 (N_3767,N_3619,N_3323);
nor U3768 (N_3768,N_3587,N_3511);
and U3769 (N_3769,N_3580,N_3464);
or U3770 (N_3770,N_3016,N_3469);
and U3771 (N_3771,N_3359,N_3245);
nor U3772 (N_3772,N_3002,N_3038);
nand U3773 (N_3773,N_3611,N_3652);
nor U3774 (N_3774,N_3338,N_3407);
nor U3775 (N_3775,N_3537,N_3432);
nor U3776 (N_3776,N_3322,N_3276);
and U3777 (N_3777,N_3305,N_3663);
and U3778 (N_3778,N_3271,N_3291);
xnor U3779 (N_3779,N_3681,N_3714);
nand U3780 (N_3780,N_3544,N_3122);
nand U3781 (N_3781,N_3749,N_3118);
or U3782 (N_3782,N_3581,N_3532);
and U3783 (N_3783,N_3410,N_3195);
or U3784 (N_3784,N_3578,N_3702);
and U3785 (N_3785,N_3157,N_3034);
xor U3786 (N_3786,N_3243,N_3411);
nand U3787 (N_3787,N_3653,N_3344);
or U3788 (N_3788,N_3185,N_3402);
and U3789 (N_3789,N_3049,N_3007);
and U3790 (N_3790,N_3232,N_3567);
and U3791 (N_3791,N_3084,N_3723);
and U3792 (N_3792,N_3427,N_3547);
nor U3793 (N_3793,N_3284,N_3146);
nor U3794 (N_3794,N_3439,N_3603);
and U3795 (N_3795,N_3492,N_3747);
nand U3796 (N_3796,N_3512,N_3334);
nand U3797 (N_3797,N_3613,N_3320);
nor U3798 (N_3798,N_3690,N_3337);
nor U3799 (N_3799,N_3301,N_3140);
and U3800 (N_3800,N_3247,N_3459);
or U3801 (N_3801,N_3623,N_3133);
nand U3802 (N_3802,N_3097,N_3566);
nand U3803 (N_3803,N_3374,N_3729);
xor U3804 (N_3804,N_3103,N_3589);
xor U3805 (N_3805,N_3229,N_3187);
and U3806 (N_3806,N_3066,N_3678);
and U3807 (N_3807,N_3599,N_3685);
nand U3808 (N_3808,N_3080,N_3482);
nor U3809 (N_3809,N_3365,N_3533);
or U3810 (N_3810,N_3008,N_3342);
and U3811 (N_3811,N_3377,N_3067);
nor U3812 (N_3812,N_3703,N_3347);
and U3813 (N_3813,N_3394,N_3264);
or U3814 (N_3814,N_3560,N_3025);
and U3815 (N_3815,N_3279,N_3233);
and U3816 (N_3816,N_3558,N_3705);
nor U3817 (N_3817,N_3349,N_3641);
nor U3818 (N_3818,N_3144,N_3015);
nand U3819 (N_3819,N_3311,N_3317);
and U3820 (N_3820,N_3501,N_3632);
nor U3821 (N_3821,N_3591,N_3708);
nor U3822 (N_3822,N_3171,N_3696);
nand U3823 (N_3823,N_3300,N_3620);
xor U3824 (N_3824,N_3078,N_3268);
nor U3825 (N_3825,N_3740,N_3330);
nor U3826 (N_3826,N_3597,N_3687);
nand U3827 (N_3827,N_3044,N_3744);
xnor U3828 (N_3828,N_3564,N_3336);
nand U3829 (N_3829,N_3092,N_3119);
nor U3830 (N_3830,N_3706,N_3403);
or U3831 (N_3831,N_3315,N_3421);
nand U3832 (N_3832,N_3333,N_3106);
nor U3833 (N_3833,N_3412,N_3590);
or U3834 (N_3834,N_3542,N_3277);
and U3835 (N_3835,N_3222,N_3104);
nor U3836 (N_3836,N_3667,N_3585);
nor U3837 (N_3837,N_3594,N_3258);
nand U3838 (N_3838,N_3463,N_3003);
or U3839 (N_3839,N_3543,N_3162);
xor U3840 (N_3840,N_3675,N_3631);
and U3841 (N_3841,N_3438,N_3425);
nand U3842 (N_3842,N_3169,N_3642);
nand U3843 (N_3843,N_3020,N_3443);
and U3844 (N_3844,N_3293,N_3075);
or U3845 (N_3845,N_3527,N_3731);
nand U3846 (N_3846,N_3040,N_3509);
and U3847 (N_3847,N_3151,N_3189);
nor U3848 (N_3848,N_3196,N_3009);
and U3849 (N_3849,N_3433,N_3064);
and U3850 (N_3850,N_3557,N_3269);
or U3851 (N_3851,N_3668,N_3312);
nand U3852 (N_3852,N_3310,N_3375);
nor U3853 (N_3853,N_3191,N_3259);
or U3854 (N_3854,N_3742,N_3689);
nand U3855 (N_3855,N_3513,N_3713);
and U3856 (N_3856,N_3304,N_3329);
nor U3857 (N_3857,N_3741,N_3252);
nor U3858 (N_3858,N_3077,N_3303);
and U3859 (N_3859,N_3528,N_3042);
nand U3860 (N_3860,N_3217,N_3664);
and U3861 (N_3861,N_3462,N_3024);
nand U3862 (N_3862,N_3110,N_3130);
and U3863 (N_3863,N_3123,N_3406);
or U3864 (N_3864,N_3691,N_3161);
and U3865 (N_3865,N_3237,N_3565);
xor U3866 (N_3866,N_3089,N_3121);
or U3867 (N_3867,N_3120,N_3444);
and U3868 (N_3868,N_3070,N_3057);
nor U3869 (N_3869,N_3460,N_3285);
and U3870 (N_3870,N_3672,N_3688);
nand U3871 (N_3871,N_3498,N_3665);
and U3872 (N_3872,N_3088,N_3554);
and U3873 (N_3873,N_3200,N_3090);
or U3874 (N_3874,N_3353,N_3506);
nand U3875 (N_3875,N_3496,N_3658);
and U3876 (N_3876,N_3137,N_3486);
xnor U3877 (N_3877,N_3112,N_3418);
nand U3878 (N_3878,N_3063,N_3056);
and U3879 (N_3879,N_3095,N_3143);
and U3880 (N_3880,N_3399,N_3419);
and U3881 (N_3881,N_3559,N_3408);
or U3882 (N_3882,N_3625,N_3027);
or U3883 (N_3883,N_3280,N_3710);
nor U3884 (N_3884,N_3052,N_3278);
nor U3885 (N_3885,N_3674,N_3636);
and U3886 (N_3886,N_3197,N_3180);
nand U3887 (N_3887,N_3686,N_3746);
and U3888 (N_3888,N_3711,N_3414);
and U3889 (N_3889,N_3286,N_3519);
and U3890 (N_3890,N_3178,N_3210);
nand U3891 (N_3891,N_3628,N_3135);
nand U3892 (N_3892,N_3199,N_3354);
nor U3893 (N_3893,N_3150,N_3129);
xor U3894 (N_3894,N_3176,N_3366);
and U3895 (N_3895,N_3473,N_3572);
nand U3896 (N_3896,N_3423,N_3014);
nand U3897 (N_3897,N_3655,N_3000);
or U3898 (N_3898,N_3649,N_3128);
and U3899 (N_3899,N_3383,N_3733);
nor U3900 (N_3900,N_3540,N_3228);
nor U3901 (N_3901,N_3417,N_3294);
nor U3902 (N_3902,N_3393,N_3577);
nand U3903 (N_3903,N_3194,N_3732);
or U3904 (N_3904,N_3182,N_3454);
xor U3905 (N_3905,N_3522,N_3607);
and U3906 (N_3906,N_3502,N_3673);
or U3907 (N_3907,N_3205,N_3530);
nand U3908 (N_3908,N_3190,N_3319);
and U3909 (N_3909,N_3539,N_3659);
and U3910 (N_3910,N_3306,N_3479);
and U3911 (N_3911,N_3545,N_3562);
or U3912 (N_3912,N_3234,N_3593);
and U3913 (N_3913,N_3270,N_3575);
and U3914 (N_3914,N_3382,N_3299);
or U3915 (N_3915,N_3013,N_3640);
nor U3916 (N_3916,N_3352,N_3721);
nand U3917 (N_3917,N_3477,N_3257);
nor U3918 (N_3918,N_3529,N_3224);
or U3919 (N_3919,N_3435,N_3332);
xor U3920 (N_3920,N_3314,N_3048);
xor U3921 (N_3921,N_3693,N_3316);
or U3922 (N_3922,N_3117,N_3221);
and U3923 (N_3923,N_3505,N_3028);
nor U3924 (N_3924,N_3508,N_3491);
and U3925 (N_3925,N_3216,N_3331);
nand U3926 (N_3926,N_3341,N_3265);
nor U3927 (N_3927,N_3437,N_3618);
xor U3928 (N_3928,N_3494,N_3204);
or U3929 (N_3929,N_3149,N_3574);
nand U3930 (N_3930,N_3029,N_3289);
and U3931 (N_3931,N_3010,N_3346);
nor U3932 (N_3932,N_3249,N_3373);
nand U3933 (N_3933,N_3541,N_3281);
and U3934 (N_3934,N_3376,N_3321);
nor U3935 (N_3935,N_3651,N_3363);
nand U3936 (N_3936,N_3163,N_3629);
xor U3937 (N_3937,N_3563,N_3475);
nor U3938 (N_3938,N_3485,N_3184);
nor U3939 (N_3939,N_3085,N_3065);
and U3940 (N_3940,N_3676,N_3388);
nor U3941 (N_3941,N_3638,N_3592);
nand U3942 (N_3942,N_3440,N_3670);
nor U3943 (N_3943,N_3476,N_3170);
and U3944 (N_3944,N_3186,N_3634);
and U3945 (N_3945,N_3356,N_3380);
nor U3946 (N_3946,N_3364,N_3083);
xnor U3947 (N_3947,N_3596,N_3630);
nand U3948 (N_3948,N_3395,N_3680);
nand U3949 (N_3949,N_3079,N_3141);
nor U3950 (N_3950,N_3134,N_3716);
or U3951 (N_3951,N_3238,N_3679);
or U3952 (N_3952,N_3308,N_3622);
and U3953 (N_3953,N_3614,N_3142);
or U3954 (N_3954,N_3449,N_3131);
and U3955 (N_3955,N_3026,N_3212);
or U3956 (N_3956,N_3017,N_3105);
nor U3957 (N_3957,N_3132,N_3646);
or U3958 (N_3958,N_3461,N_3445);
or U3959 (N_3959,N_3520,N_3521);
xnor U3960 (N_3960,N_3214,N_3692);
nand U3961 (N_3961,N_3213,N_3467);
or U3962 (N_3962,N_3136,N_3627);
xor U3963 (N_3963,N_3384,N_3579);
and U3964 (N_3964,N_3127,N_3188);
nor U3965 (N_3965,N_3236,N_3021);
or U3966 (N_3966,N_3626,N_3416);
or U3967 (N_3967,N_3072,N_3452);
or U3968 (N_3968,N_3608,N_3018);
nand U3969 (N_3969,N_3694,N_3523);
nor U3970 (N_3970,N_3495,N_3061);
nor U3971 (N_3971,N_3602,N_3242);
nand U3972 (N_3972,N_3295,N_3211);
and U3973 (N_3973,N_3173,N_3087);
and U3974 (N_3974,N_3239,N_3076);
xor U3975 (N_3975,N_3569,N_3360);
or U3976 (N_3976,N_3570,N_3071);
or U3977 (N_3977,N_3292,N_3398);
and U3978 (N_3978,N_3296,N_3043);
nand U3979 (N_3979,N_3053,N_3514);
nor U3980 (N_3980,N_3447,N_3177);
and U3981 (N_3981,N_3290,N_3719);
nor U3982 (N_3982,N_3728,N_3682);
and U3983 (N_3983,N_3114,N_3392);
and U3984 (N_3984,N_3448,N_3413);
nor U3985 (N_3985,N_3261,N_3059);
nand U3986 (N_3986,N_3734,N_3225);
and U3987 (N_3987,N_3174,N_3662);
nand U3988 (N_3988,N_3156,N_3493);
xnor U3989 (N_3989,N_3424,N_3550);
nand U3990 (N_3990,N_3643,N_3250);
nand U3991 (N_3991,N_3635,N_3724);
nor U3992 (N_3992,N_3549,N_3487);
nor U3993 (N_3993,N_3441,N_3004);
xor U3994 (N_3994,N_3111,N_3172);
nand U3995 (N_3995,N_3198,N_3039);
nand U3996 (N_3996,N_3288,N_3684);
and U3997 (N_3997,N_3736,N_3096);
nor U3998 (N_3998,N_3209,N_3109);
nand U3999 (N_3999,N_3730,N_3582);
xnor U4000 (N_4000,N_3060,N_3081);
or U4001 (N_4001,N_3046,N_3100);
or U4002 (N_4002,N_3480,N_3650);
and U4003 (N_4003,N_3517,N_3282);
nor U4004 (N_4004,N_3367,N_3094);
xnor U4005 (N_4005,N_3068,N_3241);
nor U4006 (N_4006,N_3192,N_3584);
or U4007 (N_4007,N_3218,N_3586);
nor U4008 (N_4008,N_3704,N_3720);
nand U4009 (N_4009,N_3298,N_3381);
xor U4010 (N_4010,N_3274,N_3166);
nand U4011 (N_4011,N_3255,N_3500);
nand U4012 (N_4012,N_3524,N_3556);
or U4013 (N_4013,N_3102,N_3386);
and U4014 (N_4014,N_3124,N_3054);
nand U4015 (N_4015,N_3555,N_3019);
nand U4016 (N_4016,N_3717,N_3251);
and U4017 (N_4017,N_3573,N_3159);
nand U4018 (N_4018,N_3215,N_3235);
and U4019 (N_4019,N_3051,N_3005);
or U4020 (N_4020,N_3604,N_3307);
nor U4021 (N_4021,N_3656,N_3654);
and U4022 (N_4022,N_3183,N_3260);
xor U4023 (N_4023,N_3372,N_3361);
or U4024 (N_4024,N_3645,N_3450);
and U4025 (N_4025,N_3426,N_3510);
nand U4026 (N_4026,N_3266,N_3490);
xor U4027 (N_4027,N_3516,N_3263);
nand U4028 (N_4028,N_3609,N_3011);
nand U4029 (N_4029,N_3273,N_3551);
and U4030 (N_4030,N_3526,N_3391);
nand U4031 (N_4031,N_3389,N_3203);
nand U4032 (N_4032,N_3093,N_3436);
xnor U4033 (N_4033,N_3605,N_3058);
and U4034 (N_4034,N_3219,N_3326);
nor U4035 (N_4035,N_3644,N_3610);
nand U4036 (N_4036,N_3062,N_3098);
or U4037 (N_4037,N_3154,N_3484);
or U4038 (N_4038,N_3324,N_3193);
and U4039 (N_4039,N_3488,N_3385);
and U4040 (N_4040,N_3616,N_3583);
nor U4041 (N_4041,N_3339,N_3457);
xor U4042 (N_4042,N_3738,N_3465);
and U4043 (N_4043,N_3683,N_3099);
nand U4044 (N_4044,N_3409,N_3357);
nand U4045 (N_4045,N_3006,N_3420);
or U4046 (N_4046,N_3240,N_3158);
nor U4047 (N_4047,N_3091,N_3737);
and U4048 (N_4048,N_3698,N_3576);
and U4049 (N_4049,N_3535,N_3497);
nand U4050 (N_4050,N_3715,N_3253);
or U4051 (N_4051,N_3401,N_3244);
and U4052 (N_4052,N_3726,N_3202);
nand U4053 (N_4053,N_3370,N_3328);
nand U4054 (N_4054,N_3115,N_3455);
xor U4055 (N_4055,N_3297,N_3267);
nor U4056 (N_4056,N_3223,N_3378);
or U4057 (N_4057,N_3325,N_3606);
nand U4058 (N_4058,N_3637,N_3001);
or U4059 (N_4059,N_3481,N_3397);
nor U4060 (N_4060,N_3086,N_3037);
nand U4061 (N_4061,N_3722,N_3368);
and U4062 (N_4062,N_3139,N_3126);
xor U4063 (N_4063,N_3612,N_3032);
xnor U4064 (N_4064,N_3422,N_3165);
or U4065 (N_4065,N_3700,N_3709);
nand U4066 (N_4066,N_3327,N_3335);
nand U4067 (N_4067,N_3451,N_3148);
nand U4068 (N_4068,N_3309,N_3272);
nand U4069 (N_4069,N_3152,N_3145);
nand U4070 (N_4070,N_3167,N_3246);
nor U4071 (N_4071,N_3456,N_3226);
or U4072 (N_4072,N_3400,N_3699);
nand U4073 (N_4073,N_3548,N_3248);
xor U4074 (N_4074,N_3701,N_3181);
nand U4075 (N_4075,N_3313,N_3648);
xor U4076 (N_4076,N_3598,N_3387);
and U4077 (N_4077,N_3047,N_3108);
nor U4078 (N_4078,N_3358,N_3571);
nor U4079 (N_4079,N_3446,N_3621);
and U4080 (N_4080,N_3404,N_3256);
nor U4081 (N_4081,N_3633,N_3525);
nor U4082 (N_4082,N_3262,N_3695);
nand U4083 (N_4083,N_3553,N_3069);
nand U4084 (N_4084,N_3601,N_3035);
and U4085 (N_4085,N_3030,N_3739);
xor U4086 (N_4086,N_3546,N_3478);
nor U4087 (N_4087,N_3458,N_3666);
or U4088 (N_4088,N_3472,N_3470);
nor U4089 (N_4089,N_3206,N_3125);
or U4090 (N_4090,N_3483,N_3735);
nor U4091 (N_4091,N_3405,N_3302);
nor U4092 (N_4092,N_3745,N_3287);
and U4093 (N_4093,N_3534,N_3055);
and U4094 (N_4094,N_3415,N_3022);
and U4095 (N_4095,N_3442,N_3430);
xnor U4096 (N_4096,N_3033,N_3669);
and U4097 (N_4097,N_3207,N_3113);
nor U4098 (N_4098,N_3647,N_3362);
xor U4099 (N_4099,N_3045,N_3138);
and U4100 (N_4100,N_3552,N_3657);
nand U4101 (N_4101,N_3600,N_3318);
or U4102 (N_4102,N_3012,N_3147);
and U4103 (N_4103,N_3697,N_3434);
or U4104 (N_4104,N_3082,N_3160);
xnor U4105 (N_4105,N_3275,N_3499);
nand U4106 (N_4106,N_3351,N_3283);
nand U4107 (N_4107,N_3371,N_3050);
or U4108 (N_4108,N_3615,N_3617);
nor U4109 (N_4109,N_3671,N_3507);
nand U4110 (N_4110,N_3595,N_3074);
nor U4111 (N_4111,N_3340,N_3661);
xnor U4112 (N_4112,N_3468,N_3504);
or U4113 (N_4113,N_3474,N_3036);
xor U4114 (N_4114,N_3624,N_3725);
or U4115 (N_4115,N_3536,N_3727);
nor U4116 (N_4116,N_3343,N_3471);
nor U4117 (N_4117,N_3231,N_3396);
nand U4118 (N_4118,N_3431,N_3561);
or U4119 (N_4119,N_3453,N_3031);
or U4120 (N_4120,N_3588,N_3748);
nand U4121 (N_4121,N_3503,N_3153);
or U4122 (N_4122,N_3531,N_3568);
or U4123 (N_4123,N_3107,N_3639);
nand U4124 (N_4124,N_3227,N_3379);
nand U4125 (N_4125,N_3192,N_3208);
nor U4126 (N_4126,N_3390,N_3631);
or U4127 (N_4127,N_3576,N_3690);
or U4128 (N_4128,N_3079,N_3322);
and U4129 (N_4129,N_3709,N_3679);
xnor U4130 (N_4130,N_3008,N_3688);
and U4131 (N_4131,N_3433,N_3633);
or U4132 (N_4132,N_3554,N_3445);
or U4133 (N_4133,N_3645,N_3009);
or U4134 (N_4134,N_3701,N_3344);
or U4135 (N_4135,N_3320,N_3051);
nor U4136 (N_4136,N_3411,N_3052);
or U4137 (N_4137,N_3433,N_3399);
or U4138 (N_4138,N_3236,N_3669);
or U4139 (N_4139,N_3619,N_3220);
or U4140 (N_4140,N_3413,N_3260);
nand U4141 (N_4141,N_3556,N_3430);
or U4142 (N_4142,N_3460,N_3723);
and U4143 (N_4143,N_3562,N_3313);
and U4144 (N_4144,N_3239,N_3609);
nand U4145 (N_4145,N_3430,N_3022);
xnor U4146 (N_4146,N_3596,N_3736);
and U4147 (N_4147,N_3122,N_3303);
nor U4148 (N_4148,N_3337,N_3314);
or U4149 (N_4149,N_3471,N_3286);
nor U4150 (N_4150,N_3304,N_3459);
nand U4151 (N_4151,N_3575,N_3477);
or U4152 (N_4152,N_3608,N_3702);
nor U4153 (N_4153,N_3504,N_3654);
and U4154 (N_4154,N_3181,N_3685);
nor U4155 (N_4155,N_3430,N_3193);
or U4156 (N_4156,N_3477,N_3380);
and U4157 (N_4157,N_3552,N_3043);
and U4158 (N_4158,N_3050,N_3589);
nand U4159 (N_4159,N_3361,N_3059);
nand U4160 (N_4160,N_3419,N_3692);
nor U4161 (N_4161,N_3392,N_3071);
and U4162 (N_4162,N_3695,N_3037);
and U4163 (N_4163,N_3023,N_3513);
or U4164 (N_4164,N_3331,N_3281);
and U4165 (N_4165,N_3450,N_3011);
or U4166 (N_4166,N_3289,N_3053);
nand U4167 (N_4167,N_3042,N_3114);
nor U4168 (N_4168,N_3023,N_3534);
xnor U4169 (N_4169,N_3607,N_3432);
nand U4170 (N_4170,N_3433,N_3098);
nand U4171 (N_4171,N_3436,N_3263);
and U4172 (N_4172,N_3316,N_3722);
nor U4173 (N_4173,N_3655,N_3557);
or U4174 (N_4174,N_3175,N_3207);
nor U4175 (N_4175,N_3117,N_3111);
xor U4176 (N_4176,N_3578,N_3350);
nor U4177 (N_4177,N_3589,N_3234);
or U4178 (N_4178,N_3706,N_3721);
xor U4179 (N_4179,N_3105,N_3301);
nor U4180 (N_4180,N_3581,N_3286);
nand U4181 (N_4181,N_3336,N_3692);
nand U4182 (N_4182,N_3671,N_3046);
or U4183 (N_4183,N_3489,N_3514);
and U4184 (N_4184,N_3222,N_3032);
or U4185 (N_4185,N_3374,N_3687);
or U4186 (N_4186,N_3573,N_3120);
nor U4187 (N_4187,N_3314,N_3448);
xnor U4188 (N_4188,N_3321,N_3011);
nor U4189 (N_4189,N_3561,N_3655);
nor U4190 (N_4190,N_3736,N_3473);
and U4191 (N_4191,N_3415,N_3101);
and U4192 (N_4192,N_3267,N_3440);
or U4193 (N_4193,N_3334,N_3016);
or U4194 (N_4194,N_3333,N_3125);
or U4195 (N_4195,N_3082,N_3017);
nor U4196 (N_4196,N_3200,N_3304);
and U4197 (N_4197,N_3641,N_3468);
nand U4198 (N_4198,N_3588,N_3452);
nand U4199 (N_4199,N_3363,N_3717);
and U4200 (N_4200,N_3749,N_3477);
nand U4201 (N_4201,N_3107,N_3489);
and U4202 (N_4202,N_3604,N_3516);
and U4203 (N_4203,N_3603,N_3407);
nand U4204 (N_4204,N_3293,N_3144);
or U4205 (N_4205,N_3659,N_3683);
and U4206 (N_4206,N_3101,N_3087);
nand U4207 (N_4207,N_3537,N_3388);
nor U4208 (N_4208,N_3263,N_3227);
and U4209 (N_4209,N_3608,N_3034);
or U4210 (N_4210,N_3089,N_3583);
nor U4211 (N_4211,N_3038,N_3736);
nand U4212 (N_4212,N_3550,N_3333);
nor U4213 (N_4213,N_3045,N_3645);
and U4214 (N_4214,N_3549,N_3142);
nand U4215 (N_4215,N_3296,N_3696);
and U4216 (N_4216,N_3029,N_3362);
nor U4217 (N_4217,N_3069,N_3412);
nand U4218 (N_4218,N_3565,N_3370);
or U4219 (N_4219,N_3219,N_3113);
nor U4220 (N_4220,N_3612,N_3254);
or U4221 (N_4221,N_3662,N_3113);
nor U4222 (N_4222,N_3194,N_3216);
nor U4223 (N_4223,N_3058,N_3665);
or U4224 (N_4224,N_3317,N_3148);
nand U4225 (N_4225,N_3057,N_3711);
nor U4226 (N_4226,N_3496,N_3211);
xnor U4227 (N_4227,N_3053,N_3235);
or U4228 (N_4228,N_3684,N_3734);
nor U4229 (N_4229,N_3178,N_3282);
nand U4230 (N_4230,N_3699,N_3452);
nand U4231 (N_4231,N_3186,N_3311);
nor U4232 (N_4232,N_3617,N_3231);
or U4233 (N_4233,N_3167,N_3444);
and U4234 (N_4234,N_3727,N_3281);
nand U4235 (N_4235,N_3337,N_3735);
xor U4236 (N_4236,N_3242,N_3193);
and U4237 (N_4237,N_3247,N_3117);
nand U4238 (N_4238,N_3021,N_3138);
nand U4239 (N_4239,N_3738,N_3688);
nor U4240 (N_4240,N_3524,N_3499);
or U4241 (N_4241,N_3386,N_3744);
nand U4242 (N_4242,N_3226,N_3743);
nand U4243 (N_4243,N_3276,N_3300);
nand U4244 (N_4244,N_3460,N_3576);
xnor U4245 (N_4245,N_3732,N_3330);
and U4246 (N_4246,N_3528,N_3409);
and U4247 (N_4247,N_3663,N_3419);
and U4248 (N_4248,N_3426,N_3398);
nand U4249 (N_4249,N_3085,N_3194);
and U4250 (N_4250,N_3510,N_3428);
or U4251 (N_4251,N_3234,N_3723);
nor U4252 (N_4252,N_3481,N_3688);
and U4253 (N_4253,N_3352,N_3278);
or U4254 (N_4254,N_3433,N_3525);
and U4255 (N_4255,N_3157,N_3498);
nor U4256 (N_4256,N_3298,N_3258);
nand U4257 (N_4257,N_3379,N_3084);
and U4258 (N_4258,N_3364,N_3504);
nand U4259 (N_4259,N_3438,N_3737);
nor U4260 (N_4260,N_3718,N_3294);
or U4261 (N_4261,N_3523,N_3177);
nor U4262 (N_4262,N_3423,N_3565);
nand U4263 (N_4263,N_3530,N_3655);
nor U4264 (N_4264,N_3164,N_3442);
or U4265 (N_4265,N_3242,N_3295);
or U4266 (N_4266,N_3142,N_3370);
nand U4267 (N_4267,N_3056,N_3358);
and U4268 (N_4268,N_3473,N_3043);
or U4269 (N_4269,N_3172,N_3519);
or U4270 (N_4270,N_3121,N_3351);
and U4271 (N_4271,N_3712,N_3355);
nand U4272 (N_4272,N_3107,N_3387);
nor U4273 (N_4273,N_3195,N_3070);
nand U4274 (N_4274,N_3316,N_3500);
or U4275 (N_4275,N_3587,N_3254);
nor U4276 (N_4276,N_3068,N_3065);
or U4277 (N_4277,N_3435,N_3303);
xnor U4278 (N_4278,N_3301,N_3310);
nor U4279 (N_4279,N_3338,N_3570);
nand U4280 (N_4280,N_3286,N_3544);
nand U4281 (N_4281,N_3666,N_3164);
and U4282 (N_4282,N_3179,N_3175);
and U4283 (N_4283,N_3522,N_3222);
nor U4284 (N_4284,N_3321,N_3192);
or U4285 (N_4285,N_3677,N_3393);
nor U4286 (N_4286,N_3595,N_3645);
and U4287 (N_4287,N_3599,N_3271);
nor U4288 (N_4288,N_3544,N_3451);
nor U4289 (N_4289,N_3100,N_3534);
xor U4290 (N_4290,N_3563,N_3507);
nand U4291 (N_4291,N_3730,N_3205);
nand U4292 (N_4292,N_3267,N_3527);
nor U4293 (N_4293,N_3392,N_3385);
nand U4294 (N_4294,N_3010,N_3537);
nand U4295 (N_4295,N_3551,N_3461);
and U4296 (N_4296,N_3199,N_3682);
or U4297 (N_4297,N_3597,N_3185);
nand U4298 (N_4298,N_3341,N_3268);
nand U4299 (N_4299,N_3513,N_3710);
nor U4300 (N_4300,N_3423,N_3093);
and U4301 (N_4301,N_3404,N_3214);
or U4302 (N_4302,N_3723,N_3423);
or U4303 (N_4303,N_3310,N_3175);
or U4304 (N_4304,N_3307,N_3491);
nor U4305 (N_4305,N_3180,N_3313);
or U4306 (N_4306,N_3126,N_3195);
or U4307 (N_4307,N_3380,N_3235);
xnor U4308 (N_4308,N_3393,N_3556);
or U4309 (N_4309,N_3392,N_3586);
nor U4310 (N_4310,N_3528,N_3076);
nor U4311 (N_4311,N_3251,N_3704);
or U4312 (N_4312,N_3508,N_3356);
nand U4313 (N_4313,N_3100,N_3512);
and U4314 (N_4314,N_3567,N_3010);
nor U4315 (N_4315,N_3031,N_3086);
and U4316 (N_4316,N_3692,N_3586);
and U4317 (N_4317,N_3238,N_3031);
nand U4318 (N_4318,N_3021,N_3175);
or U4319 (N_4319,N_3165,N_3544);
or U4320 (N_4320,N_3411,N_3125);
nor U4321 (N_4321,N_3444,N_3668);
nor U4322 (N_4322,N_3305,N_3525);
nor U4323 (N_4323,N_3593,N_3208);
nand U4324 (N_4324,N_3676,N_3328);
xnor U4325 (N_4325,N_3688,N_3347);
and U4326 (N_4326,N_3223,N_3595);
nor U4327 (N_4327,N_3404,N_3644);
nand U4328 (N_4328,N_3383,N_3693);
and U4329 (N_4329,N_3209,N_3096);
or U4330 (N_4330,N_3493,N_3335);
nor U4331 (N_4331,N_3613,N_3517);
nor U4332 (N_4332,N_3084,N_3198);
or U4333 (N_4333,N_3194,N_3058);
and U4334 (N_4334,N_3346,N_3729);
or U4335 (N_4335,N_3440,N_3348);
and U4336 (N_4336,N_3718,N_3414);
nand U4337 (N_4337,N_3665,N_3393);
and U4338 (N_4338,N_3541,N_3644);
and U4339 (N_4339,N_3519,N_3147);
nor U4340 (N_4340,N_3479,N_3349);
nand U4341 (N_4341,N_3017,N_3561);
or U4342 (N_4342,N_3260,N_3231);
and U4343 (N_4343,N_3422,N_3372);
and U4344 (N_4344,N_3213,N_3731);
nor U4345 (N_4345,N_3578,N_3198);
nor U4346 (N_4346,N_3328,N_3654);
nand U4347 (N_4347,N_3469,N_3349);
or U4348 (N_4348,N_3374,N_3329);
nand U4349 (N_4349,N_3590,N_3209);
nand U4350 (N_4350,N_3667,N_3352);
nor U4351 (N_4351,N_3276,N_3326);
and U4352 (N_4352,N_3466,N_3460);
nor U4353 (N_4353,N_3741,N_3054);
or U4354 (N_4354,N_3303,N_3160);
and U4355 (N_4355,N_3192,N_3644);
and U4356 (N_4356,N_3313,N_3071);
nand U4357 (N_4357,N_3418,N_3644);
xnor U4358 (N_4358,N_3692,N_3618);
xnor U4359 (N_4359,N_3459,N_3391);
nor U4360 (N_4360,N_3147,N_3388);
nand U4361 (N_4361,N_3505,N_3063);
and U4362 (N_4362,N_3164,N_3004);
and U4363 (N_4363,N_3038,N_3082);
nand U4364 (N_4364,N_3366,N_3131);
nand U4365 (N_4365,N_3359,N_3369);
or U4366 (N_4366,N_3639,N_3256);
nand U4367 (N_4367,N_3059,N_3186);
and U4368 (N_4368,N_3387,N_3392);
nor U4369 (N_4369,N_3635,N_3704);
nand U4370 (N_4370,N_3010,N_3122);
nand U4371 (N_4371,N_3547,N_3045);
and U4372 (N_4372,N_3135,N_3391);
nand U4373 (N_4373,N_3246,N_3223);
nor U4374 (N_4374,N_3739,N_3276);
and U4375 (N_4375,N_3070,N_3351);
and U4376 (N_4376,N_3560,N_3749);
nand U4377 (N_4377,N_3281,N_3473);
nor U4378 (N_4378,N_3743,N_3474);
nand U4379 (N_4379,N_3290,N_3693);
or U4380 (N_4380,N_3447,N_3435);
xnor U4381 (N_4381,N_3014,N_3424);
xor U4382 (N_4382,N_3027,N_3006);
or U4383 (N_4383,N_3239,N_3324);
or U4384 (N_4384,N_3142,N_3596);
xor U4385 (N_4385,N_3535,N_3249);
nand U4386 (N_4386,N_3245,N_3100);
and U4387 (N_4387,N_3082,N_3469);
nand U4388 (N_4388,N_3202,N_3043);
xnor U4389 (N_4389,N_3664,N_3168);
xnor U4390 (N_4390,N_3105,N_3217);
nor U4391 (N_4391,N_3622,N_3257);
nor U4392 (N_4392,N_3560,N_3307);
nand U4393 (N_4393,N_3402,N_3425);
or U4394 (N_4394,N_3504,N_3354);
nor U4395 (N_4395,N_3493,N_3101);
nor U4396 (N_4396,N_3143,N_3142);
or U4397 (N_4397,N_3348,N_3570);
xor U4398 (N_4398,N_3353,N_3015);
or U4399 (N_4399,N_3359,N_3079);
nor U4400 (N_4400,N_3695,N_3301);
or U4401 (N_4401,N_3379,N_3612);
nor U4402 (N_4402,N_3036,N_3662);
xor U4403 (N_4403,N_3272,N_3421);
and U4404 (N_4404,N_3603,N_3298);
or U4405 (N_4405,N_3196,N_3488);
xnor U4406 (N_4406,N_3626,N_3342);
nand U4407 (N_4407,N_3487,N_3680);
nand U4408 (N_4408,N_3741,N_3188);
nand U4409 (N_4409,N_3346,N_3107);
or U4410 (N_4410,N_3250,N_3455);
nand U4411 (N_4411,N_3367,N_3291);
nand U4412 (N_4412,N_3230,N_3631);
nand U4413 (N_4413,N_3532,N_3544);
or U4414 (N_4414,N_3574,N_3326);
and U4415 (N_4415,N_3173,N_3163);
nand U4416 (N_4416,N_3617,N_3627);
or U4417 (N_4417,N_3078,N_3015);
nand U4418 (N_4418,N_3237,N_3087);
nor U4419 (N_4419,N_3006,N_3073);
or U4420 (N_4420,N_3230,N_3316);
or U4421 (N_4421,N_3156,N_3548);
or U4422 (N_4422,N_3264,N_3521);
nand U4423 (N_4423,N_3022,N_3425);
nor U4424 (N_4424,N_3348,N_3494);
nand U4425 (N_4425,N_3238,N_3032);
or U4426 (N_4426,N_3549,N_3105);
nand U4427 (N_4427,N_3317,N_3617);
nor U4428 (N_4428,N_3167,N_3515);
and U4429 (N_4429,N_3574,N_3074);
nor U4430 (N_4430,N_3591,N_3005);
nand U4431 (N_4431,N_3500,N_3156);
or U4432 (N_4432,N_3625,N_3201);
and U4433 (N_4433,N_3310,N_3259);
nand U4434 (N_4434,N_3305,N_3388);
or U4435 (N_4435,N_3092,N_3326);
nor U4436 (N_4436,N_3537,N_3671);
nand U4437 (N_4437,N_3452,N_3744);
nand U4438 (N_4438,N_3748,N_3523);
nor U4439 (N_4439,N_3004,N_3741);
nor U4440 (N_4440,N_3609,N_3560);
and U4441 (N_4441,N_3012,N_3507);
nand U4442 (N_4442,N_3273,N_3605);
and U4443 (N_4443,N_3210,N_3722);
nor U4444 (N_4444,N_3485,N_3176);
xnor U4445 (N_4445,N_3482,N_3224);
nor U4446 (N_4446,N_3210,N_3361);
nand U4447 (N_4447,N_3187,N_3425);
nor U4448 (N_4448,N_3494,N_3243);
nand U4449 (N_4449,N_3293,N_3223);
and U4450 (N_4450,N_3221,N_3698);
xnor U4451 (N_4451,N_3613,N_3215);
nand U4452 (N_4452,N_3643,N_3695);
or U4453 (N_4453,N_3285,N_3104);
nand U4454 (N_4454,N_3719,N_3501);
xor U4455 (N_4455,N_3175,N_3223);
nor U4456 (N_4456,N_3225,N_3641);
and U4457 (N_4457,N_3589,N_3302);
nand U4458 (N_4458,N_3122,N_3724);
nor U4459 (N_4459,N_3209,N_3034);
or U4460 (N_4460,N_3389,N_3191);
and U4461 (N_4461,N_3157,N_3699);
and U4462 (N_4462,N_3545,N_3389);
nand U4463 (N_4463,N_3269,N_3399);
or U4464 (N_4464,N_3059,N_3615);
or U4465 (N_4465,N_3702,N_3356);
nor U4466 (N_4466,N_3133,N_3020);
nand U4467 (N_4467,N_3569,N_3242);
nand U4468 (N_4468,N_3117,N_3671);
or U4469 (N_4469,N_3435,N_3094);
and U4470 (N_4470,N_3633,N_3748);
and U4471 (N_4471,N_3565,N_3245);
nand U4472 (N_4472,N_3008,N_3202);
and U4473 (N_4473,N_3640,N_3485);
nand U4474 (N_4474,N_3523,N_3074);
or U4475 (N_4475,N_3375,N_3719);
nor U4476 (N_4476,N_3047,N_3611);
or U4477 (N_4477,N_3239,N_3469);
or U4478 (N_4478,N_3577,N_3237);
and U4479 (N_4479,N_3660,N_3108);
nand U4480 (N_4480,N_3453,N_3175);
xnor U4481 (N_4481,N_3534,N_3436);
nor U4482 (N_4482,N_3114,N_3533);
nor U4483 (N_4483,N_3587,N_3309);
nor U4484 (N_4484,N_3656,N_3489);
nand U4485 (N_4485,N_3659,N_3081);
nor U4486 (N_4486,N_3156,N_3461);
or U4487 (N_4487,N_3711,N_3596);
and U4488 (N_4488,N_3552,N_3015);
or U4489 (N_4489,N_3237,N_3169);
xnor U4490 (N_4490,N_3710,N_3229);
nor U4491 (N_4491,N_3072,N_3719);
and U4492 (N_4492,N_3359,N_3687);
or U4493 (N_4493,N_3672,N_3183);
nand U4494 (N_4494,N_3025,N_3746);
nand U4495 (N_4495,N_3646,N_3602);
nor U4496 (N_4496,N_3020,N_3360);
and U4497 (N_4497,N_3421,N_3216);
xnor U4498 (N_4498,N_3652,N_3415);
nand U4499 (N_4499,N_3234,N_3099);
nand U4500 (N_4500,N_4182,N_4436);
xnor U4501 (N_4501,N_3795,N_4209);
nand U4502 (N_4502,N_4484,N_4289);
nand U4503 (N_4503,N_4453,N_4488);
and U4504 (N_4504,N_4275,N_3937);
nor U4505 (N_4505,N_4213,N_4124);
nand U4506 (N_4506,N_3789,N_4318);
and U4507 (N_4507,N_4022,N_4199);
nor U4508 (N_4508,N_4430,N_3778);
and U4509 (N_4509,N_3934,N_4329);
nand U4510 (N_4510,N_3855,N_4399);
or U4511 (N_4511,N_3926,N_4486);
xnor U4512 (N_4512,N_3935,N_4020);
or U4513 (N_4513,N_3772,N_3792);
nand U4514 (N_4514,N_3894,N_4161);
xor U4515 (N_4515,N_4325,N_4426);
nor U4516 (N_4516,N_4025,N_4372);
nand U4517 (N_4517,N_3785,N_3886);
or U4518 (N_4518,N_4114,N_3774);
and U4519 (N_4519,N_4081,N_3864);
nor U4520 (N_4520,N_4230,N_3884);
nor U4521 (N_4521,N_4193,N_4118);
nor U4522 (N_4522,N_4190,N_4271);
or U4523 (N_4523,N_4464,N_4194);
nor U4524 (N_4524,N_4198,N_3976);
or U4525 (N_4525,N_4013,N_4374);
nor U4526 (N_4526,N_3847,N_4321);
and U4527 (N_4527,N_4274,N_4377);
and U4528 (N_4528,N_4327,N_4168);
nor U4529 (N_4529,N_4273,N_4097);
nor U4530 (N_4530,N_3911,N_3993);
nor U4531 (N_4531,N_4284,N_3907);
nor U4532 (N_4532,N_4137,N_4276);
nor U4533 (N_4533,N_4201,N_4280);
and U4534 (N_4534,N_3912,N_4225);
nor U4535 (N_4535,N_4057,N_4429);
or U4536 (N_4536,N_4195,N_4385);
or U4537 (N_4537,N_4169,N_4203);
nand U4538 (N_4538,N_3764,N_3898);
or U4539 (N_4539,N_3921,N_4078);
and U4540 (N_4540,N_3891,N_3953);
and U4541 (N_4541,N_3844,N_4497);
and U4542 (N_4542,N_4477,N_4317);
and U4543 (N_4543,N_4044,N_4040);
nand U4544 (N_4544,N_4371,N_3834);
nor U4545 (N_4545,N_3905,N_3828);
and U4546 (N_4546,N_4265,N_4499);
or U4547 (N_4547,N_3941,N_3769);
nand U4548 (N_4548,N_4476,N_4031);
and U4549 (N_4549,N_3781,N_4354);
xnor U4550 (N_4550,N_3815,N_3965);
nor U4551 (N_4551,N_3958,N_4299);
or U4552 (N_4552,N_3821,N_4469);
nor U4553 (N_4553,N_4050,N_4128);
or U4554 (N_4554,N_4316,N_4127);
nor U4555 (N_4555,N_4046,N_4247);
and U4556 (N_4556,N_3990,N_3878);
or U4557 (N_4557,N_4266,N_3945);
xnor U4558 (N_4558,N_4360,N_3827);
and U4559 (N_4559,N_3983,N_3869);
and U4560 (N_4560,N_3823,N_4176);
nor U4561 (N_4561,N_4353,N_4177);
and U4562 (N_4562,N_4009,N_4387);
or U4563 (N_4563,N_4140,N_4332);
nand U4564 (N_4564,N_4301,N_4307);
and U4565 (N_4565,N_4438,N_4378);
nor U4566 (N_4566,N_4119,N_3931);
and U4567 (N_4567,N_3752,N_3803);
nor U4568 (N_4568,N_4094,N_4216);
nor U4569 (N_4569,N_4202,N_4223);
nor U4570 (N_4570,N_4441,N_4052);
nand U4571 (N_4571,N_4397,N_3861);
or U4572 (N_4572,N_3845,N_4121);
and U4573 (N_4573,N_3784,N_4063);
xnor U4574 (N_4574,N_4033,N_4181);
nor U4575 (N_4575,N_3811,N_3768);
or U4576 (N_4576,N_4489,N_3924);
and U4577 (N_4577,N_4346,N_3765);
and U4578 (N_4578,N_4041,N_4451);
and U4579 (N_4579,N_4082,N_3751);
nand U4580 (N_4580,N_4328,N_4232);
nor U4581 (N_4581,N_4088,N_3930);
nand U4582 (N_4582,N_3885,N_3824);
nand U4583 (N_4583,N_4465,N_3760);
and U4584 (N_4584,N_4326,N_3881);
nand U4585 (N_4585,N_3996,N_4356);
or U4586 (N_4586,N_3825,N_4262);
or U4587 (N_4587,N_3813,N_3879);
or U4588 (N_4588,N_3988,N_4227);
and U4589 (N_4589,N_4023,N_4229);
nor U4590 (N_4590,N_4028,N_4269);
xor U4591 (N_4591,N_4074,N_4342);
xor U4592 (N_4592,N_4490,N_3977);
and U4593 (N_4593,N_3790,N_4466);
nand U4594 (N_4594,N_3870,N_3757);
and U4595 (N_4595,N_4285,N_4061);
nand U4596 (N_4596,N_3954,N_3853);
nor U4597 (N_4597,N_3978,N_3975);
nand U4598 (N_4598,N_4290,N_4245);
xor U4599 (N_4599,N_4086,N_4416);
nand U4600 (N_4600,N_4334,N_4395);
xor U4601 (N_4601,N_4196,N_4142);
nand U4602 (N_4602,N_4139,N_4300);
or U4603 (N_4603,N_4135,N_4043);
and U4604 (N_4604,N_4092,N_4185);
nor U4605 (N_4605,N_3793,N_3814);
nor U4606 (N_4606,N_4493,N_4107);
and U4607 (N_4607,N_4105,N_4435);
nor U4608 (N_4608,N_3797,N_4011);
and U4609 (N_4609,N_4178,N_4409);
nor U4610 (N_4610,N_4007,N_4206);
and U4611 (N_4611,N_4427,N_4117);
or U4612 (N_4612,N_3948,N_4145);
or U4613 (N_4613,N_4291,N_4143);
and U4614 (N_4614,N_4172,N_4349);
or U4615 (N_4615,N_3857,N_3974);
nand U4616 (N_4616,N_3831,N_3985);
and U4617 (N_4617,N_3997,N_4286);
and U4618 (N_4618,N_3966,N_3848);
nor U4619 (N_4619,N_3806,N_3918);
or U4620 (N_4620,N_4089,N_4101);
nand U4621 (N_4621,N_4446,N_4414);
xor U4622 (N_4622,N_4496,N_4455);
or U4623 (N_4623,N_4208,N_4217);
nand U4624 (N_4624,N_4056,N_3819);
nor U4625 (N_4625,N_4393,N_4123);
xnor U4626 (N_4626,N_4355,N_4298);
nand U4627 (N_4627,N_4174,N_3919);
nand U4628 (N_4628,N_4270,N_3961);
nor U4629 (N_4629,N_3786,N_3892);
nor U4630 (N_4630,N_4037,N_4047);
nor U4631 (N_4631,N_4204,N_4160);
or U4632 (N_4632,N_4001,N_3964);
or U4633 (N_4633,N_4084,N_4062);
nand U4634 (N_4634,N_4019,N_4015);
and U4635 (N_4635,N_4370,N_3759);
nor U4636 (N_4636,N_3807,N_4460);
xor U4637 (N_4637,N_4312,N_4320);
and U4638 (N_4638,N_4345,N_4246);
xor U4639 (N_4639,N_4150,N_3959);
nor U4640 (N_4640,N_4220,N_3908);
nor U4641 (N_4641,N_4153,N_3817);
or U4642 (N_4642,N_4002,N_4151);
nand U4643 (N_4643,N_4381,N_4402);
and U4644 (N_4644,N_4064,N_4361);
or U4645 (N_4645,N_3969,N_4308);
and U4646 (N_4646,N_4159,N_3762);
and U4647 (N_4647,N_4059,N_4167);
xor U4648 (N_4648,N_4411,N_4231);
nor U4649 (N_4649,N_4035,N_4134);
and U4650 (N_4650,N_4066,N_3841);
nand U4651 (N_4651,N_4264,N_4338);
nor U4652 (N_4652,N_4038,N_3856);
or U4653 (N_4653,N_3960,N_4241);
xor U4654 (N_4654,N_4099,N_4417);
and U4655 (N_4655,N_4113,N_4183);
nand U4656 (N_4656,N_4449,N_3780);
nor U4657 (N_4657,N_4406,N_4236);
or U4658 (N_4658,N_4358,N_4205);
nand U4659 (N_4659,N_4483,N_4297);
nor U4660 (N_4660,N_4322,N_4155);
or U4661 (N_4661,N_4122,N_3750);
nor U4662 (N_4662,N_4111,N_4392);
nand U4663 (N_4663,N_3906,N_4164);
or U4664 (N_4664,N_3865,N_4282);
xnor U4665 (N_4665,N_3850,N_4060);
nand U4666 (N_4666,N_3852,N_4260);
or U4667 (N_4667,N_4302,N_4006);
nand U4668 (N_4668,N_3777,N_4344);
nand U4669 (N_4669,N_4014,N_3917);
or U4670 (N_4670,N_3796,N_3810);
or U4671 (N_4671,N_3928,N_4067);
nor U4672 (N_4672,N_4380,N_3899);
or U4673 (N_4673,N_3770,N_3895);
or U4674 (N_4674,N_4261,N_3867);
or U4675 (N_4675,N_4186,N_4303);
or U4676 (N_4676,N_4237,N_4364);
nand U4677 (N_4677,N_4244,N_4003);
nor U4678 (N_4678,N_4224,N_3896);
or U4679 (N_4679,N_3835,N_3830);
or U4680 (N_4680,N_4373,N_4026);
nor U4681 (N_4681,N_4454,N_4382);
xor U4682 (N_4682,N_3859,N_3882);
nand U4683 (N_4683,N_4450,N_4305);
or U4684 (N_4684,N_4075,N_3956);
nor U4685 (N_4685,N_4390,N_3843);
and U4686 (N_4686,N_4173,N_3998);
xnor U4687 (N_4687,N_4422,N_3900);
or U4688 (N_4688,N_4341,N_4045);
nand U4689 (N_4689,N_4333,N_4482);
nand U4690 (N_4690,N_3876,N_3872);
nand U4691 (N_4691,N_3910,N_4188);
nor U4692 (N_4692,N_4238,N_3849);
xor U4693 (N_4693,N_4281,N_3818);
nand U4694 (N_4694,N_3913,N_4295);
or U4695 (N_4695,N_4068,N_4369);
nor U4696 (N_4696,N_4470,N_4310);
and U4697 (N_4697,N_4000,N_3922);
nor U4698 (N_4698,N_4472,N_3897);
nand U4699 (N_4699,N_4085,N_4293);
xor U4700 (N_4700,N_4268,N_4428);
and U4701 (N_4701,N_4279,N_3883);
or U4702 (N_4702,N_3787,N_4407);
nor U4703 (N_4703,N_3967,N_4218);
nor U4704 (N_4704,N_3862,N_4408);
and U4705 (N_4705,N_3950,N_4410);
and U4706 (N_4706,N_3999,N_4481);
nor U4707 (N_4707,N_4386,N_3794);
and U4708 (N_4708,N_4115,N_4027);
or U4709 (N_4709,N_4348,N_4461);
and U4710 (N_4710,N_3986,N_4219);
xor U4711 (N_4711,N_3820,N_4252);
or U4712 (N_4712,N_4263,N_4192);
nor U4713 (N_4713,N_4042,N_4313);
xnor U4714 (N_4714,N_4447,N_4309);
nor U4715 (N_4715,N_4492,N_3758);
nor U4716 (N_4716,N_3779,N_4211);
nor U4717 (N_4717,N_4331,N_4257);
xnor U4718 (N_4718,N_4100,N_4456);
and U4719 (N_4719,N_4368,N_4179);
xor U4720 (N_4720,N_4253,N_3800);
and U4721 (N_4721,N_3763,N_4158);
nor U4722 (N_4722,N_4425,N_3984);
nor U4723 (N_4723,N_4403,N_3868);
nand U4724 (N_4724,N_4288,N_4396);
or U4725 (N_4725,N_3846,N_4259);
or U4726 (N_4726,N_4180,N_3887);
and U4727 (N_4727,N_4440,N_4376);
nor U4728 (N_4728,N_4215,N_4306);
and U4729 (N_4729,N_4251,N_3914);
nand U4730 (N_4730,N_4424,N_4398);
xnor U4731 (N_4731,N_3889,N_4120);
or U4732 (N_4732,N_4383,N_3833);
or U4733 (N_4733,N_4375,N_4187);
or U4734 (N_4734,N_4171,N_4359);
or U4735 (N_4735,N_4444,N_4480);
and U4736 (N_4736,N_3936,N_4352);
nor U4737 (N_4737,N_4112,N_3880);
nor U4738 (N_4738,N_3972,N_4315);
nor U4739 (N_4739,N_4314,N_4207);
nor U4740 (N_4740,N_4255,N_3776);
xor U4741 (N_4741,N_4457,N_4391);
nand U4742 (N_4742,N_4210,N_4498);
and U4743 (N_4743,N_3771,N_4144);
and U4744 (N_4744,N_3920,N_3939);
nor U4745 (N_4745,N_4304,N_4126);
nand U4746 (N_4746,N_3952,N_4077);
or U4747 (N_4747,N_3946,N_4296);
or U4748 (N_4748,N_4110,N_3840);
nor U4749 (N_4749,N_3874,N_4479);
nor U4750 (N_4750,N_3816,N_4283);
and U4751 (N_4751,N_4362,N_3949);
xnor U4752 (N_4752,N_4434,N_4394);
nand U4753 (N_4753,N_4235,N_3863);
or U4754 (N_4754,N_4091,N_4152);
xnor U4755 (N_4755,N_4272,N_4294);
nand U4756 (N_4756,N_4054,N_4221);
or U4757 (N_4757,N_4242,N_4109);
or U4758 (N_4758,N_4175,N_3829);
nor U4759 (N_4759,N_3754,N_3970);
or U4760 (N_4760,N_4149,N_3982);
nand U4761 (N_4761,N_4350,N_3755);
nor U4762 (N_4762,N_4148,N_3812);
xor U4763 (N_4763,N_4228,N_4017);
and U4764 (N_4764,N_4049,N_3851);
nand U4765 (N_4765,N_4292,N_4189);
nor U4766 (N_4766,N_4070,N_4437);
xnor U4767 (N_4767,N_3826,N_3873);
or U4768 (N_4768,N_4065,N_4156);
and U4769 (N_4769,N_4412,N_4367);
nor U4770 (N_4770,N_4423,N_4240);
and U4771 (N_4771,N_4005,N_4039);
and U4772 (N_4772,N_4249,N_3839);
nor U4773 (N_4773,N_3989,N_4339);
nand U4774 (N_4774,N_3842,N_3971);
or U4775 (N_4775,N_4021,N_4365);
or U4776 (N_4776,N_3773,N_4448);
or U4777 (N_4777,N_4443,N_4234);
nor U4778 (N_4778,N_4491,N_4072);
nor U4779 (N_4779,N_4103,N_4384);
and U4780 (N_4780,N_3980,N_4157);
nor U4781 (N_4781,N_4474,N_3890);
and U4782 (N_4782,N_3981,N_4431);
and U4783 (N_4783,N_4467,N_3991);
xnor U4784 (N_4784,N_3963,N_3902);
nor U4785 (N_4785,N_3791,N_3877);
nor U4786 (N_4786,N_3798,N_3901);
nand U4787 (N_4787,N_4330,N_4053);
nand U4788 (N_4788,N_3836,N_4136);
xor U4789 (N_4789,N_4452,N_3909);
nand U4790 (N_4790,N_4130,N_4379);
and U4791 (N_4791,N_3940,N_4093);
nor U4792 (N_4792,N_4125,N_4102);
nor U4793 (N_4793,N_4051,N_4154);
or U4794 (N_4794,N_4404,N_4071);
xor U4795 (N_4795,N_4147,N_4048);
nor U4796 (N_4796,N_4433,N_4413);
xor U4797 (N_4797,N_4058,N_4347);
nor U4798 (N_4798,N_3979,N_4432);
and U4799 (N_4799,N_4162,N_4166);
nor U4800 (N_4800,N_4462,N_4010);
and U4801 (N_4801,N_4233,N_4250);
or U4802 (N_4802,N_3927,N_3955);
or U4803 (N_4803,N_3929,N_3915);
and U4804 (N_4804,N_3822,N_4222);
nor U4805 (N_4805,N_4277,N_4415);
or U4806 (N_4806,N_4095,N_4400);
or U4807 (N_4807,N_4463,N_4098);
or U4808 (N_4808,N_3992,N_4254);
nand U4809 (N_4809,N_3938,N_3944);
and U4810 (N_4810,N_4419,N_4200);
nand U4811 (N_4811,N_4116,N_4267);
and U4812 (N_4812,N_4343,N_3801);
nand U4813 (N_4813,N_4146,N_4494);
nor U4814 (N_4814,N_3962,N_4024);
and U4815 (N_4815,N_4141,N_3947);
and U4816 (N_4816,N_4473,N_4458);
nand U4817 (N_4817,N_4471,N_4165);
nand U4818 (N_4818,N_3957,N_4008);
or U4819 (N_4819,N_4319,N_4106);
and U4820 (N_4820,N_3893,N_4243);
or U4821 (N_4821,N_4468,N_3756);
or U4822 (N_4822,N_4073,N_3923);
or U4823 (N_4823,N_4420,N_3903);
xnor U4824 (N_4824,N_4475,N_3802);
nor U4825 (N_4825,N_4034,N_3808);
nor U4826 (N_4826,N_4018,N_4079);
nor U4827 (N_4827,N_3854,N_3987);
xnor U4828 (N_4828,N_4278,N_4029);
and U4829 (N_4829,N_4004,N_4389);
or U4830 (N_4830,N_3788,N_4340);
nor U4831 (N_4831,N_3933,N_4226);
xor U4832 (N_4832,N_4163,N_3837);
or U4833 (N_4833,N_3766,N_3942);
nor U4834 (N_4834,N_4197,N_4104);
nand U4835 (N_4835,N_3943,N_4248);
or U4836 (N_4836,N_3775,N_3968);
nand U4837 (N_4837,N_4287,N_4323);
nand U4838 (N_4838,N_3875,N_4096);
or U4839 (N_4839,N_3916,N_3871);
nand U4840 (N_4840,N_3866,N_4239);
xor U4841 (N_4841,N_4485,N_4366);
and U4842 (N_4842,N_3838,N_4442);
or U4843 (N_4843,N_4016,N_4030);
and U4844 (N_4844,N_3904,N_3995);
or U4845 (N_4845,N_3805,N_4357);
or U4846 (N_4846,N_4351,N_3761);
xnor U4847 (N_4847,N_4311,N_4214);
nand U4848 (N_4848,N_4459,N_3832);
and U4849 (N_4849,N_4191,N_3925);
or U4850 (N_4850,N_4108,N_4069);
or U4851 (N_4851,N_4401,N_3888);
nand U4852 (N_4852,N_4388,N_4487);
xnor U4853 (N_4853,N_4087,N_4184);
nand U4854 (N_4854,N_4170,N_4076);
nand U4855 (N_4855,N_4258,N_4256);
and U4856 (N_4856,N_3799,N_4036);
or U4857 (N_4857,N_4132,N_4080);
xnor U4858 (N_4858,N_3753,N_3951);
and U4859 (N_4859,N_4133,N_4418);
nand U4860 (N_4860,N_3932,N_4012);
xor U4861 (N_4861,N_3809,N_4055);
nor U4862 (N_4862,N_4131,N_4439);
and U4863 (N_4863,N_4129,N_4336);
nor U4864 (N_4864,N_3860,N_4445);
nand U4865 (N_4865,N_3973,N_4138);
nand U4866 (N_4866,N_4335,N_4212);
or U4867 (N_4867,N_3804,N_4324);
and U4868 (N_4868,N_3994,N_4478);
or U4869 (N_4869,N_3782,N_4032);
nor U4870 (N_4870,N_4405,N_4337);
nor U4871 (N_4871,N_3858,N_4363);
or U4872 (N_4872,N_4090,N_4083);
nand U4873 (N_4873,N_4495,N_3767);
nor U4874 (N_4874,N_4421,N_3783);
nand U4875 (N_4875,N_3921,N_3971);
nand U4876 (N_4876,N_4280,N_4281);
xnor U4877 (N_4877,N_4153,N_4078);
and U4878 (N_4878,N_4353,N_3806);
or U4879 (N_4879,N_4346,N_4006);
nor U4880 (N_4880,N_4392,N_3940);
nor U4881 (N_4881,N_3876,N_3750);
nand U4882 (N_4882,N_4235,N_4185);
nand U4883 (N_4883,N_4048,N_3765);
nand U4884 (N_4884,N_4347,N_4205);
nand U4885 (N_4885,N_4445,N_4383);
nor U4886 (N_4886,N_3882,N_3790);
xor U4887 (N_4887,N_4107,N_4048);
nand U4888 (N_4888,N_3856,N_3767);
or U4889 (N_4889,N_3908,N_3793);
nor U4890 (N_4890,N_3831,N_4488);
or U4891 (N_4891,N_4341,N_4232);
or U4892 (N_4892,N_4412,N_4048);
nand U4893 (N_4893,N_4175,N_3861);
nand U4894 (N_4894,N_4165,N_4259);
and U4895 (N_4895,N_3993,N_3791);
nand U4896 (N_4896,N_3940,N_4046);
xnor U4897 (N_4897,N_4248,N_4243);
nor U4898 (N_4898,N_4087,N_3887);
and U4899 (N_4899,N_3970,N_4055);
and U4900 (N_4900,N_4033,N_3894);
and U4901 (N_4901,N_4341,N_4085);
nor U4902 (N_4902,N_3914,N_4450);
or U4903 (N_4903,N_4454,N_4459);
nor U4904 (N_4904,N_4244,N_4231);
nand U4905 (N_4905,N_3862,N_4094);
or U4906 (N_4906,N_4406,N_4114);
xnor U4907 (N_4907,N_4108,N_3758);
or U4908 (N_4908,N_3880,N_4042);
nor U4909 (N_4909,N_4215,N_4263);
nand U4910 (N_4910,N_4104,N_4375);
nor U4911 (N_4911,N_3753,N_4218);
or U4912 (N_4912,N_4471,N_3940);
nor U4913 (N_4913,N_4175,N_3965);
nor U4914 (N_4914,N_3886,N_3876);
and U4915 (N_4915,N_4188,N_4057);
and U4916 (N_4916,N_4483,N_4099);
or U4917 (N_4917,N_4315,N_4386);
nand U4918 (N_4918,N_3840,N_4216);
or U4919 (N_4919,N_4379,N_4226);
nand U4920 (N_4920,N_3773,N_3942);
xnor U4921 (N_4921,N_4243,N_3910);
nor U4922 (N_4922,N_4335,N_4036);
and U4923 (N_4923,N_3876,N_4148);
and U4924 (N_4924,N_3853,N_3891);
nand U4925 (N_4925,N_3900,N_4204);
nor U4926 (N_4926,N_4203,N_4115);
and U4927 (N_4927,N_4434,N_3860);
or U4928 (N_4928,N_4202,N_4356);
xnor U4929 (N_4929,N_4324,N_4332);
and U4930 (N_4930,N_4395,N_4201);
and U4931 (N_4931,N_4240,N_3892);
or U4932 (N_4932,N_4470,N_4127);
or U4933 (N_4933,N_4298,N_4408);
and U4934 (N_4934,N_3756,N_4182);
and U4935 (N_4935,N_4108,N_4100);
nor U4936 (N_4936,N_3972,N_4137);
nand U4937 (N_4937,N_4443,N_4139);
nor U4938 (N_4938,N_3873,N_3942);
nand U4939 (N_4939,N_3994,N_4096);
nor U4940 (N_4940,N_4029,N_4096);
nor U4941 (N_4941,N_4007,N_4486);
nand U4942 (N_4942,N_4440,N_4478);
or U4943 (N_4943,N_3777,N_3948);
nand U4944 (N_4944,N_3874,N_4348);
nor U4945 (N_4945,N_3808,N_4386);
or U4946 (N_4946,N_3904,N_3932);
and U4947 (N_4947,N_3897,N_4091);
or U4948 (N_4948,N_4435,N_4078);
and U4949 (N_4949,N_3794,N_3919);
or U4950 (N_4950,N_4189,N_4279);
or U4951 (N_4951,N_4186,N_3822);
and U4952 (N_4952,N_4220,N_4363);
xor U4953 (N_4953,N_3754,N_4454);
and U4954 (N_4954,N_4039,N_3872);
nand U4955 (N_4955,N_3996,N_3828);
xor U4956 (N_4956,N_4366,N_3916);
nor U4957 (N_4957,N_4221,N_3978);
and U4958 (N_4958,N_3807,N_4408);
nand U4959 (N_4959,N_4162,N_3936);
nor U4960 (N_4960,N_3763,N_3912);
nor U4961 (N_4961,N_4123,N_4297);
xor U4962 (N_4962,N_3963,N_3898);
nor U4963 (N_4963,N_4181,N_4122);
or U4964 (N_4964,N_4038,N_4393);
xor U4965 (N_4965,N_4091,N_4246);
xnor U4966 (N_4966,N_4177,N_4242);
nor U4967 (N_4967,N_3973,N_3875);
or U4968 (N_4968,N_4154,N_4317);
xnor U4969 (N_4969,N_4141,N_3838);
xnor U4970 (N_4970,N_4238,N_4148);
xnor U4971 (N_4971,N_4445,N_4111);
and U4972 (N_4972,N_4470,N_4064);
nor U4973 (N_4973,N_4052,N_4033);
nor U4974 (N_4974,N_4330,N_3811);
nor U4975 (N_4975,N_4178,N_4300);
nand U4976 (N_4976,N_3750,N_4115);
nor U4977 (N_4977,N_4129,N_4396);
nor U4978 (N_4978,N_4479,N_4379);
nand U4979 (N_4979,N_4379,N_3755);
and U4980 (N_4980,N_4382,N_4190);
and U4981 (N_4981,N_4011,N_3790);
nand U4982 (N_4982,N_4189,N_4358);
and U4983 (N_4983,N_4357,N_3894);
nand U4984 (N_4984,N_3988,N_3899);
or U4985 (N_4985,N_4054,N_4203);
nand U4986 (N_4986,N_4205,N_4299);
or U4987 (N_4987,N_4293,N_4386);
xnor U4988 (N_4988,N_4307,N_4081);
nand U4989 (N_4989,N_4055,N_3998);
nor U4990 (N_4990,N_4211,N_4455);
and U4991 (N_4991,N_4163,N_3818);
nand U4992 (N_4992,N_4203,N_4142);
and U4993 (N_4993,N_3809,N_4133);
nand U4994 (N_4994,N_4297,N_4451);
and U4995 (N_4995,N_3999,N_4169);
or U4996 (N_4996,N_4091,N_3923);
and U4997 (N_4997,N_4152,N_3903);
and U4998 (N_4998,N_4301,N_4250);
nor U4999 (N_4999,N_4356,N_4291);
and U5000 (N_5000,N_4064,N_4439);
nand U5001 (N_5001,N_4349,N_4181);
nor U5002 (N_5002,N_3935,N_4411);
nor U5003 (N_5003,N_4356,N_3941);
xnor U5004 (N_5004,N_4445,N_4164);
or U5005 (N_5005,N_4190,N_3847);
or U5006 (N_5006,N_4098,N_3907);
xor U5007 (N_5007,N_3881,N_4151);
nor U5008 (N_5008,N_3863,N_4133);
nor U5009 (N_5009,N_4146,N_4460);
nor U5010 (N_5010,N_4208,N_3907);
nor U5011 (N_5011,N_4159,N_4481);
nor U5012 (N_5012,N_4265,N_4134);
and U5013 (N_5013,N_4196,N_4206);
or U5014 (N_5014,N_3938,N_4449);
and U5015 (N_5015,N_3956,N_3763);
and U5016 (N_5016,N_4245,N_4337);
and U5017 (N_5017,N_4038,N_4358);
or U5018 (N_5018,N_4487,N_3794);
xor U5019 (N_5019,N_4000,N_3763);
nor U5020 (N_5020,N_3792,N_4311);
xnor U5021 (N_5021,N_4226,N_3752);
xnor U5022 (N_5022,N_3947,N_3873);
and U5023 (N_5023,N_4121,N_4100);
nor U5024 (N_5024,N_4298,N_3905);
nand U5025 (N_5025,N_3954,N_4164);
xnor U5026 (N_5026,N_4166,N_3932);
nand U5027 (N_5027,N_4111,N_4118);
nor U5028 (N_5028,N_4335,N_3879);
and U5029 (N_5029,N_3760,N_4260);
or U5030 (N_5030,N_4357,N_4029);
nor U5031 (N_5031,N_4002,N_4348);
or U5032 (N_5032,N_3926,N_3782);
or U5033 (N_5033,N_4117,N_4035);
and U5034 (N_5034,N_4257,N_4036);
nand U5035 (N_5035,N_3893,N_4488);
nor U5036 (N_5036,N_4268,N_4238);
or U5037 (N_5037,N_4459,N_3905);
or U5038 (N_5038,N_4083,N_4281);
xnor U5039 (N_5039,N_4378,N_3876);
nor U5040 (N_5040,N_3857,N_4128);
and U5041 (N_5041,N_4136,N_3887);
nor U5042 (N_5042,N_3882,N_4252);
nand U5043 (N_5043,N_4209,N_4319);
or U5044 (N_5044,N_4140,N_3992);
and U5045 (N_5045,N_3761,N_4038);
nor U5046 (N_5046,N_4055,N_3764);
or U5047 (N_5047,N_3861,N_3846);
and U5048 (N_5048,N_3903,N_4482);
xnor U5049 (N_5049,N_3909,N_4427);
or U5050 (N_5050,N_3820,N_4119);
and U5051 (N_5051,N_4001,N_3890);
nand U5052 (N_5052,N_4374,N_3919);
and U5053 (N_5053,N_3848,N_4100);
or U5054 (N_5054,N_3759,N_4073);
nor U5055 (N_5055,N_4235,N_3997);
nand U5056 (N_5056,N_4002,N_4017);
and U5057 (N_5057,N_4349,N_4468);
or U5058 (N_5058,N_4384,N_4373);
nand U5059 (N_5059,N_3942,N_3937);
nor U5060 (N_5060,N_4183,N_3904);
or U5061 (N_5061,N_3780,N_4215);
and U5062 (N_5062,N_4244,N_4379);
and U5063 (N_5063,N_4289,N_4360);
nor U5064 (N_5064,N_4396,N_3899);
and U5065 (N_5065,N_3973,N_4261);
and U5066 (N_5066,N_3965,N_3946);
and U5067 (N_5067,N_4319,N_3915);
nand U5068 (N_5068,N_3983,N_3981);
nand U5069 (N_5069,N_3993,N_4149);
nor U5070 (N_5070,N_4011,N_3876);
or U5071 (N_5071,N_4430,N_4065);
and U5072 (N_5072,N_4343,N_4182);
or U5073 (N_5073,N_4215,N_3914);
nor U5074 (N_5074,N_3951,N_4198);
nor U5075 (N_5075,N_4044,N_4125);
nor U5076 (N_5076,N_4160,N_3945);
and U5077 (N_5077,N_4127,N_4267);
and U5078 (N_5078,N_4390,N_4453);
nand U5079 (N_5079,N_4032,N_4174);
nor U5080 (N_5080,N_3894,N_4097);
or U5081 (N_5081,N_4305,N_4215);
or U5082 (N_5082,N_3938,N_4079);
nand U5083 (N_5083,N_3890,N_4134);
and U5084 (N_5084,N_4025,N_3959);
nand U5085 (N_5085,N_3811,N_4058);
nand U5086 (N_5086,N_3824,N_4196);
or U5087 (N_5087,N_4078,N_3792);
xor U5088 (N_5088,N_3829,N_4136);
nor U5089 (N_5089,N_4262,N_3869);
nand U5090 (N_5090,N_3962,N_3804);
or U5091 (N_5091,N_4178,N_3799);
or U5092 (N_5092,N_4155,N_4042);
or U5093 (N_5093,N_3984,N_3888);
and U5094 (N_5094,N_4096,N_4311);
nor U5095 (N_5095,N_4003,N_4134);
and U5096 (N_5096,N_4416,N_4036);
and U5097 (N_5097,N_4231,N_3948);
and U5098 (N_5098,N_4084,N_4325);
and U5099 (N_5099,N_3804,N_4499);
or U5100 (N_5100,N_4010,N_4349);
and U5101 (N_5101,N_3936,N_4423);
and U5102 (N_5102,N_4395,N_4211);
xor U5103 (N_5103,N_4082,N_4366);
and U5104 (N_5104,N_4377,N_4099);
and U5105 (N_5105,N_4223,N_3855);
nor U5106 (N_5106,N_4025,N_4308);
and U5107 (N_5107,N_4494,N_3990);
and U5108 (N_5108,N_4165,N_4210);
nor U5109 (N_5109,N_4467,N_4264);
nand U5110 (N_5110,N_4160,N_4203);
xnor U5111 (N_5111,N_3996,N_3771);
nand U5112 (N_5112,N_4125,N_4201);
and U5113 (N_5113,N_4182,N_4109);
nor U5114 (N_5114,N_4147,N_3894);
nand U5115 (N_5115,N_4467,N_4406);
or U5116 (N_5116,N_4167,N_4285);
nand U5117 (N_5117,N_4395,N_3786);
xnor U5118 (N_5118,N_4306,N_4110);
xor U5119 (N_5119,N_4488,N_4304);
or U5120 (N_5120,N_3758,N_4247);
nand U5121 (N_5121,N_4163,N_4351);
nand U5122 (N_5122,N_3784,N_4357);
or U5123 (N_5123,N_4412,N_4465);
nand U5124 (N_5124,N_3762,N_4049);
and U5125 (N_5125,N_4201,N_4225);
xnor U5126 (N_5126,N_4377,N_4427);
nand U5127 (N_5127,N_4175,N_4298);
nand U5128 (N_5128,N_3755,N_3935);
nor U5129 (N_5129,N_3753,N_4462);
nor U5130 (N_5130,N_4367,N_4466);
or U5131 (N_5131,N_4016,N_3913);
and U5132 (N_5132,N_4363,N_3882);
nor U5133 (N_5133,N_4430,N_4241);
xor U5134 (N_5134,N_3883,N_3894);
or U5135 (N_5135,N_4392,N_4233);
nand U5136 (N_5136,N_4077,N_3921);
or U5137 (N_5137,N_3994,N_3772);
xnor U5138 (N_5138,N_4212,N_4244);
nand U5139 (N_5139,N_4197,N_3763);
xnor U5140 (N_5140,N_3871,N_4356);
nand U5141 (N_5141,N_4042,N_3764);
or U5142 (N_5142,N_4062,N_4159);
nor U5143 (N_5143,N_3943,N_3955);
nand U5144 (N_5144,N_3931,N_4022);
or U5145 (N_5145,N_3894,N_4399);
or U5146 (N_5146,N_4118,N_3805);
and U5147 (N_5147,N_3801,N_3795);
or U5148 (N_5148,N_4066,N_3976);
and U5149 (N_5149,N_4332,N_3752);
xor U5150 (N_5150,N_4141,N_3940);
nor U5151 (N_5151,N_4476,N_4235);
or U5152 (N_5152,N_3861,N_4041);
nand U5153 (N_5153,N_4360,N_3943);
nand U5154 (N_5154,N_3756,N_4494);
nand U5155 (N_5155,N_4244,N_4322);
and U5156 (N_5156,N_3999,N_4258);
nand U5157 (N_5157,N_3853,N_4217);
nand U5158 (N_5158,N_3779,N_4194);
nand U5159 (N_5159,N_4359,N_4060);
and U5160 (N_5160,N_3931,N_4042);
nor U5161 (N_5161,N_4068,N_4005);
nand U5162 (N_5162,N_4239,N_3987);
nor U5163 (N_5163,N_4288,N_4365);
nor U5164 (N_5164,N_4219,N_3990);
and U5165 (N_5165,N_4338,N_4400);
and U5166 (N_5166,N_4074,N_3930);
or U5167 (N_5167,N_4080,N_4053);
and U5168 (N_5168,N_4424,N_3780);
nand U5169 (N_5169,N_4409,N_4244);
and U5170 (N_5170,N_4142,N_4281);
nor U5171 (N_5171,N_4440,N_3812);
and U5172 (N_5172,N_3775,N_4160);
xnor U5173 (N_5173,N_3838,N_4475);
and U5174 (N_5174,N_4024,N_4265);
or U5175 (N_5175,N_3969,N_4123);
nor U5176 (N_5176,N_4243,N_3831);
nand U5177 (N_5177,N_3849,N_4143);
xnor U5178 (N_5178,N_3791,N_4074);
nor U5179 (N_5179,N_4010,N_3812);
or U5180 (N_5180,N_4351,N_4088);
nand U5181 (N_5181,N_4469,N_4028);
or U5182 (N_5182,N_4386,N_4285);
nor U5183 (N_5183,N_3996,N_4337);
and U5184 (N_5184,N_4207,N_4499);
xor U5185 (N_5185,N_3988,N_4435);
and U5186 (N_5186,N_4493,N_4245);
nor U5187 (N_5187,N_4017,N_4280);
or U5188 (N_5188,N_4132,N_4376);
xnor U5189 (N_5189,N_3766,N_4253);
nand U5190 (N_5190,N_3815,N_4074);
nand U5191 (N_5191,N_4297,N_4194);
or U5192 (N_5192,N_4275,N_4499);
nor U5193 (N_5193,N_3816,N_4245);
or U5194 (N_5194,N_4283,N_4044);
xnor U5195 (N_5195,N_4026,N_3761);
nand U5196 (N_5196,N_4159,N_4284);
or U5197 (N_5197,N_3796,N_4327);
and U5198 (N_5198,N_4294,N_4429);
nor U5199 (N_5199,N_3800,N_3769);
nor U5200 (N_5200,N_3801,N_4141);
nand U5201 (N_5201,N_4490,N_3900);
and U5202 (N_5202,N_3837,N_4363);
nand U5203 (N_5203,N_4344,N_3928);
or U5204 (N_5204,N_3764,N_3957);
or U5205 (N_5205,N_4333,N_3917);
nand U5206 (N_5206,N_3935,N_4012);
nor U5207 (N_5207,N_3911,N_3951);
xnor U5208 (N_5208,N_3833,N_4422);
nand U5209 (N_5209,N_3830,N_4459);
or U5210 (N_5210,N_3775,N_3857);
nor U5211 (N_5211,N_3798,N_3866);
or U5212 (N_5212,N_3834,N_3775);
and U5213 (N_5213,N_4412,N_4215);
or U5214 (N_5214,N_4467,N_4090);
or U5215 (N_5215,N_3816,N_4491);
or U5216 (N_5216,N_4466,N_4436);
xnor U5217 (N_5217,N_3976,N_4238);
xor U5218 (N_5218,N_3908,N_3772);
or U5219 (N_5219,N_3812,N_4437);
or U5220 (N_5220,N_4125,N_4006);
nor U5221 (N_5221,N_3853,N_4314);
and U5222 (N_5222,N_4175,N_3804);
and U5223 (N_5223,N_4208,N_4444);
nand U5224 (N_5224,N_4164,N_4452);
xor U5225 (N_5225,N_4384,N_4239);
nor U5226 (N_5226,N_4172,N_4490);
nand U5227 (N_5227,N_3892,N_4400);
nand U5228 (N_5228,N_4130,N_4351);
or U5229 (N_5229,N_4076,N_3961);
and U5230 (N_5230,N_4364,N_4388);
or U5231 (N_5231,N_3934,N_4042);
nor U5232 (N_5232,N_4322,N_4286);
or U5233 (N_5233,N_4332,N_4052);
or U5234 (N_5234,N_3886,N_4141);
nor U5235 (N_5235,N_4445,N_3968);
nand U5236 (N_5236,N_3865,N_4120);
and U5237 (N_5237,N_3836,N_4079);
xnor U5238 (N_5238,N_4291,N_3975);
nor U5239 (N_5239,N_4285,N_3794);
xor U5240 (N_5240,N_4132,N_4030);
nor U5241 (N_5241,N_3820,N_4198);
nand U5242 (N_5242,N_3781,N_4483);
and U5243 (N_5243,N_4304,N_3895);
nor U5244 (N_5244,N_4212,N_4379);
nand U5245 (N_5245,N_4224,N_3970);
or U5246 (N_5246,N_4278,N_3898);
or U5247 (N_5247,N_4258,N_4080);
and U5248 (N_5248,N_3884,N_3955);
nor U5249 (N_5249,N_3827,N_4092);
and U5250 (N_5250,N_4743,N_4919);
nor U5251 (N_5251,N_5215,N_4796);
xor U5252 (N_5252,N_4826,N_4709);
or U5253 (N_5253,N_5248,N_4902);
nand U5254 (N_5254,N_5014,N_5150);
and U5255 (N_5255,N_5249,N_5101);
nor U5256 (N_5256,N_4615,N_5038);
and U5257 (N_5257,N_4819,N_4914);
or U5258 (N_5258,N_5120,N_5035);
nand U5259 (N_5259,N_4752,N_4570);
nor U5260 (N_5260,N_5123,N_4934);
xnor U5261 (N_5261,N_5188,N_4634);
or U5262 (N_5262,N_5110,N_4917);
and U5263 (N_5263,N_4540,N_4921);
or U5264 (N_5264,N_4887,N_4771);
or U5265 (N_5265,N_5133,N_4691);
or U5266 (N_5266,N_4642,N_4616);
nand U5267 (N_5267,N_4674,N_4748);
nor U5268 (N_5268,N_4635,N_4874);
and U5269 (N_5269,N_5136,N_4682);
xnor U5270 (N_5270,N_5121,N_4918);
and U5271 (N_5271,N_5017,N_4988);
or U5272 (N_5272,N_5227,N_4942);
nor U5273 (N_5273,N_4587,N_5082);
or U5274 (N_5274,N_4516,N_5214);
nand U5275 (N_5275,N_5019,N_5238);
and U5276 (N_5276,N_4881,N_5125);
nor U5277 (N_5277,N_5045,N_4555);
nand U5278 (N_5278,N_5029,N_4529);
and U5279 (N_5279,N_5153,N_4823);
nand U5280 (N_5280,N_4590,N_4781);
nor U5281 (N_5281,N_4695,N_4738);
or U5282 (N_5282,N_4624,N_4625);
or U5283 (N_5283,N_4550,N_4611);
nand U5284 (N_5284,N_4613,N_5087);
nand U5285 (N_5285,N_4580,N_5040);
nor U5286 (N_5286,N_4524,N_4993);
or U5287 (N_5287,N_5042,N_4652);
nand U5288 (N_5288,N_5033,N_5034);
nor U5289 (N_5289,N_4564,N_4637);
nor U5290 (N_5290,N_5037,N_4766);
nand U5291 (N_5291,N_5206,N_4872);
and U5292 (N_5292,N_5068,N_5174);
and U5293 (N_5293,N_5050,N_5080);
and U5294 (N_5294,N_5200,N_4744);
nor U5295 (N_5295,N_5043,N_4729);
and U5296 (N_5296,N_4941,N_5086);
nor U5297 (N_5297,N_4757,N_5199);
or U5298 (N_5298,N_4548,N_4617);
and U5299 (N_5299,N_5139,N_4974);
nand U5300 (N_5300,N_5231,N_5218);
nor U5301 (N_5301,N_5084,N_5244);
and U5302 (N_5302,N_5162,N_4523);
nand U5303 (N_5303,N_5220,N_4777);
or U5304 (N_5304,N_5140,N_4649);
nor U5305 (N_5305,N_4556,N_5108);
and U5306 (N_5306,N_4860,N_4711);
nand U5307 (N_5307,N_4601,N_4591);
nor U5308 (N_5308,N_4506,N_4995);
or U5309 (N_5309,N_4970,N_4505);
or U5310 (N_5310,N_5069,N_4639);
and U5311 (N_5311,N_4698,N_4573);
or U5312 (N_5312,N_5224,N_4677);
nor U5313 (N_5313,N_4783,N_5073);
or U5314 (N_5314,N_4996,N_5208);
or U5315 (N_5315,N_4761,N_4673);
nand U5316 (N_5316,N_4700,N_4966);
nand U5317 (N_5317,N_5141,N_5048);
nor U5318 (N_5318,N_5064,N_4630);
or U5319 (N_5319,N_5192,N_4693);
nand U5320 (N_5320,N_4849,N_5142);
nor U5321 (N_5321,N_5147,N_4653);
xor U5322 (N_5322,N_4790,N_4913);
nor U5323 (N_5323,N_5106,N_5189);
nor U5324 (N_5324,N_4904,N_4905);
nor U5325 (N_5325,N_4575,N_4798);
xor U5326 (N_5326,N_4843,N_4769);
nand U5327 (N_5327,N_4685,N_4776);
and U5328 (N_5328,N_4515,N_5122);
xor U5329 (N_5329,N_5118,N_5180);
and U5330 (N_5330,N_4689,N_4727);
nand U5331 (N_5331,N_4560,N_5093);
nand U5332 (N_5332,N_5109,N_4861);
nand U5333 (N_5333,N_4728,N_4694);
or U5334 (N_5334,N_4566,N_4713);
and U5335 (N_5335,N_4663,N_5204);
nor U5336 (N_5336,N_4512,N_4937);
or U5337 (N_5337,N_5222,N_5072);
or U5338 (N_5338,N_5090,N_4539);
or U5339 (N_5339,N_5070,N_4609);
nand U5340 (N_5340,N_4792,N_4971);
nor U5341 (N_5341,N_4507,N_4511);
nand U5342 (N_5342,N_4562,N_4977);
and U5343 (N_5343,N_4811,N_4768);
nand U5344 (N_5344,N_4779,N_4870);
nor U5345 (N_5345,N_5155,N_4871);
nand U5346 (N_5346,N_5132,N_5098);
nor U5347 (N_5347,N_4596,N_4876);
and U5348 (N_5348,N_4712,N_4979);
nand U5349 (N_5349,N_4647,N_5113);
xor U5350 (N_5350,N_4900,N_5060);
nor U5351 (N_5351,N_4985,N_5157);
or U5352 (N_5352,N_4509,N_4845);
nor U5353 (N_5353,N_5210,N_4545);
nor U5354 (N_5354,N_4626,N_5134);
nor U5355 (N_5355,N_4950,N_4862);
nand U5356 (N_5356,N_4910,N_5236);
nand U5357 (N_5357,N_4565,N_4668);
nor U5358 (N_5358,N_4646,N_4754);
nand U5359 (N_5359,N_4620,N_5151);
nand U5360 (N_5360,N_4882,N_4621);
and U5361 (N_5361,N_5237,N_4655);
nor U5362 (N_5362,N_4670,N_5079);
and U5363 (N_5363,N_5004,N_4763);
nand U5364 (N_5364,N_5066,N_4742);
nor U5365 (N_5365,N_4662,N_4922);
nand U5366 (N_5366,N_4954,N_4983);
and U5367 (N_5367,N_5186,N_5177);
nand U5368 (N_5368,N_4561,N_5027);
or U5369 (N_5369,N_4554,N_4851);
or U5370 (N_5370,N_4707,N_4878);
or U5371 (N_5371,N_4820,N_4579);
or U5372 (N_5372,N_4852,N_4806);
nand U5373 (N_5373,N_5041,N_4794);
and U5374 (N_5374,N_5107,N_4880);
or U5375 (N_5375,N_4657,N_4961);
nor U5376 (N_5376,N_4734,N_4873);
or U5377 (N_5377,N_5225,N_5197);
or U5378 (N_5378,N_4514,N_4602);
nand U5379 (N_5379,N_5007,N_4726);
and U5380 (N_5380,N_4583,N_5239);
and U5381 (N_5381,N_4672,N_4925);
nand U5382 (N_5382,N_4931,N_4844);
nor U5383 (N_5383,N_4574,N_5124);
and U5384 (N_5384,N_4800,N_4999);
or U5385 (N_5385,N_4518,N_4740);
and U5386 (N_5386,N_5047,N_5058);
or U5387 (N_5387,N_4537,N_5053);
or U5388 (N_5388,N_4903,N_4594);
nand U5389 (N_5389,N_4853,N_4864);
nor U5390 (N_5390,N_4618,N_5002);
nand U5391 (N_5391,N_5112,N_4643);
or U5392 (N_5392,N_4830,N_4607);
or U5393 (N_5393,N_5209,N_4541);
or U5394 (N_5394,N_4708,N_4839);
and U5395 (N_5395,N_4915,N_5097);
or U5396 (N_5396,N_5039,N_4553);
nand U5397 (N_5397,N_4972,N_4586);
nor U5398 (N_5398,N_5100,N_4532);
or U5399 (N_5399,N_5005,N_5001);
or U5400 (N_5400,N_4892,N_4759);
nand U5401 (N_5401,N_4868,N_4891);
nor U5402 (N_5402,N_5078,N_4517);
nor U5403 (N_5403,N_4940,N_4821);
nand U5404 (N_5404,N_4986,N_4718);
or U5405 (N_5405,N_4831,N_4731);
and U5406 (N_5406,N_5016,N_4628);
nor U5407 (N_5407,N_4890,N_4948);
and U5408 (N_5408,N_4723,N_5051);
nand U5409 (N_5409,N_5116,N_5065);
or U5410 (N_5410,N_4536,N_5193);
xor U5411 (N_5411,N_4701,N_4837);
xor U5412 (N_5412,N_4846,N_4510);
and U5413 (N_5413,N_4982,N_4756);
or U5414 (N_5414,N_4577,N_5143);
nand U5415 (N_5415,N_4714,N_4807);
nand U5416 (N_5416,N_4725,N_5104);
nand U5417 (N_5417,N_5091,N_5171);
nor U5418 (N_5418,N_4688,N_4936);
or U5419 (N_5419,N_4829,N_4666);
and U5420 (N_5420,N_4895,N_5025);
xor U5421 (N_5421,N_5196,N_4508);
and U5422 (N_5422,N_4667,N_4664);
nor U5423 (N_5423,N_4863,N_5102);
nor U5424 (N_5424,N_4906,N_4916);
nand U5425 (N_5425,N_5096,N_5075);
nor U5426 (N_5426,N_5031,N_4824);
nor U5427 (N_5427,N_5198,N_4745);
nor U5428 (N_5428,N_5182,N_4648);
xnor U5429 (N_5429,N_4683,N_4894);
nand U5430 (N_5430,N_5088,N_5081);
nand U5431 (N_5431,N_4658,N_4981);
nand U5432 (N_5432,N_4962,N_4678);
nor U5433 (N_5433,N_4669,N_5240);
nand U5434 (N_5434,N_5063,N_5074);
and U5435 (N_5435,N_4885,N_4593);
nor U5436 (N_5436,N_5149,N_4558);
nand U5437 (N_5437,N_4651,N_4592);
or U5438 (N_5438,N_4595,N_5030);
nor U5439 (N_5439,N_4889,N_5135);
nor U5440 (N_5440,N_4793,N_4773);
or U5441 (N_5441,N_4968,N_4797);
and U5442 (N_5442,N_4912,N_4841);
xnor U5443 (N_5443,N_4681,N_4907);
nor U5444 (N_5444,N_5213,N_4526);
nand U5445 (N_5445,N_4928,N_5178);
or U5446 (N_5446,N_4898,N_4867);
xor U5447 (N_5447,N_4676,N_4959);
nand U5448 (N_5448,N_5216,N_5006);
nand U5449 (N_5449,N_5168,N_5115);
or U5450 (N_5450,N_4866,N_5181);
xor U5451 (N_5451,N_4946,N_4716);
nor U5452 (N_5452,N_4927,N_4960);
nor U5453 (N_5453,N_4782,N_5241);
and U5454 (N_5454,N_4632,N_5023);
and U5455 (N_5455,N_4786,N_4608);
nor U5456 (N_5456,N_4930,N_4998);
nand U5457 (N_5457,N_4973,N_4834);
or U5458 (N_5458,N_4569,N_5146);
or U5459 (N_5459,N_4814,N_4785);
or U5460 (N_5460,N_4772,N_5242);
nor U5461 (N_5461,N_4705,N_5137);
or U5462 (N_5462,N_4645,N_4513);
nor U5463 (N_5463,N_5011,N_4947);
or U5464 (N_5464,N_4854,N_5183);
nand U5465 (N_5465,N_5211,N_4945);
nor U5466 (N_5466,N_4546,N_4584);
nand U5467 (N_5467,N_4717,N_4957);
or U5468 (N_5468,N_4568,N_4875);
xnor U5469 (N_5469,N_5128,N_4544);
nand U5470 (N_5470,N_4893,N_5228);
nand U5471 (N_5471,N_4969,N_4578);
nand U5472 (N_5472,N_5057,N_4629);
nand U5473 (N_5473,N_4938,N_4721);
and U5474 (N_5474,N_4665,N_5169);
nand U5475 (N_5475,N_4789,N_5020);
xor U5476 (N_5476,N_4774,N_4758);
or U5477 (N_5477,N_4675,N_4877);
and U5478 (N_5478,N_5232,N_4746);
nor U5479 (N_5479,N_4987,N_5164);
and U5480 (N_5480,N_4963,N_4932);
nand U5481 (N_5481,N_4799,N_4519);
nand U5482 (N_5482,N_4636,N_4528);
nand U5483 (N_5483,N_5009,N_4585);
and U5484 (N_5484,N_4901,N_5159);
and U5485 (N_5485,N_4775,N_4842);
or U5486 (N_5486,N_5067,N_4531);
and U5487 (N_5487,N_4816,N_4989);
nand U5488 (N_5488,N_4732,N_4965);
nand U5489 (N_5489,N_4804,N_4589);
xor U5490 (N_5490,N_5148,N_4612);
or U5491 (N_5491,N_4680,N_4808);
or U5492 (N_5492,N_5233,N_4502);
or U5493 (N_5493,N_4984,N_4755);
or U5494 (N_5494,N_4690,N_4840);
and U5495 (N_5495,N_4598,N_4992);
nor U5496 (N_5496,N_5175,N_4956);
or U5497 (N_5497,N_5046,N_4503);
nor U5498 (N_5498,N_4563,N_5145);
and U5499 (N_5499,N_4627,N_4770);
and U5500 (N_5500,N_4660,N_4722);
and U5501 (N_5501,N_5000,N_4739);
nand U5502 (N_5502,N_4911,N_5117);
xnor U5503 (N_5503,N_4610,N_5217);
nand U5504 (N_5504,N_4920,N_5094);
nand U5505 (N_5505,N_5126,N_4836);
xor U5506 (N_5506,N_5187,N_4838);
nand U5507 (N_5507,N_4733,N_4538);
nand U5508 (N_5508,N_4850,N_5172);
nor U5509 (N_5509,N_4813,N_4780);
nor U5510 (N_5510,N_5201,N_4967);
nand U5511 (N_5511,N_5085,N_4525);
and U5512 (N_5512,N_5179,N_5173);
or U5513 (N_5513,N_4522,N_4958);
nor U5514 (N_5514,N_4704,N_4933);
and U5515 (N_5515,N_5076,N_5077);
nand U5516 (N_5516,N_5026,N_4926);
and U5517 (N_5517,N_5083,N_5156);
nor U5518 (N_5518,N_5203,N_4671);
and U5519 (N_5519,N_5246,N_4855);
nand U5520 (N_5520,N_4879,N_4687);
or U5521 (N_5521,N_4812,N_4869);
and U5522 (N_5522,N_4784,N_5119);
nor U5523 (N_5523,N_5158,N_5165);
xnor U5524 (N_5524,N_4848,N_4990);
xor U5525 (N_5525,N_4749,N_4500);
and U5526 (N_5526,N_4815,N_4883);
nand U5527 (N_5527,N_4659,N_4765);
or U5528 (N_5528,N_4661,N_4650);
nand U5529 (N_5529,N_4788,N_5219);
or U5530 (N_5530,N_4527,N_5221);
and U5531 (N_5531,N_5202,N_4521);
nor U5532 (N_5532,N_4778,N_4818);
nor U5533 (N_5533,N_4935,N_4571);
nor U5534 (N_5534,N_4923,N_4543);
xnor U5535 (N_5535,N_5127,N_4559);
and U5536 (N_5536,N_4994,N_4857);
and U5537 (N_5537,N_5247,N_4715);
or U5538 (N_5538,N_4787,N_5138);
nor U5539 (N_5539,N_4603,N_4640);
or U5540 (N_5540,N_4549,N_4735);
nor U5541 (N_5541,N_4805,N_4638);
nor U5542 (N_5542,N_4856,N_4547);
or U5543 (N_5543,N_5207,N_4572);
or U5544 (N_5544,N_5095,N_4817);
nand U5545 (N_5545,N_5099,N_4710);
nor U5546 (N_5546,N_4588,N_5195);
or U5547 (N_5547,N_5061,N_4750);
and U5548 (N_5548,N_5130,N_4978);
or U5549 (N_5549,N_5022,N_4832);
and U5550 (N_5550,N_5163,N_4501);
or U5551 (N_5551,N_5185,N_4767);
nand U5552 (N_5552,N_4802,N_4795);
or U5553 (N_5553,N_5028,N_4847);
xor U5554 (N_5554,N_5154,N_4741);
or U5555 (N_5555,N_4753,N_5089);
or U5556 (N_5556,N_4827,N_4614);
xnor U5557 (N_5557,N_4599,N_5167);
xor U5558 (N_5558,N_5191,N_4929);
or U5559 (N_5559,N_4896,N_4654);
or U5560 (N_5560,N_5166,N_4825);
or U5561 (N_5561,N_5036,N_4949);
nand U5562 (N_5562,N_4633,N_5092);
and U5563 (N_5563,N_4801,N_4530);
xor U5564 (N_5564,N_4909,N_4686);
and U5565 (N_5565,N_4888,N_4952);
nor U5566 (N_5566,N_4858,N_4943);
nand U5567 (N_5567,N_4809,N_5024);
nor U5568 (N_5568,N_4542,N_4597);
nor U5569 (N_5569,N_4703,N_5008);
nor U5570 (N_5570,N_4600,N_5144);
nand U5571 (N_5571,N_4697,N_5071);
or U5572 (N_5572,N_4623,N_4833);
and U5573 (N_5573,N_4533,N_4899);
nor U5574 (N_5574,N_5054,N_4656);
xor U5575 (N_5575,N_4641,N_4760);
nand U5576 (N_5576,N_5230,N_5111);
nor U5577 (N_5577,N_4803,N_4619);
or U5578 (N_5578,N_4581,N_4822);
nand U5579 (N_5579,N_4737,N_5049);
nor U5580 (N_5580,N_5184,N_4764);
xor U5581 (N_5581,N_4730,N_5161);
and U5582 (N_5582,N_5160,N_4762);
or U5583 (N_5583,N_5131,N_5235);
and U5584 (N_5584,N_5013,N_5018);
nor U5585 (N_5585,N_5176,N_4865);
or U5586 (N_5586,N_4859,N_5056);
nand U5587 (N_5587,N_4719,N_5015);
nand U5588 (N_5588,N_4751,N_4720);
nand U5589 (N_5589,N_5194,N_5234);
or U5590 (N_5590,N_4706,N_5223);
nor U5591 (N_5591,N_4828,N_4535);
nand U5592 (N_5592,N_5190,N_4810);
nand U5593 (N_5593,N_4534,N_5170);
nand U5594 (N_5594,N_4997,N_4884);
nand U5595 (N_5595,N_4897,N_4622);
and U5596 (N_5596,N_4520,N_4551);
and U5597 (N_5597,N_4953,N_4631);
or U5598 (N_5598,N_4702,N_5062);
nand U5599 (N_5599,N_4976,N_4975);
nor U5600 (N_5600,N_4576,N_5003);
or U5601 (N_5601,N_4939,N_4606);
or U5602 (N_5602,N_5044,N_4724);
and U5603 (N_5603,N_4582,N_4679);
nand U5604 (N_5604,N_5059,N_4886);
and U5605 (N_5605,N_5212,N_5103);
nand U5606 (N_5606,N_5012,N_5052);
nor U5607 (N_5607,N_4908,N_5226);
nor U5608 (N_5608,N_4991,N_4699);
nand U5609 (N_5609,N_5055,N_4504);
nor U5610 (N_5610,N_4951,N_4604);
and U5611 (N_5611,N_4964,N_4696);
or U5612 (N_5612,N_4567,N_4736);
or U5613 (N_5613,N_5021,N_5032);
and U5614 (N_5614,N_4835,N_4955);
xor U5615 (N_5615,N_4747,N_5229);
or U5616 (N_5616,N_4692,N_5105);
nor U5617 (N_5617,N_4791,N_4684);
and U5618 (N_5618,N_5114,N_5152);
xnor U5619 (N_5619,N_5010,N_5243);
nor U5620 (N_5620,N_5205,N_4980);
nand U5621 (N_5621,N_4644,N_4944);
nor U5622 (N_5622,N_4605,N_5129);
nor U5623 (N_5623,N_5245,N_4557);
and U5624 (N_5624,N_4924,N_4552);
xnor U5625 (N_5625,N_5240,N_5000);
nor U5626 (N_5626,N_5034,N_5014);
and U5627 (N_5627,N_4780,N_5086);
or U5628 (N_5628,N_5099,N_4910);
and U5629 (N_5629,N_5212,N_5055);
and U5630 (N_5630,N_4937,N_4511);
nor U5631 (N_5631,N_4672,N_5010);
nor U5632 (N_5632,N_4621,N_4676);
nand U5633 (N_5633,N_4966,N_5078);
xnor U5634 (N_5634,N_4958,N_5029);
and U5635 (N_5635,N_4561,N_4925);
and U5636 (N_5636,N_4937,N_4939);
nand U5637 (N_5637,N_4539,N_4568);
and U5638 (N_5638,N_5018,N_4732);
and U5639 (N_5639,N_4669,N_4754);
or U5640 (N_5640,N_4595,N_4644);
and U5641 (N_5641,N_4742,N_5174);
nand U5642 (N_5642,N_5230,N_4663);
nor U5643 (N_5643,N_4656,N_4566);
nand U5644 (N_5644,N_4933,N_4811);
nor U5645 (N_5645,N_4882,N_4574);
or U5646 (N_5646,N_5075,N_5128);
and U5647 (N_5647,N_4688,N_4649);
xor U5648 (N_5648,N_5190,N_5027);
or U5649 (N_5649,N_5117,N_4994);
nor U5650 (N_5650,N_4672,N_5040);
and U5651 (N_5651,N_4944,N_5026);
nor U5652 (N_5652,N_5081,N_5140);
nor U5653 (N_5653,N_4682,N_4857);
or U5654 (N_5654,N_4630,N_4979);
and U5655 (N_5655,N_5249,N_4712);
or U5656 (N_5656,N_4897,N_4953);
and U5657 (N_5657,N_4652,N_4744);
nand U5658 (N_5658,N_4643,N_4795);
xnor U5659 (N_5659,N_5220,N_5225);
and U5660 (N_5660,N_5151,N_4903);
nand U5661 (N_5661,N_5139,N_5053);
nor U5662 (N_5662,N_5243,N_4509);
xnor U5663 (N_5663,N_4523,N_5033);
and U5664 (N_5664,N_4598,N_4588);
nor U5665 (N_5665,N_4728,N_4834);
and U5666 (N_5666,N_4961,N_4621);
and U5667 (N_5667,N_4703,N_4927);
nand U5668 (N_5668,N_5239,N_5231);
and U5669 (N_5669,N_4912,N_5158);
nand U5670 (N_5670,N_5193,N_4635);
nor U5671 (N_5671,N_4939,N_4592);
nor U5672 (N_5672,N_4893,N_4625);
nand U5673 (N_5673,N_4571,N_4595);
and U5674 (N_5674,N_4956,N_4547);
and U5675 (N_5675,N_4822,N_4843);
nand U5676 (N_5676,N_4897,N_4884);
nand U5677 (N_5677,N_4558,N_4809);
or U5678 (N_5678,N_5168,N_4823);
xnor U5679 (N_5679,N_5218,N_4889);
or U5680 (N_5680,N_5125,N_4624);
nand U5681 (N_5681,N_4922,N_4897);
nand U5682 (N_5682,N_4650,N_5068);
or U5683 (N_5683,N_4690,N_4713);
nand U5684 (N_5684,N_4727,N_4730);
nor U5685 (N_5685,N_4999,N_4733);
nand U5686 (N_5686,N_5117,N_4794);
nor U5687 (N_5687,N_4990,N_4648);
xnor U5688 (N_5688,N_4914,N_4528);
or U5689 (N_5689,N_4762,N_4555);
or U5690 (N_5690,N_5056,N_5188);
nand U5691 (N_5691,N_4734,N_4905);
or U5692 (N_5692,N_5007,N_5037);
and U5693 (N_5693,N_4780,N_4686);
and U5694 (N_5694,N_5005,N_5042);
or U5695 (N_5695,N_4709,N_5059);
nor U5696 (N_5696,N_4947,N_4526);
and U5697 (N_5697,N_4655,N_4581);
or U5698 (N_5698,N_4722,N_4794);
or U5699 (N_5699,N_4992,N_4779);
nand U5700 (N_5700,N_4936,N_4831);
nand U5701 (N_5701,N_5016,N_4813);
nand U5702 (N_5702,N_4731,N_4957);
and U5703 (N_5703,N_5050,N_5161);
and U5704 (N_5704,N_4915,N_4953);
or U5705 (N_5705,N_4823,N_5154);
or U5706 (N_5706,N_5055,N_4736);
or U5707 (N_5707,N_4719,N_5082);
nand U5708 (N_5708,N_4810,N_5177);
and U5709 (N_5709,N_5226,N_4988);
nor U5710 (N_5710,N_4983,N_5147);
or U5711 (N_5711,N_5048,N_4985);
nand U5712 (N_5712,N_4793,N_4692);
xnor U5713 (N_5713,N_4981,N_5004);
and U5714 (N_5714,N_4803,N_4940);
nor U5715 (N_5715,N_5091,N_4776);
or U5716 (N_5716,N_4927,N_4800);
and U5717 (N_5717,N_5230,N_5007);
nor U5718 (N_5718,N_5010,N_4922);
xor U5719 (N_5719,N_4999,N_4707);
and U5720 (N_5720,N_4530,N_4649);
nand U5721 (N_5721,N_4621,N_5093);
nand U5722 (N_5722,N_5233,N_4622);
nor U5723 (N_5723,N_4907,N_4997);
or U5724 (N_5724,N_5092,N_4889);
or U5725 (N_5725,N_5124,N_4524);
nor U5726 (N_5726,N_5130,N_5184);
xor U5727 (N_5727,N_4937,N_4715);
or U5728 (N_5728,N_5008,N_4863);
and U5729 (N_5729,N_4607,N_4934);
or U5730 (N_5730,N_5248,N_4711);
and U5731 (N_5731,N_4773,N_4630);
or U5732 (N_5732,N_5165,N_4600);
and U5733 (N_5733,N_4999,N_5069);
or U5734 (N_5734,N_4813,N_5208);
and U5735 (N_5735,N_5067,N_5127);
nand U5736 (N_5736,N_5170,N_5092);
nand U5737 (N_5737,N_4797,N_4973);
nand U5738 (N_5738,N_5184,N_5072);
or U5739 (N_5739,N_4704,N_4731);
nor U5740 (N_5740,N_4588,N_4877);
and U5741 (N_5741,N_5043,N_5046);
or U5742 (N_5742,N_4526,N_4723);
xor U5743 (N_5743,N_4730,N_5202);
nor U5744 (N_5744,N_4883,N_4849);
and U5745 (N_5745,N_4969,N_4506);
nand U5746 (N_5746,N_5011,N_5158);
xor U5747 (N_5747,N_4734,N_5090);
and U5748 (N_5748,N_4670,N_4578);
and U5749 (N_5749,N_4652,N_4997);
nor U5750 (N_5750,N_4996,N_4924);
or U5751 (N_5751,N_5021,N_4728);
nand U5752 (N_5752,N_5087,N_5042);
nor U5753 (N_5753,N_4550,N_4904);
and U5754 (N_5754,N_4875,N_4779);
or U5755 (N_5755,N_4522,N_4524);
or U5756 (N_5756,N_5101,N_5215);
and U5757 (N_5757,N_5124,N_5155);
nor U5758 (N_5758,N_5093,N_4604);
or U5759 (N_5759,N_4807,N_5090);
and U5760 (N_5760,N_4866,N_4549);
nor U5761 (N_5761,N_4762,N_4901);
or U5762 (N_5762,N_5017,N_4634);
or U5763 (N_5763,N_5170,N_4760);
or U5764 (N_5764,N_5148,N_4705);
nand U5765 (N_5765,N_5044,N_4681);
nor U5766 (N_5766,N_5019,N_4657);
nor U5767 (N_5767,N_4629,N_5195);
and U5768 (N_5768,N_5214,N_5234);
xor U5769 (N_5769,N_5000,N_5004);
nand U5770 (N_5770,N_4865,N_4651);
or U5771 (N_5771,N_5107,N_5177);
nor U5772 (N_5772,N_5061,N_4604);
and U5773 (N_5773,N_4696,N_4516);
or U5774 (N_5774,N_5077,N_4920);
nand U5775 (N_5775,N_4755,N_5014);
nand U5776 (N_5776,N_4555,N_4571);
xor U5777 (N_5777,N_5001,N_4524);
nor U5778 (N_5778,N_4719,N_4906);
nand U5779 (N_5779,N_4544,N_5200);
nor U5780 (N_5780,N_5078,N_5088);
and U5781 (N_5781,N_4643,N_5064);
nor U5782 (N_5782,N_4540,N_4832);
nand U5783 (N_5783,N_5184,N_4969);
nor U5784 (N_5784,N_4634,N_4592);
or U5785 (N_5785,N_4592,N_5035);
nor U5786 (N_5786,N_5072,N_5189);
xor U5787 (N_5787,N_4741,N_4571);
nand U5788 (N_5788,N_5183,N_4721);
or U5789 (N_5789,N_4962,N_5218);
nor U5790 (N_5790,N_5039,N_4872);
and U5791 (N_5791,N_4870,N_5115);
and U5792 (N_5792,N_4648,N_4847);
and U5793 (N_5793,N_4879,N_5212);
and U5794 (N_5794,N_5249,N_4501);
or U5795 (N_5795,N_5085,N_4784);
and U5796 (N_5796,N_5137,N_4668);
nor U5797 (N_5797,N_4708,N_4836);
or U5798 (N_5798,N_5191,N_4991);
nand U5799 (N_5799,N_5127,N_5139);
and U5800 (N_5800,N_4969,N_5141);
or U5801 (N_5801,N_5156,N_5078);
xnor U5802 (N_5802,N_5080,N_4938);
and U5803 (N_5803,N_4738,N_4924);
nor U5804 (N_5804,N_4936,N_4648);
or U5805 (N_5805,N_4982,N_4951);
nand U5806 (N_5806,N_4700,N_5182);
or U5807 (N_5807,N_4798,N_5131);
and U5808 (N_5808,N_5150,N_4826);
nand U5809 (N_5809,N_5028,N_5197);
nor U5810 (N_5810,N_4770,N_5129);
xor U5811 (N_5811,N_5211,N_5150);
nand U5812 (N_5812,N_5235,N_4908);
nor U5813 (N_5813,N_5063,N_4906);
and U5814 (N_5814,N_4875,N_5224);
nand U5815 (N_5815,N_4945,N_4879);
nand U5816 (N_5816,N_4585,N_4936);
nor U5817 (N_5817,N_4707,N_4802);
and U5818 (N_5818,N_4509,N_4503);
and U5819 (N_5819,N_4983,N_5140);
nor U5820 (N_5820,N_4882,N_5002);
and U5821 (N_5821,N_4794,N_4553);
or U5822 (N_5822,N_4569,N_5025);
nor U5823 (N_5823,N_5056,N_4816);
and U5824 (N_5824,N_5116,N_4557);
and U5825 (N_5825,N_4606,N_5080);
and U5826 (N_5826,N_5183,N_5180);
nor U5827 (N_5827,N_4614,N_5059);
nor U5828 (N_5828,N_4542,N_5076);
or U5829 (N_5829,N_4626,N_4959);
nor U5830 (N_5830,N_4985,N_5190);
or U5831 (N_5831,N_4730,N_4948);
and U5832 (N_5832,N_5022,N_5230);
or U5833 (N_5833,N_5133,N_5124);
nand U5834 (N_5834,N_4739,N_4951);
nand U5835 (N_5835,N_4692,N_4971);
and U5836 (N_5836,N_4799,N_5117);
nand U5837 (N_5837,N_4626,N_4608);
xor U5838 (N_5838,N_4574,N_5062);
or U5839 (N_5839,N_4970,N_4834);
or U5840 (N_5840,N_5040,N_5152);
nand U5841 (N_5841,N_4704,N_4614);
xnor U5842 (N_5842,N_5148,N_4785);
xnor U5843 (N_5843,N_4791,N_4599);
and U5844 (N_5844,N_4962,N_5126);
nand U5845 (N_5845,N_4843,N_4819);
nor U5846 (N_5846,N_5198,N_4620);
or U5847 (N_5847,N_5188,N_4685);
nor U5848 (N_5848,N_4716,N_4575);
xor U5849 (N_5849,N_5129,N_4994);
nand U5850 (N_5850,N_5124,N_4689);
nor U5851 (N_5851,N_5050,N_5064);
xnor U5852 (N_5852,N_4602,N_4850);
nor U5853 (N_5853,N_4798,N_4939);
nand U5854 (N_5854,N_5108,N_5062);
nor U5855 (N_5855,N_5148,N_4971);
or U5856 (N_5856,N_4863,N_4903);
nor U5857 (N_5857,N_4582,N_5048);
and U5858 (N_5858,N_4675,N_5185);
and U5859 (N_5859,N_5080,N_4804);
nand U5860 (N_5860,N_5024,N_4879);
nor U5861 (N_5861,N_4859,N_4950);
and U5862 (N_5862,N_4867,N_4618);
or U5863 (N_5863,N_4883,N_4652);
xnor U5864 (N_5864,N_5134,N_5099);
or U5865 (N_5865,N_4886,N_4514);
nor U5866 (N_5866,N_4854,N_5221);
nor U5867 (N_5867,N_5189,N_4699);
nand U5868 (N_5868,N_4907,N_4575);
nand U5869 (N_5869,N_4662,N_5132);
nor U5870 (N_5870,N_5238,N_4750);
nand U5871 (N_5871,N_4841,N_4951);
nor U5872 (N_5872,N_4808,N_5041);
and U5873 (N_5873,N_4994,N_5204);
nand U5874 (N_5874,N_4506,N_4871);
xnor U5875 (N_5875,N_4916,N_4699);
and U5876 (N_5876,N_4813,N_5025);
and U5877 (N_5877,N_4558,N_5235);
nor U5878 (N_5878,N_4956,N_5241);
nor U5879 (N_5879,N_5109,N_4508);
or U5880 (N_5880,N_5032,N_5139);
and U5881 (N_5881,N_4771,N_4703);
nor U5882 (N_5882,N_4903,N_4530);
nand U5883 (N_5883,N_4974,N_4810);
nor U5884 (N_5884,N_5121,N_5053);
nand U5885 (N_5885,N_4786,N_4834);
nand U5886 (N_5886,N_5159,N_5168);
and U5887 (N_5887,N_5083,N_4857);
or U5888 (N_5888,N_4911,N_4616);
and U5889 (N_5889,N_4576,N_5168);
or U5890 (N_5890,N_4933,N_4902);
or U5891 (N_5891,N_4935,N_5089);
and U5892 (N_5892,N_4639,N_4653);
nand U5893 (N_5893,N_4722,N_4786);
nor U5894 (N_5894,N_5149,N_4537);
or U5895 (N_5895,N_4947,N_5224);
nor U5896 (N_5896,N_5144,N_4908);
or U5897 (N_5897,N_4931,N_4785);
nor U5898 (N_5898,N_4669,N_4522);
and U5899 (N_5899,N_4748,N_4947);
nor U5900 (N_5900,N_5246,N_4882);
nand U5901 (N_5901,N_4544,N_4791);
or U5902 (N_5902,N_4898,N_5026);
or U5903 (N_5903,N_4953,N_4973);
nand U5904 (N_5904,N_5126,N_4748);
nor U5905 (N_5905,N_5249,N_4687);
or U5906 (N_5906,N_5099,N_4584);
and U5907 (N_5907,N_5033,N_4718);
or U5908 (N_5908,N_4555,N_4584);
nor U5909 (N_5909,N_5156,N_5038);
nand U5910 (N_5910,N_5185,N_4609);
and U5911 (N_5911,N_4883,N_4504);
or U5912 (N_5912,N_4788,N_4562);
and U5913 (N_5913,N_5011,N_4886);
or U5914 (N_5914,N_5061,N_5151);
nand U5915 (N_5915,N_4755,N_4768);
or U5916 (N_5916,N_4537,N_4786);
or U5917 (N_5917,N_4660,N_4723);
and U5918 (N_5918,N_5224,N_4771);
xnor U5919 (N_5919,N_4940,N_4878);
and U5920 (N_5920,N_4927,N_4570);
nor U5921 (N_5921,N_4578,N_4510);
xor U5922 (N_5922,N_4694,N_4821);
nor U5923 (N_5923,N_4834,N_5132);
nand U5924 (N_5924,N_4628,N_4834);
nor U5925 (N_5925,N_5094,N_5201);
or U5926 (N_5926,N_4809,N_5240);
or U5927 (N_5927,N_4665,N_4761);
nand U5928 (N_5928,N_4766,N_5155);
nand U5929 (N_5929,N_4524,N_5035);
nand U5930 (N_5930,N_4872,N_4887);
and U5931 (N_5931,N_5249,N_4625);
or U5932 (N_5932,N_4602,N_5113);
or U5933 (N_5933,N_4878,N_4617);
or U5934 (N_5934,N_5128,N_4743);
nand U5935 (N_5935,N_5041,N_4596);
nand U5936 (N_5936,N_5120,N_4626);
and U5937 (N_5937,N_4621,N_4775);
nor U5938 (N_5938,N_4624,N_4800);
nor U5939 (N_5939,N_5022,N_4974);
and U5940 (N_5940,N_5139,N_5009);
nor U5941 (N_5941,N_4629,N_4756);
nor U5942 (N_5942,N_5015,N_5185);
xor U5943 (N_5943,N_4992,N_4571);
nor U5944 (N_5944,N_4821,N_5095);
or U5945 (N_5945,N_5157,N_5065);
nor U5946 (N_5946,N_4706,N_5078);
or U5947 (N_5947,N_5211,N_4768);
nand U5948 (N_5948,N_4658,N_4667);
xor U5949 (N_5949,N_4914,N_4530);
and U5950 (N_5950,N_4936,N_4996);
xnor U5951 (N_5951,N_4885,N_4773);
and U5952 (N_5952,N_4757,N_4572);
xnor U5953 (N_5953,N_4897,N_4970);
nand U5954 (N_5954,N_4889,N_4530);
and U5955 (N_5955,N_4925,N_4582);
or U5956 (N_5956,N_4541,N_4636);
nor U5957 (N_5957,N_5060,N_4747);
and U5958 (N_5958,N_4955,N_4562);
nand U5959 (N_5959,N_4895,N_4649);
or U5960 (N_5960,N_5023,N_4937);
or U5961 (N_5961,N_5091,N_4645);
or U5962 (N_5962,N_5202,N_5211);
and U5963 (N_5963,N_5074,N_4979);
and U5964 (N_5964,N_4698,N_5157);
or U5965 (N_5965,N_4986,N_4708);
or U5966 (N_5966,N_4808,N_4957);
or U5967 (N_5967,N_4829,N_4530);
nor U5968 (N_5968,N_4683,N_4910);
nor U5969 (N_5969,N_4974,N_4584);
nand U5970 (N_5970,N_4787,N_5215);
and U5971 (N_5971,N_4594,N_5234);
nor U5972 (N_5972,N_5247,N_5233);
and U5973 (N_5973,N_5213,N_5099);
and U5974 (N_5974,N_4524,N_5048);
nor U5975 (N_5975,N_4592,N_4531);
nand U5976 (N_5976,N_4523,N_4740);
and U5977 (N_5977,N_5037,N_4502);
nor U5978 (N_5978,N_5011,N_4912);
or U5979 (N_5979,N_4780,N_4601);
and U5980 (N_5980,N_4502,N_4825);
nor U5981 (N_5981,N_4575,N_5011);
xor U5982 (N_5982,N_4569,N_4515);
or U5983 (N_5983,N_4727,N_4824);
and U5984 (N_5984,N_5087,N_4643);
nor U5985 (N_5985,N_5074,N_4738);
xor U5986 (N_5986,N_4794,N_4724);
and U5987 (N_5987,N_4581,N_4964);
nand U5988 (N_5988,N_4624,N_5066);
and U5989 (N_5989,N_5050,N_4796);
nor U5990 (N_5990,N_5133,N_5243);
and U5991 (N_5991,N_4756,N_4577);
and U5992 (N_5992,N_4963,N_4907);
nor U5993 (N_5993,N_5156,N_4988);
and U5994 (N_5994,N_5008,N_4904);
nand U5995 (N_5995,N_5068,N_5178);
nor U5996 (N_5996,N_4991,N_4596);
nor U5997 (N_5997,N_4582,N_5148);
nand U5998 (N_5998,N_4616,N_5169);
or U5999 (N_5999,N_4841,N_4888);
or U6000 (N_6000,N_5289,N_5432);
and U6001 (N_6001,N_5441,N_5789);
and U6002 (N_6002,N_5829,N_5704);
or U6003 (N_6003,N_5642,N_5433);
and U6004 (N_6004,N_5611,N_5765);
or U6005 (N_6005,N_5975,N_5324);
and U6006 (N_6006,N_5830,N_5870);
or U6007 (N_6007,N_5530,N_5757);
or U6008 (N_6008,N_5454,N_5514);
nor U6009 (N_6009,N_5363,N_5339);
nor U6010 (N_6010,N_5440,N_5392);
and U6011 (N_6011,N_5863,N_5610);
xnor U6012 (N_6012,N_5472,N_5752);
or U6013 (N_6013,N_5702,N_5279);
nor U6014 (N_6014,N_5916,N_5336);
nand U6015 (N_6015,N_5853,N_5779);
or U6016 (N_6016,N_5743,N_5512);
and U6017 (N_6017,N_5971,N_5264);
nor U6018 (N_6018,N_5879,N_5891);
and U6019 (N_6019,N_5957,N_5770);
nor U6020 (N_6020,N_5535,N_5557);
or U6021 (N_6021,N_5593,N_5646);
or U6022 (N_6022,N_5873,N_5693);
nor U6023 (N_6023,N_5528,N_5526);
or U6024 (N_6024,N_5670,N_5655);
and U6025 (N_6025,N_5552,N_5768);
nand U6026 (N_6026,N_5882,N_5563);
or U6027 (N_6027,N_5660,N_5887);
and U6028 (N_6028,N_5997,N_5904);
and U6029 (N_6029,N_5272,N_5395);
nor U6030 (N_6030,N_5303,N_5658);
nor U6031 (N_6031,N_5595,N_5509);
or U6032 (N_6032,N_5826,N_5480);
nand U6033 (N_6033,N_5841,N_5974);
or U6034 (N_6034,N_5426,N_5379);
and U6035 (N_6035,N_5293,N_5403);
and U6036 (N_6036,N_5845,N_5842);
or U6037 (N_6037,N_5717,N_5321);
and U6038 (N_6038,N_5678,N_5277);
xor U6039 (N_6039,N_5527,N_5809);
xor U6040 (N_6040,N_5276,N_5946);
or U6041 (N_6041,N_5761,N_5435);
nor U6042 (N_6042,N_5894,N_5596);
nand U6043 (N_6043,N_5972,N_5382);
or U6044 (N_6044,N_5749,N_5477);
nor U6045 (N_6045,N_5418,N_5606);
nand U6046 (N_6046,N_5900,N_5544);
or U6047 (N_6047,N_5501,N_5901);
nor U6048 (N_6048,N_5281,N_5253);
nor U6049 (N_6049,N_5771,N_5333);
and U6050 (N_6050,N_5675,N_5364);
xnor U6051 (N_6051,N_5388,N_5910);
nor U6052 (N_6052,N_5663,N_5268);
or U6053 (N_6053,N_5338,N_5602);
xnor U6054 (N_6054,N_5615,N_5597);
nand U6055 (N_6055,N_5445,N_5513);
nor U6056 (N_6056,N_5381,N_5258);
nand U6057 (N_6057,N_5286,N_5627);
and U6058 (N_6058,N_5375,N_5837);
nor U6059 (N_6059,N_5412,N_5970);
nand U6060 (N_6060,N_5928,N_5929);
nand U6061 (N_6061,N_5759,N_5993);
and U6062 (N_6062,N_5455,N_5899);
xnor U6063 (N_6063,N_5995,N_5843);
and U6064 (N_6064,N_5958,N_5547);
or U6065 (N_6065,N_5346,N_5621);
or U6066 (N_6066,N_5943,N_5963);
nand U6067 (N_6067,N_5591,N_5653);
xnor U6068 (N_6068,N_5878,N_5780);
or U6069 (N_6069,N_5319,N_5612);
and U6070 (N_6070,N_5959,N_5951);
or U6071 (N_6071,N_5518,N_5636);
nand U6072 (N_6072,N_5483,N_5764);
nor U6073 (N_6073,N_5795,N_5648);
xor U6074 (N_6074,N_5603,N_5256);
or U6075 (N_6075,N_5792,N_5534);
nor U6076 (N_6076,N_5654,N_5462);
and U6077 (N_6077,N_5340,N_5589);
or U6078 (N_6078,N_5681,N_5685);
or U6079 (N_6079,N_5417,N_5793);
nand U6080 (N_6080,N_5730,N_5976);
nor U6081 (N_6081,N_5927,N_5955);
nor U6082 (N_6082,N_5539,N_5817);
nand U6083 (N_6083,N_5430,N_5605);
xnor U6084 (N_6084,N_5502,N_5920);
or U6085 (N_6085,N_5291,N_5868);
xnor U6086 (N_6086,N_5748,N_5851);
or U6087 (N_6087,N_5444,N_5821);
nand U6088 (N_6088,N_5991,N_5383);
xor U6089 (N_6089,N_5989,N_5687);
or U6090 (N_6090,N_5747,N_5849);
nor U6091 (N_6091,N_5738,N_5896);
or U6092 (N_6092,N_5923,N_5564);
and U6093 (N_6093,N_5292,N_5366);
or U6094 (N_6094,N_5827,N_5871);
or U6095 (N_6095,N_5525,N_5760);
xor U6096 (N_6096,N_5949,N_5549);
or U6097 (N_6097,N_5798,N_5332);
xnor U6098 (N_6098,N_5372,N_5697);
nor U6099 (N_6099,N_5778,N_5890);
nand U6100 (N_6100,N_5574,N_5608);
nand U6101 (N_6101,N_5977,N_5296);
nor U6102 (N_6102,N_5688,N_5695);
or U6103 (N_6103,N_5712,N_5618);
nand U6104 (N_6104,N_5847,N_5425);
and U6105 (N_6105,N_5408,N_5573);
nand U6106 (N_6106,N_5616,N_5952);
nand U6107 (N_6107,N_5893,N_5945);
and U6108 (N_6108,N_5607,N_5800);
nor U6109 (N_6109,N_5968,N_5885);
or U6110 (N_6110,N_5632,N_5302);
and U6111 (N_6111,N_5938,N_5576);
nand U6112 (N_6112,N_5950,N_5263);
and U6113 (N_6113,N_5369,N_5703);
and U6114 (N_6114,N_5569,N_5742);
nor U6115 (N_6115,N_5781,N_5400);
xor U6116 (N_6116,N_5884,N_5325);
and U6117 (N_6117,N_5541,N_5815);
nor U6118 (N_6118,N_5337,N_5583);
and U6119 (N_6119,N_5719,N_5909);
xor U6120 (N_6120,N_5796,N_5553);
nor U6121 (N_6121,N_5915,N_5650);
nand U6122 (N_6122,N_5314,N_5620);
nand U6123 (N_6123,N_5838,N_5278);
or U6124 (N_6124,N_5311,N_5990);
nand U6125 (N_6125,N_5373,N_5932);
and U6126 (N_6126,N_5404,N_5588);
xnor U6127 (N_6127,N_5814,N_5758);
nor U6128 (N_6128,N_5808,N_5753);
nand U6129 (N_6129,N_5722,N_5714);
or U6130 (N_6130,N_5736,N_5511);
nand U6131 (N_6131,N_5460,N_5832);
nand U6132 (N_6132,N_5331,N_5427);
nor U6133 (N_6133,N_5255,N_5361);
and U6134 (N_6134,N_5546,N_5860);
or U6135 (N_6135,N_5266,N_5516);
or U6136 (N_6136,N_5844,N_5506);
or U6137 (N_6137,N_5741,N_5305);
and U6138 (N_6138,N_5297,N_5327);
nor U6139 (N_6139,N_5385,N_5594);
nand U6140 (N_6140,N_5579,N_5592);
or U6141 (N_6141,N_5755,N_5967);
nor U6142 (N_6142,N_5848,N_5405);
nand U6143 (N_6143,N_5399,N_5707);
and U6144 (N_6144,N_5565,N_5250);
or U6145 (N_6145,N_5275,N_5496);
and U6146 (N_6146,N_5876,N_5918);
and U6147 (N_6147,N_5861,N_5322);
nor U6148 (N_6148,N_5877,N_5811);
nand U6149 (N_6149,N_5582,N_5323);
and U6150 (N_6150,N_5914,N_5874);
and U6151 (N_6151,N_5485,N_5396);
nand U6152 (N_6152,N_5746,N_5422);
nand U6153 (N_6153,N_5862,N_5543);
and U6154 (N_6154,N_5922,N_5280);
xor U6155 (N_6155,N_5442,N_5601);
nor U6156 (N_6156,N_5452,N_5710);
nor U6157 (N_6157,N_5451,N_5407);
nand U6158 (N_6158,N_5898,N_5684);
nand U6159 (N_6159,N_5691,N_5739);
and U6160 (N_6160,N_5356,N_5969);
or U6161 (N_6161,N_5931,N_5803);
nor U6162 (N_6162,N_5482,N_5822);
nand U6163 (N_6163,N_5810,N_5799);
and U6164 (N_6164,N_5661,N_5816);
and U6165 (N_6165,N_5791,N_5619);
nand U6166 (N_6166,N_5668,N_5756);
nand U6167 (N_6167,N_5499,N_5584);
and U6168 (N_6168,N_5979,N_5343);
nand U6169 (N_6169,N_5744,N_5492);
nor U6170 (N_6170,N_5585,N_5686);
and U6171 (N_6171,N_5365,N_5902);
or U6172 (N_6172,N_5575,N_5812);
and U6173 (N_6173,N_5358,N_5913);
nor U6174 (N_6174,N_5329,N_5802);
nand U6175 (N_6175,N_5473,N_5348);
nand U6176 (N_6176,N_5732,N_5907);
and U6177 (N_6177,N_5628,N_5315);
nor U6178 (N_6178,N_5858,N_5353);
nand U6179 (N_6179,N_5897,N_5423);
nand U6180 (N_6180,N_5466,N_5437);
xnor U6181 (N_6181,N_5572,N_5490);
and U6182 (N_6182,N_5623,N_5669);
and U6183 (N_6183,N_5652,N_5370);
or U6184 (N_6184,N_5458,N_5984);
nand U6185 (N_6185,N_5820,N_5921);
nand U6186 (N_6186,N_5298,N_5637);
nand U6187 (N_6187,N_5443,N_5368);
nand U6188 (N_6188,N_5804,N_5320);
nand U6189 (N_6189,N_5677,N_5698);
or U6190 (N_6190,N_5386,N_5998);
nand U6191 (N_6191,N_5420,N_5726);
or U6192 (N_6192,N_5304,N_5510);
and U6193 (N_6193,N_5538,N_5282);
or U6194 (N_6194,N_5474,N_5252);
and U6195 (N_6195,N_5888,N_5359);
xnor U6196 (N_6196,N_5641,N_5580);
nand U6197 (N_6197,N_5469,N_5766);
nor U6198 (N_6198,N_5834,N_5631);
nor U6199 (N_6199,N_5560,N_5926);
nand U6200 (N_6200,N_5797,N_5775);
nand U6201 (N_6201,N_5447,N_5475);
xnor U6202 (N_6202,N_5886,N_5416);
or U6203 (N_6203,N_5629,N_5288);
nand U6204 (N_6204,N_5529,N_5413);
and U6205 (N_6205,N_5507,N_5309);
and U6206 (N_6206,N_5783,N_5270);
or U6207 (N_6207,N_5590,N_5371);
or U6208 (N_6208,N_5831,N_5568);
nor U6209 (N_6209,N_5828,N_5721);
nand U6210 (N_6210,N_5767,N_5694);
nor U6211 (N_6211,N_5545,N_5456);
nand U6212 (N_6212,N_5470,N_5428);
nand U6213 (N_6213,N_5318,N_5344);
or U6214 (N_6214,N_5776,N_5777);
nor U6215 (N_6215,N_5942,N_5273);
and U6216 (N_6216,N_5561,N_5349);
nor U6217 (N_6217,N_5788,N_5479);
or U6218 (N_6218,N_5617,N_5699);
xnor U6219 (N_6219,N_5727,N_5493);
nor U6220 (N_6220,N_5645,N_5450);
and U6221 (N_6221,N_5737,N_5941);
and U6222 (N_6222,N_5377,N_5638);
xnor U6223 (N_6223,N_5762,N_5944);
nor U6224 (N_6224,N_5639,N_5733);
nand U6225 (N_6225,N_5978,N_5672);
or U6226 (N_6226,N_5785,N_5833);
nor U6227 (N_6227,N_5310,N_5287);
nor U6228 (N_6228,N_5328,N_5351);
and U6229 (N_6229,N_5986,N_5414);
or U6230 (N_6230,N_5503,N_5463);
nand U6231 (N_6231,N_5763,N_5720);
nand U6232 (N_6232,N_5647,N_5786);
xor U6233 (N_6233,N_5341,N_5936);
or U6234 (N_6234,N_5892,N_5505);
nor U6235 (N_6235,N_5740,N_5262);
xor U6236 (N_6236,N_5662,N_5419);
or U6237 (N_6237,N_5495,N_5784);
or U6238 (N_6238,N_5352,N_5981);
nand U6239 (N_6239,N_5824,N_5259);
nor U6240 (N_6240,N_5536,N_5261);
xor U6241 (N_6241,N_5912,N_5634);
nor U6242 (N_6242,N_5285,N_5532);
or U6243 (N_6243,N_5599,N_5850);
or U6244 (N_6244,N_5855,N_5269);
nand U6245 (N_6245,N_5614,N_5586);
nor U6246 (N_6246,N_5992,N_5515);
or U6247 (N_6247,N_5271,N_5836);
nand U6248 (N_6248,N_5609,N_5644);
nand U6249 (N_6249,N_5446,N_5643);
or U6250 (N_6250,N_5478,N_5805);
nand U6251 (N_6251,N_5659,N_5999);
nand U6252 (N_6252,N_5774,N_5376);
xnor U6253 (N_6253,N_5713,N_5581);
and U6254 (N_6254,N_5772,N_5571);
xnor U6255 (N_6255,N_5718,N_5360);
nor U6256 (N_6256,N_5924,N_5531);
xnor U6257 (N_6257,N_5961,N_5604);
or U6258 (N_6258,N_5988,N_5983);
nor U6259 (N_6259,N_5705,N_5947);
or U6260 (N_6260,N_5731,N_5554);
or U6261 (N_6261,N_5925,N_5389);
nor U6262 (N_6262,N_5709,N_5267);
xor U6263 (N_6263,N_5251,N_5728);
or U6264 (N_6264,N_5347,N_5700);
nor U6265 (N_6265,N_5857,N_5937);
nor U6266 (N_6266,N_5839,N_5613);
nor U6267 (N_6267,N_5881,N_5725);
nand U6268 (N_6268,N_5489,N_5939);
xor U6269 (N_6269,N_5835,N_5708);
nand U6270 (N_6270,N_5980,N_5819);
and U6271 (N_6271,N_5449,N_5504);
or U6272 (N_6272,N_5872,N_5459);
xor U6273 (N_6273,N_5859,N_5933);
nor U6274 (N_6274,N_5265,N_5556);
nand U6275 (N_6275,N_5402,N_5434);
nor U6276 (N_6276,N_5486,N_5962);
xor U6277 (N_6277,N_5550,N_5484);
or U6278 (N_6278,N_5313,N_5558);
nor U6279 (N_6279,N_5295,N_5378);
nor U6280 (N_6280,N_5517,N_5956);
nor U6281 (N_6281,N_5551,N_5674);
nor U6282 (N_6282,N_5421,N_5683);
or U6283 (N_6283,N_5567,N_5671);
nor U6284 (N_6284,N_5665,N_5716);
and U6285 (N_6285,N_5431,N_5640);
xor U6286 (N_6286,N_5335,N_5257);
nor U6287 (N_6287,N_5308,N_5657);
nand U6288 (N_6288,N_5555,N_5867);
and U6289 (N_6289,N_5317,N_5494);
and U6290 (N_6290,N_5301,N_5578);
nand U6291 (N_6291,N_5488,N_5656);
nor U6292 (N_6292,N_5806,N_5491);
nand U6293 (N_6293,N_5626,N_5439);
nor U6294 (N_6294,N_5520,N_5935);
or U6295 (N_6295,N_5953,N_5880);
nor U6296 (N_6296,N_5409,N_5985);
or U6297 (N_6297,N_5846,N_5715);
nor U6298 (N_6298,N_5476,N_5326);
xnor U6299 (N_6299,N_5919,N_5689);
nor U6300 (N_6300,N_5342,N_5498);
or U6301 (N_6301,N_5312,N_5745);
nand U6302 (N_6302,N_5696,N_5673);
nor U6303 (N_6303,N_5401,N_5410);
or U6304 (N_6304,N_5587,N_5598);
nor U6305 (N_6305,N_5682,N_5316);
or U6306 (N_6306,N_5254,N_5782);
nor U6307 (N_6307,N_5667,N_5711);
or U6308 (N_6308,N_5300,N_5415);
nand U6309 (N_6309,N_5911,N_5274);
xnor U6310 (N_6310,N_5865,N_5866);
nand U6311 (N_6311,N_5468,N_5453);
or U6312 (N_6312,N_5290,N_5464);
xor U6313 (N_6313,N_5905,N_5906);
and U6314 (N_6314,N_5651,N_5630);
or U6315 (N_6315,N_5773,N_5790);
nor U6316 (N_6316,N_5436,N_5367);
xor U6317 (N_6317,N_5299,N_5701);
nor U6318 (N_6318,N_5982,N_5622);
and U6319 (N_6319,N_5750,N_5624);
nand U6320 (N_6320,N_5965,N_5948);
and U6321 (N_6321,N_5334,N_5559);
nand U6322 (N_6322,N_5869,N_5537);
and U6323 (N_6323,N_5649,N_5883);
and U6324 (N_6324,N_5706,N_5954);
and U6325 (N_6325,N_5570,N_5519);
nor U6326 (N_6326,N_5397,N_5438);
and U6327 (N_6327,N_5680,N_5394);
nand U6328 (N_6328,N_5524,N_5330);
or U6329 (N_6329,N_5917,N_5735);
nand U6330 (N_6330,N_5635,N_5964);
nand U6331 (N_6331,N_5889,N_5723);
and U6332 (N_6332,N_5350,N_5856);
and U6333 (N_6333,N_5448,N_5406);
nand U6334 (N_6334,N_5676,N_5294);
nand U6335 (N_6335,N_5903,N_5345);
and U6336 (N_6336,N_5487,N_5875);
and U6337 (N_6337,N_5306,N_5429);
or U6338 (N_6338,N_5908,N_5751);
nand U6339 (N_6339,N_5825,N_5283);
nand U6340 (N_6340,N_5996,N_5497);
or U6341 (N_6341,N_5754,N_5522);
or U6342 (N_6342,N_5966,N_5940);
and U6343 (N_6343,N_5818,N_5533);
nand U6344 (N_6344,N_5508,N_5633);
nor U6345 (N_6345,N_5387,N_5724);
or U6346 (N_6346,N_5354,N_5362);
nor U6347 (N_6347,N_5457,N_5374);
nor U6348 (N_6348,N_5461,N_5577);
and U6349 (N_6349,N_5540,N_5523);
and U6350 (N_6350,N_5729,N_5852);
nor U6351 (N_6351,N_5794,N_5424);
nand U6352 (N_6352,N_5471,N_5769);
nor U6353 (N_6353,N_5854,N_5973);
nand U6354 (N_6354,N_5562,N_5411);
nor U6355 (N_6355,N_5284,N_5355);
nand U6356 (N_6356,N_5692,N_5548);
and U6357 (N_6357,N_5864,N_5566);
nand U6358 (N_6358,N_5393,N_5664);
and U6359 (N_6359,N_5807,N_5934);
or U6360 (N_6360,N_5823,N_5467);
and U6361 (N_6361,N_5895,N_5391);
and U6362 (N_6362,N_5398,N_5679);
nand U6363 (N_6363,N_5465,N_5500);
xnor U6364 (N_6364,N_5625,N_5840);
nor U6365 (N_6365,N_5390,N_5801);
nand U6366 (N_6366,N_5521,N_5600);
and U6367 (N_6367,N_5481,N_5994);
xor U6368 (N_6368,N_5930,N_5260);
nor U6369 (N_6369,N_5384,N_5380);
nand U6370 (N_6370,N_5960,N_5357);
nor U6371 (N_6371,N_5987,N_5542);
or U6372 (N_6372,N_5734,N_5666);
or U6373 (N_6373,N_5787,N_5307);
nor U6374 (N_6374,N_5690,N_5813);
nand U6375 (N_6375,N_5783,N_5258);
nand U6376 (N_6376,N_5367,N_5304);
and U6377 (N_6377,N_5341,N_5899);
nor U6378 (N_6378,N_5996,N_5562);
nand U6379 (N_6379,N_5908,N_5609);
and U6380 (N_6380,N_5527,N_5347);
and U6381 (N_6381,N_5703,N_5904);
nor U6382 (N_6382,N_5483,N_5356);
nor U6383 (N_6383,N_5503,N_5331);
nor U6384 (N_6384,N_5472,N_5546);
nor U6385 (N_6385,N_5614,N_5521);
and U6386 (N_6386,N_5642,N_5750);
or U6387 (N_6387,N_5529,N_5559);
or U6388 (N_6388,N_5464,N_5405);
xnor U6389 (N_6389,N_5876,N_5861);
nor U6390 (N_6390,N_5736,N_5636);
nor U6391 (N_6391,N_5641,N_5314);
xor U6392 (N_6392,N_5733,N_5522);
nand U6393 (N_6393,N_5481,N_5564);
or U6394 (N_6394,N_5325,N_5594);
nand U6395 (N_6395,N_5256,N_5290);
xor U6396 (N_6396,N_5604,N_5477);
nor U6397 (N_6397,N_5732,N_5542);
nor U6398 (N_6398,N_5996,N_5293);
or U6399 (N_6399,N_5722,N_5284);
nor U6400 (N_6400,N_5549,N_5761);
or U6401 (N_6401,N_5783,N_5719);
nand U6402 (N_6402,N_5284,N_5671);
nor U6403 (N_6403,N_5780,N_5690);
xnor U6404 (N_6404,N_5311,N_5552);
nor U6405 (N_6405,N_5625,N_5780);
xor U6406 (N_6406,N_5691,N_5487);
xnor U6407 (N_6407,N_5525,N_5560);
xnor U6408 (N_6408,N_5652,N_5923);
xor U6409 (N_6409,N_5988,N_5859);
or U6410 (N_6410,N_5491,N_5873);
nor U6411 (N_6411,N_5287,N_5370);
nand U6412 (N_6412,N_5301,N_5660);
and U6413 (N_6413,N_5875,N_5833);
nand U6414 (N_6414,N_5945,N_5914);
and U6415 (N_6415,N_5618,N_5760);
nand U6416 (N_6416,N_5267,N_5445);
or U6417 (N_6417,N_5912,N_5485);
xor U6418 (N_6418,N_5340,N_5780);
nor U6419 (N_6419,N_5932,N_5836);
nor U6420 (N_6420,N_5686,N_5544);
nand U6421 (N_6421,N_5497,N_5975);
nand U6422 (N_6422,N_5677,N_5748);
and U6423 (N_6423,N_5953,N_5391);
nand U6424 (N_6424,N_5362,N_5923);
xor U6425 (N_6425,N_5288,N_5926);
or U6426 (N_6426,N_5635,N_5544);
xnor U6427 (N_6427,N_5979,N_5406);
nand U6428 (N_6428,N_5567,N_5709);
nor U6429 (N_6429,N_5953,N_5409);
nand U6430 (N_6430,N_5425,N_5531);
nor U6431 (N_6431,N_5615,N_5735);
nor U6432 (N_6432,N_5765,N_5265);
nor U6433 (N_6433,N_5781,N_5865);
or U6434 (N_6434,N_5874,N_5324);
nand U6435 (N_6435,N_5515,N_5412);
nor U6436 (N_6436,N_5365,N_5762);
nand U6437 (N_6437,N_5736,N_5323);
nor U6438 (N_6438,N_5668,N_5919);
or U6439 (N_6439,N_5300,N_5596);
nor U6440 (N_6440,N_5886,N_5575);
nor U6441 (N_6441,N_5281,N_5987);
nand U6442 (N_6442,N_5549,N_5528);
nand U6443 (N_6443,N_5515,N_5659);
and U6444 (N_6444,N_5333,N_5970);
nor U6445 (N_6445,N_5664,N_5569);
nor U6446 (N_6446,N_5432,N_5287);
and U6447 (N_6447,N_5372,N_5964);
and U6448 (N_6448,N_5421,N_5758);
nor U6449 (N_6449,N_5494,N_5966);
nand U6450 (N_6450,N_5965,N_5597);
nor U6451 (N_6451,N_5268,N_5801);
nor U6452 (N_6452,N_5358,N_5985);
or U6453 (N_6453,N_5958,N_5846);
and U6454 (N_6454,N_5300,N_5716);
or U6455 (N_6455,N_5516,N_5306);
and U6456 (N_6456,N_5487,N_5432);
or U6457 (N_6457,N_5483,N_5668);
or U6458 (N_6458,N_5667,N_5831);
nand U6459 (N_6459,N_5735,N_5322);
nand U6460 (N_6460,N_5930,N_5866);
or U6461 (N_6461,N_5756,N_5959);
and U6462 (N_6462,N_5349,N_5435);
nand U6463 (N_6463,N_5645,N_5268);
xnor U6464 (N_6464,N_5965,N_5935);
or U6465 (N_6465,N_5979,N_5747);
and U6466 (N_6466,N_5323,N_5324);
nor U6467 (N_6467,N_5930,N_5864);
nand U6468 (N_6468,N_5334,N_5767);
or U6469 (N_6469,N_5391,N_5860);
nor U6470 (N_6470,N_5811,N_5328);
xor U6471 (N_6471,N_5555,N_5695);
nand U6472 (N_6472,N_5597,N_5642);
nor U6473 (N_6473,N_5266,N_5508);
nor U6474 (N_6474,N_5657,N_5290);
or U6475 (N_6475,N_5471,N_5565);
nand U6476 (N_6476,N_5525,N_5283);
xnor U6477 (N_6477,N_5631,N_5820);
nand U6478 (N_6478,N_5278,N_5662);
xnor U6479 (N_6479,N_5488,N_5267);
nor U6480 (N_6480,N_5800,N_5693);
nor U6481 (N_6481,N_5646,N_5729);
xor U6482 (N_6482,N_5309,N_5619);
or U6483 (N_6483,N_5693,N_5399);
xor U6484 (N_6484,N_5588,N_5550);
nand U6485 (N_6485,N_5278,N_5510);
nand U6486 (N_6486,N_5659,N_5716);
nand U6487 (N_6487,N_5623,N_5730);
or U6488 (N_6488,N_5910,N_5838);
and U6489 (N_6489,N_5250,N_5276);
or U6490 (N_6490,N_5955,N_5498);
nor U6491 (N_6491,N_5264,N_5550);
nor U6492 (N_6492,N_5376,N_5841);
nor U6493 (N_6493,N_5982,N_5734);
or U6494 (N_6494,N_5510,N_5936);
nor U6495 (N_6495,N_5351,N_5870);
and U6496 (N_6496,N_5540,N_5257);
xnor U6497 (N_6497,N_5250,N_5987);
nor U6498 (N_6498,N_5528,N_5836);
nand U6499 (N_6499,N_5581,N_5776);
nand U6500 (N_6500,N_5753,N_5657);
and U6501 (N_6501,N_5499,N_5514);
xnor U6502 (N_6502,N_5709,N_5635);
xor U6503 (N_6503,N_5253,N_5267);
or U6504 (N_6504,N_5716,N_5411);
or U6505 (N_6505,N_5358,N_5574);
xor U6506 (N_6506,N_5269,N_5856);
nand U6507 (N_6507,N_5440,N_5873);
nand U6508 (N_6508,N_5650,N_5906);
or U6509 (N_6509,N_5556,N_5774);
nand U6510 (N_6510,N_5621,N_5608);
or U6511 (N_6511,N_5861,N_5393);
nand U6512 (N_6512,N_5742,N_5591);
and U6513 (N_6513,N_5419,N_5334);
xor U6514 (N_6514,N_5563,N_5491);
or U6515 (N_6515,N_5734,N_5811);
and U6516 (N_6516,N_5516,N_5337);
and U6517 (N_6517,N_5283,N_5270);
or U6518 (N_6518,N_5595,N_5936);
or U6519 (N_6519,N_5499,N_5400);
nand U6520 (N_6520,N_5526,N_5659);
nor U6521 (N_6521,N_5379,N_5815);
and U6522 (N_6522,N_5730,N_5589);
nand U6523 (N_6523,N_5928,N_5618);
nor U6524 (N_6524,N_5721,N_5510);
nor U6525 (N_6525,N_5311,N_5345);
or U6526 (N_6526,N_5551,N_5455);
nor U6527 (N_6527,N_5744,N_5875);
and U6528 (N_6528,N_5529,N_5783);
or U6529 (N_6529,N_5664,N_5753);
xor U6530 (N_6530,N_5865,N_5698);
and U6531 (N_6531,N_5806,N_5942);
nand U6532 (N_6532,N_5509,N_5758);
or U6533 (N_6533,N_5547,N_5477);
xnor U6534 (N_6534,N_5479,N_5625);
or U6535 (N_6535,N_5927,N_5865);
nor U6536 (N_6536,N_5876,N_5270);
or U6537 (N_6537,N_5796,N_5801);
nor U6538 (N_6538,N_5368,N_5549);
nor U6539 (N_6539,N_5291,N_5779);
xnor U6540 (N_6540,N_5355,N_5751);
nor U6541 (N_6541,N_5341,N_5466);
and U6542 (N_6542,N_5939,N_5494);
and U6543 (N_6543,N_5495,N_5568);
and U6544 (N_6544,N_5851,N_5991);
and U6545 (N_6545,N_5864,N_5402);
nand U6546 (N_6546,N_5634,N_5922);
and U6547 (N_6547,N_5371,N_5470);
and U6548 (N_6548,N_5835,N_5804);
and U6549 (N_6549,N_5612,N_5461);
nand U6550 (N_6550,N_5796,N_5755);
nand U6551 (N_6551,N_5451,N_5313);
nor U6552 (N_6552,N_5656,N_5466);
nand U6553 (N_6553,N_5930,N_5285);
or U6554 (N_6554,N_5268,N_5399);
and U6555 (N_6555,N_5959,N_5526);
or U6556 (N_6556,N_5796,N_5863);
nor U6557 (N_6557,N_5817,N_5585);
or U6558 (N_6558,N_5713,N_5284);
or U6559 (N_6559,N_5534,N_5355);
nand U6560 (N_6560,N_5415,N_5983);
and U6561 (N_6561,N_5850,N_5999);
xor U6562 (N_6562,N_5306,N_5468);
or U6563 (N_6563,N_5922,N_5967);
nand U6564 (N_6564,N_5787,N_5280);
nand U6565 (N_6565,N_5926,N_5913);
nor U6566 (N_6566,N_5564,N_5354);
and U6567 (N_6567,N_5462,N_5759);
nor U6568 (N_6568,N_5853,N_5436);
and U6569 (N_6569,N_5276,N_5299);
or U6570 (N_6570,N_5322,N_5775);
nor U6571 (N_6571,N_5432,N_5614);
nand U6572 (N_6572,N_5937,N_5538);
and U6573 (N_6573,N_5806,N_5465);
nor U6574 (N_6574,N_5309,N_5744);
nor U6575 (N_6575,N_5402,N_5651);
nand U6576 (N_6576,N_5703,N_5889);
nand U6577 (N_6577,N_5771,N_5614);
or U6578 (N_6578,N_5402,N_5457);
and U6579 (N_6579,N_5655,N_5718);
and U6580 (N_6580,N_5324,N_5255);
nor U6581 (N_6581,N_5409,N_5750);
or U6582 (N_6582,N_5350,N_5531);
nand U6583 (N_6583,N_5436,N_5262);
nand U6584 (N_6584,N_5708,N_5626);
nor U6585 (N_6585,N_5702,N_5461);
nor U6586 (N_6586,N_5804,N_5936);
nand U6587 (N_6587,N_5418,N_5645);
xor U6588 (N_6588,N_5858,N_5653);
or U6589 (N_6589,N_5463,N_5269);
nand U6590 (N_6590,N_5724,N_5297);
or U6591 (N_6591,N_5560,N_5409);
and U6592 (N_6592,N_5802,N_5904);
and U6593 (N_6593,N_5995,N_5931);
and U6594 (N_6594,N_5913,N_5566);
nor U6595 (N_6595,N_5340,N_5866);
nor U6596 (N_6596,N_5890,N_5557);
and U6597 (N_6597,N_5320,N_5704);
nand U6598 (N_6598,N_5938,N_5608);
and U6599 (N_6599,N_5575,N_5471);
nor U6600 (N_6600,N_5629,N_5363);
xnor U6601 (N_6601,N_5564,N_5927);
xor U6602 (N_6602,N_5352,N_5731);
or U6603 (N_6603,N_5628,N_5694);
and U6604 (N_6604,N_5362,N_5395);
or U6605 (N_6605,N_5907,N_5608);
xnor U6606 (N_6606,N_5816,N_5440);
nand U6607 (N_6607,N_5766,N_5876);
and U6608 (N_6608,N_5930,N_5845);
nand U6609 (N_6609,N_5354,N_5801);
nor U6610 (N_6610,N_5717,N_5391);
nand U6611 (N_6611,N_5976,N_5660);
and U6612 (N_6612,N_5555,N_5717);
nand U6613 (N_6613,N_5520,N_5667);
or U6614 (N_6614,N_5755,N_5656);
or U6615 (N_6615,N_5873,N_5609);
nor U6616 (N_6616,N_5738,N_5539);
nor U6617 (N_6617,N_5538,N_5728);
nor U6618 (N_6618,N_5521,N_5658);
nand U6619 (N_6619,N_5879,N_5632);
xnor U6620 (N_6620,N_5512,N_5919);
nor U6621 (N_6621,N_5853,N_5415);
nor U6622 (N_6622,N_5794,N_5526);
and U6623 (N_6623,N_5581,N_5292);
nor U6624 (N_6624,N_5255,N_5422);
xor U6625 (N_6625,N_5410,N_5435);
nand U6626 (N_6626,N_5799,N_5406);
nand U6627 (N_6627,N_5793,N_5478);
or U6628 (N_6628,N_5866,N_5416);
nand U6629 (N_6629,N_5985,N_5590);
and U6630 (N_6630,N_5916,N_5629);
and U6631 (N_6631,N_5665,N_5872);
and U6632 (N_6632,N_5592,N_5702);
xnor U6633 (N_6633,N_5827,N_5969);
and U6634 (N_6634,N_5338,N_5917);
or U6635 (N_6635,N_5745,N_5870);
nor U6636 (N_6636,N_5390,N_5335);
and U6637 (N_6637,N_5944,N_5682);
and U6638 (N_6638,N_5365,N_5452);
or U6639 (N_6639,N_5641,N_5786);
xnor U6640 (N_6640,N_5796,N_5772);
nor U6641 (N_6641,N_5689,N_5614);
nand U6642 (N_6642,N_5610,N_5846);
nand U6643 (N_6643,N_5558,N_5947);
or U6644 (N_6644,N_5910,N_5853);
nor U6645 (N_6645,N_5785,N_5475);
nand U6646 (N_6646,N_5626,N_5555);
nor U6647 (N_6647,N_5624,N_5915);
nor U6648 (N_6648,N_5407,N_5748);
nand U6649 (N_6649,N_5302,N_5534);
nand U6650 (N_6650,N_5736,N_5953);
nor U6651 (N_6651,N_5820,N_5675);
and U6652 (N_6652,N_5564,N_5501);
or U6653 (N_6653,N_5852,N_5722);
or U6654 (N_6654,N_5313,N_5699);
or U6655 (N_6655,N_5758,N_5598);
or U6656 (N_6656,N_5480,N_5312);
xnor U6657 (N_6657,N_5429,N_5847);
or U6658 (N_6658,N_5782,N_5356);
and U6659 (N_6659,N_5781,N_5822);
nand U6660 (N_6660,N_5321,N_5520);
nand U6661 (N_6661,N_5853,N_5549);
or U6662 (N_6662,N_5883,N_5708);
nand U6663 (N_6663,N_5746,N_5976);
and U6664 (N_6664,N_5780,N_5594);
nor U6665 (N_6665,N_5350,N_5788);
or U6666 (N_6666,N_5859,N_5251);
xnor U6667 (N_6667,N_5768,N_5563);
or U6668 (N_6668,N_5740,N_5571);
nor U6669 (N_6669,N_5629,N_5822);
xor U6670 (N_6670,N_5970,N_5613);
nor U6671 (N_6671,N_5392,N_5821);
and U6672 (N_6672,N_5714,N_5362);
nand U6673 (N_6673,N_5399,N_5569);
nor U6674 (N_6674,N_5725,N_5611);
and U6675 (N_6675,N_5826,N_5309);
nand U6676 (N_6676,N_5782,N_5886);
nand U6677 (N_6677,N_5400,N_5442);
or U6678 (N_6678,N_5810,N_5515);
nor U6679 (N_6679,N_5856,N_5311);
nand U6680 (N_6680,N_5779,N_5693);
and U6681 (N_6681,N_5614,N_5541);
nand U6682 (N_6682,N_5564,N_5779);
or U6683 (N_6683,N_5321,N_5727);
or U6684 (N_6684,N_5255,N_5281);
nor U6685 (N_6685,N_5846,N_5964);
nand U6686 (N_6686,N_5481,N_5417);
nand U6687 (N_6687,N_5727,N_5775);
xnor U6688 (N_6688,N_5881,N_5624);
or U6689 (N_6689,N_5458,N_5490);
or U6690 (N_6690,N_5315,N_5970);
nand U6691 (N_6691,N_5854,N_5481);
and U6692 (N_6692,N_5440,N_5496);
nor U6693 (N_6693,N_5354,N_5740);
and U6694 (N_6694,N_5446,N_5285);
nor U6695 (N_6695,N_5721,N_5475);
nand U6696 (N_6696,N_5411,N_5987);
and U6697 (N_6697,N_5932,N_5413);
nand U6698 (N_6698,N_5788,N_5495);
nor U6699 (N_6699,N_5735,N_5686);
or U6700 (N_6700,N_5962,N_5974);
or U6701 (N_6701,N_5556,N_5725);
and U6702 (N_6702,N_5344,N_5646);
xnor U6703 (N_6703,N_5700,N_5916);
nand U6704 (N_6704,N_5558,N_5353);
nor U6705 (N_6705,N_5900,N_5926);
or U6706 (N_6706,N_5339,N_5872);
nand U6707 (N_6707,N_5930,N_5629);
or U6708 (N_6708,N_5253,N_5771);
xor U6709 (N_6709,N_5660,N_5874);
and U6710 (N_6710,N_5627,N_5320);
and U6711 (N_6711,N_5622,N_5957);
nor U6712 (N_6712,N_5586,N_5588);
nand U6713 (N_6713,N_5821,N_5555);
and U6714 (N_6714,N_5346,N_5780);
xor U6715 (N_6715,N_5559,N_5707);
nor U6716 (N_6716,N_5895,N_5620);
and U6717 (N_6717,N_5302,N_5682);
nor U6718 (N_6718,N_5630,N_5613);
xnor U6719 (N_6719,N_5263,N_5850);
nand U6720 (N_6720,N_5791,N_5269);
nand U6721 (N_6721,N_5478,N_5828);
xor U6722 (N_6722,N_5565,N_5966);
or U6723 (N_6723,N_5528,N_5432);
nor U6724 (N_6724,N_5733,N_5549);
xnor U6725 (N_6725,N_5420,N_5865);
nand U6726 (N_6726,N_5924,N_5554);
or U6727 (N_6727,N_5268,N_5313);
or U6728 (N_6728,N_5702,N_5571);
or U6729 (N_6729,N_5965,N_5599);
or U6730 (N_6730,N_5422,N_5426);
or U6731 (N_6731,N_5310,N_5644);
or U6732 (N_6732,N_5502,N_5295);
nand U6733 (N_6733,N_5574,N_5840);
and U6734 (N_6734,N_5835,N_5318);
nand U6735 (N_6735,N_5453,N_5338);
or U6736 (N_6736,N_5781,N_5871);
or U6737 (N_6737,N_5705,N_5796);
and U6738 (N_6738,N_5673,N_5908);
and U6739 (N_6739,N_5413,N_5276);
and U6740 (N_6740,N_5911,N_5881);
or U6741 (N_6741,N_5977,N_5780);
or U6742 (N_6742,N_5546,N_5972);
nand U6743 (N_6743,N_5754,N_5616);
nor U6744 (N_6744,N_5994,N_5897);
nor U6745 (N_6745,N_5549,N_5658);
or U6746 (N_6746,N_5343,N_5621);
nand U6747 (N_6747,N_5304,N_5336);
and U6748 (N_6748,N_5788,N_5345);
or U6749 (N_6749,N_5866,N_5983);
nor U6750 (N_6750,N_6232,N_6076);
nand U6751 (N_6751,N_6263,N_6516);
or U6752 (N_6752,N_6186,N_6414);
nand U6753 (N_6753,N_6624,N_6269);
nor U6754 (N_6754,N_6506,N_6339);
nor U6755 (N_6755,N_6373,N_6551);
and U6756 (N_6756,N_6268,N_6111);
nor U6757 (N_6757,N_6068,N_6161);
nand U6758 (N_6758,N_6655,N_6073);
or U6759 (N_6759,N_6172,N_6081);
nor U6760 (N_6760,N_6157,N_6703);
nand U6761 (N_6761,N_6147,N_6710);
and U6762 (N_6762,N_6140,N_6517);
nand U6763 (N_6763,N_6208,N_6451);
or U6764 (N_6764,N_6440,N_6283);
nor U6765 (N_6765,N_6088,N_6329);
xor U6766 (N_6766,N_6652,N_6118);
nor U6767 (N_6767,N_6654,N_6555);
and U6768 (N_6768,N_6303,N_6742);
nand U6769 (N_6769,N_6052,N_6615);
or U6770 (N_6770,N_6291,N_6385);
or U6771 (N_6771,N_6025,N_6488);
nand U6772 (N_6772,N_6336,N_6252);
nor U6773 (N_6773,N_6535,N_6564);
nor U6774 (N_6774,N_6350,N_6097);
nor U6775 (N_6775,N_6162,N_6332);
nor U6776 (N_6776,N_6279,N_6374);
and U6777 (N_6777,N_6197,N_6204);
or U6778 (N_6778,N_6302,N_6433);
or U6779 (N_6779,N_6563,N_6594);
nand U6780 (N_6780,N_6155,N_6523);
nand U6781 (N_6781,N_6454,N_6595);
and U6782 (N_6782,N_6665,N_6477);
and U6783 (N_6783,N_6249,N_6711);
or U6784 (N_6784,N_6632,N_6643);
or U6785 (N_6785,N_6103,N_6337);
or U6786 (N_6786,N_6014,N_6008);
nand U6787 (N_6787,N_6188,N_6436);
and U6788 (N_6788,N_6457,N_6091);
nor U6789 (N_6789,N_6254,N_6178);
or U6790 (N_6790,N_6098,N_6031);
or U6791 (N_6791,N_6005,N_6158);
and U6792 (N_6792,N_6420,N_6275);
and U6793 (N_6793,N_6018,N_6587);
xor U6794 (N_6794,N_6276,N_6050);
or U6795 (N_6795,N_6554,N_6738);
or U6796 (N_6796,N_6273,N_6530);
and U6797 (N_6797,N_6514,N_6138);
and U6798 (N_6798,N_6307,N_6467);
or U6799 (N_6799,N_6601,N_6362);
or U6800 (N_6800,N_6460,N_6203);
nor U6801 (N_6801,N_6537,N_6439);
and U6802 (N_6802,N_6109,N_6065);
and U6803 (N_6803,N_6745,N_6657);
nor U6804 (N_6804,N_6735,N_6424);
nor U6805 (N_6805,N_6707,N_6349);
or U6806 (N_6806,N_6412,N_6744);
and U6807 (N_6807,N_6270,N_6720);
and U6808 (N_6808,N_6661,N_6653);
nand U6809 (N_6809,N_6588,N_6258);
and U6810 (N_6810,N_6628,N_6251);
nand U6811 (N_6811,N_6437,N_6305);
and U6812 (N_6812,N_6331,N_6583);
nand U6813 (N_6813,N_6061,N_6714);
and U6814 (N_6814,N_6579,N_6070);
and U6815 (N_6815,N_6681,N_6569);
nand U6816 (N_6816,N_6019,N_6104);
and U6817 (N_6817,N_6450,N_6567);
and U6818 (N_6818,N_6280,N_6132);
nand U6819 (N_6819,N_6730,N_6447);
nand U6820 (N_6820,N_6430,N_6009);
xor U6821 (N_6821,N_6641,N_6465);
nand U6822 (N_6822,N_6190,N_6668);
nand U6823 (N_6823,N_6473,N_6692);
nand U6824 (N_6824,N_6020,N_6046);
nor U6825 (N_6825,N_6380,N_6156);
nor U6826 (N_6826,N_6746,N_6266);
or U6827 (N_6827,N_6059,N_6577);
xor U6828 (N_6828,N_6574,N_6542);
xor U6829 (N_6829,N_6146,N_6194);
nor U6830 (N_6830,N_6029,N_6401);
and U6831 (N_6831,N_6464,N_6407);
nor U6832 (N_6832,N_6358,N_6598);
nand U6833 (N_6833,N_6347,N_6013);
and U6834 (N_6834,N_6066,N_6067);
nor U6835 (N_6835,N_6313,N_6035);
nand U6836 (N_6836,N_6130,N_6548);
and U6837 (N_6837,N_6037,N_6578);
xor U6838 (N_6838,N_6558,N_6051);
nand U6839 (N_6839,N_6443,N_6151);
or U6840 (N_6840,N_6021,N_6573);
or U6841 (N_6841,N_6345,N_6584);
nand U6842 (N_6842,N_6235,N_6087);
nor U6843 (N_6843,N_6028,N_6344);
nand U6844 (N_6844,N_6671,N_6141);
and U6845 (N_6845,N_6731,N_6304);
nor U6846 (N_6846,N_6078,N_6187);
or U6847 (N_6847,N_6055,N_6480);
and U6848 (N_6848,N_6015,N_6502);
nand U6849 (N_6849,N_6122,N_6474);
nor U6850 (N_6850,N_6136,N_6384);
nand U6851 (N_6851,N_6640,N_6402);
or U6852 (N_6852,N_6072,N_6196);
nand U6853 (N_6853,N_6165,N_6348);
and U6854 (N_6854,N_6164,N_6160);
or U6855 (N_6855,N_6701,N_6369);
or U6856 (N_6856,N_6333,N_6697);
nand U6857 (N_6857,N_6298,N_6647);
nor U6858 (N_6858,N_6000,N_6328);
nand U6859 (N_6859,N_6603,N_6127);
nor U6860 (N_6860,N_6521,N_6475);
and U6861 (N_6861,N_6518,N_6452);
xnor U6862 (N_6862,N_6716,N_6192);
xor U6863 (N_6863,N_6054,N_6565);
and U6864 (N_6864,N_6079,N_6642);
nor U6865 (N_6865,N_6680,N_6561);
nand U6866 (N_6866,N_6592,N_6179);
and U6867 (N_6867,N_6117,N_6288);
nand U6868 (N_6868,N_6515,N_6580);
and U6869 (N_6869,N_6543,N_6379);
nor U6870 (N_6870,N_6609,N_6060);
xnor U6871 (N_6871,N_6256,N_6429);
nor U6872 (N_6872,N_6743,N_6610);
or U6873 (N_6873,N_6685,N_6495);
xnor U6874 (N_6874,N_6717,N_6063);
and U6875 (N_6875,N_6570,N_6618);
or U6876 (N_6876,N_6623,N_6531);
nand U6877 (N_6877,N_6572,N_6282);
nor U6878 (N_6878,N_6651,N_6293);
nor U6879 (N_6879,N_6704,N_6544);
and U6880 (N_6880,N_6511,N_6696);
xnor U6881 (N_6881,N_6434,N_6575);
xnor U6882 (N_6882,N_6231,N_6619);
nand U6883 (N_6883,N_6327,N_6239);
xnor U6884 (N_6884,N_6033,N_6694);
and U6885 (N_6885,N_6485,N_6597);
or U6886 (N_6886,N_6686,N_6023);
and U6887 (N_6887,N_6360,N_6687);
or U6888 (N_6888,N_6128,N_6416);
nand U6889 (N_6889,N_6223,N_6453);
nand U6890 (N_6890,N_6290,N_6620);
nor U6891 (N_6891,N_6142,N_6176);
nand U6892 (N_6892,N_6581,N_6183);
and U6893 (N_6893,N_6189,N_6016);
xor U6894 (N_6894,N_6718,N_6113);
nand U6895 (N_6895,N_6472,N_6728);
or U6896 (N_6896,N_6041,N_6427);
nor U6897 (N_6897,N_6227,N_6108);
and U6898 (N_6898,N_6706,N_6483);
and U6899 (N_6899,N_6378,N_6342);
nor U6900 (N_6900,N_6324,N_6422);
or U6901 (N_6901,N_6116,N_6636);
and U6902 (N_6902,N_6367,N_6505);
nor U6903 (N_6903,N_6124,N_6670);
and U6904 (N_6904,N_6074,N_6616);
nand U6905 (N_6905,N_6556,N_6519);
or U6906 (N_6906,N_6482,N_6012);
nor U6907 (N_6907,N_6094,N_6368);
nor U6908 (N_6908,N_6526,N_6528);
and U6909 (N_6909,N_6214,N_6481);
xor U6910 (N_6910,N_6295,N_6330);
nor U6911 (N_6911,N_6418,N_6391);
and U6912 (N_6912,N_6411,N_6672);
xnor U6913 (N_6913,N_6207,N_6226);
nor U6914 (N_6914,N_6287,N_6137);
and U6915 (N_6915,N_6712,N_6247);
nor U6916 (N_6916,N_6622,N_6101);
and U6917 (N_6917,N_6026,N_6599);
nor U6918 (N_6918,N_6497,N_6634);
nand U6919 (N_6919,N_6646,N_6510);
nor U6920 (N_6920,N_6719,N_6110);
nand U6921 (N_6921,N_6677,N_6082);
and U6922 (N_6922,N_6377,N_6590);
or U6923 (N_6923,N_6382,N_6487);
and U6924 (N_6924,N_6191,N_6708);
nand U6925 (N_6925,N_6351,N_6312);
and U6926 (N_6926,N_6359,N_6679);
and U6927 (N_6927,N_6170,N_6501);
nand U6928 (N_6928,N_6229,N_6478);
and U6929 (N_6929,N_6106,N_6343);
nor U6930 (N_6930,N_6205,N_6727);
or U6931 (N_6931,N_6648,N_6354);
and U6932 (N_6932,N_6455,N_6027);
nor U6933 (N_6933,N_6498,N_6315);
nand U6934 (N_6934,N_6722,N_6356);
or U6935 (N_6935,N_6408,N_6419);
and U6936 (N_6936,N_6093,N_6089);
nor U6937 (N_6937,N_6319,N_6096);
and U6938 (N_6938,N_6185,N_6370);
nand U6939 (N_6939,N_6639,N_6394);
and U6940 (N_6940,N_6484,N_6237);
nand U6941 (N_6941,N_6123,N_6198);
and U6942 (N_6942,N_6702,N_6209);
or U6943 (N_6943,N_6689,N_6213);
and U6944 (N_6944,N_6586,N_6119);
or U6945 (N_6945,N_6663,N_6086);
or U6946 (N_6946,N_6285,N_6371);
or U6947 (N_6947,N_6316,N_6202);
or U6948 (N_6948,N_6605,N_6084);
nor U6949 (N_6949,N_6099,N_6272);
nand U6950 (N_6950,N_6614,N_6168);
and U6951 (N_6951,N_6080,N_6524);
or U6952 (N_6952,N_6318,N_6236);
and U6953 (N_6953,N_6201,N_6666);
nor U6954 (N_6954,N_6069,N_6660);
nor U6955 (N_6955,N_6238,N_6612);
and U6956 (N_6956,N_6107,N_6077);
and U6957 (N_6957,N_6267,N_6010);
or U6958 (N_6958,N_6507,N_6695);
and U6959 (N_6959,N_6734,N_6644);
nor U6960 (N_6960,N_6011,N_6334);
nand U6961 (N_6961,N_6150,N_6326);
or U6962 (N_6962,N_6662,N_6406);
nor U6963 (N_6963,N_6626,N_6725);
nor U6964 (N_6964,N_6534,N_6220);
or U6965 (N_6965,N_6700,N_6489);
nand U6966 (N_6966,N_6723,N_6085);
nor U6967 (N_6967,N_6071,N_6134);
or U6968 (N_6968,N_6233,N_6423);
or U6969 (N_6969,N_6396,N_6314);
and U6970 (N_6970,N_6007,N_6729);
and U6971 (N_6971,N_6259,N_6678);
nand U6972 (N_6972,N_6540,N_6715);
nor U6973 (N_6973,N_6043,N_6320);
nand U6974 (N_6974,N_6365,N_6552);
or U6975 (N_6975,N_6001,N_6322);
nand U6976 (N_6976,N_6635,N_6277);
nor U6977 (N_6977,N_6039,N_6265);
nand U6978 (N_6978,N_6264,N_6173);
and U6979 (N_6979,N_6449,N_6664);
nand U6980 (N_6980,N_6533,N_6306);
or U6981 (N_6981,N_6159,N_6244);
xor U6982 (N_6982,N_6056,N_6499);
nor U6983 (N_6983,N_6390,N_6600);
or U6984 (N_6984,N_6032,N_6549);
or U6985 (N_6985,N_6121,N_6181);
xnor U6986 (N_6986,N_6346,N_6248);
nor U6987 (N_6987,N_6299,N_6112);
xnor U6988 (N_6988,N_6102,N_6174);
nand U6989 (N_6989,N_6645,N_6149);
xor U6990 (N_6990,N_6053,N_6486);
and U6991 (N_6991,N_6426,N_6625);
nor U6992 (N_6992,N_6047,N_6144);
xor U6993 (N_6993,N_6748,N_6741);
or U6994 (N_6994,N_6493,N_6260);
and U6995 (N_6995,N_6338,N_6215);
nor U6996 (N_6996,N_6309,N_6462);
nand U6997 (N_6997,N_6576,N_6323);
nand U6998 (N_6998,N_6361,N_6566);
nand U6999 (N_6999,N_6463,N_6199);
and U7000 (N_7000,N_6064,N_6513);
or U7001 (N_7001,N_6177,N_6432);
nor U7002 (N_7002,N_6532,N_6428);
and U7003 (N_7003,N_6659,N_6057);
nand U7004 (N_7004,N_6040,N_6739);
and U7005 (N_7005,N_6292,N_6490);
xor U7006 (N_7006,N_6496,N_6568);
or U7007 (N_7007,N_6261,N_6355);
nand U7008 (N_7008,N_6656,N_6049);
nand U7009 (N_7009,N_6509,N_6296);
nor U7010 (N_7010,N_6195,N_6404);
nor U7011 (N_7011,N_6669,N_6243);
nand U7012 (N_7012,N_6317,N_6441);
and U7013 (N_7013,N_6629,N_6250);
nand U7014 (N_7014,N_6550,N_6733);
nand U7015 (N_7015,N_6658,N_6002);
nand U7016 (N_7016,N_6503,N_6271);
nand U7017 (N_7017,N_6732,N_6274);
and U7018 (N_7018,N_6456,N_6633);
xor U7019 (N_7019,N_6425,N_6504);
and U7020 (N_7020,N_6684,N_6352);
xnor U7021 (N_7021,N_6397,N_6675);
nand U7022 (N_7022,N_6289,N_6152);
nand U7023 (N_7023,N_6163,N_6593);
nor U7024 (N_7024,N_6448,N_6638);
nand U7025 (N_7025,N_6224,N_6421);
and U7026 (N_7026,N_6726,N_6310);
or U7027 (N_7027,N_6721,N_6120);
and U7028 (N_7028,N_6126,N_6649);
or U7029 (N_7029,N_6253,N_6212);
and U7030 (N_7030,N_6562,N_6627);
nand U7031 (N_7031,N_6479,N_6539);
nand U7032 (N_7032,N_6491,N_6699);
and U7033 (N_7033,N_6105,N_6153);
or U7034 (N_7034,N_6022,N_6713);
nand U7035 (N_7035,N_6747,N_6637);
nor U7036 (N_7036,N_6353,N_6459);
nand U7037 (N_7037,N_6621,N_6557);
or U7038 (N_7038,N_6284,N_6737);
or U7039 (N_7039,N_6222,N_6048);
nor U7040 (N_7040,N_6241,N_6547);
nand U7041 (N_7041,N_6321,N_6300);
or U7042 (N_7042,N_6038,N_6682);
nand U7043 (N_7043,N_6042,N_6230);
or U7044 (N_7044,N_6006,N_6184);
nor U7045 (N_7045,N_6045,N_6129);
nor U7046 (N_7046,N_6145,N_6278);
xor U7047 (N_7047,N_6257,N_6115);
or U7048 (N_7048,N_6468,N_6591);
and U7049 (N_7049,N_6133,N_6400);
nand U7050 (N_7050,N_6438,N_6431);
and U7051 (N_7051,N_6596,N_6034);
and U7052 (N_7052,N_6262,N_6180);
or U7053 (N_7053,N_6674,N_6245);
nand U7054 (N_7054,N_6175,N_6210);
nor U7055 (N_7055,N_6617,N_6469);
nand U7056 (N_7056,N_6325,N_6169);
or U7057 (N_7057,N_6494,N_6240);
or U7058 (N_7058,N_6286,N_6386);
nor U7059 (N_7059,N_6709,N_6090);
nand U7060 (N_7060,N_6083,N_6376);
nor U7061 (N_7061,N_6415,N_6221);
xor U7062 (N_7062,N_6387,N_6017);
xor U7063 (N_7063,N_6604,N_6749);
xor U7064 (N_7064,N_6389,N_6559);
nor U7065 (N_7065,N_6435,N_6470);
nor U7066 (N_7066,N_6357,N_6442);
nand U7067 (N_7067,N_6044,N_6395);
nor U7068 (N_7068,N_6611,N_6512);
or U7069 (N_7069,N_6375,N_6536);
nand U7070 (N_7070,N_6405,N_6381);
nand U7071 (N_7071,N_6058,N_6246);
and U7072 (N_7072,N_6698,N_6538);
nor U7073 (N_7073,N_6606,N_6004);
or U7074 (N_7074,N_6667,N_6541);
or U7075 (N_7075,N_6154,N_6585);
and U7076 (N_7076,N_6148,N_6030);
nor U7077 (N_7077,N_6399,N_6690);
nor U7078 (N_7078,N_6413,N_6392);
and U7079 (N_7079,N_6693,N_6508);
and U7080 (N_7080,N_6143,N_6705);
nand U7081 (N_7081,N_6242,N_6545);
and U7082 (N_7082,N_6341,N_6092);
or U7083 (N_7083,N_6630,N_6131);
or U7084 (N_7084,N_6571,N_6075);
or U7085 (N_7085,N_6492,N_6217);
nand U7086 (N_7086,N_6553,N_6476);
xor U7087 (N_7087,N_6281,N_6114);
nor U7088 (N_7088,N_6546,N_6100);
nand U7089 (N_7089,N_6417,N_6294);
and U7090 (N_7090,N_6255,N_6383);
nor U7091 (N_7091,N_6676,N_6461);
nor U7092 (N_7092,N_6398,N_6135);
nor U7093 (N_7093,N_6216,N_6409);
nand U7094 (N_7094,N_6631,N_6311);
nor U7095 (N_7095,N_6650,N_6206);
xor U7096 (N_7096,N_6003,N_6166);
nand U7097 (N_7097,N_6062,N_6182);
nand U7098 (N_7098,N_6167,N_6218);
and U7099 (N_7099,N_6525,N_6366);
nand U7100 (N_7100,N_6529,N_6024);
or U7101 (N_7101,N_6527,N_6471);
or U7102 (N_7102,N_6613,N_6740);
and U7103 (N_7103,N_6458,N_6393);
or U7104 (N_7104,N_6335,N_6301);
or U7105 (N_7105,N_6364,N_6520);
nand U7106 (N_7106,N_6410,N_6193);
nor U7107 (N_7107,N_6688,N_6522);
nor U7108 (N_7108,N_6446,N_6219);
nor U7109 (N_7109,N_6297,N_6691);
nor U7110 (N_7110,N_6683,N_6234);
xor U7111 (N_7111,N_6372,N_6171);
nand U7112 (N_7112,N_6582,N_6388);
or U7113 (N_7113,N_6095,N_6445);
or U7114 (N_7114,N_6608,N_6500);
and U7115 (N_7115,N_6403,N_6602);
nor U7116 (N_7116,N_6607,N_6211);
nand U7117 (N_7117,N_6225,N_6139);
nand U7118 (N_7118,N_6724,N_6673);
or U7119 (N_7119,N_6466,N_6200);
xnor U7120 (N_7120,N_6363,N_6228);
nand U7121 (N_7121,N_6308,N_6444);
xnor U7122 (N_7122,N_6036,N_6560);
nor U7123 (N_7123,N_6589,N_6125);
nor U7124 (N_7124,N_6736,N_6340);
nand U7125 (N_7125,N_6017,N_6236);
nand U7126 (N_7126,N_6167,N_6567);
or U7127 (N_7127,N_6146,N_6417);
nor U7128 (N_7128,N_6341,N_6199);
xor U7129 (N_7129,N_6571,N_6744);
nand U7130 (N_7130,N_6139,N_6209);
or U7131 (N_7131,N_6349,N_6382);
or U7132 (N_7132,N_6378,N_6360);
nor U7133 (N_7133,N_6366,N_6192);
or U7134 (N_7134,N_6346,N_6633);
xor U7135 (N_7135,N_6085,N_6617);
and U7136 (N_7136,N_6481,N_6388);
nor U7137 (N_7137,N_6398,N_6120);
and U7138 (N_7138,N_6454,N_6652);
nand U7139 (N_7139,N_6010,N_6330);
nand U7140 (N_7140,N_6319,N_6511);
or U7141 (N_7141,N_6244,N_6041);
or U7142 (N_7142,N_6315,N_6344);
or U7143 (N_7143,N_6258,N_6016);
nor U7144 (N_7144,N_6285,N_6167);
and U7145 (N_7145,N_6654,N_6392);
nand U7146 (N_7146,N_6236,N_6544);
nand U7147 (N_7147,N_6661,N_6549);
nor U7148 (N_7148,N_6113,N_6493);
and U7149 (N_7149,N_6735,N_6562);
xor U7150 (N_7150,N_6534,N_6703);
or U7151 (N_7151,N_6168,N_6286);
nand U7152 (N_7152,N_6432,N_6458);
nand U7153 (N_7153,N_6145,N_6153);
nor U7154 (N_7154,N_6178,N_6250);
nand U7155 (N_7155,N_6722,N_6650);
nor U7156 (N_7156,N_6599,N_6076);
or U7157 (N_7157,N_6491,N_6032);
nor U7158 (N_7158,N_6462,N_6725);
nand U7159 (N_7159,N_6289,N_6728);
nor U7160 (N_7160,N_6641,N_6342);
nor U7161 (N_7161,N_6398,N_6064);
nor U7162 (N_7162,N_6480,N_6397);
and U7163 (N_7163,N_6198,N_6692);
nor U7164 (N_7164,N_6023,N_6682);
xnor U7165 (N_7165,N_6246,N_6182);
nor U7166 (N_7166,N_6083,N_6304);
nor U7167 (N_7167,N_6504,N_6568);
nor U7168 (N_7168,N_6589,N_6349);
xnor U7169 (N_7169,N_6708,N_6247);
or U7170 (N_7170,N_6039,N_6436);
nor U7171 (N_7171,N_6555,N_6689);
and U7172 (N_7172,N_6381,N_6139);
nand U7173 (N_7173,N_6644,N_6027);
nand U7174 (N_7174,N_6374,N_6734);
or U7175 (N_7175,N_6545,N_6139);
nor U7176 (N_7176,N_6631,N_6336);
nand U7177 (N_7177,N_6425,N_6393);
nand U7178 (N_7178,N_6274,N_6024);
and U7179 (N_7179,N_6712,N_6666);
nand U7180 (N_7180,N_6587,N_6534);
nand U7181 (N_7181,N_6238,N_6226);
xnor U7182 (N_7182,N_6487,N_6536);
nand U7183 (N_7183,N_6007,N_6008);
nor U7184 (N_7184,N_6597,N_6173);
and U7185 (N_7185,N_6641,N_6018);
nor U7186 (N_7186,N_6359,N_6245);
or U7187 (N_7187,N_6391,N_6140);
xor U7188 (N_7188,N_6134,N_6666);
nand U7189 (N_7189,N_6431,N_6715);
or U7190 (N_7190,N_6106,N_6668);
nand U7191 (N_7191,N_6285,N_6033);
or U7192 (N_7192,N_6601,N_6212);
nand U7193 (N_7193,N_6741,N_6223);
and U7194 (N_7194,N_6476,N_6166);
or U7195 (N_7195,N_6598,N_6659);
nand U7196 (N_7196,N_6025,N_6102);
nand U7197 (N_7197,N_6583,N_6264);
and U7198 (N_7198,N_6255,N_6451);
nor U7199 (N_7199,N_6599,N_6038);
xnor U7200 (N_7200,N_6042,N_6125);
nor U7201 (N_7201,N_6531,N_6003);
nand U7202 (N_7202,N_6036,N_6233);
nand U7203 (N_7203,N_6722,N_6573);
and U7204 (N_7204,N_6103,N_6396);
nor U7205 (N_7205,N_6748,N_6461);
nor U7206 (N_7206,N_6683,N_6200);
nor U7207 (N_7207,N_6523,N_6543);
or U7208 (N_7208,N_6522,N_6188);
nor U7209 (N_7209,N_6165,N_6494);
or U7210 (N_7210,N_6268,N_6383);
and U7211 (N_7211,N_6513,N_6610);
nor U7212 (N_7212,N_6320,N_6240);
and U7213 (N_7213,N_6217,N_6597);
nor U7214 (N_7214,N_6498,N_6480);
nand U7215 (N_7215,N_6617,N_6654);
nand U7216 (N_7216,N_6108,N_6659);
and U7217 (N_7217,N_6215,N_6225);
or U7218 (N_7218,N_6366,N_6306);
nor U7219 (N_7219,N_6643,N_6343);
or U7220 (N_7220,N_6476,N_6255);
or U7221 (N_7221,N_6517,N_6646);
xor U7222 (N_7222,N_6324,N_6136);
nor U7223 (N_7223,N_6417,N_6522);
or U7224 (N_7224,N_6597,N_6338);
and U7225 (N_7225,N_6297,N_6414);
nand U7226 (N_7226,N_6529,N_6721);
and U7227 (N_7227,N_6308,N_6089);
nor U7228 (N_7228,N_6407,N_6104);
and U7229 (N_7229,N_6650,N_6454);
xnor U7230 (N_7230,N_6165,N_6187);
nand U7231 (N_7231,N_6523,N_6489);
nand U7232 (N_7232,N_6231,N_6635);
and U7233 (N_7233,N_6300,N_6552);
nor U7234 (N_7234,N_6480,N_6596);
xnor U7235 (N_7235,N_6319,N_6351);
nand U7236 (N_7236,N_6240,N_6124);
nand U7237 (N_7237,N_6724,N_6197);
nor U7238 (N_7238,N_6731,N_6471);
and U7239 (N_7239,N_6007,N_6498);
nand U7240 (N_7240,N_6208,N_6020);
and U7241 (N_7241,N_6434,N_6236);
xnor U7242 (N_7242,N_6219,N_6270);
nor U7243 (N_7243,N_6570,N_6342);
nor U7244 (N_7244,N_6626,N_6272);
nor U7245 (N_7245,N_6279,N_6268);
xnor U7246 (N_7246,N_6426,N_6583);
nor U7247 (N_7247,N_6703,N_6051);
and U7248 (N_7248,N_6223,N_6215);
or U7249 (N_7249,N_6536,N_6514);
and U7250 (N_7250,N_6437,N_6459);
nand U7251 (N_7251,N_6150,N_6059);
or U7252 (N_7252,N_6547,N_6292);
or U7253 (N_7253,N_6596,N_6036);
or U7254 (N_7254,N_6097,N_6517);
nor U7255 (N_7255,N_6598,N_6713);
nor U7256 (N_7256,N_6006,N_6407);
or U7257 (N_7257,N_6305,N_6039);
and U7258 (N_7258,N_6066,N_6044);
nor U7259 (N_7259,N_6701,N_6185);
or U7260 (N_7260,N_6507,N_6198);
and U7261 (N_7261,N_6167,N_6321);
or U7262 (N_7262,N_6682,N_6097);
nor U7263 (N_7263,N_6020,N_6303);
and U7264 (N_7264,N_6195,N_6366);
xnor U7265 (N_7265,N_6427,N_6101);
and U7266 (N_7266,N_6437,N_6618);
or U7267 (N_7267,N_6040,N_6501);
and U7268 (N_7268,N_6519,N_6390);
nor U7269 (N_7269,N_6324,N_6155);
nand U7270 (N_7270,N_6745,N_6587);
nor U7271 (N_7271,N_6010,N_6456);
nand U7272 (N_7272,N_6383,N_6642);
xnor U7273 (N_7273,N_6027,N_6229);
nand U7274 (N_7274,N_6710,N_6700);
xor U7275 (N_7275,N_6636,N_6499);
or U7276 (N_7276,N_6147,N_6568);
xor U7277 (N_7277,N_6182,N_6455);
xnor U7278 (N_7278,N_6020,N_6168);
or U7279 (N_7279,N_6289,N_6552);
and U7280 (N_7280,N_6556,N_6474);
nor U7281 (N_7281,N_6736,N_6584);
and U7282 (N_7282,N_6307,N_6102);
nor U7283 (N_7283,N_6662,N_6497);
or U7284 (N_7284,N_6191,N_6472);
or U7285 (N_7285,N_6393,N_6278);
and U7286 (N_7286,N_6654,N_6098);
nor U7287 (N_7287,N_6259,N_6586);
or U7288 (N_7288,N_6609,N_6126);
and U7289 (N_7289,N_6463,N_6236);
nor U7290 (N_7290,N_6249,N_6338);
or U7291 (N_7291,N_6116,N_6330);
nor U7292 (N_7292,N_6029,N_6000);
or U7293 (N_7293,N_6561,N_6094);
and U7294 (N_7294,N_6519,N_6379);
and U7295 (N_7295,N_6543,N_6022);
or U7296 (N_7296,N_6104,N_6224);
xor U7297 (N_7297,N_6577,N_6612);
or U7298 (N_7298,N_6153,N_6305);
or U7299 (N_7299,N_6337,N_6542);
nand U7300 (N_7300,N_6424,N_6334);
or U7301 (N_7301,N_6141,N_6615);
nand U7302 (N_7302,N_6584,N_6738);
nor U7303 (N_7303,N_6499,N_6179);
or U7304 (N_7304,N_6081,N_6523);
nand U7305 (N_7305,N_6084,N_6128);
or U7306 (N_7306,N_6506,N_6403);
nor U7307 (N_7307,N_6028,N_6620);
nor U7308 (N_7308,N_6056,N_6568);
or U7309 (N_7309,N_6062,N_6692);
nand U7310 (N_7310,N_6728,N_6324);
and U7311 (N_7311,N_6701,N_6239);
nand U7312 (N_7312,N_6323,N_6724);
and U7313 (N_7313,N_6377,N_6251);
or U7314 (N_7314,N_6068,N_6199);
and U7315 (N_7315,N_6553,N_6556);
or U7316 (N_7316,N_6620,N_6097);
nor U7317 (N_7317,N_6117,N_6215);
or U7318 (N_7318,N_6395,N_6426);
or U7319 (N_7319,N_6517,N_6128);
and U7320 (N_7320,N_6393,N_6436);
nand U7321 (N_7321,N_6533,N_6231);
xnor U7322 (N_7322,N_6388,N_6344);
nor U7323 (N_7323,N_6658,N_6540);
nand U7324 (N_7324,N_6346,N_6520);
xor U7325 (N_7325,N_6064,N_6036);
nand U7326 (N_7326,N_6416,N_6067);
nand U7327 (N_7327,N_6392,N_6085);
and U7328 (N_7328,N_6711,N_6085);
nor U7329 (N_7329,N_6593,N_6531);
nand U7330 (N_7330,N_6681,N_6073);
and U7331 (N_7331,N_6352,N_6305);
nor U7332 (N_7332,N_6007,N_6734);
nor U7333 (N_7333,N_6647,N_6511);
and U7334 (N_7334,N_6503,N_6733);
and U7335 (N_7335,N_6173,N_6350);
or U7336 (N_7336,N_6205,N_6075);
nor U7337 (N_7337,N_6684,N_6034);
and U7338 (N_7338,N_6559,N_6483);
or U7339 (N_7339,N_6110,N_6002);
nor U7340 (N_7340,N_6238,N_6081);
nand U7341 (N_7341,N_6616,N_6331);
or U7342 (N_7342,N_6585,N_6453);
nand U7343 (N_7343,N_6455,N_6691);
nand U7344 (N_7344,N_6582,N_6042);
xnor U7345 (N_7345,N_6340,N_6543);
or U7346 (N_7346,N_6694,N_6292);
or U7347 (N_7347,N_6644,N_6500);
nand U7348 (N_7348,N_6647,N_6152);
nand U7349 (N_7349,N_6431,N_6255);
and U7350 (N_7350,N_6304,N_6180);
xnor U7351 (N_7351,N_6429,N_6372);
xor U7352 (N_7352,N_6526,N_6155);
or U7353 (N_7353,N_6403,N_6383);
nand U7354 (N_7354,N_6058,N_6489);
nand U7355 (N_7355,N_6745,N_6066);
and U7356 (N_7356,N_6747,N_6744);
or U7357 (N_7357,N_6699,N_6157);
nand U7358 (N_7358,N_6426,N_6393);
nor U7359 (N_7359,N_6399,N_6084);
nand U7360 (N_7360,N_6092,N_6323);
nor U7361 (N_7361,N_6523,N_6690);
nand U7362 (N_7362,N_6043,N_6559);
and U7363 (N_7363,N_6147,N_6145);
and U7364 (N_7364,N_6698,N_6018);
or U7365 (N_7365,N_6634,N_6234);
or U7366 (N_7366,N_6000,N_6209);
nor U7367 (N_7367,N_6507,N_6105);
nand U7368 (N_7368,N_6123,N_6368);
nor U7369 (N_7369,N_6698,N_6435);
and U7370 (N_7370,N_6198,N_6444);
nor U7371 (N_7371,N_6601,N_6701);
and U7372 (N_7372,N_6377,N_6387);
nor U7373 (N_7373,N_6607,N_6074);
or U7374 (N_7374,N_6015,N_6471);
or U7375 (N_7375,N_6474,N_6528);
and U7376 (N_7376,N_6554,N_6183);
or U7377 (N_7377,N_6379,N_6021);
and U7378 (N_7378,N_6321,N_6558);
nand U7379 (N_7379,N_6359,N_6643);
nand U7380 (N_7380,N_6118,N_6382);
nand U7381 (N_7381,N_6741,N_6593);
nand U7382 (N_7382,N_6626,N_6134);
nor U7383 (N_7383,N_6545,N_6405);
or U7384 (N_7384,N_6107,N_6693);
or U7385 (N_7385,N_6146,N_6218);
or U7386 (N_7386,N_6662,N_6743);
nand U7387 (N_7387,N_6219,N_6351);
xnor U7388 (N_7388,N_6308,N_6665);
nand U7389 (N_7389,N_6333,N_6309);
and U7390 (N_7390,N_6190,N_6715);
nand U7391 (N_7391,N_6471,N_6611);
nand U7392 (N_7392,N_6126,N_6578);
xor U7393 (N_7393,N_6476,N_6068);
nor U7394 (N_7394,N_6451,N_6717);
and U7395 (N_7395,N_6469,N_6044);
and U7396 (N_7396,N_6029,N_6184);
nand U7397 (N_7397,N_6600,N_6682);
and U7398 (N_7398,N_6178,N_6221);
and U7399 (N_7399,N_6134,N_6432);
and U7400 (N_7400,N_6328,N_6380);
or U7401 (N_7401,N_6205,N_6322);
or U7402 (N_7402,N_6464,N_6717);
nor U7403 (N_7403,N_6693,N_6314);
nand U7404 (N_7404,N_6387,N_6227);
nand U7405 (N_7405,N_6624,N_6359);
and U7406 (N_7406,N_6061,N_6114);
and U7407 (N_7407,N_6417,N_6454);
and U7408 (N_7408,N_6748,N_6736);
and U7409 (N_7409,N_6012,N_6658);
nand U7410 (N_7410,N_6121,N_6164);
nand U7411 (N_7411,N_6272,N_6461);
nand U7412 (N_7412,N_6325,N_6569);
and U7413 (N_7413,N_6132,N_6034);
nor U7414 (N_7414,N_6186,N_6734);
xnor U7415 (N_7415,N_6011,N_6447);
nor U7416 (N_7416,N_6184,N_6577);
and U7417 (N_7417,N_6149,N_6140);
or U7418 (N_7418,N_6599,N_6120);
xor U7419 (N_7419,N_6190,N_6391);
nand U7420 (N_7420,N_6581,N_6437);
and U7421 (N_7421,N_6215,N_6126);
or U7422 (N_7422,N_6570,N_6094);
and U7423 (N_7423,N_6398,N_6153);
xor U7424 (N_7424,N_6353,N_6482);
nor U7425 (N_7425,N_6341,N_6179);
nor U7426 (N_7426,N_6511,N_6635);
nand U7427 (N_7427,N_6642,N_6017);
or U7428 (N_7428,N_6662,N_6071);
or U7429 (N_7429,N_6110,N_6458);
nor U7430 (N_7430,N_6029,N_6285);
nand U7431 (N_7431,N_6052,N_6561);
nor U7432 (N_7432,N_6565,N_6292);
or U7433 (N_7433,N_6402,N_6005);
and U7434 (N_7434,N_6134,N_6260);
or U7435 (N_7435,N_6281,N_6621);
nor U7436 (N_7436,N_6422,N_6703);
or U7437 (N_7437,N_6295,N_6451);
or U7438 (N_7438,N_6272,N_6335);
and U7439 (N_7439,N_6195,N_6270);
or U7440 (N_7440,N_6155,N_6204);
and U7441 (N_7441,N_6055,N_6739);
and U7442 (N_7442,N_6677,N_6162);
nor U7443 (N_7443,N_6070,N_6109);
nor U7444 (N_7444,N_6166,N_6271);
nand U7445 (N_7445,N_6540,N_6476);
and U7446 (N_7446,N_6116,N_6241);
and U7447 (N_7447,N_6022,N_6726);
or U7448 (N_7448,N_6241,N_6076);
nor U7449 (N_7449,N_6612,N_6515);
and U7450 (N_7450,N_6431,N_6199);
nor U7451 (N_7451,N_6035,N_6397);
and U7452 (N_7452,N_6118,N_6419);
and U7453 (N_7453,N_6701,N_6119);
or U7454 (N_7454,N_6131,N_6115);
or U7455 (N_7455,N_6340,N_6192);
nor U7456 (N_7456,N_6195,N_6575);
nor U7457 (N_7457,N_6187,N_6307);
and U7458 (N_7458,N_6738,N_6370);
nand U7459 (N_7459,N_6621,N_6017);
nor U7460 (N_7460,N_6460,N_6534);
and U7461 (N_7461,N_6466,N_6360);
xor U7462 (N_7462,N_6042,N_6611);
nor U7463 (N_7463,N_6055,N_6379);
and U7464 (N_7464,N_6344,N_6437);
or U7465 (N_7465,N_6049,N_6323);
and U7466 (N_7466,N_6221,N_6590);
xor U7467 (N_7467,N_6484,N_6026);
or U7468 (N_7468,N_6682,N_6374);
nand U7469 (N_7469,N_6371,N_6108);
or U7470 (N_7470,N_6526,N_6402);
nand U7471 (N_7471,N_6167,N_6612);
and U7472 (N_7472,N_6598,N_6480);
nor U7473 (N_7473,N_6725,N_6599);
nand U7474 (N_7474,N_6108,N_6174);
xnor U7475 (N_7475,N_6236,N_6621);
nor U7476 (N_7476,N_6484,N_6294);
and U7477 (N_7477,N_6183,N_6713);
nor U7478 (N_7478,N_6356,N_6327);
and U7479 (N_7479,N_6016,N_6056);
xor U7480 (N_7480,N_6346,N_6011);
nor U7481 (N_7481,N_6513,N_6442);
nor U7482 (N_7482,N_6556,N_6280);
xnor U7483 (N_7483,N_6323,N_6154);
or U7484 (N_7484,N_6446,N_6086);
or U7485 (N_7485,N_6592,N_6664);
nand U7486 (N_7486,N_6170,N_6303);
nand U7487 (N_7487,N_6198,N_6517);
nor U7488 (N_7488,N_6568,N_6293);
xor U7489 (N_7489,N_6433,N_6493);
nor U7490 (N_7490,N_6659,N_6101);
nor U7491 (N_7491,N_6533,N_6639);
nor U7492 (N_7492,N_6022,N_6050);
or U7493 (N_7493,N_6681,N_6041);
nand U7494 (N_7494,N_6505,N_6027);
nor U7495 (N_7495,N_6570,N_6617);
nand U7496 (N_7496,N_6157,N_6602);
and U7497 (N_7497,N_6648,N_6475);
nor U7498 (N_7498,N_6512,N_6428);
nor U7499 (N_7499,N_6277,N_6347);
and U7500 (N_7500,N_7290,N_7438);
or U7501 (N_7501,N_7393,N_7368);
nor U7502 (N_7502,N_7214,N_6842);
xor U7503 (N_7503,N_7338,N_6835);
nand U7504 (N_7504,N_7392,N_7359);
nand U7505 (N_7505,N_7265,N_6757);
and U7506 (N_7506,N_7286,N_7135);
and U7507 (N_7507,N_7361,N_7482);
and U7508 (N_7508,N_7322,N_6862);
nand U7509 (N_7509,N_6929,N_7232);
xor U7510 (N_7510,N_7484,N_6807);
or U7511 (N_7511,N_6993,N_7164);
nor U7512 (N_7512,N_7189,N_6819);
or U7513 (N_7513,N_7496,N_7159);
or U7514 (N_7514,N_7384,N_6755);
nor U7515 (N_7515,N_7009,N_7326);
or U7516 (N_7516,N_6945,N_7269);
or U7517 (N_7517,N_7068,N_7288);
nand U7518 (N_7518,N_7455,N_6784);
nor U7519 (N_7519,N_7499,N_7071);
xor U7520 (N_7520,N_6833,N_7405);
nand U7521 (N_7521,N_7031,N_6778);
or U7522 (N_7522,N_7398,N_7349);
nand U7523 (N_7523,N_7430,N_6915);
nor U7524 (N_7524,N_7259,N_7397);
and U7525 (N_7525,N_7495,N_6900);
nand U7526 (N_7526,N_7126,N_6793);
nor U7527 (N_7527,N_7419,N_7321);
nor U7528 (N_7528,N_7471,N_7141);
or U7529 (N_7529,N_7457,N_7001);
nor U7530 (N_7530,N_7012,N_7435);
and U7531 (N_7531,N_7160,N_6760);
or U7532 (N_7532,N_7025,N_6973);
or U7533 (N_7533,N_6999,N_6931);
and U7534 (N_7534,N_7400,N_6939);
xor U7535 (N_7535,N_6856,N_6913);
or U7536 (N_7536,N_7078,N_7377);
and U7537 (N_7537,N_7351,N_6919);
nand U7538 (N_7538,N_7032,N_7454);
or U7539 (N_7539,N_7390,N_7289);
and U7540 (N_7540,N_6866,N_6986);
and U7541 (N_7541,N_7373,N_7412);
nand U7542 (N_7542,N_7003,N_7328);
nand U7543 (N_7543,N_7313,N_7221);
and U7544 (N_7544,N_6927,N_6896);
and U7545 (N_7545,N_7305,N_6974);
nand U7546 (N_7546,N_7143,N_7279);
and U7547 (N_7547,N_7493,N_7278);
nand U7548 (N_7548,N_7169,N_7465);
or U7549 (N_7549,N_7103,N_6920);
nand U7550 (N_7550,N_7404,N_6924);
or U7551 (N_7551,N_7145,N_7040);
or U7552 (N_7552,N_7357,N_6858);
or U7553 (N_7553,N_7070,N_7415);
xor U7554 (N_7554,N_7249,N_7231);
and U7555 (N_7555,N_7475,N_6877);
nand U7556 (N_7556,N_7139,N_6957);
and U7557 (N_7557,N_7242,N_7476);
and U7558 (N_7558,N_7258,N_6911);
nor U7559 (N_7559,N_7191,N_7117);
nor U7560 (N_7560,N_7329,N_6841);
or U7561 (N_7561,N_7345,N_6815);
or U7562 (N_7562,N_7150,N_7355);
nand U7563 (N_7563,N_6776,N_6846);
xor U7564 (N_7564,N_7335,N_7367);
nor U7565 (N_7565,N_7051,N_6855);
nor U7566 (N_7566,N_7294,N_7134);
nor U7567 (N_7567,N_7247,N_6795);
nor U7568 (N_7568,N_7195,N_7101);
xnor U7569 (N_7569,N_7196,N_7156);
or U7570 (N_7570,N_7459,N_7488);
or U7571 (N_7571,N_6770,N_7133);
or U7572 (N_7572,N_6802,N_7203);
nand U7573 (N_7573,N_7206,N_6800);
nand U7574 (N_7574,N_7007,N_6948);
nor U7575 (N_7575,N_7467,N_7014);
or U7576 (N_7576,N_6863,N_7217);
nor U7577 (N_7577,N_7181,N_6792);
nand U7578 (N_7578,N_7152,N_7116);
and U7579 (N_7579,N_7030,N_7396);
or U7580 (N_7580,N_7386,N_7084);
and U7581 (N_7581,N_7416,N_6859);
and U7582 (N_7582,N_7016,N_7029);
xnor U7583 (N_7583,N_7251,N_6799);
nor U7584 (N_7584,N_6774,N_7082);
nor U7585 (N_7585,N_7244,N_6960);
and U7586 (N_7586,N_7375,N_6892);
nand U7587 (N_7587,N_7445,N_6910);
nor U7588 (N_7588,N_6798,N_7420);
nand U7589 (N_7589,N_6972,N_6752);
or U7590 (N_7590,N_7486,N_7093);
and U7591 (N_7591,N_7019,N_6830);
and U7592 (N_7592,N_7260,N_7151);
and U7593 (N_7593,N_7446,N_7055);
or U7594 (N_7594,N_7175,N_6959);
nand U7595 (N_7595,N_7287,N_7180);
xnor U7596 (N_7596,N_7474,N_7241);
and U7597 (N_7597,N_7198,N_7108);
and U7598 (N_7598,N_7276,N_6767);
or U7599 (N_7599,N_7268,N_6909);
nor U7600 (N_7600,N_6926,N_6982);
and U7601 (N_7601,N_7158,N_6963);
nor U7602 (N_7602,N_7077,N_7006);
nor U7603 (N_7603,N_6946,N_7118);
nand U7604 (N_7604,N_6822,N_7194);
nor U7605 (N_7605,N_6902,N_7138);
and U7606 (N_7606,N_7469,N_7312);
xnor U7607 (N_7607,N_7492,N_7490);
or U7608 (N_7608,N_6838,N_6994);
nand U7609 (N_7609,N_7215,N_7418);
nor U7610 (N_7610,N_7155,N_6810);
nor U7611 (N_7611,N_7255,N_7429);
and U7612 (N_7612,N_6895,N_7114);
xor U7613 (N_7613,N_7017,N_7491);
or U7614 (N_7614,N_7202,N_7046);
nor U7615 (N_7615,N_7171,N_7274);
or U7616 (N_7616,N_7065,N_7207);
nand U7617 (N_7617,N_6843,N_7240);
or U7618 (N_7618,N_6874,N_6906);
or U7619 (N_7619,N_6912,N_7256);
and U7620 (N_7620,N_7449,N_7153);
nor U7621 (N_7621,N_7154,N_7186);
nand U7622 (N_7622,N_7401,N_7026);
nor U7623 (N_7623,N_6780,N_7498);
nand U7624 (N_7624,N_6989,N_7324);
nor U7625 (N_7625,N_6901,N_6861);
and U7626 (N_7626,N_6781,N_6849);
nor U7627 (N_7627,N_7410,N_6873);
nor U7628 (N_7628,N_6857,N_6918);
or U7629 (N_7629,N_6992,N_6851);
nor U7630 (N_7630,N_7140,N_7450);
nor U7631 (N_7631,N_7489,N_6865);
nand U7632 (N_7632,N_7344,N_7237);
nor U7633 (N_7633,N_7443,N_7352);
nand U7634 (N_7634,N_6979,N_7226);
or U7635 (N_7635,N_7076,N_6949);
nand U7636 (N_7636,N_7297,N_7275);
and U7637 (N_7637,N_6821,N_6867);
and U7638 (N_7638,N_6935,N_7110);
nand U7639 (N_7639,N_7383,N_7057);
xnor U7640 (N_7640,N_7038,N_6875);
xnor U7641 (N_7641,N_6839,N_6816);
nor U7642 (N_7642,N_7147,N_7165);
nor U7643 (N_7643,N_6933,N_7044);
nand U7644 (N_7644,N_6758,N_7102);
nand U7645 (N_7645,N_7334,N_7358);
nand U7646 (N_7646,N_7075,N_6785);
or U7647 (N_7647,N_7130,N_7252);
nand U7648 (N_7648,N_7222,N_6951);
and U7649 (N_7649,N_7109,N_7376);
and U7650 (N_7650,N_6996,N_7149);
nor U7651 (N_7651,N_6884,N_7323);
xnor U7652 (N_7652,N_7127,N_7295);
nand U7653 (N_7653,N_7235,N_6970);
nor U7654 (N_7654,N_6832,N_7319);
nor U7655 (N_7655,N_7441,N_6987);
and U7656 (N_7656,N_6831,N_7122);
and U7657 (N_7657,N_7406,N_6940);
or U7658 (N_7658,N_7172,N_7049);
or U7659 (N_7659,N_6783,N_6947);
or U7660 (N_7660,N_7285,N_7059);
or U7661 (N_7661,N_7119,N_7088);
and U7662 (N_7662,N_7188,N_7060);
xor U7663 (N_7663,N_7485,N_6768);
xnor U7664 (N_7664,N_7021,N_7477);
nand U7665 (N_7665,N_6791,N_7052);
xnor U7666 (N_7666,N_6932,N_7472);
nor U7667 (N_7667,N_6789,N_7163);
or U7668 (N_7668,N_6847,N_7316);
nand U7669 (N_7669,N_7142,N_7374);
nor U7670 (N_7670,N_7079,N_6983);
xor U7671 (N_7671,N_7183,N_7028);
and U7672 (N_7672,N_6864,N_7098);
and U7673 (N_7673,N_7096,N_7364);
xor U7674 (N_7674,N_7131,N_6990);
nor U7675 (N_7675,N_7456,N_7213);
or U7676 (N_7676,N_6897,N_6828);
nand U7677 (N_7677,N_7094,N_6890);
nor U7678 (N_7678,N_7166,N_6905);
nor U7679 (N_7679,N_7440,N_6881);
xnor U7680 (N_7680,N_6790,N_7085);
or U7681 (N_7681,N_7092,N_7487);
nand U7682 (N_7682,N_7343,N_7434);
or U7683 (N_7683,N_6891,N_7437);
nor U7684 (N_7684,N_7327,N_7246);
or U7685 (N_7685,N_7107,N_7233);
nor U7686 (N_7686,N_7023,N_7378);
nand U7687 (N_7687,N_6981,N_6808);
xnor U7688 (N_7688,N_7366,N_7413);
and U7689 (N_7689,N_6812,N_7080);
nand U7690 (N_7690,N_6777,N_6955);
and U7691 (N_7691,N_6950,N_6764);
or U7692 (N_7692,N_7005,N_6942);
nand U7693 (N_7693,N_7381,N_7033);
nor U7694 (N_7694,N_7045,N_7043);
xor U7695 (N_7695,N_7190,N_7220);
and U7696 (N_7696,N_7199,N_7011);
or U7697 (N_7697,N_7216,N_7425);
nand U7698 (N_7698,N_7253,N_6888);
nor U7699 (N_7699,N_7168,N_6977);
nand U7700 (N_7700,N_6882,N_7053);
nor U7701 (N_7701,N_7004,N_6907);
nand U7702 (N_7702,N_7162,N_6969);
or U7703 (N_7703,N_7185,N_7097);
and U7704 (N_7704,N_7061,N_7081);
and U7705 (N_7705,N_7270,N_7447);
or U7706 (N_7706,N_7174,N_7090);
nand U7707 (N_7707,N_7058,N_7308);
xnor U7708 (N_7708,N_7315,N_7365);
nor U7709 (N_7709,N_6925,N_6968);
or U7710 (N_7710,N_7144,N_7362);
xor U7711 (N_7711,N_7264,N_7304);
nor U7712 (N_7712,N_7218,N_7111);
nor U7713 (N_7713,N_7320,N_7099);
xnor U7714 (N_7714,N_6965,N_7219);
nand U7715 (N_7715,N_6876,N_7347);
nand U7716 (N_7716,N_7027,N_7243);
nand U7717 (N_7717,N_7042,N_6756);
nand U7718 (N_7718,N_7238,N_7481);
nor U7719 (N_7719,N_7192,N_7224);
nand U7720 (N_7720,N_6854,N_6850);
nand U7721 (N_7721,N_7035,N_7281);
and U7722 (N_7722,N_6872,N_7010);
nand U7723 (N_7723,N_6771,N_7337);
and U7724 (N_7724,N_7262,N_7466);
and U7725 (N_7725,N_7372,N_7056);
or U7726 (N_7726,N_7125,N_6887);
or U7727 (N_7727,N_6788,N_6765);
nor U7728 (N_7728,N_7248,N_6811);
or U7729 (N_7729,N_7123,N_7385);
nand U7730 (N_7730,N_7417,N_7064);
nor U7731 (N_7731,N_6952,N_7179);
or U7732 (N_7732,N_7483,N_7271);
xor U7733 (N_7733,N_6796,N_7066);
xor U7734 (N_7734,N_7132,N_7228);
nor U7735 (N_7735,N_6904,N_6797);
nand U7736 (N_7736,N_7414,N_7409);
or U7737 (N_7737,N_6984,N_7239);
or U7738 (N_7738,N_6769,N_6880);
or U7739 (N_7739,N_6921,N_7301);
xnor U7740 (N_7740,N_7284,N_6786);
and U7741 (N_7741,N_6885,N_6825);
nand U7742 (N_7742,N_7353,N_7054);
or U7743 (N_7743,N_7048,N_6988);
nand U7744 (N_7744,N_7015,N_7382);
or U7745 (N_7745,N_6967,N_7293);
nand U7746 (N_7746,N_6916,N_7310);
xnor U7747 (N_7747,N_7148,N_6953);
and U7748 (N_7748,N_7176,N_6943);
and U7749 (N_7749,N_6827,N_7037);
and U7750 (N_7750,N_6848,N_6779);
nand U7751 (N_7751,N_7369,N_7105);
and U7752 (N_7752,N_7212,N_7480);
or U7753 (N_7753,N_7063,N_7451);
nand U7754 (N_7754,N_6844,N_7403);
or U7755 (N_7755,N_7340,N_7177);
nor U7756 (N_7756,N_6868,N_7356);
or U7757 (N_7757,N_6813,N_7234);
xnor U7758 (N_7758,N_6934,N_7047);
and U7759 (N_7759,N_7291,N_7432);
or U7760 (N_7760,N_7000,N_6995);
nor U7761 (N_7761,N_7250,N_7433);
or U7762 (N_7762,N_7436,N_7354);
and U7763 (N_7763,N_6908,N_7086);
and U7764 (N_7764,N_7205,N_6878);
or U7765 (N_7765,N_6894,N_7442);
nor U7766 (N_7766,N_7298,N_6936);
and U7767 (N_7767,N_6775,N_7089);
or U7768 (N_7768,N_7245,N_6930);
or U7769 (N_7769,N_6903,N_6870);
or U7770 (N_7770,N_6823,N_7204);
nor U7771 (N_7771,N_6818,N_6751);
and U7772 (N_7772,N_7306,N_7303);
nand U7773 (N_7773,N_6966,N_7309);
xor U7774 (N_7774,N_7399,N_7494);
and U7775 (N_7775,N_7339,N_7193);
and U7776 (N_7776,N_7113,N_7273);
and U7777 (N_7777,N_7106,N_7261);
nand U7778 (N_7778,N_7277,N_7227);
or U7779 (N_7779,N_7104,N_7464);
or U7780 (N_7780,N_7317,N_6820);
nand U7781 (N_7781,N_6997,N_6845);
nor U7782 (N_7782,N_7318,N_6879);
nand U7783 (N_7783,N_6923,N_7091);
nor U7784 (N_7784,N_6886,N_6893);
xor U7785 (N_7785,N_7333,N_7041);
and U7786 (N_7786,N_7209,N_7395);
xor U7787 (N_7787,N_7254,N_7002);
nor U7788 (N_7788,N_7167,N_7008);
nor U7789 (N_7789,N_7307,N_7391);
and U7790 (N_7790,N_7330,N_6998);
nor U7791 (N_7791,N_7427,N_7263);
nand U7792 (N_7792,N_7020,N_6817);
and U7793 (N_7793,N_6917,N_7407);
or U7794 (N_7794,N_7095,N_7311);
nor U7795 (N_7795,N_7426,N_7266);
and U7796 (N_7796,N_6824,N_7100);
nand U7797 (N_7797,N_6961,N_6883);
and U7798 (N_7798,N_6871,N_6801);
or U7799 (N_7799,N_7453,N_6809);
nor U7800 (N_7800,N_7423,N_7018);
nor U7801 (N_7801,N_6899,N_7282);
or U7802 (N_7802,N_6938,N_6826);
and U7803 (N_7803,N_7341,N_7034);
and U7804 (N_7804,N_7013,N_7473);
and U7805 (N_7805,N_7348,N_7074);
xor U7806 (N_7806,N_6852,N_6836);
xor U7807 (N_7807,N_7115,N_6944);
and U7808 (N_7808,N_7463,N_7036);
nor U7809 (N_7809,N_6853,N_7422);
xnor U7810 (N_7810,N_7112,N_7230);
nor U7811 (N_7811,N_7267,N_7050);
and U7812 (N_7812,N_7462,N_7121);
nor U7813 (N_7813,N_6834,N_7363);
and U7814 (N_7814,N_7039,N_6772);
nand U7815 (N_7815,N_7137,N_7411);
nor U7816 (N_7816,N_7073,N_6787);
nor U7817 (N_7817,N_7087,N_6928);
or U7818 (N_7818,N_7452,N_7302);
and U7819 (N_7819,N_6803,N_6889);
or U7820 (N_7820,N_7062,N_6761);
and U7821 (N_7821,N_7182,N_7439);
nor U7822 (N_7822,N_7072,N_7370);
nand U7823 (N_7823,N_7200,N_7067);
and U7824 (N_7824,N_7211,N_7187);
and U7825 (N_7825,N_6860,N_6922);
nor U7826 (N_7826,N_7283,N_7325);
nor U7827 (N_7827,N_7342,N_7428);
nor U7828 (N_7828,N_7458,N_7360);
or U7829 (N_7829,N_6958,N_7387);
and U7830 (N_7830,N_6898,N_7022);
nand U7831 (N_7831,N_6773,N_7146);
xnor U7832 (N_7832,N_6941,N_6763);
nand U7833 (N_7833,N_7300,N_7346);
or U7834 (N_7834,N_7157,N_6980);
xor U7835 (N_7835,N_6991,N_6766);
or U7836 (N_7836,N_6829,N_6806);
or U7837 (N_7837,N_6937,N_7479);
nor U7838 (N_7838,N_7083,N_6975);
nand U7839 (N_7839,N_6754,N_7379);
and U7840 (N_7840,N_7394,N_7208);
and U7841 (N_7841,N_7460,N_6804);
nor U7842 (N_7842,N_6753,N_7184);
nand U7843 (N_7843,N_6976,N_7350);
or U7844 (N_7844,N_6985,N_6794);
or U7845 (N_7845,N_7229,N_7448);
or U7846 (N_7846,N_7402,N_7331);
and U7847 (N_7847,N_7332,N_7424);
or U7848 (N_7848,N_7136,N_7421);
xnor U7849 (N_7849,N_6956,N_6869);
nor U7850 (N_7850,N_7124,N_6782);
and U7851 (N_7851,N_6840,N_6914);
or U7852 (N_7852,N_7444,N_7225);
nor U7853 (N_7853,N_7408,N_7178);
and U7854 (N_7854,N_7371,N_7296);
or U7855 (N_7855,N_6954,N_7299);
xnor U7856 (N_7856,N_7170,N_7257);
nand U7857 (N_7857,N_7431,N_7380);
or U7858 (N_7858,N_7336,N_6814);
nand U7859 (N_7859,N_6759,N_6762);
or U7860 (N_7860,N_7210,N_7292);
nor U7861 (N_7861,N_6837,N_6964);
nor U7862 (N_7862,N_7129,N_7120);
or U7863 (N_7863,N_7478,N_7470);
or U7864 (N_7864,N_6750,N_7128);
and U7865 (N_7865,N_7223,N_7161);
or U7866 (N_7866,N_6971,N_6962);
and U7867 (N_7867,N_7069,N_7197);
and U7868 (N_7868,N_7389,N_7280);
nand U7869 (N_7869,N_6805,N_7468);
and U7870 (N_7870,N_7024,N_7236);
xor U7871 (N_7871,N_7461,N_7388);
or U7872 (N_7872,N_7272,N_7314);
and U7873 (N_7873,N_7201,N_6978);
nor U7874 (N_7874,N_7173,N_7497);
and U7875 (N_7875,N_6927,N_7106);
nand U7876 (N_7876,N_7134,N_6919);
nand U7877 (N_7877,N_7427,N_6920);
or U7878 (N_7878,N_7054,N_7016);
nor U7879 (N_7879,N_6780,N_6806);
or U7880 (N_7880,N_7135,N_7456);
and U7881 (N_7881,N_7033,N_6770);
nor U7882 (N_7882,N_7038,N_7219);
or U7883 (N_7883,N_7391,N_7356);
or U7884 (N_7884,N_7101,N_7379);
and U7885 (N_7885,N_6764,N_7238);
nor U7886 (N_7886,N_7215,N_7269);
and U7887 (N_7887,N_7023,N_7178);
nand U7888 (N_7888,N_6786,N_7243);
nor U7889 (N_7889,N_6828,N_7038);
nor U7890 (N_7890,N_6943,N_6816);
nor U7891 (N_7891,N_7164,N_7369);
nor U7892 (N_7892,N_7360,N_7075);
or U7893 (N_7893,N_7307,N_7056);
or U7894 (N_7894,N_6933,N_7448);
or U7895 (N_7895,N_7160,N_6974);
and U7896 (N_7896,N_7376,N_7424);
and U7897 (N_7897,N_7447,N_7260);
nor U7898 (N_7898,N_6750,N_7187);
xor U7899 (N_7899,N_6997,N_7487);
and U7900 (N_7900,N_7433,N_6985);
and U7901 (N_7901,N_7270,N_6785);
xnor U7902 (N_7902,N_6813,N_7381);
nor U7903 (N_7903,N_6768,N_7442);
and U7904 (N_7904,N_6950,N_7089);
nor U7905 (N_7905,N_7222,N_7415);
nor U7906 (N_7906,N_7033,N_7142);
xnor U7907 (N_7907,N_6788,N_7406);
or U7908 (N_7908,N_7295,N_7181);
xnor U7909 (N_7909,N_6942,N_6800);
xnor U7910 (N_7910,N_7393,N_6877);
or U7911 (N_7911,N_6801,N_7413);
nor U7912 (N_7912,N_7407,N_6760);
nor U7913 (N_7913,N_7167,N_7111);
or U7914 (N_7914,N_7485,N_7247);
nand U7915 (N_7915,N_7345,N_7074);
nor U7916 (N_7916,N_6795,N_7024);
or U7917 (N_7917,N_7495,N_7197);
nor U7918 (N_7918,N_7236,N_7144);
nand U7919 (N_7919,N_7379,N_7196);
and U7920 (N_7920,N_6961,N_7177);
nor U7921 (N_7921,N_7169,N_6859);
nor U7922 (N_7922,N_6792,N_6897);
xnor U7923 (N_7923,N_7438,N_7471);
nor U7924 (N_7924,N_6765,N_6895);
nor U7925 (N_7925,N_7399,N_7286);
nor U7926 (N_7926,N_7411,N_7060);
xnor U7927 (N_7927,N_6892,N_6761);
xor U7928 (N_7928,N_7415,N_7206);
nand U7929 (N_7929,N_7140,N_7059);
or U7930 (N_7930,N_7230,N_7149);
nor U7931 (N_7931,N_7095,N_6926);
nor U7932 (N_7932,N_7069,N_7477);
or U7933 (N_7933,N_6781,N_7265);
and U7934 (N_7934,N_6858,N_7298);
nand U7935 (N_7935,N_7223,N_7041);
nor U7936 (N_7936,N_7472,N_6840);
and U7937 (N_7937,N_7158,N_7170);
nand U7938 (N_7938,N_6892,N_7120);
nor U7939 (N_7939,N_7206,N_7081);
and U7940 (N_7940,N_7313,N_6813);
xnor U7941 (N_7941,N_6823,N_6959);
or U7942 (N_7942,N_6820,N_6922);
and U7943 (N_7943,N_7104,N_7099);
nand U7944 (N_7944,N_6911,N_7003);
or U7945 (N_7945,N_6848,N_7488);
and U7946 (N_7946,N_7103,N_7100);
nor U7947 (N_7947,N_6986,N_7403);
nor U7948 (N_7948,N_7424,N_7483);
nand U7949 (N_7949,N_7413,N_7337);
or U7950 (N_7950,N_6916,N_7391);
nand U7951 (N_7951,N_7152,N_6773);
nand U7952 (N_7952,N_7305,N_6964);
nor U7953 (N_7953,N_6789,N_7470);
nor U7954 (N_7954,N_6800,N_7259);
and U7955 (N_7955,N_6930,N_6912);
or U7956 (N_7956,N_7295,N_6854);
nor U7957 (N_7957,N_6916,N_6965);
nor U7958 (N_7958,N_7013,N_7162);
nor U7959 (N_7959,N_7181,N_7006);
and U7960 (N_7960,N_6842,N_7108);
and U7961 (N_7961,N_7406,N_6965);
nand U7962 (N_7962,N_6756,N_7219);
nor U7963 (N_7963,N_6975,N_6758);
xor U7964 (N_7964,N_7217,N_6759);
nor U7965 (N_7965,N_7400,N_7036);
and U7966 (N_7966,N_7319,N_7442);
nor U7967 (N_7967,N_7319,N_7315);
or U7968 (N_7968,N_6825,N_7404);
nand U7969 (N_7969,N_7304,N_6979);
nor U7970 (N_7970,N_7307,N_7285);
and U7971 (N_7971,N_6902,N_7445);
or U7972 (N_7972,N_7137,N_7339);
nor U7973 (N_7973,N_7285,N_7366);
and U7974 (N_7974,N_7353,N_7245);
and U7975 (N_7975,N_7215,N_6903);
nand U7976 (N_7976,N_6840,N_7494);
or U7977 (N_7977,N_7478,N_7037);
and U7978 (N_7978,N_6763,N_7153);
or U7979 (N_7979,N_6882,N_7247);
nor U7980 (N_7980,N_7481,N_6929);
nor U7981 (N_7981,N_7167,N_7228);
or U7982 (N_7982,N_7201,N_7432);
or U7983 (N_7983,N_7320,N_7234);
nand U7984 (N_7984,N_6902,N_6839);
and U7985 (N_7985,N_6760,N_7208);
nand U7986 (N_7986,N_7293,N_6919);
and U7987 (N_7987,N_7121,N_6921);
and U7988 (N_7988,N_7085,N_7496);
or U7989 (N_7989,N_7238,N_7212);
nor U7990 (N_7990,N_7231,N_7243);
or U7991 (N_7991,N_6984,N_7106);
nor U7992 (N_7992,N_6926,N_7284);
nor U7993 (N_7993,N_7473,N_6951);
nor U7994 (N_7994,N_7086,N_7392);
xnor U7995 (N_7995,N_6870,N_7114);
xor U7996 (N_7996,N_6953,N_6863);
and U7997 (N_7997,N_7246,N_7115);
nand U7998 (N_7998,N_7391,N_7207);
nor U7999 (N_7999,N_7013,N_7232);
and U8000 (N_8000,N_7301,N_7381);
xor U8001 (N_8001,N_7298,N_7238);
or U8002 (N_8002,N_7262,N_7260);
or U8003 (N_8003,N_7341,N_6848);
and U8004 (N_8004,N_7363,N_7445);
or U8005 (N_8005,N_6978,N_7427);
nor U8006 (N_8006,N_7147,N_7471);
and U8007 (N_8007,N_6861,N_6956);
nor U8008 (N_8008,N_7301,N_6959);
nor U8009 (N_8009,N_7379,N_7075);
xor U8010 (N_8010,N_7179,N_6997);
nand U8011 (N_8011,N_7096,N_7226);
or U8012 (N_8012,N_7346,N_7033);
and U8013 (N_8013,N_6952,N_7273);
or U8014 (N_8014,N_7334,N_6902);
or U8015 (N_8015,N_7162,N_7133);
nand U8016 (N_8016,N_6833,N_7019);
and U8017 (N_8017,N_6809,N_7145);
nor U8018 (N_8018,N_7128,N_7389);
and U8019 (N_8019,N_6916,N_7209);
and U8020 (N_8020,N_6977,N_7467);
nand U8021 (N_8021,N_7004,N_7211);
and U8022 (N_8022,N_6774,N_7258);
and U8023 (N_8023,N_6929,N_7428);
nand U8024 (N_8024,N_6919,N_7230);
nor U8025 (N_8025,N_7043,N_7048);
or U8026 (N_8026,N_6758,N_7442);
nand U8027 (N_8027,N_6775,N_7273);
nand U8028 (N_8028,N_6879,N_6861);
xnor U8029 (N_8029,N_7483,N_6825);
or U8030 (N_8030,N_7168,N_7023);
nand U8031 (N_8031,N_6988,N_6816);
nor U8032 (N_8032,N_6830,N_7084);
and U8033 (N_8033,N_6988,N_7341);
xor U8034 (N_8034,N_7401,N_7147);
and U8035 (N_8035,N_7466,N_7175);
or U8036 (N_8036,N_7170,N_7268);
or U8037 (N_8037,N_6780,N_7107);
nor U8038 (N_8038,N_7489,N_6778);
nand U8039 (N_8039,N_6820,N_7017);
nand U8040 (N_8040,N_6986,N_7188);
nor U8041 (N_8041,N_7175,N_7001);
and U8042 (N_8042,N_7126,N_7217);
nor U8043 (N_8043,N_7339,N_7040);
or U8044 (N_8044,N_7256,N_7443);
nand U8045 (N_8045,N_7086,N_7085);
nand U8046 (N_8046,N_7459,N_7417);
nor U8047 (N_8047,N_6850,N_6897);
xnor U8048 (N_8048,N_6803,N_7276);
nand U8049 (N_8049,N_6769,N_7079);
nor U8050 (N_8050,N_7368,N_6759);
xnor U8051 (N_8051,N_6800,N_7113);
or U8052 (N_8052,N_6833,N_7295);
nor U8053 (N_8053,N_7210,N_7155);
nand U8054 (N_8054,N_7487,N_7420);
and U8055 (N_8055,N_7161,N_7257);
nor U8056 (N_8056,N_6916,N_7424);
or U8057 (N_8057,N_7475,N_7415);
nor U8058 (N_8058,N_6930,N_7285);
and U8059 (N_8059,N_7362,N_6865);
nor U8060 (N_8060,N_7044,N_7442);
or U8061 (N_8061,N_7099,N_6895);
nor U8062 (N_8062,N_7292,N_6933);
xnor U8063 (N_8063,N_7047,N_7439);
or U8064 (N_8064,N_6838,N_7165);
or U8065 (N_8065,N_7413,N_7487);
and U8066 (N_8066,N_7343,N_6845);
and U8067 (N_8067,N_7202,N_7015);
nor U8068 (N_8068,N_6922,N_7028);
nor U8069 (N_8069,N_7205,N_6774);
and U8070 (N_8070,N_7401,N_6792);
nor U8071 (N_8071,N_7245,N_7495);
and U8072 (N_8072,N_6984,N_7488);
nand U8073 (N_8073,N_6870,N_6850);
nand U8074 (N_8074,N_7407,N_6957);
and U8075 (N_8075,N_7426,N_7128);
nor U8076 (N_8076,N_6819,N_7150);
xor U8077 (N_8077,N_7335,N_6893);
or U8078 (N_8078,N_6947,N_7243);
or U8079 (N_8079,N_7153,N_7439);
xor U8080 (N_8080,N_7059,N_7159);
and U8081 (N_8081,N_7136,N_7449);
nor U8082 (N_8082,N_7088,N_7056);
or U8083 (N_8083,N_7232,N_7168);
xnor U8084 (N_8084,N_7173,N_7215);
and U8085 (N_8085,N_7326,N_6851);
nand U8086 (N_8086,N_6978,N_6963);
or U8087 (N_8087,N_7162,N_7328);
or U8088 (N_8088,N_7103,N_6935);
or U8089 (N_8089,N_7324,N_6934);
and U8090 (N_8090,N_6886,N_7497);
nor U8091 (N_8091,N_7115,N_7181);
nor U8092 (N_8092,N_6931,N_6911);
or U8093 (N_8093,N_7471,N_6979);
and U8094 (N_8094,N_7446,N_7004);
nand U8095 (N_8095,N_7382,N_7355);
or U8096 (N_8096,N_7074,N_7337);
and U8097 (N_8097,N_7157,N_7442);
nand U8098 (N_8098,N_6933,N_7391);
and U8099 (N_8099,N_7016,N_6853);
nor U8100 (N_8100,N_7164,N_7411);
xnor U8101 (N_8101,N_7268,N_7252);
nor U8102 (N_8102,N_6870,N_6822);
and U8103 (N_8103,N_7086,N_7379);
nor U8104 (N_8104,N_6769,N_7453);
or U8105 (N_8105,N_7454,N_7216);
nor U8106 (N_8106,N_6802,N_7284);
nand U8107 (N_8107,N_7250,N_7397);
xnor U8108 (N_8108,N_7026,N_7174);
nor U8109 (N_8109,N_6896,N_6905);
and U8110 (N_8110,N_6948,N_7365);
and U8111 (N_8111,N_6802,N_7491);
xor U8112 (N_8112,N_7473,N_6971);
nand U8113 (N_8113,N_7041,N_7113);
and U8114 (N_8114,N_7181,N_7042);
or U8115 (N_8115,N_7478,N_7388);
or U8116 (N_8116,N_7245,N_6999);
or U8117 (N_8117,N_7468,N_7015);
or U8118 (N_8118,N_6803,N_7484);
and U8119 (N_8119,N_7400,N_7321);
nand U8120 (N_8120,N_6933,N_7100);
nor U8121 (N_8121,N_6977,N_6765);
or U8122 (N_8122,N_6802,N_6919);
nand U8123 (N_8123,N_7474,N_7021);
or U8124 (N_8124,N_6767,N_6877);
or U8125 (N_8125,N_6778,N_6998);
nand U8126 (N_8126,N_6980,N_7144);
nor U8127 (N_8127,N_6791,N_7037);
or U8128 (N_8128,N_7171,N_6955);
and U8129 (N_8129,N_7390,N_7292);
xnor U8130 (N_8130,N_7341,N_7089);
and U8131 (N_8131,N_7303,N_7410);
nand U8132 (N_8132,N_7095,N_7387);
nand U8133 (N_8133,N_7112,N_7141);
nor U8134 (N_8134,N_6857,N_7390);
nand U8135 (N_8135,N_7199,N_7270);
xnor U8136 (N_8136,N_7079,N_6874);
nor U8137 (N_8137,N_7488,N_7362);
nor U8138 (N_8138,N_7133,N_7273);
nor U8139 (N_8139,N_7148,N_6921);
and U8140 (N_8140,N_6887,N_7307);
or U8141 (N_8141,N_7389,N_6973);
or U8142 (N_8142,N_7283,N_6831);
nand U8143 (N_8143,N_6815,N_6989);
xnor U8144 (N_8144,N_6876,N_7320);
nand U8145 (N_8145,N_6866,N_7498);
nor U8146 (N_8146,N_6785,N_6837);
nand U8147 (N_8147,N_7118,N_6764);
xnor U8148 (N_8148,N_7083,N_7244);
nand U8149 (N_8149,N_7449,N_6879);
xnor U8150 (N_8150,N_7137,N_7445);
nand U8151 (N_8151,N_7339,N_6962);
and U8152 (N_8152,N_7116,N_7320);
and U8153 (N_8153,N_7466,N_7000);
or U8154 (N_8154,N_7220,N_7399);
and U8155 (N_8155,N_6777,N_7173);
nand U8156 (N_8156,N_6798,N_7342);
or U8157 (N_8157,N_6901,N_7227);
nand U8158 (N_8158,N_7129,N_7350);
or U8159 (N_8159,N_7413,N_7499);
nand U8160 (N_8160,N_7101,N_7332);
or U8161 (N_8161,N_7286,N_7390);
nand U8162 (N_8162,N_6842,N_7250);
and U8163 (N_8163,N_6909,N_7165);
nor U8164 (N_8164,N_6962,N_7077);
xnor U8165 (N_8165,N_7148,N_7213);
nand U8166 (N_8166,N_7396,N_6920);
or U8167 (N_8167,N_7336,N_6987);
nor U8168 (N_8168,N_7260,N_7431);
and U8169 (N_8169,N_7409,N_6793);
nand U8170 (N_8170,N_6896,N_7102);
nor U8171 (N_8171,N_6768,N_7480);
nor U8172 (N_8172,N_6756,N_6979);
nor U8173 (N_8173,N_7350,N_7330);
nor U8174 (N_8174,N_7343,N_7054);
and U8175 (N_8175,N_7203,N_7074);
or U8176 (N_8176,N_6806,N_7134);
nand U8177 (N_8177,N_7343,N_6823);
nor U8178 (N_8178,N_6815,N_7012);
nand U8179 (N_8179,N_6813,N_7409);
or U8180 (N_8180,N_7272,N_6854);
or U8181 (N_8181,N_6960,N_7119);
and U8182 (N_8182,N_7213,N_7299);
or U8183 (N_8183,N_7382,N_7484);
nand U8184 (N_8184,N_6896,N_6783);
nor U8185 (N_8185,N_7082,N_7320);
and U8186 (N_8186,N_7041,N_7427);
and U8187 (N_8187,N_7071,N_7177);
nor U8188 (N_8188,N_7247,N_7374);
or U8189 (N_8189,N_7396,N_6879);
nor U8190 (N_8190,N_7079,N_7287);
or U8191 (N_8191,N_7436,N_7432);
nand U8192 (N_8192,N_7272,N_6924);
nor U8193 (N_8193,N_6809,N_7061);
nand U8194 (N_8194,N_7091,N_7116);
nor U8195 (N_8195,N_7196,N_7402);
nor U8196 (N_8196,N_7486,N_6927);
and U8197 (N_8197,N_7208,N_7379);
nor U8198 (N_8198,N_7028,N_7053);
or U8199 (N_8199,N_6836,N_7236);
or U8200 (N_8200,N_6954,N_6995);
and U8201 (N_8201,N_7172,N_6928);
and U8202 (N_8202,N_6778,N_6770);
and U8203 (N_8203,N_7253,N_7428);
and U8204 (N_8204,N_7312,N_6913);
xnor U8205 (N_8205,N_7376,N_6832);
nand U8206 (N_8206,N_6978,N_7113);
nand U8207 (N_8207,N_7439,N_6983);
nor U8208 (N_8208,N_7223,N_7436);
nor U8209 (N_8209,N_6901,N_6946);
nor U8210 (N_8210,N_6880,N_7016);
xor U8211 (N_8211,N_6845,N_7124);
nand U8212 (N_8212,N_7091,N_7199);
nand U8213 (N_8213,N_7372,N_7356);
nor U8214 (N_8214,N_7143,N_7383);
nor U8215 (N_8215,N_6818,N_7130);
nand U8216 (N_8216,N_7174,N_7397);
nor U8217 (N_8217,N_7262,N_7467);
xnor U8218 (N_8218,N_7194,N_6903);
and U8219 (N_8219,N_7130,N_6900);
nor U8220 (N_8220,N_7286,N_7275);
nor U8221 (N_8221,N_7118,N_7202);
xor U8222 (N_8222,N_7342,N_6917);
or U8223 (N_8223,N_7347,N_6753);
and U8224 (N_8224,N_7238,N_6916);
and U8225 (N_8225,N_6855,N_6951);
and U8226 (N_8226,N_7427,N_7348);
and U8227 (N_8227,N_6930,N_6829);
and U8228 (N_8228,N_7128,N_7173);
nor U8229 (N_8229,N_7469,N_6851);
nor U8230 (N_8230,N_7093,N_7020);
or U8231 (N_8231,N_6805,N_7332);
or U8232 (N_8232,N_7297,N_6900);
xor U8233 (N_8233,N_6835,N_6792);
or U8234 (N_8234,N_7061,N_7176);
nand U8235 (N_8235,N_7046,N_6870);
nand U8236 (N_8236,N_7435,N_7383);
and U8237 (N_8237,N_6960,N_6801);
nor U8238 (N_8238,N_7460,N_6873);
nand U8239 (N_8239,N_7080,N_7479);
or U8240 (N_8240,N_7393,N_6820);
xor U8241 (N_8241,N_7433,N_7498);
nor U8242 (N_8242,N_7314,N_7304);
and U8243 (N_8243,N_7403,N_7471);
or U8244 (N_8244,N_7362,N_7083);
nor U8245 (N_8245,N_7368,N_6755);
nand U8246 (N_8246,N_7394,N_6861);
nand U8247 (N_8247,N_6854,N_6832);
nor U8248 (N_8248,N_7161,N_7059);
nand U8249 (N_8249,N_6861,N_7257);
nand U8250 (N_8250,N_8069,N_7533);
xnor U8251 (N_8251,N_8132,N_7686);
nor U8252 (N_8252,N_7811,N_8074);
xnor U8253 (N_8253,N_7973,N_7831);
and U8254 (N_8254,N_7992,N_7613);
nand U8255 (N_8255,N_7968,N_7738);
nand U8256 (N_8256,N_7753,N_7893);
and U8257 (N_8257,N_7796,N_7855);
xor U8258 (N_8258,N_8025,N_7710);
nor U8259 (N_8259,N_7772,N_7592);
or U8260 (N_8260,N_7816,N_8052);
or U8261 (N_8261,N_7912,N_7777);
or U8262 (N_8262,N_8080,N_8200);
nor U8263 (N_8263,N_7630,N_8182);
nand U8264 (N_8264,N_8057,N_8042);
nor U8265 (N_8265,N_8210,N_7746);
nand U8266 (N_8266,N_8249,N_8140);
nand U8267 (N_8267,N_7733,N_8135);
nor U8268 (N_8268,N_8183,N_7515);
nor U8269 (N_8269,N_7940,N_7875);
nand U8270 (N_8270,N_7953,N_7759);
nand U8271 (N_8271,N_8102,N_8227);
nor U8272 (N_8272,N_7619,N_8173);
or U8273 (N_8273,N_7558,N_7654);
nor U8274 (N_8274,N_7503,N_7891);
or U8275 (N_8275,N_7775,N_8056);
nand U8276 (N_8276,N_8141,N_7703);
nand U8277 (N_8277,N_7516,N_8213);
nor U8278 (N_8278,N_7776,N_8201);
and U8279 (N_8279,N_7827,N_7945);
nand U8280 (N_8280,N_7795,N_7878);
nand U8281 (N_8281,N_8167,N_7697);
or U8282 (N_8282,N_7907,N_7844);
or U8283 (N_8283,N_7798,N_8158);
xnor U8284 (N_8284,N_8126,N_7652);
or U8285 (N_8285,N_7958,N_8022);
nor U8286 (N_8286,N_7648,N_8187);
or U8287 (N_8287,N_7994,N_7614);
nand U8288 (N_8288,N_7846,N_7562);
and U8289 (N_8289,N_8136,N_7505);
or U8290 (N_8290,N_7514,N_7821);
nand U8291 (N_8291,N_7814,N_7991);
and U8292 (N_8292,N_7695,N_7799);
or U8293 (N_8293,N_8021,N_8010);
or U8294 (N_8294,N_7681,N_8230);
and U8295 (N_8295,N_7770,N_7598);
nor U8296 (N_8296,N_7883,N_7886);
or U8297 (N_8297,N_7895,N_7944);
nand U8298 (N_8298,N_8092,N_7930);
and U8299 (N_8299,N_8191,N_7576);
xnor U8300 (N_8300,N_7732,N_7610);
nor U8301 (N_8301,N_7773,N_7760);
or U8302 (N_8302,N_7588,N_7726);
nor U8303 (N_8303,N_8111,N_7651);
nand U8304 (N_8304,N_8202,N_7602);
nand U8305 (N_8305,N_7699,N_8225);
and U8306 (N_8306,N_7828,N_8030);
and U8307 (N_8307,N_8186,N_7571);
and U8308 (N_8308,N_7673,N_8081);
nand U8309 (N_8309,N_7584,N_7669);
nor U8310 (N_8310,N_7823,N_7802);
or U8311 (N_8311,N_7641,N_7877);
and U8312 (N_8312,N_7579,N_7764);
and U8313 (N_8313,N_8134,N_8151);
or U8314 (N_8314,N_7500,N_7555);
or U8315 (N_8315,N_7986,N_7911);
nor U8316 (N_8316,N_7859,N_7763);
nor U8317 (N_8317,N_7692,N_7573);
xnor U8318 (N_8318,N_7727,N_8164);
or U8319 (N_8319,N_7964,N_8205);
nand U8320 (N_8320,N_7590,N_8168);
xnor U8321 (N_8321,N_7554,N_7910);
and U8322 (N_8322,N_7946,N_8098);
xor U8323 (N_8323,N_7658,N_7966);
or U8324 (N_8324,N_7624,N_7595);
or U8325 (N_8325,N_8090,N_7841);
nor U8326 (N_8326,N_7633,N_7606);
and U8327 (N_8327,N_8162,N_7631);
xnor U8328 (N_8328,N_8181,N_7525);
or U8329 (N_8329,N_8246,N_8223);
or U8330 (N_8330,N_7801,N_8059);
or U8331 (N_8331,N_7677,N_7626);
nand U8332 (N_8332,N_8019,N_7593);
and U8333 (N_8333,N_8247,N_7700);
nor U8334 (N_8334,N_7863,N_8082);
and U8335 (N_8335,N_7840,N_8094);
or U8336 (N_8336,N_7939,N_8107);
nor U8337 (N_8337,N_8128,N_7596);
and U8338 (N_8338,N_7664,N_7548);
nand U8339 (N_8339,N_7531,N_7847);
nand U8340 (N_8340,N_8076,N_7949);
nor U8341 (N_8341,N_7605,N_7611);
nand U8342 (N_8342,N_8043,N_7933);
xor U8343 (N_8343,N_7993,N_7524);
nand U8344 (N_8344,N_7998,N_8119);
nor U8345 (N_8345,N_7540,N_7979);
or U8346 (N_8346,N_7952,N_7976);
and U8347 (N_8347,N_7919,N_7922);
xnor U8348 (N_8348,N_8089,N_7679);
and U8349 (N_8349,N_8045,N_7999);
xnor U8350 (N_8350,N_7905,N_7898);
and U8351 (N_8351,N_7668,N_7815);
or U8352 (N_8352,N_8160,N_8017);
nor U8353 (N_8353,N_7935,N_8122);
nor U8354 (N_8354,N_7767,N_8003);
and U8355 (N_8355,N_7586,N_7983);
or U8356 (N_8356,N_8127,N_7961);
and U8357 (N_8357,N_8156,N_7774);
and U8358 (N_8358,N_8189,N_8245);
nor U8359 (N_8359,N_8097,N_8023);
nand U8360 (N_8360,N_8207,N_7559);
nand U8361 (N_8361,N_8063,N_7527);
nor U8362 (N_8362,N_8058,N_7532);
or U8363 (N_8363,N_8064,N_8037);
or U8364 (N_8364,N_8006,N_7545);
and U8365 (N_8365,N_7591,N_7781);
nor U8366 (N_8366,N_7535,N_8234);
xnor U8367 (N_8367,N_8159,N_8112);
xor U8368 (N_8368,N_8077,N_7685);
or U8369 (N_8369,N_7716,N_7707);
and U8370 (N_8370,N_8060,N_7825);
nand U8371 (N_8371,N_7659,N_7849);
or U8372 (N_8372,N_7556,N_7587);
nand U8373 (N_8373,N_7861,N_7519);
nor U8374 (N_8374,N_8196,N_8242);
and U8375 (N_8375,N_8055,N_7885);
xnor U8376 (N_8376,N_7601,N_7520);
and U8377 (N_8377,N_8009,N_7561);
nand U8378 (N_8378,N_7742,N_7636);
or U8379 (N_8379,N_7938,N_7536);
nor U8380 (N_8380,N_8114,N_8026);
or U8381 (N_8381,N_7783,N_8216);
nand U8382 (N_8382,N_7529,N_7736);
nor U8383 (N_8383,N_7534,N_7644);
and U8384 (N_8384,N_7580,N_8143);
nand U8385 (N_8385,N_8012,N_8229);
or U8386 (N_8386,N_7780,N_8075);
nor U8387 (N_8387,N_7768,N_7889);
or U8388 (N_8388,N_7622,N_8149);
nor U8389 (N_8389,N_7955,N_8174);
nor U8390 (N_8390,N_7918,N_8120);
nor U8391 (N_8391,N_7927,N_7517);
xor U8392 (N_8392,N_7680,N_7567);
nor U8393 (N_8393,N_7510,N_8088);
or U8394 (N_8394,N_7609,N_8235);
nand U8395 (N_8395,N_8068,N_7565);
and U8396 (N_8396,N_7676,N_7739);
nand U8397 (N_8397,N_8038,N_8222);
or U8398 (N_8398,N_7879,N_8214);
and U8399 (N_8399,N_7936,N_8199);
xnor U8400 (N_8400,N_7671,N_8220);
and U8401 (N_8401,N_7714,N_8138);
nor U8402 (N_8402,N_7807,N_7719);
nand U8403 (N_8403,N_7954,N_7537);
and U8404 (N_8404,N_7741,N_8150);
nor U8405 (N_8405,N_8050,N_7959);
and U8406 (N_8406,N_7523,N_7972);
and U8407 (N_8407,N_7544,N_8031);
and U8408 (N_8408,N_7706,N_8175);
or U8409 (N_8409,N_7574,N_7766);
or U8410 (N_8410,N_7645,N_8071);
and U8411 (N_8411,N_7805,N_8121);
and U8412 (N_8412,N_8095,N_7789);
nor U8413 (N_8413,N_7778,N_7720);
nor U8414 (N_8414,N_7518,N_7755);
nor U8415 (N_8415,N_8035,N_7984);
nor U8416 (N_8416,N_8113,N_8061);
and U8417 (N_8417,N_7583,N_7832);
nor U8418 (N_8418,N_8169,N_8033);
nor U8419 (N_8419,N_8165,N_8016);
and U8420 (N_8420,N_8192,N_8190);
or U8421 (N_8421,N_7876,N_7657);
nand U8422 (N_8422,N_7818,N_7600);
and U8423 (N_8423,N_7747,N_7978);
nor U8424 (N_8424,N_7694,N_7674);
and U8425 (N_8425,N_7608,N_7868);
nand U8426 (N_8426,N_7634,N_7808);
or U8427 (N_8427,N_8116,N_8243);
and U8428 (N_8428,N_7987,N_8139);
nor U8429 (N_8429,N_7552,N_7717);
xnor U8430 (N_8430,N_7512,N_7572);
and U8431 (N_8431,N_8212,N_8203);
or U8432 (N_8432,N_7838,N_7585);
xnor U8433 (N_8433,N_8041,N_7996);
and U8434 (N_8434,N_7678,N_8194);
nor U8435 (N_8435,N_8040,N_7744);
nand U8436 (N_8436,N_8130,N_7923);
nand U8437 (N_8437,N_7752,N_8099);
or U8438 (N_8438,N_7509,N_7803);
or U8439 (N_8439,N_7734,N_7672);
nand U8440 (N_8440,N_7908,N_7790);
or U8441 (N_8441,N_7543,N_8231);
nor U8442 (N_8442,N_7771,N_8087);
and U8443 (N_8443,N_7682,N_7542);
or U8444 (N_8444,N_7743,N_7860);
xor U8445 (N_8445,N_8125,N_7570);
or U8446 (N_8446,N_7950,N_7662);
nor U8447 (N_8447,N_7513,N_7712);
or U8448 (N_8448,N_7862,N_7963);
and U8449 (N_8449,N_8008,N_7691);
or U8450 (N_8450,N_7621,N_7675);
nand U8451 (N_8451,N_7581,N_7728);
or U8452 (N_8452,N_7553,N_7757);
nor U8453 (N_8453,N_8176,N_8148);
nand U8454 (N_8454,N_7575,N_8015);
nor U8455 (N_8455,N_7835,N_8157);
xnor U8456 (N_8456,N_8248,N_7965);
nand U8457 (N_8457,N_8096,N_7792);
and U8458 (N_8458,N_8171,N_7563);
nor U8459 (N_8459,N_8144,N_7639);
nand U8460 (N_8460,N_8154,N_7618);
xor U8461 (N_8461,N_8219,N_7696);
nand U8462 (N_8462,N_7812,N_7826);
nand U8463 (N_8463,N_7722,N_8228);
nand U8464 (N_8464,N_7990,N_7926);
nand U8465 (N_8465,N_7615,N_7962);
or U8466 (N_8466,N_7948,N_7845);
nand U8467 (N_8467,N_7892,N_8027);
and U8468 (N_8468,N_7701,N_8195);
or U8469 (N_8469,N_7568,N_7989);
nor U8470 (N_8470,N_7506,N_7689);
xnor U8471 (N_8471,N_7830,N_7873);
nor U8472 (N_8472,N_8101,N_8067);
nor U8473 (N_8473,N_7937,N_8197);
and U8474 (N_8474,N_7920,N_8044);
or U8475 (N_8475,N_7715,N_7745);
nor U8476 (N_8476,N_8211,N_8240);
xor U8477 (N_8477,N_7934,N_7848);
nand U8478 (N_8478,N_8185,N_7909);
nor U8479 (N_8479,N_8218,N_7882);
nand U8480 (N_8480,N_8123,N_8085);
nand U8481 (N_8481,N_7971,N_7906);
nand U8482 (N_8482,N_7507,N_7723);
nand U8483 (N_8483,N_7667,N_7748);
nand U8484 (N_8484,N_8054,N_8002);
and U8485 (N_8485,N_8103,N_8078);
or U8486 (N_8486,N_7837,N_7929);
or U8487 (N_8487,N_7858,N_7985);
and U8488 (N_8488,N_7737,N_7538);
nand U8489 (N_8489,N_8244,N_7599);
or U8490 (N_8490,N_7521,N_8053);
xor U8491 (N_8491,N_7819,N_7511);
and U8492 (N_8492,N_7903,N_8118);
nand U8493 (N_8493,N_7688,N_8047);
or U8494 (N_8494,N_8237,N_8170);
xnor U8495 (N_8495,N_7617,N_7566);
nand U8496 (N_8496,N_8152,N_8028);
and U8497 (N_8497,N_7791,N_7725);
and U8498 (N_8498,N_7967,N_8048);
nor U8499 (N_8499,N_7684,N_7632);
nand U8500 (N_8500,N_7800,N_7751);
nor U8501 (N_8501,N_7833,N_7502);
xor U8502 (N_8502,N_7541,N_7547);
nor U8503 (N_8503,N_8070,N_7779);
or U8504 (N_8504,N_7637,N_7756);
nor U8505 (N_8505,N_8188,N_8072);
nand U8506 (N_8506,N_8100,N_7897);
or U8507 (N_8507,N_7836,N_7607);
and U8508 (N_8508,N_7915,N_7917);
nand U8509 (N_8509,N_8106,N_7951);
or U8510 (N_8510,N_7942,N_7932);
nor U8511 (N_8511,N_7822,N_7550);
nand U8512 (N_8512,N_7501,N_7888);
nor U8513 (N_8513,N_7749,N_7661);
xnor U8514 (N_8514,N_8206,N_7642);
and U8515 (N_8515,N_8163,N_7627);
and U8516 (N_8516,N_8145,N_7941);
or U8517 (N_8517,N_8013,N_7730);
and U8518 (N_8518,N_8153,N_8109);
and U8519 (N_8519,N_8020,N_8146);
nand U8520 (N_8520,N_7647,N_7890);
nand U8521 (N_8521,N_8131,N_7975);
nor U8522 (N_8522,N_7857,N_7709);
and U8523 (N_8523,N_7980,N_8198);
and U8524 (N_8524,N_7969,N_8036);
and U8525 (N_8525,N_8104,N_7522);
nor U8526 (N_8526,N_7564,N_7569);
nand U8527 (N_8527,N_7539,N_7718);
and U8528 (N_8528,N_7977,N_7867);
nand U8529 (N_8529,N_8224,N_8051);
nor U8530 (N_8530,N_7797,N_8024);
and U8531 (N_8531,N_7761,N_7549);
and U8532 (N_8532,N_8001,N_8193);
xor U8533 (N_8533,N_7850,N_8093);
or U8534 (N_8534,N_8065,N_7809);
nor U8535 (N_8535,N_8034,N_8147);
nor U8536 (N_8536,N_7702,N_7735);
xor U8537 (N_8537,N_8179,N_7902);
and U8538 (N_8538,N_7869,N_7865);
nor U8539 (N_8539,N_7834,N_7872);
or U8540 (N_8540,N_7981,N_7899);
nor U8541 (N_8541,N_7784,N_7504);
nand U8542 (N_8542,N_7731,N_8018);
nor U8543 (N_8543,N_7794,N_7787);
nand U8544 (N_8544,N_8105,N_8032);
nand U8545 (N_8545,N_7650,N_7925);
and U8546 (N_8546,N_7900,N_7653);
nand U8547 (N_8547,N_7704,N_7616);
xor U8548 (N_8548,N_7729,N_7995);
and U8549 (N_8549,N_7638,N_8091);
and U8550 (N_8550,N_7649,N_7643);
nor U8551 (N_8551,N_7880,N_8011);
and U8552 (N_8552,N_8232,N_7557);
nand U8553 (N_8553,N_7901,N_7666);
or U8554 (N_8554,N_7974,N_7612);
nand U8555 (N_8555,N_8086,N_7546);
nor U8556 (N_8556,N_7829,N_8221);
or U8557 (N_8557,N_7721,N_7884);
or U8558 (N_8558,N_7646,N_7788);
and U8559 (N_8559,N_7793,N_7625);
nor U8560 (N_8560,N_8046,N_8217);
or U8561 (N_8561,N_7824,N_7629);
and U8562 (N_8562,N_8108,N_7693);
nand U8563 (N_8563,N_7690,N_7960);
xor U8564 (N_8564,N_7594,N_8177);
nor U8565 (N_8565,N_8137,N_8115);
or U8566 (N_8566,N_8209,N_7804);
or U8567 (N_8567,N_7750,N_7853);
xnor U8568 (N_8568,N_7871,N_7683);
nand U8569 (N_8569,N_7874,N_7852);
or U8570 (N_8570,N_7916,N_8005);
nor U8571 (N_8571,N_7839,N_7724);
nor U8572 (N_8572,N_7656,N_7663);
and U8573 (N_8573,N_7843,N_7758);
and U8574 (N_8574,N_8215,N_7687);
nor U8575 (N_8575,N_7577,N_8226);
xnor U8576 (N_8576,N_7956,N_8049);
or U8577 (N_8577,N_7970,N_7660);
nand U8578 (N_8578,N_7896,N_7782);
nor U8579 (N_8579,N_7603,N_7817);
nor U8580 (N_8580,N_8204,N_7914);
or U8581 (N_8581,N_7708,N_7597);
nor U8582 (N_8582,N_8073,N_7740);
nand U8583 (N_8583,N_7887,N_7620);
nor U8584 (N_8584,N_7813,N_8233);
or U8585 (N_8585,N_7665,N_7870);
nor U8586 (N_8586,N_7508,N_8014);
or U8587 (N_8587,N_8142,N_8208);
nand U8588 (N_8588,N_7528,N_8110);
nor U8589 (N_8589,N_8161,N_7894);
nand U8590 (N_8590,N_7810,N_7866);
and U8591 (N_8591,N_7806,N_7854);
and U8592 (N_8592,N_7769,N_8166);
or U8593 (N_8593,N_8236,N_8238);
xor U8594 (N_8594,N_8062,N_7705);
nor U8595 (N_8595,N_8079,N_7924);
nor U8596 (N_8596,N_7754,N_7698);
xnor U8597 (N_8597,N_7864,N_7765);
and U8598 (N_8598,N_8172,N_8066);
nand U8599 (N_8599,N_8239,N_7711);
or U8600 (N_8600,N_7928,N_8241);
nor U8601 (N_8601,N_8180,N_8155);
and U8602 (N_8602,N_8129,N_7526);
nand U8603 (N_8603,N_7947,N_7820);
nand U8604 (N_8604,N_7785,N_7670);
nor U8605 (N_8605,N_8007,N_7921);
or U8606 (N_8606,N_7931,N_7713);
and U8607 (N_8607,N_8000,N_7842);
xnor U8608 (N_8608,N_7530,N_7551);
or U8609 (N_8609,N_8117,N_7988);
nand U8610 (N_8610,N_8178,N_7982);
nor U8611 (N_8611,N_7628,N_7560);
nor U8612 (N_8612,N_8084,N_7997);
or U8613 (N_8613,N_7762,N_8029);
or U8614 (N_8614,N_7635,N_7957);
or U8615 (N_8615,N_7655,N_7582);
nor U8616 (N_8616,N_7943,N_7786);
or U8617 (N_8617,N_8133,N_7589);
nand U8618 (N_8618,N_7851,N_8124);
or U8619 (N_8619,N_8083,N_7904);
or U8620 (N_8620,N_8184,N_7881);
or U8621 (N_8621,N_7578,N_7913);
and U8622 (N_8622,N_8039,N_8004);
nand U8623 (N_8623,N_7623,N_7856);
or U8624 (N_8624,N_7640,N_7604);
nor U8625 (N_8625,N_7685,N_8029);
and U8626 (N_8626,N_8079,N_7679);
and U8627 (N_8627,N_8211,N_8115);
or U8628 (N_8628,N_7600,N_8041);
and U8629 (N_8629,N_7970,N_7743);
or U8630 (N_8630,N_7559,N_7976);
nor U8631 (N_8631,N_7871,N_7891);
or U8632 (N_8632,N_7556,N_7797);
nor U8633 (N_8633,N_7927,N_7812);
or U8634 (N_8634,N_7878,N_7587);
or U8635 (N_8635,N_7874,N_8163);
nor U8636 (N_8636,N_8082,N_7948);
and U8637 (N_8637,N_8119,N_8157);
nor U8638 (N_8638,N_7946,N_7921);
and U8639 (N_8639,N_8111,N_7811);
nand U8640 (N_8640,N_7946,N_7787);
and U8641 (N_8641,N_8030,N_7614);
nor U8642 (N_8642,N_7926,N_7669);
or U8643 (N_8643,N_8005,N_8119);
nor U8644 (N_8644,N_7719,N_7823);
or U8645 (N_8645,N_8114,N_8007);
nand U8646 (N_8646,N_8063,N_7603);
or U8647 (N_8647,N_8097,N_7799);
or U8648 (N_8648,N_7852,N_8213);
and U8649 (N_8649,N_8021,N_7841);
and U8650 (N_8650,N_7819,N_7841);
and U8651 (N_8651,N_7954,N_7568);
and U8652 (N_8652,N_7681,N_7773);
or U8653 (N_8653,N_7504,N_7745);
nor U8654 (N_8654,N_7626,N_8007);
or U8655 (N_8655,N_8180,N_7699);
and U8656 (N_8656,N_8022,N_7738);
nand U8657 (N_8657,N_7621,N_8220);
nor U8658 (N_8658,N_7690,N_8012);
xor U8659 (N_8659,N_8107,N_7520);
and U8660 (N_8660,N_7688,N_7510);
nor U8661 (N_8661,N_7764,N_7874);
nand U8662 (N_8662,N_7595,N_7955);
nor U8663 (N_8663,N_7903,N_7885);
nor U8664 (N_8664,N_7563,N_7625);
and U8665 (N_8665,N_8229,N_8042);
or U8666 (N_8666,N_7825,N_7659);
nand U8667 (N_8667,N_7571,N_8071);
or U8668 (N_8668,N_7715,N_7875);
and U8669 (N_8669,N_8174,N_7502);
xor U8670 (N_8670,N_7632,N_8173);
xor U8671 (N_8671,N_7901,N_7648);
and U8672 (N_8672,N_8118,N_8214);
nand U8673 (N_8673,N_7514,N_7701);
or U8674 (N_8674,N_7708,N_8215);
nor U8675 (N_8675,N_8080,N_7617);
and U8676 (N_8676,N_8112,N_7630);
and U8677 (N_8677,N_7735,N_7602);
nor U8678 (N_8678,N_8177,N_7539);
xnor U8679 (N_8679,N_8235,N_8150);
or U8680 (N_8680,N_8037,N_8188);
nand U8681 (N_8681,N_8031,N_7510);
nand U8682 (N_8682,N_8157,N_7941);
and U8683 (N_8683,N_7966,N_8068);
nor U8684 (N_8684,N_7810,N_7732);
or U8685 (N_8685,N_7842,N_7596);
nand U8686 (N_8686,N_7702,N_8236);
nor U8687 (N_8687,N_7722,N_7654);
nand U8688 (N_8688,N_7584,N_7995);
nor U8689 (N_8689,N_7833,N_7955);
nand U8690 (N_8690,N_7770,N_7562);
or U8691 (N_8691,N_7572,N_7756);
and U8692 (N_8692,N_8149,N_8216);
nand U8693 (N_8693,N_7891,N_7899);
nand U8694 (N_8694,N_8113,N_8004);
nand U8695 (N_8695,N_7646,N_7744);
and U8696 (N_8696,N_8175,N_8181);
nor U8697 (N_8697,N_7756,N_7919);
and U8698 (N_8698,N_8065,N_7812);
nor U8699 (N_8699,N_7965,N_7936);
nand U8700 (N_8700,N_7524,N_8155);
or U8701 (N_8701,N_7686,N_7706);
and U8702 (N_8702,N_7514,N_8003);
or U8703 (N_8703,N_8232,N_8052);
nand U8704 (N_8704,N_7610,N_8086);
or U8705 (N_8705,N_7674,N_7984);
nand U8706 (N_8706,N_8145,N_7757);
nor U8707 (N_8707,N_7832,N_8124);
or U8708 (N_8708,N_7766,N_8216);
nand U8709 (N_8709,N_7757,N_8170);
and U8710 (N_8710,N_7900,N_7714);
and U8711 (N_8711,N_7679,N_7542);
nand U8712 (N_8712,N_7747,N_7743);
nand U8713 (N_8713,N_7995,N_7577);
or U8714 (N_8714,N_7783,N_7651);
or U8715 (N_8715,N_7852,N_7720);
and U8716 (N_8716,N_7726,N_7751);
or U8717 (N_8717,N_7996,N_7758);
and U8718 (N_8718,N_7610,N_7541);
xor U8719 (N_8719,N_8081,N_7795);
and U8720 (N_8720,N_8116,N_8107);
and U8721 (N_8721,N_7769,N_7864);
and U8722 (N_8722,N_7607,N_7840);
and U8723 (N_8723,N_8158,N_7508);
nand U8724 (N_8724,N_7738,N_8127);
or U8725 (N_8725,N_8018,N_7725);
nor U8726 (N_8726,N_8113,N_7963);
nor U8727 (N_8727,N_7862,N_7607);
nor U8728 (N_8728,N_7623,N_7648);
nand U8729 (N_8729,N_8053,N_7538);
or U8730 (N_8730,N_8137,N_7878);
or U8731 (N_8731,N_8077,N_7837);
or U8732 (N_8732,N_7801,N_7803);
nor U8733 (N_8733,N_7965,N_7586);
nand U8734 (N_8734,N_7961,N_7740);
and U8735 (N_8735,N_7938,N_7530);
or U8736 (N_8736,N_8036,N_7587);
or U8737 (N_8737,N_7901,N_8090);
or U8738 (N_8738,N_7589,N_7790);
or U8739 (N_8739,N_7819,N_8072);
nand U8740 (N_8740,N_8170,N_8055);
nor U8741 (N_8741,N_8082,N_8056);
nor U8742 (N_8742,N_8109,N_7507);
or U8743 (N_8743,N_7698,N_7683);
nor U8744 (N_8744,N_7884,N_7634);
xnor U8745 (N_8745,N_7588,N_7797);
nor U8746 (N_8746,N_7833,N_8194);
and U8747 (N_8747,N_7882,N_7816);
or U8748 (N_8748,N_7596,N_8009);
nand U8749 (N_8749,N_7516,N_7664);
and U8750 (N_8750,N_7649,N_7886);
and U8751 (N_8751,N_8062,N_8034);
nor U8752 (N_8752,N_8007,N_8175);
nor U8753 (N_8753,N_8132,N_7653);
and U8754 (N_8754,N_7639,N_7942);
nand U8755 (N_8755,N_8066,N_8213);
or U8756 (N_8756,N_7713,N_8056);
nor U8757 (N_8757,N_7783,N_8175);
nand U8758 (N_8758,N_7654,N_7643);
and U8759 (N_8759,N_7744,N_7803);
and U8760 (N_8760,N_7877,N_8188);
nor U8761 (N_8761,N_7656,N_7630);
and U8762 (N_8762,N_8172,N_8126);
and U8763 (N_8763,N_7864,N_7799);
and U8764 (N_8764,N_8142,N_7860);
xor U8765 (N_8765,N_8221,N_8045);
and U8766 (N_8766,N_7881,N_7618);
nor U8767 (N_8767,N_7826,N_7707);
nand U8768 (N_8768,N_8008,N_8044);
and U8769 (N_8769,N_7667,N_7655);
or U8770 (N_8770,N_7842,N_7697);
nor U8771 (N_8771,N_7557,N_8059);
nand U8772 (N_8772,N_8012,N_7564);
nand U8773 (N_8773,N_7776,N_8009);
or U8774 (N_8774,N_7785,N_7886);
nand U8775 (N_8775,N_8068,N_8158);
and U8776 (N_8776,N_7530,N_8213);
or U8777 (N_8777,N_7598,N_7612);
and U8778 (N_8778,N_7681,N_8241);
nor U8779 (N_8779,N_8111,N_7927);
and U8780 (N_8780,N_8015,N_7845);
nand U8781 (N_8781,N_7503,N_7518);
nand U8782 (N_8782,N_8092,N_8133);
or U8783 (N_8783,N_7797,N_7533);
xnor U8784 (N_8784,N_7699,N_7904);
nand U8785 (N_8785,N_7658,N_8007);
nor U8786 (N_8786,N_8039,N_7765);
xnor U8787 (N_8787,N_7588,N_7578);
nand U8788 (N_8788,N_7894,N_8092);
and U8789 (N_8789,N_8067,N_7789);
nor U8790 (N_8790,N_7832,N_7548);
xnor U8791 (N_8791,N_8028,N_7984);
xnor U8792 (N_8792,N_7576,N_7596);
nor U8793 (N_8793,N_7818,N_7553);
or U8794 (N_8794,N_7717,N_7757);
nor U8795 (N_8795,N_7717,N_8175);
xor U8796 (N_8796,N_8123,N_7763);
nand U8797 (N_8797,N_7687,N_7704);
and U8798 (N_8798,N_7832,N_8024);
nand U8799 (N_8799,N_8004,N_8211);
and U8800 (N_8800,N_8028,N_8129);
and U8801 (N_8801,N_7724,N_7534);
xor U8802 (N_8802,N_7953,N_7617);
or U8803 (N_8803,N_8002,N_8218);
nand U8804 (N_8804,N_7818,N_7663);
and U8805 (N_8805,N_8116,N_7566);
nand U8806 (N_8806,N_7870,N_8193);
or U8807 (N_8807,N_7804,N_7732);
xor U8808 (N_8808,N_7765,N_8214);
and U8809 (N_8809,N_7859,N_7784);
nand U8810 (N_8810,N_7576,N_7999);
nand U8811 (N_8811,N_8123,N_7628);
nor U8812 (N_8812,N_7732,N_8091);
nand U8813 (N_8813,N_8184,N_7917);
nor U8814 (N_8814,N_7915,N_7675);
nor U8815 (N_8815,N_8073,N_7613);
or U8816 (N_8816,N_7589,N_7884);
xor U8817 (N_8817,N_7684,N_8135);
nor U8818 (N_8818,N_8011,N_8206);
and U8819 (N_8819,N_8143,N_7866);
xor U8820 (N_8820,N_7643,N_7672);
nor U8821 (N_8821,N_7973,N_7515);
nor U8822 (N_8822,N_8131,N_8048);
nand U8823 (N_8823,N_7594,N_8083);
nand U8824 (N_8824,N_7741,N_8222);
nand U8825 (N_8825,N_7853,N_7543);
or U8826 (N_8826,N_7891,N_7629);
nor U8827 (N_8827,N_7601,N_7949);
nor U8828 (N_8828,N_8134,N_7935);
nand U8829 (N_8829,N_7757,N_7827);
xnor U8830 (N_8830,N_7971,N_8068);
and U8831 (N_8831,N_8075,N_7732);
nor U8832 (N_8832,N_7808,N_7748);
and U8833 (N_8833,N_8030,N_7785);
or U8834 (N_8834,N_7614,N_7885);
or U8835 (N_8835,N_8015,N_7520);
nand U8836 (N_8836,N_7869,N_7890);
nor U8837 (N_8837,N_7538,N_7898);
xnor U8838 (N_8838,N_7554,N_7652);
and U8839 (N_8839,N_7520,N_8179);
nor U8840 (N_8840,N_8223,N_7623);
nor U8841 (N_8841,N_7670,N_7775);
or U8842 (N_8842,N_8102,N_7573);
or U8843 (N_8843,N_7869,N_7690);
nor U8844 (N_8844,N_7916,N_8045);
nand U8845 (N_8845,N_7711,N_7528);
and U8846 (N_8846,N_7997,N_7506);
and U8847 (N_8847,N_8134,N_7934);
and U8848 (N_8848,N_8241,N_7694);
nand U8849 (N_8849,N_7956,N_7797);
xor U8850 (N_8850,N_7983,N_8117);
and U8851 (N_8851,N_7507,N_7844);
nor U8852 (N_8852,N_7609,N_8185);
and U8853 (N_8853,N_7838,N_7644);
or U8854 (N_8854,N_7646,N_7732);
or U8855 (N_8855,N_7773,N_7902);
or U8856 (N_8856,N_7780,N_7889);
xor U8857 (N_8857,N_7994,N_7977);
and U8858 (N_8858,N_8064,N_7973);
nand U8859 (N_8859,N_8112,N_8187);
xor U8860 (N_8860,N_7995,N_8123);
xnor U8861 (N_8861,N_7919,N_7765);
nand U8862 (N_8862,N_8168,N_7963);
nor U8863 (N_8863,N_7535,N_7516);
xor U8864 (N_8864,N_7915,N_8021);
nand U8865 (N_8865,N_7876,N_8000);
and U8866 (N_8866,N_7692,N_7602);
nor U8867 (N_8867,N_8147,N_7803);
nor U8868 (N_8868,N_7790,N_7634);
nor U8869 (N_8869,N_7977,N_7639);
or U8870 (N_8870,N_7764,N_8009);
nand U8871 (N_8871,N_7969,N_7924);
and U8872 (N_8872,N_8115,N_8099);
and U8873 (N_8873,N_7846,N_7927);
or U8874 (N_8874,N_7539,N_7744);
nor U8875 (N_8875,N_8157,N_7511);
or U8876 (N_8876,N_7993,N_7515);
and U8877 (N_8877,N_7585,N_7529);
and U8878 (N_8878,N_7595,N_7814);
nand U8879 (N_8879,N_7692,N_7966);
and U8880 (N_8880,N_8171,N_8054);
nand U8881 (N_8881,N_7519,N_7612);
or U8882 (N_8882,N_8114,N_7510);
or U8883 (N_8883,N_8127,N_8047);
nand U8884 (N_8884,N_7928,N_8243);
nor U8885 (N_8885,N_8228,N_7525);
and U8886 (N_8886,N_8078,N_7747);
and U8887 (N_8887,N_8110,N_8126);
nand U8888 (N_8888,N_7808,N_7792);
nor U8889 (N_8889,N_8053,N_8012);
or U8890 (N_8890,N_7532,N_8002);
nand U8891 (N_8891,N_7663,N_8192);
nand U8892 (N_8892,N_7642,N_8059);
nor U8893 (N_8893,N_7931,N_8130);
or U8894 (N_8894,N_7787,N_8128);
nand U8895 (N_8895,N_7629,N_8071);
nand U8896 (N_8896,N_7830,N_8089);
nor U8897 (N_8897,N_8108,N_8009);
or U8898 (N_8898,N_7697,N_8134);
and U8899 (N_8899,N_7775,N_8050);
nand U8900 (N_8900,N_8097,N_7678);
or U8901 (N_8901,N_7720,N_7849);
nand U8902 (N_8902,N_7723,N_7815);
or U8903 (N_8903,N_8107,N_7754);
nand U8904 (N_8904,N_7989,N_8036);
or U8905 (N_8905,N_8135,N_8136);
nor U8906 (N_8906,N_8160,N_7649);
or U8907 (N_8907,N_8194,N_7686);
nor U8908 (N_8908,N_7675,N_7903);
or U8909 (N_8909,N_8155,N_8120);
nand U8910 (N_8910,N_7866,N_8009);
nand U8911 (N_8911,N_7520,N_8137);
nor U8912 (N_8912,N_7531,N_7870);
nand U8913 (N_8913,N_7614,N_8187);
nor U8914 (N_8914,N_7813,N_8175);
or U8915 (N_8915,N_8062,N_7993);
or U8916 (N_8916,N_7730,N_8160);
nand U8917 (N_8917,N_8032,N_7819);
or U8918 (N_8918,N_7648,N_7774);
or U8919 (N_8919,N_7646,N_7927);
nor U8920 (N_8920,N_7942,N_8137);
nand U8921 (N_8921,N_7703,N_7592);
nor U8922 (N_8922,N_7700,N_7514);
nand U8923 (N_8923,N_7825,N_7931);
nor U8924 (N_8924,N_7685,N_7582);
and U8925 (N_8925,N_7905,N_8198);
nand U8926 (N_8926,N_7814,N_7775);
nor U8927 (N_8927,N_7952,N_8042);
and U8928 (N_8928,N_8159,N_7600);
nor U8929 (N_8929,N_8105,N_7795);
and U8930 (N_8930,N_7891,N_7849);
and U8931 (N_8931,N_7873,N_8173);
nor U8932 (N_8932,N_8186,N_7908);
nand U8933 (N_8933,N_7775,N_7649);
or U8934 (N_8934,N_7502,N_7696);
and U8935 (N_8935,N_7586,N_7570);
nand U8936 (N_8936,N_7893,N_7659);
nand U8937 (N_8937,N_7925,N_8030);
and U8938 (N_8938,N_7796,N_8172);
nor U8939 (N_8939,N_7882,N_8194);
nor U8940 (N_8940,N_7662,N_7505);
nand U8941 (N_8941,N_8062,N_7816);
nand U8942 (N_8942,N_8096,N_7698);
nor U8943 (N_8943,N_8075,N_8020);
or U8944 (N_8944,N_7762,N_7526);
and U8945 (N_8945,N_8191,N_7643);
nor U8946 (N_8946,N_7904,N_7917);
nand U8947 (N_8947,N_8087,N_7784);
nand U8948 (N_8948,N_7768,N_7518);
nor U8949 (N_8949,N_7738,N_7912);
nand U8950 (N_8950,N_8239,N_7531);
or U8951 (N_8951,N_7836,N_7691);
nor U8952 (N_8952,N_7791,N_7836);
or U8953 (N_8953,N_7658,N_8217);
nor U8954 (N_8954,N_8138,N_8020);
nand U8955 (N_8955,N_7874,N_7671);
and U8956 (N_8956,N_8137,N_8130);
or U8957 (N_8957,N_7994,N_8070);
nor U8958 (N_8958,N_8114,N_7709);
xnor U8959 (N_8959,N_7577,N_8092);
and U8960 (N_8960,N_7630,N_7703);
nor U8961 (N_8961,N_7689,N_7741);
and U8962 (N_8962,N_7554,N_7580);
and U8963 (N_8963,N_8025,N_7831);
xor U8964 (N_8964,N_7656,N_7892);
nand U8965 (N_8965,N_7533,N_7745);
nand U8966 (N_8966,N_8220,N_7858);
nand U8967 (N_8967,N_7893,N_8061);
nor U8968 (N_8968,N_7585,N_7853);
nor U8969 (N_8969,N_7713,N_7909);
and U8970 (N_8970,N_7959,N_7506);
nand U8971 (N_8971,N_7745,N_7920);
or U8972 (N_8972,N_8101,N_7640);
nand U8973 (N_8973,N_7761,N_8140);
nor U8974 (N_8974,N_7501,N_8134);
or U8975 (N_8975,N_8109,N_8001);
and U8976 (N_8976,N_8020,N_7781);
or U8977 (N_8977,N_8104,N_7756);
nor U8978 (N_8978,N_7724,N_7941);
or U8979 (N_8979,N_7921,N_7829);
and U8980 (N_8980,N_7916,N_7975);
nor U8981 (N_8981,N_7772,N_8205);
nor U8982 (N_8982,N_8094,N_7519);
nand U8983 (N_8983,N_7867,N_7997);
nand U8984 (N_8984,N_7957,N_7670);
nor U8985 (N_8985,N_7784,N_7955);
nor U8986 (N_8986,N_7616,N_8201);
nor U8987 (N_8987,N_7656,N_7661);
or U8988 (N_8988,N_8168,N_8019);
or U8989 (N_8989,N_7652,N_7900);
nor U8990 (N_8990,N_7954,N_8060);
nor U8991 (N_8991,N_7917,N_7857);
or U8992 (N_8992,N_7787,N_8188);
or U8993 (N_8993,N_8231,N_7590);
nand U8994 (N_8994,N_7873,N_7599);
or U8995 (N_8995,N_7599,N_7822);
nand U8996 (N_8996,N_7620,N_7689);
or U8997 (N_8997,N_8209,N_8231);
and U8998 (N_8998,N_8156,N_8026);
nand U8999 (N_8999,N_8163,N_7599);
nand U9000 (N_9000,N_8665,N_8687);
nand U9001 (N_9001,N_8768,N_8622);
nor U9002 (N_9002,N_8600,N_8696);
and U9003 (N_9003,N_8461,N_8787);
nand U9004 (N_9004,N_8816,N_8976);
or U9005 (N_9005,N_8440,N_8486);
nand U9006 (N_9006,N_8459,N_8915);
and U9007 (N_9007,N_8711,N_8849);
or U9008 (N_9008,N_8760,N_8263);
xnor U9009 (N_9009,N_8605,N_8356);
or U9010 (N_9010,N_8380,N_8564);
nor U9011 (N_9011,N_8551,N_8612);
nand U9012 (N_9012,N_8691,N_8791);
or U9013 (N_9013,N_8530,N_8950);
nor U9014 (N_9014,N_8286,N_8826);
and U9015 (N_9015,N_8875,N_8435);
or U9016 (N_9016,N_8429,N_8424);
nand U9017 (N_9017,N_8666,N_8702);
nand U9018 (N_9018,N_8788,N_8761);
and U9019 (N_9019,N_8673,N_8796);
xor U9020 (N_9020,N_8689,N_8954);
and U9021 (N_9021,N_8303,N_8872);
or U9022 (N_9022,N_8784,N_8740);
nand U9023 (N_9023,N_8864,N_8458);
nand U9024 (N_9024,N_8621,N_8928);
nor U9025 (N_9025,N_8755,N_8643);
nor U9026 (N_9026,N_8683,N_8619);
and U9027 (N_9027,N_8722,N_8443);
nand U9028 (N_9028,N_8721,N_8972);
nor U9029 (N_9029,N_8542,N_8822);
nand U9030 (N_9030,N_8569,N_8865);
nand U9031 (N_9031,N_8715,N_8771);
or U9032 (N_9032,N_8631,N_8640);
and U9033 (N_9033,N_8739,N_8521);
nand U9034 (N_9034,N_8331,N_8975);
and U9035 (N_9035,N_8897,N_8328);
xor U9036 (N_9036,N_8795,N_8828);
nand U9037 (N_9037,N_8686,N_8746);
xor U9038 (N_9038,N_8276,N_8322);
xor U9039 (N_9039,N_8381,N_8388);
or U9040 (N_9040,N_8995,N_8676);
nor U9041 (N_9041,N_8283,N_8310);
nand U9042 (N_9042,N_8448,N_8273);
xnor U9043 (N_9043,N_8939,N_8730);
xor U9044 (N_9044,N_8814,N_8378);
and U9045 (N_9045,N_8359,N_8329);
nor U9046 (N_9046,N_8653,N_8978);
nor U9047 (N_9047,N_8602,N_8894);
or U9048 (N_9048,N_8874,N_8471);
nand U9049 (N_9049,N_8667,N_8473);
nor U9050 (N_9050,N_8425,N_8825);
and U9051 (N_9051,N_8457,N_8520);
or U9052 (N_9052,N_8367,N_8346);
or U9053 (N_9053,N_8983,N_8743);
or U9054 (N_9054,N_8922,N_8365);
nand U9055 (N_9055,N_8581,N_8349);
or U9056 (N_9056,N_8762,N_8731);
xnor U9057 (N_9057,N_8835,N_8748);
or U9058 (N_9058,N_8566,N_8971);
nand U9059 (N_9059,N_8422,N_8499);
and U9060 (N_9060,N_8675,N_8908);
or U9061 (N_9061,N_8452,N_8268);
or U9062 (N_9062,N_8627,N_8963);
xnor U9063 (N_9063,N_8688,N_8280);
and U9064 (N_9064,N_8586,N_8684);
and U9065 (N_9065,N_8753,N_8384);
nand U9066 (N_9066,N_8831,N_8759);
nor U9067 (N_9067,N_8379,N_8668);
or U9068 (N_9068,N_8254,N_8638);
nor U9069 (N_9069,N_8817,N_8271);
and U9070 (N_9070,N_8538,N_8964);
nand U9071 (N_9071,N_8999,N_8574);
nand U9072 (N_9072,N_8652,N_8832);
nand U9073 (N_9073,N_8301,N_8726);
or U9074 (N_9074,N_8355,N_8576);
and U9075 (N_9075,N_8636,N_8981);
and U9076 (N_9076,N_8483,N_8557);
nor U9077 (N_9077,N_8855,N_8515);
nor U9078 (N_9078,N_8315,N_8871);
nor U9079 (N_9079,N_8464,N_8754);
and U9080 (N_9080,N_8590,N_8779);
xor U9081 (N_9081,N_8386,N_8518);
and U9082 (N_9082,N_8769,N_8930);
and U9083 (N_9083,N_8973,N_8392);
and U9084 (N_9084,N_8757,N_8660);
nor U9085 (N_9085,N_8509,N_8906);
nand U9086 (N_9086,N_8377,N_8732);
or U9087 (N_9087,N_8742,N_8827);
and U9088 (N_9088,N_8823,N_8998);
nor U9089 (N_9089,N_8878,N_8713);
xnor U9090 (N_9090,N_8617,N_8848);
xor U9091 (N_9091,N_8733,N_8709);
or U9092 (N_9092,N_8965,N_8588);
nor U9093 (N_9093,N_8707,N_8592);
nor U9094 (N_9094,N_8727,N_8843);
nand U9095 (N_9095,N_8750,N_8423);
nand U9096 (N_9096,N_8396,N_8919);
nand U9097 (N_9097,N_8401,N_8413);
xor U9098 (N_9098,N_8993,N_8992);
and U9099 (N_9099,N_8775,N_8411);
nand U9100 (N_9100,N_8360,N_8312);
or U9101 (N_9101,N_8320,N_8647);
and U9102 (N_9102,N_8902,N_8867);
and U9103 (N_9103,N_8970,N_8945);
nor U9104 (N_9104,N_8598,N_8275);
and U9105 (N_9105,N_8336,N_8904);
nand U9106 (N_9106,N_8737,N_8561);
or U9107 (N_9107,N_8299,N_8445);
nand U9108 (N_9108,N_8968,N_8745);
and U9109 (N_9109,N_8559,N_8671);
and U9110 (N_9110,N_8670,N_8723);
and U9111 (N_9111,N_8255,N_8880);
or U9112 (N_9112,N_8813,N_8535);
nand U9113 (N_9113,N_8962,N_8808);
nand U9114 (N_9114,N_8747,N_8434);
or U9115 (N_9115,N_8293,N_8372);
nand U9116 (N_9116,N_8390,N_8446);
nor U9117 (N_9117,N_8261,N_8785);
and U9118 (N_9118,N_8318,N_8585);
nand U9119 (N_9119,N_8541,N_8794);
nand U9120 (N_9120,N_8432,N_8931);
nor U9121 (N_9121,N_8869,N_8568);
nor U9122 (N_9122,N_8385,N_8948);
and U9123 (N_9123,N_8735,N_8571);
or U9124 (N_9124,N_8302,N_8252);
nand U9125 (N_9125,N_8540,N_8756);
or U9126 (N_9126,N_8637,N_8433);
xnor U9127 (N_9127,N_8916,N_8801);
and U9128 (N_9128,N_8833,N_8421);
and U9129 (N_9129,N_8606,N_8265);
and U9130 (N_9130,N_8701,N_8489);
nor U9131 (N_9131,N_8654,N_8497);
xnor U9132 (N_9132,N_8669,N_8951);
or U9133 (N_9133,N_8543,N_8342);
or U9134 (N_9134,N_8466,N_8933);
xor U9135 (N_9135,N_8887,N_8890);
and U9136 (N_9136,N_8475,N_8719);
nand U9137 (N_9137,N_8967,N_8615);
nor U9138 (N_9138,N_8498,N_8526);
xor U9139 (N_9139,N_8623,N_8339);
and U9140 (N_9140,N_8921,N_8681);
nand U9141 (N_9141,N_8815,N_8343);
nor U9142 (N_9142,N_8389,N_8692);
nor U9143 (N_9143,N_8896,N_8929);
xnor U9144 (N_9144,N_8257,N_8484);
or U9145 (N_9145,N_8527,N_8752);
nor U9146 (N_9146,N_8524,N_8829);
nor U9147 (N_9147,N_8758,N_8682);
or U9148 (N_9148,N_8593,N_8469);
or U9149 (N_9149,N_8853,N_8382);
nor U9150 (N_9150,N_8279,N_8420);
nor U9151 (N_9151,N_8662,N_8493);
nor U9152 (N_9152,N_8934,N_8258);
nor U9153 (N_9153,N_8391,N_8632);
nor U9154 (N_9154,N_8729,N_8845);
and U9155 (N_9155,N_8861,N_8531);
or U9156 (N_9156,N_8313,N_8259);
nand U9157 (N_9157,N_8468,N_8399);
or U9158 (N_9158,N_8834,N_8905);
and U9159 (N_9159,N_8725,N_8626);
nand U9160 (N_9160,N_8441,N_8810);
nand U9161 (N_9161,N_8304,N_8899);
or U9162 (N_9162,N_8393,N_8327);
nor U9163 (N_9163,N_8503,N_8570);
nor U9164 (N_9164,N_8495,N_8272);
nor U9165 (N_9165,N_8514,N_8348);
or U9166 (N_9166,N_8376,N_8639);
nor U9167 (N_9167,N_8923,N_8982);
and U9168 (N_9168,N_8886,N_8837);
nor U9169 (N_9169,N_8749,N_8482);
or U9170 (N_9170,N_8262,N_8937);
nand U9171 (N_9171,N_8251,N_8942);
nor U9172 (N_9172,N_8935,N_8918);
nand U9173 (N_9173,N_8604,N_8809);
xor U9174 (N_9174,N_8596,N_8405);
and U9175 (N_9175,N_8644,N_8984);
nor U9176 (N_9176,N_8465,N_8502);
nand U9177 (N_9177,N_8901,N_8717);
nor U9178 (N_9178,N_8319,N_8920);
nand U9179 (N_9179,N_8578,N_8690);
xor U9180 (N_9180,N_8885,N_8513);
nor U9181 (N_9181,N_8591,N_8764);
nand U9182 (N_9182,N_8549,N_8851);
and U9183 (N_9183,N_8672,N_8558);
and U9184 (N_9184,N_8341,N_8633);
or U9185 (N_9185,N_8804,N_8987);
nor U9186 (N_9186,N_8295,N_8517);
xnor U9187 (N_9187,N_8625,N_8510);
nor U9188 (N_9188,N_8364,N_8988);
or U9189 (N_9189,N_8986,N_8294);
nor U9190 (N_9190,N_8895,N_8353);
xor U9191 (N_9191,N_8693,N_8567);
or U9192 (N_9192,N_8783,N_8694);
or U9193 (N_9193,N_8577,N_8716);
or U9194 (N_9194,N_8680,N_8789);
and U9195 (N_9195,N_8395,N_8264);
and U9196 (N_9196,N_8402,N_8373);
nand U9197 (N_9197,N_8888,N_8534);
and U9198 (N_9198,N_8774,N_8846);
nand U9199 (N_9199,N_8989,N_8278);
nand U9200 (N_9200,N_8481,N_8253);
nand U9201 (N_9201,N_8428,N_8351);
nand U9202 (N_9202,N_8354,N_8324);
nand U9203 (N_9203,N_8778,N_8338);
nor U9204 (N_9204,N_8790,N_8357);
or U9205 (N_9205,N_8881,N_8679);
nand U9206 (N_9206,N_8601,N_8607);
and U9207 (N_9207,N_8734,N_8439);
xnor U9208 (N_9208,N_8418,N_8546);
xor U9209 (N_9209,N_8620,N_8494);
nor U9210 (N_9210,N_8800,N_8641);
or U9211 (N_9211,N_8649,N_8474);
nand U9212 (N_9212,N_8798,N_8580);
nor U9213 (N_9213,N_8563,N_8587);
nand U9214 (N_9214,N_8917,N_8720);
and U9215 (N_9215,N_8932,N_8589);
and U9216 (N_9216,N_8956,N_8250);
nand U9217 (N_9217,N_8595,N_8335);
nand U9218 (N_9218,N_8565,N_8609);
nand U9219 (N_9219,N_8806,N_8270);
xnor U9220 (N_9220,N_8485,N_8281);
or U9221 (N_9221,N_8957,N_8496);
nor U9222 (N_9222,N_8488,N_8553);
or U9223 (N_9223,N_8959,N_8859);
or U9224 (N_9224,N_8907,N_8480);
nand U9225 (N_9225,N_8579,N_8997);
and U9226 (N_9226,N_8462,N_8751);
nand U9227 (N_9227,N_8892,N_8700);
nor U9228 (N_9228,N_8802,N_8290);
nand U9229 (N_9229,N_8856,N_8415);
or U9230 (N_9230,N_8560,N_8333);
xor U9231 (N_9231,N_8269,N_8436);
and U9232 (N_9232,N_8614,N_8642);
nor U9233 (N_9233,N_8736,N_8765);
or U9234 (N_9234,N_8599,N_8799);
nor U9235 (N_9235,N_8476,N_8697);
nor U9236 (N_9236,N_8447,N_8508);
and U9237 (N_9237,N_8532,N_8528);
and U9238 (N_9238,N_8285,N_8877);
and U9239 (N_9239,N_8613,N_8979);
nand U9240 (N_9240,N_8410,N_8961);
and U9241 (N_9241,N_8852,N_8883);
nand U9242 (N_9242,N_8334,N_8903);
and U9243 (N_9243,N_8345,N_8925);
nor U9244 (N_9244,N_8635,N_8347);
or U9245 (N_9245,N_8426,N_8974);
nand U9246 (N_9246,N_8891,N_8451);
nand U9247 (N_9247,N_8479,N_8504);
and U9248 (N_9248,N_8830,N_8298);
nand U9249 (N_9249,N_8512,N_8330);
nand U9250 (N_9250,N_8317,N_8844);
nor U9251 (N_9251,N_8927,N_8572);
nor U9252 (N_9252,N_8400,N_8501);
nor U9253 (N_9253,N_8430,N_8936);
and U9254 (N_9254,N_8416,N_8898);
or U9255 (N_9255,N_8966,N_8492);
or U9256 (N_9256,N_8664,N_8548);
nand U9257 (N_9257,N_8912,N_8383);
xnor U9258 (N_9258,N_8550,N_8363);
nor U9259 (N_9259,N_8511,N_8792);
nand U9260 (N_9260,N_8340,N_8407);
nand U9261 (N_9261,N_8884,N_8659);
or U9262 (N_9262,N_8704,N_8763);
nand U9263 (N_9263,N_8952,N_8554);
nor U9264 (N_9264,N_8944,N_8332);
or U9265 (N_9265,N_8807,N_8374);
and U9266 (N_9266,N_8417,N_8767);
and U9267 (N_9267,N_8695,N_8926);
nor U9268 (N_9268,N_8824,N_8487);
or U9269 (N_9269,N_8337,N_8685);
nor U9270 (N_9270,N_8724,N_8953);
nor U9271 (N_9271,N_8544,N_8977);
or U9272 (N_9272,N_8584,N_8710);
nor U9273 (N_9273,N_8900,N_8868);
xor U9274 (N_9274,N_8780,N_8708);
nand U9275 (N_9275,N_8914,N_8398);
or U9276 (N_9276,N_8876,N_8292);
and U9277 (N_9277,N_8661,N_8362);
and U9278 (N_9278,N_8366,N_8409);
or U9279 (N_9279,N_8924,N_8256);
and U9280 (N_9280,N_8525,N_8841);
xnor U9281 (N_9281,N_8387,N_8350);
or U9282 (N_9282,N_8323,N_8656);
xnor U9283 (N_9283,N_8836,N_8523);
nor U9284 (N_9284,N_8994,N_8996);
nor U9285 (N_9285,N_8533,N_8478);
nand U9286 (N_9286,N_8412,N_8985);
or U9287 (N_9287,N_8805,N_8352);
and U9288 (N_9288,N_8857,N_8536);
and U9289 (N_9289,N_8913,N_8819);
nor U9290 (N_9290,N_8506,N_8776);
or U9291 (N_9291,N_8949,N_8547);
nor U9292 (N_9292,N_8960,N_8705);
xor U9293 (N_9293,N_8943,N_8529);
or U9294 (N_9294,N_8616,N_8624);
and U9295 (N_9295,N_8594,N_8990);
xor U9296 (N_9296,N_8490,N_8545);
xor U9297 (N_9297,N_8893,N_8555);
nor U9298 (N_9298,N_8408,N_8296);
nand U9299 (N_9299,N_8860,N_8838);
nand U9300 (N_9300,N_8404,N_8882);
nor U9301 (N_9301,N_8463,N_8406);
nor U9302 (N_9302,N_8854,N_8611);
nor U9303 (N_9303,N_8911,N_8870);
and U9304 (N_9304,N_8358,N_8454);
or U9305 (N_9305,N_8797,N_8738);
and U9306 (N_9306,N_8307,N_8812);
nand U9307 (N_9307,N_8698,N_8840);
xnor U9308 (N_9308,N_8842,N_8274);
nor U9309 (N_9309,N_8821,N_8427);
or U9310 (N_9310,N_8397,N_8282);
xnor U9311 (N_9311,N_8291,N_8326);
xor U9312 (N_9312,N_8862,N_8793);
and U9313 (N_9313,N_8267,N_8909);
or U9314 (N_9314,N_8403,N_8414);
nand U9315 (N_9315,N_8575,N_8657);
nand U9316 (N_9316,N_8958,N_8314);
nand U9317 (N_9317,N_8618,N_8368);
and U9318 (N_9318,N_8453,N_8678);
and U9319 (N_9319,N_8782,N_8266);
nand U9320 (N_9320,N_8450,N_8889);
or U9321 (N_9321,N_8718,N_8308);
nand U9322 (N_9322,N_8562,N_8629);
and U9323 (N_9323,N_8477,N_8449);
nand U9324 (N_9324,N_8500,N_8820);
nand U9325 (N_9325,N_8773,N_8300);
or U9326 (N_9326,N_8552,N_8277);
or U9327 (N_9327,N_8610,N_8516);
and U9328 (N_9328,N_8699,N_8309);
or U9329 (N_9329,N_8786,N_8288);
nand U9330 (N_9330,N_8940,N_8879);
or U9331 (N_9331,N_8369,N_8645);
nor U9332 (N_9332,N_8603,N_8941);
and U9333 (N_9333,N_8646,N_8634);
nor U9334 (N_9334,N_8573,N_8938);
nand U9335 (N_9335,N_8284,N_8437);
nand U9336 (N_9336,N_8651,N_8419);
xor U9337 (N_9337,N_8655,N_8847);
and U9338 (N_9338,N_8955,N_8522);
nor U9339 (N_9339,N_8582,N_8777);
nor U9340 (N_9340,N_8781,N_8537);
or U9341 (N_9341,N_8714,N_8811);
nand U9342 (N_9342,N_8839,N_8728);
nand U9343 (N_9343,N_8287,N_8766);
or U9344 (N_9344,N_8969,N_8703);
nor U9345 (N_9345,N_8630,N_8431);
nor U9346 (N_9346,N_8910,N_8344);
and U9347 (N_9347,N_8260,N_8456);
or U9348 (N_9348,N_8650,N_8306);
nor U9349 (N_9349,N_8305,N_8394);
or U9350 (N_9350,N_8628,N_8370);
xnor U9351 (N_9351,N_8706,N_8491);
or U9352 (N_9352,N_8505,N_8311);
nand U9353 (N_9353,N_8507,N_8980);
or U9354 (N_9354,N_8297,N_8556);
and U9355 (N_9355,N_8858,N_8539);
and U9356 (N_9356,N_8375,N_8442);
or U9357 (N_9357,N_8361,N_8316);
and U9358 (N_9358,N_8519,N_8470);
or U9359 (N_9359,N_8455,N_8677);
nand U9360 (N_9360,N_8818,N_8873);
or U9361 (N_9361,N_8946,N_8289);
nand U9362 (N_9362,N_8712,N_8850);
or U9363 (N_9363,N_8770,N_8371);
xnor U9364 (N_9364,N_8444,N_8597);
nand U9365 (N_9365,N_8472,N_8866);
xnor U9366 (N_9366,N_8991,N_8325);
and U9367 (N_9367,N_8663,N_8803);
nand U9368 (N_9368,N_8321,N_8863);
or U9369 (N_9369,N_8741,N_8658);
and U9370 (N_9370,N_8772,N_8438);
nand U9371 (N_9371,N_8467,N_8744);
and U9372 (N_9372,N_8648,N_8674);
nor U9373 (N_9373,N_8608,N_8460);
and U9374 (N_9374,N_8583,N_8947);
nor U9375 (N_9375,N_8427,N_8360);
nor U9376 (N_9376,N_8414,N_8280);
or U9377 (N_9377,N_8427,N_8523);
nor U9378 (N_9378,N_8504,N_8804);
nand U9379 (N_9379,N_8735,N_8298);
or U9380 (N_9380,N_8832,N_8667);
xnor U9381 (N_9381,N_8625,N_8691);
nand U9382 (N_9382,N_8836,N_8573);
nor U9383 (N_9383,N_8327,N_8492);
and U9384 (N_9384,N_8516,N_8343);
and U9385 (N_9385,N_8330,N_8924);
and U9386 (N_9386,N_8700,N_8592);
nor U9387 (N_9387,N_8934,N_8621);
or U9388 (N_9388,N_8604,N_8327);
nand U9389 (N_9389,N_8377,N_8642);
nand U9390 (N_9390,N_8509,N_8993);
and U9391 (N_9391,N_8853,N_8772);
nand U9392 (N_9392,N_8757,N_8429);
nor U9393 (N_9393,N_8630,N_8339);
nand U9394 (N_9394,N_8863,N_8532);
or U9395 (N_9395,N_8938,N_8879);
or U9396 (N_9396,N_8801,N_8881);
xor U9397 (N_9397,N_8695,N_8479);
xnor U9398 (N_9398,N_8638,N_8463);
and U9399 (N_9399,N_8891,N_8740);
nor U9400 (N_9400,N_8953,N_8902);
nand U9401 (N_9401,N_8326,N_8599);
and U9402 (N_9402,N_8571,N_8558);
nor U9403 (N_9403,N_8433,N_8865);
or U9404 (N_9404,N_8548,N_8291);
nand U9405 (N_9405,N_8967,N_8844);
xnor U9406 (N_9406,N_8494,N_8913);
or U9407 (N_9407,N_8686,N_8472);
and U9408 (N_9408,N_8293,N_8479);
or U9409 (N_9409,N_8694,N_8949);
xnor U9410 (N_9410,N_8915,N_8394);
or U9411 (N_9411,N_8255,N_8307);
and U9412 (N_9412,N_8854,N_8304);
nand U9413 (N_9413,N_8316,N_8687);
nand U9414 (N_9414,N_8629,N_8860);
and U9415 (N_9415,N_8968,N_8695);
or U9416 (N_9416,N_8336,N_8602);
nand U9417 (N_9417,N_8381,N_8822);
nor U9418 (N_9418,N_8446,N_8874);
or U9419 (N_9419,N_8571,N_8827);
nor U9420 (N_9420,N_8909,N_8924);
xnor U9421 (N_9421,N_8273,N_8616);
or U9422 (N_9422,N_8263,N_8875);
nand U9423 (N_9423,N_8418,N_8703);
xor U9424 (N_9424,N_8520,N_8836);
nand U9425 (N_9425,N_8327,N_8894);
nand U9426 (N_9426,N_8296,N_8984);
nor U9427 (N_9427,N_8303,N_8511);
and U9428 (N_9428,N_8905,N_8378);
nor U9429 (N_9429,N_8479,N_8812);
nand U9430 (N_9430,N_8689,N_8570);
nand U9431 (N_9431,N_8443,N_8731);
nor U9432 (N_9432,N_8467,N_8377);
xnor U9433 (N_9433,N_8792,N_8503);
nor U9434 (N_9434,N_8872,N_8725);
nor U9435 (N_9435,N_8902,N_8819);
xor U9436 (N_9436,N_8655,N_8395);
nor U9437 (N_9437,N_8724,N_8627);
and U9438 (N_9438,N_8339,N_8695);
and U9439 (N_9439,N_8451,N_8960);
nand U9440 (N_9440,N_8828,N_8979);
nor U9441 (N_9441,N_8469,N_8791);
xnor U9442 (N_9442,N_8436,N_8250);
or U9443 (N_9443,N_8278,N_8612);
or U9444 (N_9444,N_8542,N_8278);
nand U9445 (N_9445,N_8748,N_8342);
nor U9446 (N_9446,N_8374,N_8265);
nand U9447 (N_9447,N_8651,N_8805);
and U9448 (N_9448,N_8458,N_8712);
nand U9449 (N_9449,N_8537,N_8963);
or U9450 (N_9450,N_8940,N_8536);
or U9451 (N_9451,N_8896,N_8788);
nor U9452 (N_9452,N_8933,N_8732);
nor U9453 (N_9453,N_8723,N_8293);
or U9454 (N_9454,N_8809,N_8497);
and U9455 (N_9455,N_8268,N_8532);
nor U9456 (N_9456,N_8447,N_8363);
and U9457 (N_9457,N_8805,N_8452);
and U9458 (N_9458,N_8990,N_8267);
and U9459 (N_9459,N_8406,N_8319);
or U9460 (N_9460,N_8466,N_8563);
nor U9461 (N_9461,N_8912,N_8789);
nor U9462 (N_9462,N_8300,N_8951);
and U9463 (N_9463,N_8741,N_8591);
and U9464 (N_9464,N_8881,N_8962);
xor U9465 (N_9465,N_8480,N_8537);
nand U9466 (N_9466,N_8976,N_8610);
nor U9467 (N_9467,N_8574,N_8791);
and U9468 (N_9468,N_8773,N_8605);
and U9469 (N_9469,N_8374,N_8700);
nor U9470 (N_9470,N_8297,N_8969);
xor U9471 (N_9471,N_8437,N_8422);
or U9472 (N_9472,N_8673,N_8584);
nand U9473 (N_9473,N_8398,N_8289);
or U9474 (N_9474,N_8267,N_8612);
and U9475 (N_9475,N_8780,N_8973);
nor U9476 (N_9476,N_8779,N_8508);
nand U9477 (N_9477,N_8507,N_8359);
nand U9478 (N_9478,N_8481,N_8649);
and U9479 (N_9479,N_8592,N_8422);
nor U9480 (N_9480,N_8430,N_8292);
nand U9481 (N_9481,N_8733,N_8354);
or U9482 (N_9482,N_8755,N_8349);
xor U9483 (N_9483,N_8250,N_8696);
nor U9484 (N_9484,N_8661,N_8983);
or U9485 (N_9485,N_8585,N_8942);
and U9486 (N_9486,N_8696,N_8907);
and U9487 (N_9487,N_8598,N_8907);
xnor U9488 (N_9488,N_8283,N_8331);
nor U9489 (N_9489,N_8859,N_8792);
or U9490 (N_9490,N_8960,N_8980);
xor U9491 (N_9491,N_8534,N_8337);
nand U9492 (N_9492,N_8326,N_8383);
nand U9493 (N_9493,N_8800,N_8779);
and U9494 (N_9494,N_8485,N_8260);
nand U9495 (N_9495,N_8472,N_8282);
nor U9496 (N_9496,N_8587,N_8750);
nand U9497 (N_9497,N_8979,N_8409);
xnor U9498 (N_9498,N_8934,N_8854);
and U9499 (N_9499,N_8691,N_8391);
nand U9500 (N_9500,N_8832,N_8671);
or U9501 (N_9501,N_8653,N_8588);
nand U9502 (N_9502,N_8891,N_8851);
or U9503 (N_9503,N_8375,N_8948);
nor U9504 (N_9504,N_8739,N_8917);
or U9505 (N_9505,N_8738,N_8886);
xnor U9506 (N_9506,N_8671,N_8492);
nor U9507 (N_9507,N_8741,N_8523);
nand U9508 (N_9508,N_8839,N_8844);
nor U9509 (N_9509,N_8779,N_8541);
and U9510 (N_9510,N_8541,N_8781);
or U9511 (N_9511,N_8504,N_8513);
or U9512 (N_9512,N_8591,N_8606);
and U9513 (N_9513,N_8830,N_8463);
nand U9514 (N_9514,N_8793,N_8613);
or U9515 (N_9515,N_8716,N_8766);
xor U9516 (N_9516,N_8287,N_8325);
nor U9517 (N_9517,N_8654,N_8759);
nand U9518 (N_9518,N_8812,N_8518);
or U9519 (N_9519,N_8605,N_8626);
nor U9520 (N_9520,N_8261,N_8431);
or U9521 (N_9521,N_8920,N_8772);
and U9522 (N_9522,N_8323,N_8794);
or U9523 (N_9523,N_8399,N_8758);
and U9524 (N_9524,N_8901,N_8614);
nand U9525 (N_9525,N_8891,N_8379);
nand U9526 (N_9526,N_8667,N_8774);
nor U9527 (N_9527,N_8425,N_8314);
xor U9528 (N_9528,N_8811,N_8683);
and U9529 (N_9529,N_8923,N_8827);
xor U9530 (N_9530,N_8467,N_8461);
and U9531 (N_9531,N_8730,N_8396);
or U9532 (N_9532,N_8752,N_8265);
nand U9533 (N_9533,N_8856,N_8387);
or U9534 (N_9534,N_8663,N_8485);
nor U9535 (N_9535,N_8615,N_8873);
nor U9536 (N_9536,N_8376,N_8989);
nor U9537 (N_9537,N_8823,N_8435);
nand U9538 (N_9538,N_8501,N_8849);
nand U9539 (N_9539,N_8335,N_8532);
nor U9540 (N_9540,N_8950,N_8536);
and U9541 (N_9541,N_8405,N_8717);
and U9542 (N_9542,N_8862,N_8953);
nand U9543 (N_9543,N_8983,N_8579);
and U9544 (N_9544,N_8358,N_8918);
nand U9545 (N_9545,N_8415,N_8431);
or U9546 (N_9546,N_8888,N_8920);
nor U9547 (N_9547,N_8975,N_8933);
nand U9548 (N_9548,N_8820,N_8942);
nand U9549 (N_9549,N_8742,N_8431);
or U9550 (N_9550,N_8714,N_8935);
and U9551 (N_9551,N_8291,N_8559);
and U9552 (N_9552,N_8582,N_8933);
and U9553 (N_9553,N_8307,N_8965);
and U9554 (N_9554,N_8989,N_8847);
and U9555 (N_9555,N_8759,N_8933);
nor U9556 (N_9556,N_8871,N_8642);
nor U9557 (N_9557,N_8801,N_8729);
nand U9558 (N_9558,N_8914,N_8747);
or U9559 (N_9559,N_8828,N_8539);
nand U9560 (N_9560,N_8458,N_8443);
and U9561 (N_9561,N_8269,N_8764);
or U9562 (N_9562,N_8292,N_8883);
xor U9563 (N_9563,N_8481,N_8963);
and U9564 (N_9564,N_8889,N_8693);
and U9565 (N_9565,N_8380,N_8833);
and U9566 (N_9566,N_8859,N_8498);
xnor U9567 (N_9567,N_8348,N_8550);
and U9568 (N_9568,N_8893,N_8877);
nand U9569 (N_9569,N_8700,N_8915);
and U9570 (N_9570,N_8913,N_8680);
and U9571 (N_9571,N_8626,N_8364);
or U9572 (N_9572,N_8975,N_8864);
or U9573 (N_9573,N_8600,N_8415);
xor U9574 (N_9574,N_8432,N_8250);
nand U9575 (N_9575,N_8959,N_8427);
nor U9576 (N_9576,N_8763,N_8746);
and U9577 (N_9577,N_8872,N_8320);
and U9578 (N_9578,N_8972,N_8617);
or U9579 (N_9579,N_8660,N_8971);
and U9580 (N_9580,N_8323,N_8552);
and U9581 (N_9581,N_8998,N_8989);
nand U9582 (N_9582,N_8484,N_8425);
or U9583 (N_9583,N_8914,N_8994);
and U9584 (N_9584,N_8726,N_8511);
nand U9585 (N_9585,N_8444,N_8779);
and U9586 (N_9586,N_8860,N_8522);
or U9587 (N_9587,N_8744,N_8853);
and U9588 (N_9588,N_8572,N_8531);
nand U9589 (N_9589,N_8969,N_8746);
nor U9590 (N_9590,N_8284,N_8413);
nor U9591 (N_9591,N_8486,N_8813);
or U9592 (N_9592,N_8741,N_8284);
nand U9593 (N_9593,N_8564,N_8546);
nand U9594 (N_9594,N_8399,N_8972);
nor U9595 (N_9595,N_8614,N_8667);
or U9596 (N_9596,N_8636,N_8879);
xor U9597 (N_9597,N_8303,N_8980);
or U9598 (N_9598,N_8750,N_8645);
and U9599 (N_9599,N_8963,N_8938);
nor U9600 (N_9600,N_8890,N_8598);
nand U9601 (N_9601,N_8280,N_8270);
and U9602 (N_9602,N_8572,N_8767);
or U9603 (N_9603,N_8756,N_8327);
nor U9604 (N_9604,N_8623,N_8913);
and U9605 (N_9605,N_8763,N_8728);
or U9606 (N_9606,N_8313,N_8996);
and U9607 (N_9607,N_8703,N_8384);
and U9608 (N_9608,N_8537,N_8873);
and U9609 (N_9609,N_8290,N_8351);
nand U9610 (N_9610,N_8524,N_8984);
nor U9611 (N_9611,N_8689,N_8622);
and U9612 (N_9612,N_8971,N_8869);
and U9613 (N_9613,N_8378,N_8960);
and U9614 (N_9614,N_8257,N_8699);
and U9615 (N_9615,N_8571,N_8625);
xor U9616 (N_9616,N_8756,N_8801);
and U9617 (N_9617,N_8390,N_8591);
nand U9618 (N_9618,N_8797,N_8835);
nand U9619 (N_9619,N_8782,N_8814);
nor U9620 (N_9620,N_8754,N_8925);
or U9621 (N_9621,N_8409,N_8753);
or U9622 (N_9622,N_8635,N_8351);
and U9623 (N_9623,N_8554,N_8963);
xnor U9624 (N_9624,N_8780,N_8667);
or U9625 (N_9625,N_8254,N_8956);
or U9626 (N_9626,N_8682,N_8530);
nor U9627 (N_9627,N_8345,N_8387);
or U9628 (N_9628,N_8738,N_8781);
nand U9629 (N_9629,N_8451,N_8346);
nor U9630 (N_9630,N_8706,N_8373);
and U9631 (N_9631,N_8978,N_8301);
and U9632 (N_9632,N_8586,N_8762);
and U9633 (N_9633,N_8983,N_8936);
or U9634 (N_9634,N_8962,N_8860);
nor U9635 (N_9635,N_8755,N_8672);
and U9636 (N_9636,N_8426,N_8291);
and U9637 (N_9637,N_8380,N_8626);
nor U9638 (N_9638,N_8629,N_8877);
nor U9639 (N_9639,N_8870,N_8676);
or U9640 (N_9640,N_8734,N_8408);
and U9641 (N_9641,N_8424,N_8885);
or U9642 (N_9642,N_8974,N_8896);
and U9643 (N_9643,N_8769,N_8330);
nand U9644 (N_9644,N_8440,N_8362);
or U9645 (N_9645,N_8836,N_8642);
xnor U9646 (N_9646,N_8938,N_8993);
and U9647 (N_9647,N_8464,N_8899);
nor U9648 (N_9648,N_8284,N_8795);
and U9649 (N_9649,N_8372,N_8652);
and U9650 (N_9650,N_8612,N_8261);
nor U9651 (N_9651,N_8832,N_8299);
nand U9652 (N_9652,N_8964,N_8280);
xnor U9653 (N_9653,N_8409,N_8887);
xor U9654 (N_9654,N_8878,N_8334);
nand U9655 (N_9655,N_8841,N_8787);
or U9656 (N_9656,N_8377,N_8518);
nand U9657 (N_9657,N_8303,N_8403);
nand U9658 (N_9658,N_8639,N_8695);
or U9659 (N_9659,N_8377,N_8433);
nor U9660 (N_9660,N_8940,N_8380);
or U9661 (N_9661,N_8842,N_8650);
or U9662 (N_9662,N_8576,N_8319);
xor U9663 (N_9663,N_8793,N_8795);
nand U9664 (N_9664,N_8869,N_8982);
or U9665 (N_9665,N_8837,N_8858);
nand U9666 (N_9666,N_8608,N_8797);
or U9667 (N_9667,N_8518,N_8627);
xor U9668 (N_9668,N_8264,N_8391);
or U9669 (N_9669,N_8373,N_8427);
or U9670 (N_9670,N_8779,N_8536);
and U9671 (N_9671,N_8442,N_8286);
xor U9672 (N_9672,N_8755,N_8576);
nor U9673 (N_9673,N_8569,N_8990);
nor U9674 (N_9674,N_8550,N_8698);
nand U9675 (N_9675,N_8341,N_8263);
nor U9676 (N_9676,N_8509,N_8613);
xor U9677 (N_9677,N_8874,N_8601);
xor U9678 (N_9678,N_8666,N_8707);
nand U9679 (N_9679,N_8303,N_8483);
or U9680 (N_9680,N_8681,N_8571);
or U9681 (N_9681,N_8297,N_8506);
and U9682 (N_9682,N_8904,N_8768);
nor U9683 (N_9683,N_8883,N_8615);
or U9684 (N_9684,N_8252,N_8289);
or U9685 (N_9685,N_8645,N_8478);
nand U9686 (N_9686,N_8650,N_8315);
nor U9687 (N_9687,N_8622,N_8792);
or U9688 (N_9688,N_8539,N_8949);
nor U9689 (N_9689,N_8347,N_8393);
or U9690 (N_9690,N_8684,N_8987);
xor U9691 (N_9691,N_8987,N_8989);
nand U9692 (N_9692,N_8553,N_8339);
nand U9693 (N_9693,N_8604,N_8820);
or U9694 (N_9694,N_8882,N_8563);
nor U9695 (N_9695,N_8742,N_8493);
nand U9696 (N_9696,N_8366,N_8633);
or U9697 (N_9697,N_8812,N_8677);
or U9698 (N_9698,N_8625,N_8914);
or U9699 (N_9699,N_8959,N_8424);
or U9700 (N_9700,N_8919,N_8810);
and U9701 (N_9701,N_8924,N_8959);
nor U9702 (N_9702,N_8721,N_8798);
nor U9703 (N_9703,N_8837,N_8316);
and U9704 (N_9704,N_8508,N_8996);
nand U9705 (N_9705,N_8967,N_8453);
nor U9706 (N_9706,N_8972,N_8678);
nor U9707 (N_9707,N_8663,N_8970);
or U9708 (N_9708,N_8343,N_8909);
xnor U9709 (N_9709,N_8355,N_8919);
xnor U9710 (N_9710,N_8254,N_8619);
or U9711 (N_9711,N_8782,N_8655);
and U9712 (N_9712,N_8641,N_8391);
nand U9713 (N_9713,N_8822,N_8306);
nand U9714 (N_9714,N_8718,N_8949);
or U9715 (N_9715,N_8881,N_8893);
nand U9716 (N_9716,N_8853,N_8606);
and U9717 (N_9717,N_8488,N_8437);
nor U9718 (N_9718,N_8586,N_8265);
and U9719 (N_9719,N_8829,N_8393);
nor U9720 (N_9720,N_8671,N_8350);
and U9721 (N_9721,N_8996,N_8390);
xor U9722 (N_9722,N_8659,N_8704);
xnor U9723 (N_9723,N_8969,N_8818);
xor U9724 (N_9724,N_8914,N_8968);
or U9725 (N_9725,N_8948,N_8877);
nor U9726 (N_9726,N_8658,N_8875);
nor U9727 (N_9727,N_8552,N_8734);
or U9728 (N_9728,N_8680,N_8278);
nor U9729 (N_9729,N_8991,N_8764);
xor U9730 (N_9730,N_8455,N_8768);
and U9731 (N_9731,N_8336,N_8761);
nor U9732 (N_9732,N_8287,N_8569);
or U9733 (N_9733,N_8858,N_8606);
nor U9734 (N_9734,N_8408,N_8719);
nor U9735 (N_9735,N_8829,N_8406);
or U9736 (N_9736,N_8311,N_8389);
nor U9737 (N_9737,N_8835,N_8761);
nor U9738 (N_9738,N_8603,N_8371);
or U9739 (N_9739,N_8449,N_8734);
xnor U9740 (N_9740,N_8999,N_8572);
nand U9741 (N_9741,N_8883,N_8385);
nand U9742 (N_9742,N_8982,N_8662);
nor U9743 (N_9743,N_8761,N_8533);
and U9744 (N_9744,N_8340,N_8659);
or U9745 (N_9745,N_8309,N_8700);
and U9746 (N_9746,N_8417,N_8298);
and U9747 (N_9747,N_8616,N_8330);
or U9748 (N_9748,N_8597,N_8551);
and U9749 (N_9749,N_8786,N_8628);
and U9750 (N_9750,N_9061,N_9486);
nand U9751 (N_9751,N_9736,N_9400);
nand U9752 (N_9752,N_9244,N_9650);
or U9753 (N_9753,N_9673,N_9266);
xnor U9754 (N_9754,N_9341,N_9638);
nand U9755 (N_9755,N_9725,N_9472);
nor U9756 (N_9756,N_9058,N_9492);
xor U9757 (N_9757,N_9134,N_9221);
or U9758 (N_9758,N_9245,N_9576);
nor U9759 (N_9759,N_9352,N_9347);
nor U9760 (N_9760,N_9585,N_9099);
nor U9761 (N_9761,N_9697,N_9672);
nor U9762 (N_9762,N_9278,N_9542);
and U9763 (N_9763,N_9212,N_9493);
nand U9764 (N_9764,N_9327,N_9277);
nand U9765 (N_9765,N_9595,N_9251);
nand U9766 (N_9766,N_9398,N_9580);
and U9767 (N_9767,N_9622,N_9391);
xor U9768 (N_9768,N_9397,N_9282);
nor U9769 (N_9769,N_9551,N_9142);
nand U9770 (N_9770,N_9183,N_9406);
and U9771 (N_9771,N_9315,N_9586);
nor U9772 (N_9772,N_9129,N_9163);
or U9773 (N_9773,N_9598,N_9021);
and U9774 (N_9774,N_9373,N_9228);
nor U9775 (N_9775,N_9111,N_9197);
nor U9776 (N_9776,N_9178,N_9574);
nor U9777 (N_9777,N_9036,N_9258);
nand U9778 (N_9778,N_9479,N_9507);
and U9779 (N_9779,N_9057,N_9363);
and U9780 (N_9780,N_9646,N_9381);
or U9781 (N_9781,N_9648,N_9149);
and U9782 (N_9782,N_9601,N_9417);
and U9783 (N_9783,N_9426,N_9664);
or U9784 (N_9784,N_9560,N_9686);
or U9785 (N_9785,N_9103,N_9465);
nor U9786 (N_9786,N_9074,N_9699);
and U9787 (N_9787,N_9559,N_9056);
or U9788 (N_9788,N_9035,N_9467);
or U9789 (N_9789,N_9466,N_9067);
nand U9790 (N_9790,N_9550,N_9105);
nand U9791 (N_9791,N_9308,N_9174);
nor U9792 (N_9792,N_9191,N_9563);
nand U9793 (N_9793,N_9445,N_9006);
or U9794 (N_9794,N_9716,N_9351);
nand U9795 (N_9795,N_9041,N_9541);
nand U9796 (N_9796,N_9499,N_9692);
or U9797 (N_9797,N_9602,N_9296);
nor U9798 (N_9798,N_9700,N_9032);
nand U9799 (N_9799,N_9185,N_9123);
xnor U9800 (N_9800,N_9038,N_9702);
nor U9801 (N_9801,N_9225,N_9167);
or U9802 (N_9802,N_9546,N_9500);
xor U9803 (N_9803,N_9484,N_9357);
and U9804 (N_9804,N_9524,N_9243);
xor U9805 (N_9805,N_9722,N_9442);
xnor U9806 (N_9806,N_9687,N_9085);
nor U9807 (N_9807,N_9179,N_9677);
and U9808 (N_9808,N_9594,N_9530);
or U9809 (N_9809,N_9195,N_9135);
nand U9810 (N_9810,N_9469,N_9659);
nand U9811 (N_9811,N_9423,N_9114);
or U9812 (N_9812,N_9124,N_9495);
xor U9813 (N_9813,N_9115,N_9512);
or U9814 (N_9814,N_9079,N_9414);
or U9815 (N_9815,N_9269,N_9411);
and U9816 (N_9816,N_9305,N_9353);
or U9817 (N_9817,N_9667,N_9377);
nor U9818 (N_9818,N_9077,N_9583);
and U9819 (N_9819,N_9342,N_9435);
or U9820 (N_9820,N_9713,N_9360);
or U9821 (N_9821,N_9177,N_9651);
nor U9822 (N_9822,N_9165,N_9140);
nor U9823 (N_9823,N_9072,N_9248);
nor U9824 (N_9824,N_9131,N_9476);
or U9825 (N_9825,N_9012,N_9297);
and U9826 (N_9826,N_9071,N_9535);
and U9827 (N_9827,N_9480,N_9421);
and U9828 (N_9828,N_9169,N_9196);
nand U9829 (N_9829,N_9683,N_9365);
and U9830 (N_9830,N_9572,N_9705);
and U9831 (N_9831,N_9506,N_9270);
or U9832 (N_9832,N_9022,N_9017);
nand U9833 (N_9833,N_9275,N_9468);
nor U9834 (N_9834,N_9049,N_9428);
nor U9835 (N_9835,N_9289,N_9592);
or U9836 (N_9836,N_9382,N_9189);
or U9837 (N_9837,N_9749,N_9656);
and U9838 (N_9838,N_9520,N_9090);
nor U9839 (N_9839,N_9652,N_9273);
or U9840 (N_9840,N_9561,N_9358);
nand U9841 (N_9841,N_9660,N_9604);
nand U9842 (N_9842,N_9459,N_9047);
nor U9843 (N_9843,N_9075,N_9742);
or U9844 (N_9844,N_9511,N_9577);
and U9845 (N_9845,N_9238,N_9141);
or U9846 (N_9846,N_9732,N_9587);
nand U9847 (N_9847,N_9211,N_9291);
or U9848 (N_9848,N_9657,N_9116);
and U9849 (N_9849,N_9402,N_9454);
or U9850 (N_9850,N_9457,N_9614);
and U9851 (N_9851,N_9002,N_9707);
nor U9852 (N_9852,N_9706,N_9582);
nand U9853 (N_9853,N_9219,N_9117);
nor U9854 (N_9854,N_9300,N_9101);
and U9855 (N_9855,N_9125,N_9098);
nor U9856 (N_9856,N_9139,N_9525);
or U9857 (N_9857,N_9218,N_9120);
nor U9858 (N_9858,N_9655,N_9444);
nor U9859 (N_9859,N_9171,N_9376);
or U9860 (N_9860,N_9069,N_9470);
nor U9861 (N_9861,N_9431,N_9724);
or U9862 (N_9862,N_9073,N_9362);
nand U9863 (N_9863,N_9184,N_9051);
or U9864 (N_9864,N_9094,N_9045);
or U9865 (N_9865,N_9625,N_9523);
nor U9866 (N_9866,N_9048,N_9663);
nor U9867 (N_9867,N_9538,N_9126);
nand U9868 (N_9868,N_9256,N_9557);
or U9869 (N_9869,N_9581,N_9158);
xnor U9870 (N_9870,N_9746,N_9693);
nand U9871 (N_9871,N_9611,N_9387);
nor U9872 (N_9872,N_9681,N_9146);
or U9873 (N_9873,N_9737,N_9691);
and U9874 (N_9874,N_9534,N_9626);
xnor U9875 (N_9875,N_9393,N_9010);
or U9876 (N_9876,N_9145,N_9319);
xor U9877 (N_9877,N_9740,N_9689);
and U9878 (N_9878,N_9276,N_9320);
nand U9879 (N_9879,N_9175,N_9734);
nand U9880 (N_9880,N_9159,N_9436);
or U9881 (N_9881,N_9517,N_9224);
and U9882 (N_9882,N_9739,N_9370);
nor U9883 (N_9883,N_9422,N_9588);
or U9884 (N_9884,N_9122,N_9003);
nor U9885 (N_9885,N_9569,N_9412);
or U9886 (N_9886,N_9433,N_9247);
and U9887 (N_9887,N_9407,N_9513);
and U9888 (N_9888,N_9324,N_9043);
xor U9889 (N_9889,N_9578,N_9025);
nor U9890 (N_9890,N_9425,N_9223);
and U9891 (N_9891,N_9390,N_9237);
nor U9892 (N_9892,N_9590,N_9503);
xnor U9893 (N_9893,N_9232,N_9635);
nand U9894 (N_9894,N_9458,N_9579);
nor U9895 (N_9895,N_9264,N_9628);
or U9896 (N_9896,N_9285,N_9063);
or U9897 (N_9897,N_9555,N_9000);
or U9898 (N_9898,N_9645,N_9632);
xnor U9899 (N_9899,N_9509,N_9093);
nand U9900 (N_9900,N_9344,N_9603);
or U9901 (N_9901,N_9318,N_9610);
nand U9902 (N_9902,N_9455,N_9389);
and U9903 (N_9903,N_9272,N_9182);
nand U9904 (N_9904,N_9483,N_9662);
or U9905 (N_9905,N_9494,N_9214);
nor U9906 (N_9906,N_9015,N_9331);
nand U9907 (N_9907,N_9521,N_9157);
and U9908 (N_9908,N_9311,N_9104);
nand U9909 (N_9909,N_9137,N_9649);
and U9910 (N_9910,N_9384,N_9263);
xnor U9911 (N_9911,N_9250,N_9338);
or U9912 (N_9912,N_9661,N_9288);
or U9913 (N_9913,N_9350,N_9679);
xnor U9914 (N_9914,N_9037,N_9597);
and U9915 (N_9915,N_9392,N_9526);
nand U9916 (N_9916,N_9226,N_9441);
and U9917 (N_9917,N_9078,N_9418);
nor U9918 (N_9918,N_9631,N_9127);
nor U9919 (N_9919,N_9608,N_9514);
and U9920 (N_9920,N_9685,N_9385);
or U9921 (N_9921,N_9473,N_9231);
nand U9922 (N_9922,N_9440,N_9055);
nor U9923 (N_9923,N_9354,N_9086);
or U9924 (N_9924,N_9034,N_9607);
xnor U9925 (N_9925,N_9533,N_9676);
and U9926 (N_9926,N_9430,N_9497);
and U9927 (N_9927,N_9540,N_9719);
xor U9928 (N_9928,N_9147,N_9314);
nand U9929 (N_9929,N_9170,N_9206);
xnor U9930 (N_9930,N_9684,N_9102);
and U9931 (N_9931,N_9748,N_9284);
nor U9932 (N_9932,N_9408,N_9304);
or U9933 (N_9933,N_9227,N_9532);
xnor U9934 (N_9934,N_9571,N_9720);
nor U9935 (N_9935,N_9419,N_9570);
and U9936 (N_9936,N_9089,N_9505);
nand U9937 (N_9937,N_9715,N_9153);
or U9938 (N_9938,N_9543,N_9413);
nand U9939 (N_9939,N_9404,N_9229);
and U9940 (N_9940,N_9348,N_9088);
or U9941 (N_9941,N_9704,N_9738);
xor U9942 (N_9942,N_9567,N_9312);
nand U9943 (N_9943,N_9302,N_9138);
and U9944 (N_9944,N_9031,N_9013);
nand U9945 (N_9945,N_9463,N_9005);
nand U9946 (N_9946,N_9584,N_9680);
nand U9947 (N_9947,N_9081,N_9011);
nand U9948 (N_9948,N_9053,N_9420);
xor U9949 (N_9949,N_9029,N_9027);
nor U9950 (N_9950,N_9380,N_9236);
nand U9951 (N_9951,N_9447,N_9675);
nand U9952 (N_9952,N_9489,N_9144);
nor U9953 (N_9953,N_9213,N_9233);
and U9954 (N_9954,N_9016,N_9471);
xnor U9955 (N_9955,N_9207,N_9204);
nand U9956 (N_9956,N_9456,N_9621);
xor U9957 (N_9957,N_9334,N_9453);
xor U9958 (N_9958,N_9059,N_9537);
nor U9959 (N_9959,N_9619,N_9708);
and U9960 (N_9960,N_9162,N_9620);
xnor U9961 (N_9961,N_9670,N_9694);
or U9962 (N_9962,N_9313,N_9554);
xnor U9963 (N_9963,N_9432,N_9019);
or U9964 (N_9964,N_9379,N_9014);
or U9965 (N_9965,N_9084,N_9293);
and U9966 (N_9966,N_9295,N_9399);
and U9967 (N_9967,N_9405,N_9630);
nor U9968 (N_9968,N_9415,N_9642);
nor U9969 (N_9969,N_9064,N_9150);
or U9970 (N_9970,N_9361,N_9695);
nor U9971 (N_9971,N_9599,N_9616);
and U9972 (N_9972,N_9508,N_9332);
and U9973 (N_9973,N_9046,N_9726);
and U9974 (N_9974,N_9188,N_9292);
or U9975 (N_9975,N_9222,N_9666);
or U9976 (N_9976,N_9255,N_9378);
nor U9977 (N_9977,N_9623,N_9148);
and U9978 (N_9978,N_9464,N_9596);
or U9979 (N_9979,N_9488,N_9346);
nor U9980 (N_9980,N_9460,N_9065);
and U9981 (N_9981,N_9100,N_9249);
or U9982 (N_9982,N_9136,N_9593);
and U9983 (N_9983,N_9703,N_9723);
or U9984 (N_9984,N_9186,N_9082);
and U9985 (N_9985,N_9443,N_9491);
nand U9986 (N_9986,N_9682,N_9710);
xnor U9987 (N_9987,N_9409,N_9629);
nor U9988 (N_9988,N_9092,N_9234);
or U9989 (N_9989,N_9688,N_9155);
nand U9990 (N_9990,N_9539,N_9640);
nand U9991 (N_9991,N_9235,N_9589);
or U9992 (N_9992,N_9427,N_9173);
and U9993 (N_9993,N_9033,N_9368);
and U9994 (N_9994,N_9439,N_9083);
nand U9995 (N_9995,N_9070,N_9556);
nor U9996 (N_9996,N_9307,N_9118);
or U9997 (N_9997,N_9565,N_9267);
and U9998 (N_9998,N_9215,N_9558);
nand U9999 (N_9999,N_9097,N_9653);
and U10000 (N_10000,N_9452,N_9612);
or U10001 (N_10001,N_9239,N_9449);
or U10002 (N_10002,N_9210,N_9450);
nand U10003 (N_10003,N_9375,N_9383);
xor U10004 (N_10004,N_9330,N_9545);
nor U10005 (N_10005,N_9271,N_9437);
or U10006 (N_10006,N_9333,N_9721);
or U10007 (N_10007,N_9299,N_9709);
and U10008 (N_10008,N_9575,N_9429);
nor U10009 (N_10009,N_9253,N_9388);
or U10010 (N_10010,N_9156,N_9529);
or U10011 (N_10011,N_9477,N_9080);
or U10012 (N_10012,N_9605,N_9403);
nor U10013 (N_10013,N_9128,N_9042);
nor U10014 (N_10014,N_9424,N_9259);
nor U10015 (N_10015,N_9714,N_9478);
nand U10016 (N_10016,N_9246,N_9260);
nand U10017 (N_10017,N_9108,N_9161);
nand U10018 (N_10018,N_9257,N_9743);
xnor U10019 (N_10019,N_9600,N_9335);
and U10020 (N_10020,N_9730,N_9050);
or U10021 (N_10021,N_9690,N_9096);
or U10022 (N_10022,N_9321,N_9181);
nor U10023 (N_10023,N_9696,N_9166);
xor U10024 (N_10024,N_9735,N_9323);
nand U10025 (N_10025,N_9202,N_9252);
nor U10026 (N_10026,N_9240,N_9728);
or U10027 (N_10027,N_9194,N_9281);
nand U10028 (N_10028,N_9192,N_9671);
or U10029 (N_10029,N_9242,N_9668);
or U10030 (N_10030,N_9474,N_9634);
xor U10031 (N_10031,N_9717,N_9698);
and U10032 (N_10032,N_9522,N_9254);
nand U10033 (N_10033,N_9023,N_9369);
or U10034 (N_10034,N_9669,N_9180);
and U10035 (N_10035,N_9008,N_9109);
nand U10036 (N_10036,N_9303,N_9261);
and U10037 (N_10037,N_9609,N_9310);
nand U10038 (N_10038,N_9451,N_9168);
nand U10039 (N_10039,N_9265,N_9639);
and U10040 (N_10040,N_9279,N_9618);
and U10041 (N_10041,N_9396,N_9544);
nand U10042 (N_10042,N_9340,N_9328);
nor U10043 (N_10043,N_9110,N_9615);
and U10044 (N_10044,N_9367,N_9501);
or U10045 (N_10045,N_9203,N_9658);
and U10046 (N_10046,N_9054,N_9654);
or U10047 (N_10047,N_9549,N_9198);
nand U10048 (N_10048,N_9268,N_9510);
nand U10049 (N_10049,N_9386,N_9306);
nand U10050 (N_10050,N_9107,N_9741);
or U10051 (N_10051,N_9401,N_9633);
nand U10052 (N_10052,N_9502,N_9349);
or U10053 (N_10053,N_9481,N_9193);
nor U10054 (N_10054,N_9356,N_9009);
nand U10055 (N_10055,N_9712,N_9026);
or U10056 (N_10056,N_9066,N_9644);
or U10057 (N_10057,N_9290,N_9566);
nand U10058 (N_10058,N_9372,N_9280);
nor U10059 (N_10059,N_9241,N_9498);
nand U10060 (N_10060,N_9744,N_9325);
and U10061 (N_10061,N_9317,N_9143);
nor U10062 (N_10062,N_9217,N_9573);
nand U10063 (N_10063,N_9643,N_9462);
xor U10064 (N_10064,N_9637,N_9665);
xor U10065 (N_10065,N_9030,N_9617);
nand U10066 (N_10066,N_9007,N_9087);
nor U10067 (N_10067,N_9062,N_9152);
xor U10068 (N_10068,N_9286,N_9040);
nand U10069 (N_10069,N_9641,N_9519);
nor U10070 (N_10070,N_9106,N_9515);
or U10071 (N_10071,N_9496,N_9337);
nand U10072 (N_10072,N_9187,N_9461);
nand U10073 (N_10073,N_9701,N_9119);
nor U10074 (N_10074,N_9627,N_9316);
or U10075 (N_10075,N_9130,N_9287);
nand U10076 (N_10076,N_9091,N_9283);
and U10077 (N_10077,N_9164,N_9060);
nand U10078 (N_10078,N_9678,N_9018);
or U10079 (N_10079,N_9718,N_9547);
xor U10080 (N_10080,N_9371,N_9624);
nor U10081 (N_10081,N_9674,N_9216);
or U10082 (N_10082,N_9095,N_9729);
nand U10083 (N_10083,N_9294,N_9438);
and U10084 (N_10084,N_9446,N_9200);
and U10085 (N_10085,N_9044,N_9343);
nand U10086 (N_10086,N_9132,N_9024);
nor U10087 (N_10087,N_9395,N_9208);
or U10088 (N_10088,N_9274,N_9004);
or U10089 (N_10089,N_9504,N_9199);
nor U10090 (N_10090,N_9366,N_9531);
and U10091 (N_10091,N_9355,N_9548);
and U10092 (N_10092,N_9482,N_9113);
nor U10093 (N_10093,N_9606,N_9326);
and U10094 (N_10094,N_9490,N_9731);
and U10095 (N_10095,N_9727,N_9364);
nand U10096 (N_10096,N_9190,N_9711);
xor U10097 (N_10097,N_9154,N_9564);
xor U10098 (N_10098,N_9733,N_9518);
nand U10099 (N_10099,N_9121,N_9528);
nor U10100 (N_10100,N_9475,N_9485);
nor U10101 (N_10101,N_9172,N_9591);
nand U10102 (N_10102,N_9552,N_9052);
and U10103 (N_10103,N_9028,N_9747);
xnor U10104 (N_10104,N_9039,N_9336);
xor U10105 (N_10105,N_9448,N_9068);
and U10106 (N_10106,N_9133,N_9209);
nor U10107 (N_10107,N_9020,N_9076);
nor U10108 (N_10108,N_9160,N_9345);
and U10109 (N_10109,N_9205,N_9394);
or U10110 (N_10110,N_9322,N_9516);
nor U10111 (N_10111,N_9309,N_9339);
and U10112 (N_10112,N_9201,N_9527);
nand U10113 (N_10113,N_9230,N_9359);
or U10114 (N_10114,N_9416,N_9568);
or U10115 (N_10115,N_9553,N_9536);
nand U10116 (N_10116,N_9112,N_9262);
nand U10117 (N_10117,N_9176,N_9151);
or U10118 (N_10118,N_9636,N_9410);
nor U10119 (N_10119,N_9001,N_9434);
nand U10120 (N_10120,N_9562,N_9301);
nand U10121 (N_10121,N_9298,N_9745);
xnor U10122 (N_10122,N_9374,N_9487);
nand U10123 (N_10123,N_9329,N_9647);
and U10124 (N_10124,N_9613,N_9220);
or U10125 (N_10125,N_9257,N_9599);
or U10126 (N_10126,N_9015,N_9672);
nor U10127 (N_10127,N_9023,N_9679);
xor U10128 (N_10128,N_9171,N_9168);
nor U10129 (N_10129,N_9717,N_9357);
nor U10130 (N_10130,N_9681,N_9127);
nand U10131 (N_10131,N_9715,N_9051);
or U10132 (N_10132,N_9219,N_9511);
nand U10133 (N_10133,N_9605,N_9687);
and U10134 (N_10134,N_9119,N_9711);
nor U10135 (N_10135,N_9042,N_9472);
nor U10136 (N_10136,N_9140,N_9004);
nand U10137 (N_10137,N_9072,N_9018);
nand U10138 (N_10138,N_9398,N_9731);
and U10139 (N_10139,N_9221,N_9548);
and U10140 (N_10140,N_9173,N_9267);
and U10141 (N_10141,N_9628,N_9499);
and U10142 (N_10142,N_9678,N_9374);
nor U10143 (N_10143,N_9720,N_9341);
nor U10144 (N_10144,N_9589,N_9625);
and U10145 (N_10145,N_9058,N_9396);
or U10146 (N_10146,N_9560,N_9321);
and U10147 (N_10147,N_9470,N_9039);
nand U10148 (N_10148,N_9266,N_9236);
xnor U10149 (N_10149,N_9338,N_9026);
nand U10150 (N_10150,N_9561,N_9117);
nor U10151 (N_10151,N_9147,N_9565);
or U10152 (N_10152,N_9315,N_9067);
or U10153 (N_10153,N_9179,N_9156);
nand U10154 (N_10154,N_9680,N_9741);
or U10155 (N_10155,N_9009,N_9566);
or U10156 (N_10156,N_9139,N_9431);
and U10157 (N_10157,N_9548,N_9376);
and U10158 (N_10158,N_9613,N_9748);
and U10159 (N_10159,N_9347,N_9561);
or U10160 (N_10160,N_9488,N_9459);
or U10161 (N_10161,N_9072,N_9179);
or U10162 (N_10162,N_9567,N_9324);
and U10163 (N_10163,N_9504,N_9009);
or U10164 (N_10164,N_9377,N_9598);
nand U10165 (N_10165,N_9658,N_9451);
nor U10166 (N_10166,N_9591,N_9185);
nor U10167 (N_10167,N_9414,N_9355);
xnor U10168 (N_10168,N_9499,N_9022);
xor U10169 (N_10169,N_9227,N_9422);
nor U10170 (N_10170,N_9471,N_9659);
nand U10171 (N_10171,N_9264,N_9205);
or U10172 (N_10172,N_9644,N_9155);
or U10173 (N_10173,N_9322,N_9212);
nor U10174 (N_10174,N_9284,N_9317);
xnor U10175 (N_10175,N_9520,N_9594);
xor U10176 (N_10176,N_9101,N_9678);
or U10177 (N_10177,N_9099,N_9206);
or U10178 (N_10178,N_9700,N_9039);
or U10179 (N_10179,N_9729,N_9385);
nor U10180 (N_10180,N_9746,N_9627);
nand U10181 (N_10181,N_9246,N_9397);
nand U10182 (N_10182,N_9293,N_9273);
or U10183 (N_10183,N_9199,N_9229);
or U10184 (N_10184,N_9547,N_9064);
or U10185 (N_10185,N_9624,N_9399);
and U10186 (N_10186,N_9385,N_9384);
nand U10187 (N_10187,N_9349,N_9599);
or U10188 (N_10188,N_9291,N_9558);
nand U10189 (N_10189,N_9433,N_9157);
and U10190 (N_10190,N_9649,N_9516);
nor U10191 (N_10191,N_9454,N_9521);
and U10192 (N_10192,N_9369,N_9648);
xor U10193 (N_10193,N_9522,N_9572);
nor U10194 (N_10194,N_9044,N_9632);
nor U10195 (N_10195,N_9422,N_9721);
or U10196 (N_10196,N_9454,N_9619);
nor U10197 (N_10197,N_9734,N_9129);
and U10198 (N_10198,N_9423,N_9033);
nand U10199 (N_10199,N_9188,N_9060);
and U10200 (N_10200,N_9279,N_9616);
nand U10201 (N_10201,N_9198,N_9635);
xnor U10202 (N_10202,N_9358,N_9575);
nor U10203 (N_10203,N_9073,N_9187);
or U10204 (N_10204,N_9683,N_9744);
and U10205 (N_10205,N_9672,N_9434);
nor U10206 (N_10206,N_9609,N_9200);
nor U10207 (N_10207,N_9494,N_9203);
or U10208 (N_10208,N_9354,N_9689);
nand U10209 (N_10209,N_9060,N_9636);
or U10210 (N_10210,N_9491,N_9039);
nand U10211 (N_10211,N_9706,N_9276);
or U10212 (N_10212,N_9493,N_9597);
xnor U10213 (N_10213,N_9603,N_9725);
nand U10214 (N_10214,N_9013,N_9640);
xor U10215 (N_10215,N_9325,N_9130);
nand U10216 (N_10216,N_9367,N_9228);
nand U10217 (N_10217,N_9102,N_9518);
xor U10218 (N_10218,N_9329,N_9620);
xnor U10219 (N_10219,N_9188,N_9277);
nand U10220 (N_10220,N_9009,N_9326);
and U10221 (N_10221,N_9142,N_9728);
nand U10222 (N_10222,N_9709,N_9520);
nor U10223 (N_10223,N_9459,N_9432);
and U10224 (N_10224,N_9503,N_9615);
or U10225 (N_10225,N_9180,N_9452);
nand U10226 (N_10226,N_9487,N_9288);
nand U10227 (N_10227,N_9047,N_9574);
or U10228 (N_10228,N_9486,N_9594);
xnor U10229 (N_10229,N_9370,N_9178);
and U10230 (N_10230,N_9085,N_9036);
and U10231 (N_10231,N_9589,N_9117);
xor U10232 (N_10232,N_9358,N_9224);
and U10233 (N_10233,N_9154,N_9437);
or U10234 (N_10234,N_9423,N_9699);
or U10235 (N_10235,N_9425,N_9515);
nor U10236 (N_10236,N_9516,N_9409);
nand U10237 (N_10237,N_9093,N_9468);
and U10238 (N_10238,N_9250,N_9314);
nand U10239 (N_10239,N_9653,N_9146);
or U10240 (N_10240,N_9073,N_9702);
xnor U10241 (N_10241,N_9334,N_9232);
nor U10242 (N_10242,N_9370,N_9500);
and U10243 (N_10243,N_9122,N_9544);
nand U10244 (N_10244,N_9315,N_9663);
or U10245 (N_10245,N_9568,N_9014);
nor U10246 (N_10246,N_9613,N_9234);
and U10247 (N_10247,N_9271,N_9552);
and U10248 (N_10248,N_9662,N_9745);
nor U10249 (N_10249,N_9237,N_9629);
nor U10250 (N_10250,N_9151,N_9060);
and U10251 (N_10251,N_9091,N_9698);
nor U10252 (N_10252,N_9227,N_9594);
xnor U10253 (N_10253,N_9729,N_9637);
or U10254 (N_10254,N_9450,N_9438);
nor U10255 (N_10255,N_9321,N_9521);
and U10256 (N_10256,N_9149,N_9637);
or U10257 (N_10257,N_9674,N_9354);
nand U10258 (N_10258,N_9494,N_9646);
and U10259 (N_10259,N_9475,N_9061);
or U10260 (N_10260,N_9042,N_9737);
nor U10261 (N_10261,N_9713,N_9099);
nand U10262 (N_10262,N_9271,N_9225);
or U10263 (N_10263,N_9038,N_9390);
or U10264 (N_10264,N_9530,N_9378);
nand U10265 (N_10265,N_9444,N_9545);
and U10266 (N_10266,N_9193,N_9689);
and U10267 (N_10267,N_9170,N_9493);
nor U10268 (N_10268,N_9265,N_9246);
xor U10269 (N_10269,N_9132,N_9519);
nand U10270 (N_10270,N_9488,N_9149);
nor U10271 (N_10271,N_9075,N_9288);
nand U10272 (N_10272,N_9162,N_9388);
and U10273 (N_10273,N_9527,N_9069);
xnor U10274 (N_10274,N_9304,N_9102);
nand U10275 (N_10275,N_9132,N_9223);
nand U10276 (N_10276,N_9227,N_9019);
or U10277 (N_10277,N_9687,N_9444);
xnor U10278 (N_10278,N_9418,N_9017);
nand U10279 (N_10279,N_9170,N_9069);
or U10280 (N_10280,N_9044,N_9175);
nand U10281 (N_10281,N_9651,N_9068);
nand U10282 (N_10282,N_9728,N_9273);
and U10283 (N_10283,N_9703,N_9461);
and U10284 (N_10284,N_9236,N_9387);
or U10285 (N_10285,N_9138,N_9612);
nor U10286 (N_10286,N_9515,N_9434);
xor U10287 (N_10287,N_9443,N_9374);
and U10288 (N_10288,N_9137,N_9317);
nor U10289 (N_10289,N_9327,N_9687);
nor U10290 (N_10290,N_9087,N_9675);
and U10291 (N_10291,N_9217,N_9064);
nand U10292 (N_10292,N_9643,N_9359);
nand U10293 (N_10293,N_9130,N_9566);
and U10294 (N_10294,N_9223,N_9468);
and U10295 (N_10295,N_9573,N_9041);
nor U10296 (N_10296,N_9187,N_9632);
or U10297 (N_10297,N_9514,N_9431);
nand U10298 (N_10298,N_9038,N_9532);
and U10299 (N_10299,N_9462,N_9146);
and U10300 (N_10300,N_9606,N_9129);
xnor U10301 (N_10301,N_9589,N_9662);
or U10302 (N_10302,N_9542,N_9687);
or U10303 (N_10303,N_9003,N_9746);
nor U10304 (N_10304,N_9377,N_9457);
and U10305 (N_10305,N_9676,N_9459);
or U10306 (N_10306,N_9041,N_9614);
xnor U10307 (N_10307,N_9198,N_9523);
nor U10308 (N_10308,N_9351,N_9059);
nand U10309 (N_10309,N_9652,N_9432);
or U10310 (N_10310,N_9165,N_9185);
or U10311 (N_10311,N_9174,N_9177);
nor U10312 (N_10312,N_9734,N_9003);
or U10313 (N_10313,N_9559,N_9095);
and U10314 (N_10314,N_9016,N_9177);
nand U10315 (N_10315,N_9207,N_9081);
xnor U10316 (N_10316,N_9348,N_9469);
xnor U10317 (N_10317,N_9579,N_9366);
or U10318 (N_10318,N_9347,N_9503);
nand U10319 (N_10319,N_9356,N_9370);
xor U10320 (N_10320,N_9550,N_9375);
and U10321 (N_10321,N_9474,N_9184);
and U10322 (N_10322,N_9081,N_9529);
xor U10323 (N_10323,N_9600,N_9312);
nor U10324 (N_10324,N_9722,N_9205);
nand U10325 (N_10325,N_9652,N_9425);
and U10326 (N_10326,N_9186,N_9518);
nor U10327 (N_10327,N_9730,N_9339);
nor U10328 (N_10328,N_9362,N_9156);
nor U10329 (N_10329,N_9240,N_9446);
xnor U10330 (N_10330,N_9255,N_9576);
nor U10331 (N_10331,N_9441,N_9186);
nor U10332 (N_10332,N_9603,N_9667);
or U10333 (N_10333,N_9745,N_9169);
xnor U10334 (N_10334,N_9170,N_9176);
nand U10335 (N_10335,N_9660,N_9300);
or U10336 (N_10336,N_9517,N_9550);
or U10337 (N_10337,N_9745,N_9551);
and U10338 (N_10338,N_9692,N_9391);
xor U10339 (N_10339,N_9241,N_9208);
xnor U10340 (N_10340,N_9338,N_9655);
and U10341 (N_10341,N_9630,N_9207);
nand U10342 (N_10342,N_9530,N_9452);
nand U10343 (N_10343,N_9167,N_9453);
and U10344 (N_10344,N_9294,N_9432);
xnor U10345 (N_10345,N_9668,N_9223);
xor U10346 (N_10346,N_9339,N_9027);
nor U10347 (N_10347,N_9202,N_9003);
xnor U10348 (N_10348,N_9070,N_9466);
or U10349 (N_10349,N_9212,N_9144);
nand U10350 (N_10350,N_9570,N_9241);
and U10351 (N_10351,N_9380,N_9704);
or U10352 (N_10352,N_9165,N_9526);
or U10353 (N_10353,N_9464,N_9166);
nand U10354 (N_10354,N_9030,N_9229);
nor U10355 (N_10355,N_9458,N_9158);
nor U10356 (N_10356,N_9570,N_9306);
nor U10357 (N_10357,N_9675,N_9028);
nor U10358 (N_10358,N_9286,N_9673);
nand U10359 (N_10359,N_9476,N_9401);
nand U10360 (N_10360,N_9081,N_9298);
nor U10361 (N_10361,N_9076,N_9427);
nor U10362 (N_10362,N_9484,N_9693);
or U10363 (N_10363,N_9370,N_9042);
or U10364 (N_10364,N_9100,N_9559);
and U10365 (N_10365,N_9715,N_9682);
nor U10366 (N_10366,N_9015,N_9492);
nor U10367 (N_10367,N_9428,N_9116);
xnor U10368 (N_10368,N_9564,N_9463);
nor U10369 (N_10369,N_9346,N_9610);
nor U10370 (N_10370,N_9418,N_9012);
and U10371 (N_10371,N_9611,N_9727);
nand U10372 (N_10372,N_9438,N_9399);
and U10373 (N_10373,N_9715,N_9334);
xnor U10374 (N_10374,N_9420,N_9475);
or U10375 (N_10375,N_9586,N_9355);
nand U10376 (N_10376,N_9039,N_9693);
or U10377 (N_10377,N_9702,N_9672);
or U10378 (N_10378,N_9718,N_9300);
and U10379 (N_10379,N_9670,N_9259);
and U10380 (N_10380,N_9668,N_9537);
nand U10381 (N_10381,N_9400,N_9273);
or U10382 (N_10382,N_9485,N_9463);
nand U10383 (N_10383,N_9483,N_9520);
and U10384 (N_10384,N_9510,N_9428);
nor U10385 (N_10385,N_9149,N_9169);
or U10386 (N_10386,N_9013,N_9411);
or U10387 (N_10387,N_9093,N_9412);
nand U10388 (N_10388,N_9242,N_9532);
and U10389 (N_10389,N_9397,N_9584);
or U10390 (N_10390,N_9126,N_9367);
nand U10391 (N_10391,N_9249,N_9465);
nor U10392 (N_10392,N_9370,N_9112);
xnor U10393 (N_10393,N_9697,N_9548);
nand U10394 (N_10394,N_9403,N_9005);
xor U10395 (N_10395,N_9456,N_9074);
nand U10396 (N_10396,N_9260,N_9570);
or U10397 (N_10397,N_9300,N_9020);
or U10398 (N_10398,N_9017,N_9643);
and U10399 (N_10399,N_9237,N_9042);
or U10400 (N_10400,N_9304,N_9653);
and U10401 (N_10401,N_9400,N_9093);
nand U10402 (N_10402,N_9388,N_9079);
nor U10403 (N_10403,N_9354,N_9387);
nor U10404 (N_10404,N_9004,N_9357);
or U10405 (N_10405,N_9344,N_9054);
nand U10406 (N_10406,N_9439,N_9272);
and U10407 (N_10407,N_9164,N_9731);
and U10408 (N_10408,N_9525,N_9741);
nor U10409 (N_10409,N_9719,N_9605);
nand U10410 (N_10410,N_9076,N_9575);
xor U10411 (N_10411,N_9059,N_9307);
nand U10412 (N_10412,N_9455,N_9332);
nor U10413 (N_10413,N_9243,N_9151);
nand U10414 (N_10414,N_9435,N_9526);
nor U10415 (N_10415,N_9737,N_9097);
or U10416 (N_10416,N_9625,N_9509);
and U10417 (N_10417,N_9580,N_9413);
and U10418 (N_10418,N_9626,N_9414);
or U10419 (N_10419,N_9179,N_9465);
and U10420 (N_10420,N_9119,N_9334);
and U10421 (N_10421,N_9483,N_9456);
and U10422 (N_10422,N_9621,N_9229);
or U10423 (N_10423,N_9547,N_9310);
or U10424 (N_10424,N_9506,N_9674);
nor U10425 (N_10425,N_9359,N_9029);
or U10426 (N_10426,N_9447,N_9739);
nor U10427 (N_10427,N_9329,N_9706);
nor U10428 (N_10428,N_9563,N_9547);
or U10429 (N_10429,N_9422,N_9118);
or U10430 (N_10430,N_9169,N_9110);
nor U10431 (N_10431,N_9523,N_9740);
or U10432 (N_10432,N_9232,N_9198);
nand U10433 (N_10433,N_9254,N_9397);
xnor U10434 (N_10434,N_9113,N_9509);
nor U10435 (N_10435,N_9592,N_9683);
and U10436 (N_10436,N_9668,N_9209);
nor U10437 (N_10437,N_9135,N_9010);
xnor U10438 (N_10438,N_9400,N_9040);
and U10439 (N_10439,N_9163,N_9490);
and U10440 (N_10440,N_9505,N_9071);
xor U10441 (N_10441,N_9317,N_9201);
or U10442 (N_10442,N_9556,N_9421);
and U10443 (N_10443,N_9295,N_9492);
nand U10444 (N_10444,N_9519,N_9585);
nor U10445 (N_10445,N_9272,N_9462);
nand U10446 (N_10446,N_9109,N_9557);
nand U10447 (N_10447,N_9571,N_9587);
nor U10448 (N_10448,N_9072,N_9744);
and U10449 (N_10449,N_9124,N_9551);
nor U10450 (N_10450,N_9636,N_9037);
xor U10451 (N_10451,N_9539,N_9419);
or U10452 (N_10452,N_9692,N_9085);
nand U10453 (N_10453,N_9362,N_9545);
and U10454 (N_10454,N_9498,N_9662);
nand U10455 (N_10455,N_9649,N_9171);
nor U10456 (N_10456,N_9396,N_9702);
xor U10457 (N_10457,N_9669,N_9400);
nand U10458 (N_10458,N_9646,N_9559);
nor U10459 (N_10459,N_9576,N_9117);
or U10460 (N_10460,N_9658,N_9555);
or U10461 (N_10461,N_9648,N_9337);
nand U10462 (N_10462,N_9684,N_9113);
and U10463 (N_10463,N_9537,N_9456);
or U10464 (N_10464,N_9720,N_9120);
nand U10465 (N_10465,N_9454,N_9268);
xnor U10466 (N_10466,N_9304,N_9522);
or U10467 (N_10467,N_9286,N_9015);
nor U10468 (N_10468,N_9523,N_9219);
or U10469 (N_10469,N_9082,N_9720);
and U10470 (N_10470,N_9396,N_9641);
and U10471 (N_10471,N_9118,N_9494);
and U10472 (N_10472,N_9109,N_9660);
and U10473 (N_10473,N_9053,N_9196);
nand U10474 (N_10474,N_9081,N_9353);
and U10475 (N_10475,N_9103,N_9439);
or U10476 (N_10476,N_9454,N_9490);
and U10477 (N_10477,N_9665,N_9155);
and U10478 (N_10478,N_9329,N_9698);
or U10479 (N_10479,N_9562,N_9577);
nand U10480 (N_10480,N_9317,N_9711);
or U10481 (N_10481,N_9259,N_9180);
nand U10482 (N_10482,N_9617,N_9457);
nand U10483 (N_10483,N_9601,N_9278);
or U10484 (N_10484,N_9319,N_9645);
and U10485 (N_10485,N_9413,N_9402);
xor U10486 (N_10486,N_9568,N_9477);
nor U10487 (N_10487,N_9494,N_9518);
or U10488 (N_10488,N_9200,N_9132);
nor U10489 (N_10489,N_9647,N_9499);
or U10490 (N_10490,N_9327,N_9038);
nand U10491 (N_10491,N_9621,N_9057);
nand U10492 (N_10492,N_9749,N_9455);
nor U10493 (N_10493,N_9300,N_9175);
nand U10494 (N_10494,N_9376,N_9356);
xor U10495 (N_10495,N_9617,N_9696);
or U10496 (N_10496,N_9081,N_9033);
nand U10497 (N_10497,N_9410,N_9176);
and U10498 (N_10498,N_9011,N_9197);
nor U10499 (N_10499,N_9592,N_9572);
nand U10500 (N_10500,N_10205,N_10278);
nor U10501 (N_10501,N_10105,N_10144);
nand U10502 (N_10502,N_10159,N_10294);
nor U10503 (N_10503,N_10177,N_10235);
and U10504 (N_10504,N_9817,N_10348);
nor U10505 (N_10505,N_9779,N_10484);
nor U10506 (N_10506,N_10377,N_9838);
nand U10507 (N_10507,N_9768,N_10085);
or U10508 (N_10508,N_10417,N_10028);
xor U10509 (N_10509,N_10126,N_9769);
or U10510 (N_10510,N_10449,N_10232);
nor U10511 (N_10511,N_9765,N_10053);
and U10512 (N_10512,N_9940,N_10258);
or U10513 (N_10513,N_10179,N_10213);
or U10514 (N_10514,N_10451,N_9926);
xnor U10515 (N_10515,N_9952,N_9843);
and U10516 (N_10516,N_10151,N_9849);
or U10517 (N_10517,N_10009,N_9937);
or U10518 (N_10518,N_9785,N_10345);
nand U10519 (N_10519,N_10314,N_9879);
and U10520 (N_10520,N_10383,N_9798);
nand U10521 (N_10521,N_9840,N_9772);
nand U10522 (N_10522,N_9985,N_10471);
nor U10523 (N_10523,N_10243,N_10200);
or U10524 (N_10524,N_9869,N_9992);
or U10525 (N_10525,N_9999,N_9927);
nor U10526 (N_10526,N_10236,N_10171);
nand U10527 (N_10527,N_10251,N_10344);
nand U10528 (N_10528,N_10107,N_9880);
and U10529 (N_10529,N_10161,N_9812);
and U10530 (N_10530,N_9947,N_9872);
and U10531 (N_10531,N_10439,N_10296);
or U10532 (N_10532,N_9924,N_10066);
and U10533 (N_10533,N_10195,N_10096);
and U10534 (N_10534,N_10368,N_10190);
nand U10535 (N_10535,N_10478,N_10095);
and U10536 (N_10536,N_10413,N_10091);
xnor U10537 (N_10537,N_10142,N_10005);
nor U10538 (N_10538,N_9990,N_9891);
nand U10539 (N_10539,N_9784,N_10070);
or U10540 (N_10540,N_10396,N_10322);
or U10541 (N_10541,N_10412,N_9809);
and U10542 (N_10542,N_10360,N_10194);
or U10543 (N_10543,N_10046,N_10189);
and U10544 (N_10544,N_10361,N_10365);
nor U10545 (N_10545,N_10264,N_10160);
or U10546 (N_10546,N_10440,N_10332);
nand U10547 (N_10547,N_10485,N_9896);
and U10548 (N_10548,N_10188,N_9877);
nor U10549 (N_10549,N_9903,N_10068);
nor U10550 (N_10550,N_9839,N_9908);
nand U10551 (N_10551,N_10252,N_10434);
nand U10552 (N_10552,N_10473,N_10209);
xor U10553 (N_10553,N_9954,N_9808);
nand U10554 (N_10554,N_10287,N_9868);
nand U10555 (N_10555,N_10398,N_10409);
or U10556 (N_10556,N_10271,N_9942);
nand U10557 (N_10557,N_10386,N_10077);
and U10558 (N_10558,N_10459,N_10312);
nand U10559 (N_10559,N_10430,N_10115);
and U10560 (N_10560,N_10432,N_10134);
xnor U10561 (N_10561,N_10109,N_10220);
nor U10562 (N_10562,N_10221,N_9805);
nor U10563 (N_10563,N_9958,N_10491);
or U10564 (N_10564,N_9885,N_9864);
nor U10565 (N_10565,N_10114,N_9964);
nor U10566 (N_10566,N_10423,N_9807);
nor U10567 (N_10567,N_10438,N_10495);
nand U10568 (N_10568,N_10058,N_10355);
nand U10569 (N_10569,N_10364,N_10204);
and U10570 (N_10570,N_9874,N_10445);
nor U10571 (N_10571,N_10320,N_9944);
nand U10572 (N_10572,N_10101,N_10457);
nor U10573 (N_10573,N_10039,N_10162);
nand U10574 (N_10574,N_10133,N_9984);
nor U10575 (N_10575,N_9789,N_9901);
xnor U10576 (N_10576,N_9788,N_10152);
and U10577 (N_10577,N_10427,N_9821);
and U10578 (N_10578,N_10196,N_10444);
nand U10579 (N_10579,N_10489,N_10158);
xnor U10580 (N_10580,N_10167,N_10022);
nand U10581 (N_10581,N_9753,N_10197);
or U10582 (N_10582,N_10141,N_9887);
xor U10583 (N_10583,N_10276,N_10044);
or U10584 (N_10584,N_10388,N_10234);
or U10585 (N_10585,N_10352,N_10420);
nor U10586 (N_10586,N_9776,N_10029);
nor U10587 (N_10587,N_9801,N_10291);
xor U10588 (N_10588,N_10048,N_10443);
nand U10589 (N_10589,N_10260,N_9799);
and U10590 (N_10590,N_10326,N_10173);
xnor U10591 (N_10591,N_9888,N_10037);
nand U10592 (N_10592,N_10008,N_10049);
and U10593 (N_10593,N_9850,N_10230);
nor U10594 (N_10594,N_9794,N_10042);
nand U10595 (N_10595,N_10324,N_9921);
or U10596 (N_10596,N_10238,N_9906);
and U10597 (N_10597,N_10191,N_10001);
nand U10598 (N_10598,N_10273,N_10131);
nand U10599 (N_10599,N_10168,N_10269);
xnor U10600 (N_10600,N_9957,N_9848);
nand U10601 (N_10601,N_9894,N_10328);
and U10602 (N_10602,N_10429,N_10202);
and U10603 (N_10603,N_9963,N_9970);
nor U10604 (N_10604,N_9875,N_10498);
or U10605 (N_10605,N_10071,N_10309);
and U10606 (N_10606,N_9950,N_10392);
or U10607 (N_10607,N_9841,N_10353);
nand U10608 (N_10608,N_10004,N_10479);
and U10609 (N_10609,N_9866,N_10208);
or U10610 (N_10610,N_10362,N_9978);
nor U10611 (N_10611,N_9831,N_10482);
or U10612 (N_10612,N_10329,N_10062);
nor U10613 (N_10613,N_10032,N_9960);
nor U10614 (N_10614,N_9910,N_10100);
and U10615 (N_10615,N_10020,N_10285);
nor U10616 (N_10616,N_9777,N_10120);
or U10617 (N_10617,N_10448,N_10371);
and U10618 (N_10618,N_10033,N_10303);
xor U10619 (N_10619,N_10082,N_9827);
nand U10620 (N_10620,N_10358,N_9905);
or U10621 (N_10621,N_10246,N_9844);
or U10622 (N_10622,N_10336,N_10316);
and U10623 (N_10623,N_10376,N_9948);
and U10624 (N_10624,N_9792,N_10227);
nand U10625 (N_10625,N_10424,N_10415);
nand U10626 (N_10626,N_10452,N_9916);
nand U10627 (N_10627,N_10181,N_10472);
or U10628 (N_10628,N_10229,N_10405);
or U10629 (N_10629,N_9800,N_9969);
nor U10630 (N_10630,N_10488,N_9878);
nor U10631 (N_10631,N_10057,N_10119);
or U10632 (N_10632,N_10241,N_9846);
or U10633 (N_10633,N_10225,N_9857);
nand U10634 (N_10634,N_10040,N_10325);
nand U10635 (N_10635,N_9783,N_9802);
xor U10636 (N_10636,N_10043,N_10143);
nor U10637 (N_10637,N_10047,N_9778);
nand U10638 (N_10638,N_10006,N_9912);
or U10639 (N_10639,N_10308,N_10318);
nor U10640 (N_10640,N_10223,N_9833);
nor U10641 (N_10641,N_10447,N_10180);
nor U10642 (N_10642,N_9959,N_10468);
and U10643 (N_10643,N_10395,N_10099);
nand U10644 (N_10644,N_9949,N_10342);
and U10645 (N_10645,N_9980,N_10455);
xor U10646 (N_10646,N_10384,N_10450);
nand U10647 (N_10647,N_10215,N_9867);
and U10648 (N_10648,N_10261,N_10397);
and U10649 (N_10649,N_10127,N_10201);
or U10650 (N_10650,N_10274,N_10295);
nand U10651 (N_10651,N_10340,N_10497);
or U10652 (N_10652,N_9917,N_10380);
and U10653 (N_10653,N_9832,N_10017);
and U10654 (N_10654,N_10078,N_9972);
and U10655 (N_10655,N_10083,N_10061);
nand U10656 (N_10656,N_10321,N_10080);
or U10657 (N_10657,N_10074,N_10374);
or U10658 (N_10658,N_10060,N_10437);
nand U10659 (N_10659,N_10165,N_9935);
or U10660 (N_10660,N_10469,N_10277);
nor U10661 (N_10661,N_10351,N_10354);
nor U10662 (N_10662,N_10249,N_10012);
xor U10663 (N_10663,N_10418,N_10065);
xor U10664 (N_10664,N_9892,N_9813);
nor U10665 (N_10665,N_10301,N_10268);
nor U10666 (N_10666,N_10063,N_10297);
and U10667 (N_10667,N_10199,N_9781);
nor U10668 (N_10668,N_10050,N_9923);
nand U10669 (N_10669,N_9943,N_9767);
and U10670 (N_10670,N_10132,N_10406);
nand U10671 (N_10671,N_10334,N_9981);
and U10672 (N_10672,N_9967,N_10490);
and U10673 (N_10673,N_10094,N_10442);
nand U10674 (N_10674,N_10248,N_10300);
and U10675 (N_10675,N_10394,N_10129);
and U10676 (N_10676,N_10024,N_10462);
and U10677 (N_10677,N_10335,N_9899);
nand U10678 (N_10678,N_10346,N_10084);
nor U10679 (N_10679,N_10390,N_10319);
nor U10680 (N_10680,N_9824,N_9835);
nand U10681 (N_10681,N_9863,N_10186);
and U10682 (N_10682,N_10150,N_9876);
or U10683 (N_10683,N_10460,N_9871);
or U10684 (N_10684,N_10426,N_9818);
nor U10685 (N_10685,N_9830,N_9974);
or U10686 (N_10686,N_10370,N_10403);
nand U10687 (N_10687,N_10454,N_9902);
nand U10688 (N_10688,N_9825,N_10428);
or U10689 (N_10689,N_9847,N_10212);
nand U10690 (N_10690,N_10156,N_9815);
and U10691 (N_10691,N_9762,N_10292);
nor U10692 (N_10692,N_9962,N_10250);
nor U10693 (N_10693,N_9965,N_10014);
and U10694 (N_10694,N_9983,N_10128);
and U10695 (N_10695,N_9966,N_10140);
xnor U10696 (N_10696,N_10481,N_10339);
nand U10697 (N_10697,N_9856,N_10389);
or U10698 (N_10698,N_10216,N_9929);
xnor U10699 (N_10699,N_10494,N_10123);
nor U10700 (N_10700,N_10217,N_9811);
or U10701 (N_10701,N_9938,N_9911);
nor U10702 (N_10702,N_10337,N_9986);
or U10703 (N_10703,N_9975,N_10002);
or U10704 (N_10704,N_10456,N_9861);
and U10705 (N_10705,N_10496,N_10385);
and U10706 (N_10706,N_9837,N_10366);
xor U10707 (N_10707,N_10102,N_10486);
nand U10708 (N_10708,N_9836,N_9760);
nor U10709 (N_10709,N_9771,N_9754);
nor U10710 (N_10710,N_10372,N_10493);
nor U10711 (N_10711,N_9982,N_10193);
or U10712 (N_10712,N_9907,N_10175);
and U10713 (N_10713,N_9791,N_10011);
nor U10714 (N_10714,N_10356,N_10087);
xnor U10715 (N_10715,N_10419,N_9997);
and U10716 (N_10716,N_10067,N_10282);
nand U10717 (N_10717,N_10408,N_10147);
nor U10718 (N_10718,N_10476,N_10045);
and U10719 (N_10719,N_9763,N_9823);
and U10720 (N_10720,N_10214,N_10130);
or U10721 (N_10721,N_9774,N_10219);
or U10722 (N_10722,N_10313,N_9851);
nor U10723 (N_10723,N_10228,N_10453);
and U10724 (N_10724,N_10035,N_9826);
or U10725 (N_10725,N_10170,N_10184);
or U10726 (N_10726,N_10203,N_10064);
nand U10727 (N_10727,N_10155,N_10375);
xnor U10728 (N_10728,N_9852,N_10436);
or U10729 (N_10729,N_10373,N_9855);
or U10730 (N_10730,N_10330,N_10266);
and U10731 (N_10731,N_10183,N_10010);
or U10732 (N_10732,N_9803,N_10139);
nand U10733 (N_10733,N_9820,N_10174);
nand U10734 (N_10734,N_10108,N_10092);
and U10735 (N_10735,N_9883,N_10247);
nand U10736 (N_10736,N_10369,N_10036);
and U10737 (N_10737,N_9936,N_9755);
xor U10738 (N_10738,N_9932,N_10027);
or U10739 (N_10739,N_9764,N_10347);
xnor U10740 (N_10740,N_10079,N_10145);
nor U10741 (N_10741,N_10000,N_9773);
nor U10742 (N_10742,N_10149,N_10304);
or U10743 (N_10743,N_10007,N_10331);
and U10744 (N_10744,N_10477,N_9928);
nand U10745 (N_10745,N_10237,N_10192);
nand U10746 (N_10746,N_10317,N_10272);
nand U10747 (N_10747,N_10176,N_10410);
xnor U10748 (N_10748,N_10016,N_10302);
nor U10749 (N_10749,N_10441,N_10379);
nor U10750 (N_10750,N_9858,N_9787);
or U10751 (N_10751,N_10465,N_10431);
nand U10752 (N_10752,N_10466,N_9961);
nand U10753 (N_10753,N_9918,N_9895);
nor U10754 (N_10754,N_10169,N_10135);
or U10755 (N_10755,N_10148,N_10030);
nand U10756 (N_10756,N_10224,N_10402);
and U10757 (N_10757,N_10433,N_10327);
nor U10758 (N_10758,N_9786,N_9925);
nor U10759 (N_10759,N_10172,N_9909);
or U10760 (N_10760,N_10088,N_10233);
xnor U10761 (N_10761,N_10111,N_10343);
nand U10762 (N_10762,N_10122,N_10298);
or U10763 (N_10763,N_10367,N_9761);
nand U10764 (N_10764,N_9989,N_9759);
or U10765 (N_10765,N_10023,N_10019);
nand U10766 (N_10766,N_10182,N_9976);
and U10767 (N_10767,N_10178,N_10113);
or U10768 (N_10768,N_9904,N_10422);
nand U10769 (N_10769,N_10106,N_10446);
nand U10770 (N_10770,N_10210,N_10401);
nor U10771 (N_10771,N_9893,N_9933);
nor U10772 (N_10772,N_9956,N_9987);
or U10773 (N_10773,N_10306,N_10474);
nand U10774 (N_10774,N_9915,N_10110);
and U10775 (N_10775,N_10055,N_9993);
nor U10776 (N_10776,N_10041,N_9797);
xor U10777 (N_10777,N_10255,N_9971);
xnor U10778 (N_10778,N_9750,N_10254);
nor U10779 (N_10779,N_10279,N_9816);
nand U10780 (N_10780,N_10359,N_10015);
nor U10781 (N_10781,N_9941,N_10026);
and U10782 (N_10782,N_10121,N_9920);
nor U10783 (N_10783,N_10499,N_10226);
and U10784 (N_10784,N_10052,N_10307);
and U10785 (N_10785,N_9930,N_9790);
nand U10786 (N_10786,N_9860,N_9810);
xor U10787 (N_10787,N_10073,N_9796);
xor U10788 (N_10788,N_10054,N_10137);
nand U10789 (N_10789,N_10104,N_9853);
and U10790 (N_10790,N_10117,N_10076);
and U10791 (N_10791,N_9806,N_10198);
nor U10792 (N_10792,N_10378,N_10283);
and U10793 (N_10793,N_10086,N_10245);
or U10794 (N_10794,N_10414,N_10393);
and U10795 (N_10795,N_9919,N_10310);
nor U10796 (N_10796,N_10492,N_9994);
nand U10797 (N_10797,N_10341,N_10265);
or U10798 (N_10798,N_10338,N_9758);
nor U10799 (N_10799,N_9991,N_9782);
and U10800 (N_10800,N_9898,N_9854);
or U10801 (N_10801,N_10480,N_10425);
nor U10802 (N_10802,N_9819,N_9890);
and U10803 (N_10803,N_10146,N_9834);
nand U10804 (N_10804,N_10464,N_10242);
nand U10805 (N_10805,N_10289,N_9793);
nor U10806 (N_10806,N_10103,N_10034);
nand U10807 (N_10807,N_9889,N_10185);
or U10808 (N_10808,N_10038,N_9955);
or U10809 (N_10809,N_9795,N_9996);
or U10810 (N_10810,N_9751,N_10069);
or U10811 (N_10811,N_10267,N_9934);
nand U10812 (N_10812,N_10299,N_10125);
nor U10813 (N_10813,N_10056,N_10239);
and U10814 (N_10814,N_10421,N_9914);
nand U10815 (N_10815,N_10013,N_10458);
or U10816 (N_10816,N_9931,N_9953);
or U10817 (N_10817,N_9951,N_9939);
nor U10818 (N_10818,N_10311,N_9922);
nor U10819 (N_10819,N_10098,N_9973);
nand U10820 (N_10820,N_10118,N_10270);
nand U10821 (N_10821,N_10089,N_10259);
nor U10822 (N_10822,N_9886,N_9766);
nor U10823 (N_10823,N_9913,N_10124);
nor U10824 (N_10824,N_10263,N_10470);
or U10825 (N_10825,N_10157,N_9998);
or U10826 (N_10826,N_10404,N_10240);
nand U10827 (N_10827,N_10059,N_10483);
and U10828 (N_10828,N_10391,N_10323);
nand U10829 (N_10829,N_10093,N_9752);
nor U10830 (N_10830,N_10387,N_9829);
nand U10831 (N_10831,N_10075,N_9828);
nor U10832 (N_10832,N_10275,N_9945);
and U10833 (N_10833,N_10218,N_10051);
nand U10834 (N_10834,N_10435,N_10333);
xnor U10835 (N_10835,N_10257,N_9900);
xnor U10836 (N_10836,N_9884,N_9881);
or U10837 (N_10837,N_10411,N_9865);
or U10838 (N_10838,N_10138,N_10284);
xor U10839 (N_10839,N_10280,N_10382);
and U10840 (N_10840,N_10072,N_10305);
and U10841 (N_10841,N_10349,N_10136);
or U10842 (N_10842,N_10407,N_10262);
or U10843 (N_10843,N_10281,N_10211);
or U10844 (N_10844,N_9988,N_9946);
nor U10845 (N_10845,N_10467,N_10315);
and U10846 (N_10846,N_10461,N_10222);
nor U10847 (N_10847,N_9842,N_10416);
or U10848 (N_10848,N_10164,N_9814);
and U10849 (N_10849,N_10097,N_10154);
and U10850 (N_10850,N_9757,N_10399);
and U10851 (N_10851,N_10350,N_10025);
nand U10852 (N_10852,N_10381,N_10400);
nand U10853 (N_10853,N_10163,N_9775);
or U10854 (N_10854,N_9770,N_9979);
nor U10855 (N_10855,N_9882,N_10018);
and U10856 (N_10856,N_9862,N_9756);
nor U10857 (N_10857,N_9859,N_9977);
nor U10858 (N_10858,N_10231,N_10363);
nand U10859 (N_10859,N_10153,N_10286);
xor U10860 (N_10860,N_10206,N_9995);
and U10861 (N_10861,N_10116,N_10207);
and U10862 (N_10862,N_10081,N_10112);
and U10863 (N_10863,N_10166,N_10487);
nor U10864 (N_10864,N_9897,N_10187);
nor U10865 (N_10865,N_9822,N_9873);
nand U10866 (N_10866,N_10244,N_10003);
and U10867 (N_10867,N_9804,N_10288);
nand U10868 (N_10868,N_9845,N_10256);
nand U10869 (N_10869,N_10463,N_9780);
nand U10870 (N_10870,N_10293,N_10021);
nor U10871 (N_10871,N_10031,N_10253);
and U10872 (N_10872,N_10290,N_10090);
or U10873 (N_10873,N_9968,N_10475);
and U10874 (N_10874,N_9870,N_10357);
nor U10875 (N_10875,N_9889,N_9793);
or U10876 (N_10876,N_10133,N_10477);
and U10877 (N_10877,N_10208,N_10286);
and U10878 (N_10878,N_10347,N_9773);
or U10879 (N_10879,N_10466,N_9940);
nor U10880 (N_10880,N_10155,N_10127);
nand U10881 (N_10881,N_10222,N_10345);
nand U10882 (N_10882,N_10322,N_10405);
and U10883 (N_10883,N_10075,N_9920);
or U10884 (N_10884,N_10156,N_9957);
and U10885 (N_10885,N_9766,N_9798);
nor U10886 (N_10886,N_9947,N_10086);
xnor U10887 (N_10887,N_10361,N_10096);
xnor U10888 (N_10888,N_10270,N_10267);
xor U10889 (N_10889,N_10165,N_10166);
nor U10890 (N_10890,N_10142,N_10216);
nor U10891 (N_10891,N_10228,N_9993);
and U10892 (N_10892,N_10455,N_9984);
nor U10893 (N_10893,N_10466,N_10036);
xor U10894 (N_10894,N_10049,N_10323);
nand U10895 (N_10895,N_10324,N_10412);
nand U10896 (N_10896,N_10234,N_10082);
nor U10897 (N_10897,N_9857,N_10258);
nor U10898 (N_10898,N_9944,N_10152);
and U10899 (N_10899,N_10475,N_9824);
or U10900 (N_10900,N_10035,N_10060);
nand U10901 (N_10901,N_10194,N_9909);
or U10902 (N_10902,N_10419,N_10452);
or U10903 (N_10903,N_10205,N_9923);
and U10904 (N_10904,N_9968,N_10309);
or U10905 (N_10905,N_10082,N_10038);
nor U10906 (N_10906,N_9892,N_10484);
and U10907 (N_10907,N_10312,N_9860);
nor U10908 (N_10908,N_9781,N_10019);
xnor U10909 (N_10909,N_10481,N_9779);
and U10910 (N_10910,N_10019,N_10436);
or U10911 (N_10911,N_9923,N_10094);
xor U10912 (N_10912,N_10295,N_10363);
or U10913 (N_10913,N_10351,N_10410);
or U10914 (N_10914,N_9813,N_9967);
and U10915 (N_10915,N_10448,N_10374);
or U10916 (N_10916,N_10236,N_10487);
and U10917 (N_10917,N_10451,N_10498);
nor U10918 (N_10918,N_10335,N_10455);
nor U10919 (N_10919,N_10285,N_10174);
nor U10920 (N_10920,N_10415,N_9966);
and U10921 (N_10921,N_10321,N_10448);
and U10922 (N_10922,N_9947,N_10050);
nand U10923 (N_10923,N_9790,N_10049);
nor U10924 (N_10924,N_10063,N_10080);
nand U10925 (N_10925,N_10115,N_10495);
nand U10926 (N_10926,N_10126,N_9985);
nor U10927 (N_10927,N_10497,N_10217);
or U10928 (N_10928,N_9854,N_10266);
nand U10929 (N_10929,N_9860,N_9981);
nor U10930 (N_10930,N_10107,N_9938);
or U10931 (N_10931,N_10220,N_10406);
or U10932 (N_10932,N_9957,N_9760);
nand U10933 (N_10933,N_10158,N_9874);
nor U10934 (N_10934,N_10309,N_9929);
nor U10935 (N_10935,N_10205,N_9898);
xnor U10936 (N_10936,N_9931,N_9865);
xnor U10937 (N_10937,N_10205,N_10294);
nor U10938 (N_10938,N_10139,N_10477);
nand U10939 (N_10939,N_10435,N_9911);
and U10940 (N_10940,N_10215,N_10163);
nand U10941 (N_10941,N_10002,N_10383);
nand U10942 (N_10942,N_10393,N_9854);
and U10943 (N_10943,N_9947,N_9876);
or U10944 (N_10944,N_10022,N_9938);
and U10945 (N_10945,N_9763,N_10128);
and U10946 (N_10946,N_10348,N_10168);
nand U10947 (N_10947,N_10453,N_10398);
nor U10948 (N_10948,N_10283,N_9992);
nand U10949 (N_10949,N_9967,N_10046);
nand U10950 (N_10950,N_9997,N_10090);
and U10951 (N_10951,N_9934,N_10481);
nand U10952 (N_10952,N_10052,N_9921);
xnor U10953 (N_10953,N_10444,N_10080);
nor U10954 (N_10954,N_10195,N_10050);
or U10955 (N_10955,N_10062,N_10375);
nor U10956 (N_10956,N_9799,N_10224);
xor U10957 (N_10957,N_10013,N_10496);
and U10958 (N_10958,N_9861,N_10344);
nand U10959 (N_10959,N_10359,N_10000);
xor U10960 (N_10960,N_10113,N_10182);
or U10961 (N_10961,N_10458,N_10288);
xor U10962 (N_10962,N_10277,N_9759);
nand U10963 (N_10963,N_10167,N_10421);
or U10964 (N_10964,N_9841,N_10490);
nor U10965 (N_10965,N_10280,N_9921);
and U10966 (N_10966,N_10243,N_9762);
or U10967 (N_10967,N_10272,N_10187);
or U10968 (N_10968,N_10255,N_10037);
and U10969 (N_10969,N_10000,N_10353);
nand U10970 (N_10970,N_10309,N_10453);
nor U10971 (N_10971,N_10080,N_9989);
nand U10972 (N_10972,N_9940,N_10447);
nand U10973 (N_10973,N_10487,N_9791);
and U10974 (N_10974,N_10148,N_10032);
and U10975 (N_10975,N_9902,N_10163);
nand U10976 (N_10976,N_10088,N_10122);
or U10977 (N_10977,N_9840,N_10185);
or U10978 (N_10978,N_10189,N_9903);
xor U10979 (N_10979,N_10218,N_10003);
nor U10980 (N_10980,N_9891,N_9964);
nand U10981 (N_10981,N_9802,N_9807);
or U10982 (N_10982,N_10268,N_10488);
and U10983 (N_10983,N_10153,N_9838);
and U10984 (N_10984,N_10142,N_9836);
nand U10985 (N_10985,N_10153,N_10287);
or U10986 (N_10986,N_10188,N_10481);
nand U10987 (N_10987,N_9918,N_10017);
nand U10988 (N_10988,N_9840,N_10081);
or U10989 (N_10989,N_10117,N_9753);
xnor U10990 (N_10990,N_9925,N_9928);
xnor U10991 (N_10991,N_10353,N_10215);
and U10992 (N_10992,N_9943,N_10208);
or U10993 (N_10993,N_10468,N_9851);
or U10994 (N_10994,N_10049,N_10100);
nor U10995 (N_10995,N_10264,N_10097);
nand U10996 (N_10996,N_10346,N_9826);
or U10997 (N_10997,N_9887,N_9933);
nor U10998 (N_10998,N_10120,N_10426);
or U10999 (N_10999,N_10222,N_9939);
or U11000 (N_11000,N_10323,N_10091);
xor U11001 (N_11001,N_9890,N_10084);
and U11002 (N_11002,N_10070,N_10432);
nand U11003 (N_11003,N_9775,N_9956);
nand U11004 (N_11004,N_10495,N_10009);
and U11005 (N_11005,N_10192,N_10194);
nor U11006 (N_11006,N_10478,N_10456);
xor U11007 (N_11007,N_10368,N_9751);
nor U11008 (N_11008,N_10056,N_9974);
nand U11009 (N_11009,N_10319,N_9828);
nand U11010 (N_11010,N_10096,N_9800);
xnor U11011 (N_11011,N_10225,N_9822);
xor U11012 (N_11012,N_10326,N_10137);
nand U11013 (N_11013,N_9758,N_10116);
nand U11014 (N_11014,N_10202,N_10406);
or U11015 (N_11015,N_10213,N_10440);
nor U11016 (N_11016,N_10329,N_9851);
xor U11017 (N_11017,N_10266,N_9784);
nand U11018 (N_11018,N_10359,N_9861);
and U11019 (N_11019,N_10133,N_10462);
and U11020 (N_11020,N_10286,N_10023);
or U11021 (N_11021,N_10308,N_9756);
nand U11022 (N_11022,N_10272,N_10111);
xor U11023 (N_11023,N_10244,N_9972);
or U11024 (N_11024,N_9781,N_10302);
and U11025 (N_11025,N_9792,N_10013);
nand U11026 (N_11026,N_10176,N_10306);
nor U11027 (N_11027,N_9839,N_10225);
nand U11028 (N_11028,N_9756,N_10246);
nor U11029 (N_11029,N_9773,N_9966);
nor U11030 (N_11030,N_9991,N_10122);
nand U11031 (N_11031,N_10040,N_10450);
nor U11032 (N_11032,N_10260,N_10254);
and U11033 (N_11033,N_10454,N_9910);
nand U11034 (N_11034,N_10116,N_10353);
nand U11035 (N_11035,N_10074,N_10433);
nand U11036 (N_11036,N_9837,N_9988);
nand U11037 (N_11037,N_10239,N_10271);
and U11038 (N_11038,N_10337,N_10282);
or U11039 (N_11039,N_10186,N_9788);
or U11040 (N_11040,N_10125,N_10234);
and U11041 (N_11041,N_10019,N_9985);
or U11042 (N_11042,N_10047,N_10077);
nor U11043 (N_11043,N_9952,N_10320);
nor U11044 (N_11044,N_9805,N_9807);
and U11045 (N_11045,N_10098,N_9759);
and U11046 (N_11046,N_10452,N_9850);
or U11047 (N_11047,N_10081,N_10411);
nor U11048 (N_11048,N_10058,N_10408);
nor U11049 (N_11049,N_10097,N_9781);
and U11050 (N_11050,N_9910,N_10083);
and U11051 (N_11051,N_9884,N_10134);
or U11052 (N_11052,N_9865,N_9756);
xor U11053 (N_11053,N_10303,N_10148);
or U11054 (N_11054,N_9913,N_9908);
or U11055 (N_11055,N_10303,N_10302);
nand U11056 (N_11056,N_10355,N_10199);
and U11057 (N_11057,N_10037,N_9809);
and U11058 (N_11058,N_9853,N_10299);
or U11059 (N_11059,N_9752,N_9879);
or U11060 (N_11060,N_9935,N_9980);
nor U11061 (N_11061,N_9805,N_10344);
nand U11062 (N_11062,N_9789,N_9770);
nor U11063 (N_11063,N_9967,N_9793);
or U11064 (N_11064,N_9773,N_10375);
nand U11065 (N_11065,N_9865,N_10231);
nand U11066 (N_11066,N_9936,N_10377);
nand U11067 (N_11067,N_10465,N_10194);
and U11068 (N_11068,N_10133,N_9966);
nor U11069 (N_11069,N_10044,N_10266);
nand U11070 (N_11070,N_10062,N_10344);
nand U11071 (N_11071,N_9954,N_10092);
or U11072 (N_11072,N_10197,N_9770);
nand U11073 (N_11073,N_9931,N_10472);
nand U11074 (N_11074,N_10002,N_10305);
and U11075 (N_11075,N_9833,N_10004);
or U11076 (N_11076,N_10161,N_10018);
or U11077 (N_11077,N_10049,N_9787);
or U11078 (N_11078,N_10433,N_10369);
and U11079 (N_11079,N_9775,N_10443);
nor U11080 (N_11080,N_9842,N_10286);
nor U11081 (N_11081,N_10048,N_9789);
nor U11082 (N_11082,N_10262,N_9806);
or U11083 (N_11083,N_10274,N_9803);
or U11084 (N_11084,N_10126,N_9819);
nand U11085 (N_11085,N_10495,N_10428);
nor U11086 (N_11086,N_10089,N_10314);
nor U11087 (N_11087,N_10014,N_9779);
and U11088 (N_11088,N_10471,N_10490);
nand U11089 (N_11089,N_9840,N_10102);
nand U11090 (N_11090,N_10230,N_9890);
nor U11091 (N_11091,N_10388,N_10204);
and U11092 (N_11092,N_10051,N_10124);
or U11093 (N_11093,N_10137,N_10095);
xor U11094 (N_11094,N_10084,N_10310);
nor U11095 (N_11095,N_10340,N_9930);
xor U11096 (N_11096,N_10033,N_10030);
or U11097 (N_11097,N_9985,N_9837);
and U11098 (N_11098,N_9804,N_9960);
nand U11099 (N_11099,N_9933,N_10206);
nand U11100 (N_11100,N_9776,N_10335);
and U11101 (N_11101,N_10059,N_10157);
xor U11102 (N_11102,N_9870,N_9948);
or U11103 (N_11103,N_10020,N_10425);
and U11104 (N_11104,N_9853,N_9803);
and U11105 (N_11105,N_10475,N_10312);
and U11106 (N_11106,N_10365,N_9989);
or U11107 (N_11107,N_10484,N_9989);
nor U11108 (N_11108,N_9853,N_9962);
nor U11109 (N_11109,N_10172,N_10299);
or U11110 (N_11110,N_10204,N_9902);
nor U11111 (N_11111,N_10274,N_10112);
or U11112 (N_11112,N_10334,N_10415);
or U11113 (N_11113,N_10114,N_10459);
or U11114 (N_11114,N_10389,N_10258);
nor U11115 (N_11115,N_10384,N_10345);
xor U11116 (N_11116,N_9806,N_9830);
nand U11117 (N_11117,N_10149,N_10323);
nor U11118 (N_11118,N_9887,N_10488);
or U11119 (N_11119,N_10212,N_9853);
xor U11120 (N_11120,N_10130,N_10354);
nand U11121 (N_11121,N_10314,N_10452);
xnor U11122 (N_11122,N_9875,N_10414);
nor U11123 (N_11123,N_9901,N_10205);
nand U11124 (N_11124,N_10432,N_10485);
or U11125 (N_11125,N_10057,N_10180);
and U11126 (N_11126,N_10464,N_10309);
or U11127 (N_11127,N_10459,N_9851);
and U11128 (N_11128,N_10225,N_10160);
nor U11129 (N_11129,N_9944,N_10148);
nor U11130 (N_11130,N_9885,N_10200);
nor U11131 (N_11131,N_10412,N_10462);
or U11132 (N_11132,N_10473,N_10001);
nand U11133 (N_11133,N_9882,N_10324);
nand U11134 (N_11134,N_9924,N_10303);
nor U11135 (N_11135,N_10048,N_9908);
or U11136 (N_11136,N_9909,N_10085);
or U11137 (N_11137,N_9828,N_10137);
nor U11138 (N_11138,N_10150,N_10226);
xor U11139 (N_11139,N_10301,N_10125);
or U11140 (N_11140,N_10328,N_10073);
nand U11141 (N_11141,N_9965,N_9898);
or U11142 (N_11142,N_9800,N_10040);
and U11143 (N_11143,N_10320,N_10007);
nor U11144 (N_11144,N_9752,N_9903);
or U11145 (N_11145,N_10234,N_9876);
nor U11146 (N_11146,N_10016,N_9800);
and U11147 (N_11147,N_10188,N_10382);
and U11148 (N_11148,N_10339,N_9795);
nand U11149 (N_11149,N_10280,N_9839);
or U11150 (N_11150,N_10306,N_10295);
and U11151 (N_11151,N_10425,N_10470);
nand U11152 (N_11152,N_10069,N_10398);
and U11153 (N_11153,N_10139,N_10138);
and U11154 (N_11154,N_10136,N_10235);
and U11155 (N_11155,N_10069,N_10156);
xor U11156 (N_11156,N_10465,N_9789);
nand U11157 (N_11157,N_10431,N_9918);
nor U11158 (N_11158,N_9839,N_10076);
nor U11159 (N_11159,N_10422,N_10131);
nor U11160 (N_11160,N_10094,N_9881);
or U11161 (N_11161,N_10263,N_10173);
or U11162 (N_11162,N_10478,N_10299);
or U11163 (N_11163,N_9917,N_9766);
nand U11164 (N_11164,N_9784,N_10363);
and U11165 (N_11165,N_10366,N_10119);
nor U11166 (N_11166,N_9754,N_10427);
or U11167 (N_11167,N_9767,N_10351);
or U11168 (N_11168,N_10408,N_10364);
nor U11169 (N_11169,N_10245,N_10217);
and U11170 (N_11170,N_10220,N_10056);
or U11171 (N_11171,N_10193,N_9873);
nand U11172 (N_11172,N_9974,N_10437);
xor U11173 (N_11173,N_9886,N_9773);
or U11174 (N_11174,N_10402,N_10257);
nor U11175 (N_11175,N_10011,N_9917);
nand U11176 (N_11176,N_10287,N_10279);
and U11177 (N_11177,N_10496,N_10405);
and U11178 (N_11178,N_9853,N_9987);
and U11179 (N_11179,N_10185,N_9878);
nand U11180 (N_11180,N_9999,N_10325);
nor U11181 (N_11181,N_10446,N_10121);
nor U11182 (N_11182,N_10383,N_10448);
nand U11183 (N_11183,N_10235,N_9879);
or U11184 (N_11184,N_10291,N_10301);
nand U11185 (N_11185,N_9990,N_9788);
and U11186 (N_11186,N_10489,N_10241);
and U11187 (N_11187,N_10272,N_10487);
nand U11188 (N_11188,N_10371,N_9943);
and U11189 (N_11189,N_10194,N_10027);
nor U11190 (N_11190,N_10347,N_10343);
nor U11191 (N_11191,N_10473,N_10372);
nor U11192 (N_11192,N_10360,N_10175);
or U11193 (N_11193,N_10139,N_10416);
and U11194 (N_11194,N_9900,N_10363);
and U11195 (N_11195,N_10198,N_10019);
nand U11196 (N_11196,N_9792,N_10065);
nand U11197 (N_11197,N_10099,N_10205);
nand U11198 (N_11198,N_9922,N_9765);
and U11199 (N_11199,N_9953,N_9783);
or U11200 (N_11200,N_9852,N_10135);
or U11201 (N_11201,N_10337,N_9765);
and U11202 (N_11202,N_9880,N_10012);
or U11203 (N_11203,N_10230,N_9948);
and U11204 (N_11204,N_10221,N_10179);
or U11205 (N_11205,N_9877,N_9784);
nand U11206 (N_11206,N_10254,N_10270);
nand U11207 (N_11207,N_10150,N_10085);
nand U11208 (N_11208,N_10300,N_10148);
xor U11209 (N_11209,N_10453,N_10444);
nand U11210 (N_11210,N_10347,N_10309);
nand U11211 (N_11211,N_10450,N_10349);
or U11212 (N_11212,N_10035,N_9954);
nor U11213 (N_11213,N_10406,N_10407);
or U11214 (N_11214,N_9980,N_10497);
or U11215 (N_11215,N_9988,N_10139);
and U11216 (N_11216,N_9866,N_9923);
nor U11217 (N_11217,N_10401,N_10267);
and U11218 (N_11218,N_9894,N_9960);
and U11219 (N_11219,N_10483,N_9873);
nand U11220 (N_11220,N_9754,N_9988);
xnor U11221 (N_11221,N_10228,N_10122);
nor U11222 (N_11222,N_9901,N_10160);
nor U11223 (N_11223,N_10024,N_9776);
and U11224 (N_11224,N_10285,N_10370);
and U11225 (N_11225,N_9925,N_10092);
or U11226 (N_11226,N_10199,N_10221);
nor U11227 (N_11227,N_10065,N_10468);
or U11228 (N_11228,N_10291,N_10244);
nand U11229 (N_11229,N_10390,N_10191);
nand U11230 (N_11230,N_10121,N_9791);
nor U11231 (N_11231,N_10069,N_10260);
nor U11232 (N_11232,N_10443,N_10152);
and U11233 (N_11233,N_10014,N_10485);
and U11234 (N_11234,N_10059,N_10046);
nand U11235 (N_11235,N_10382,N_10215);
or U11236 (N_11236,N_10408,N_9999);
or U11237 (N_11237,N_10109,N_9978);
or U11238 (N_11238,N_9862,N_10388);
or U11239 (N_11239,N_10253,N_10387);
nor U11240 (N_11240,N_10064,N_9980);
and U11241 (N_11241,N_9835,N_10140);
nor U11242 (N_11242,N_10200,N_9952);
nand U11243 (N_11243,N_10428,N_10195);
and U11244 (N_11244,N_9771,N_10188);
and U11245 (N_11245,N_10307,N_9816);
and U11246 (N_11246,N_10008,N_10170);
nor U11247 (N_11247,N_10409,N_10379);
or U11248 (N_11248,N_9856,N_10112);
nor U11249 (N_11249,N_9952,N_9953);
and U11250 (N_11250,N_10767,N_10626);
nand U11251 (N_11251,N_10682,N_11082);
nand U11252 (N_11252,N_10867,N_10727);
and U11253 (N_11253,N_10689,N_10528);
nand U11254 (N_11254,N_11247,N_10893);
and U11255 (N_11255,N_10668,N_10806);
nor U11256 (N_11256,N_10914,N_10765);
nor U11257 (N_11257,N_10809,N_10699);
nand U11258 (N_11258,N_10812,N_10583);
and U11259 (N_11259,N_10625,N_11199);
and U11260 (N_11260,N_10850,N_10522);
and U11261 (N_11261,N_10684,N_11213);
nor U11262 (N_11262,N_10779,N_10603);
and U11263 (N_11263,N_11016,N_11165);
nor U11264 (N_11264,N_10995,N_11019);
or U11265 (N_11265,N_11054,N_11201);
and U11266 (N_11266,N_10550,N_10660);
and U11267 (N_11267,N_11242,N_11109);
and U11268 (N_11268,N_10553,N_11227);
nand U11269 (N_11269,N_11230,N_11013);
or U11270 (N_11270,N_10944,N_10665);
or U11271 (N_11271,N_11212,N_11145);
and U11272 (N_11272,N_11080,N_11192);
nor U11273 (N_11273,N_10957,N_10711);
nand U11274 (N_11274,N_11166,N_11138);
nand U11275 (N_11275,N_10904,N_11141);
and U11276 (N_11276,N_10916,N_11134);
xnor U11277 (N_11277,N_11170,N_11036);
nand U11278 (N_11278,N_10956,N_10620);
and U11279 (N_11279,N_10892,N_10577);
nand U11280 (N_11280,N_11030,N_10718);
nand U11281 (N_11281,N_11221,N_10931);
nor U11282 (N_11282,N_10630,N_10647);
or U11283 (N_11283,N_11225,N_10876);
nand U11284 (N_11284,N_10961,N_10586);
nand U11285 (N_11285,N_10955,N_10905);
and U11286 (N_11286,N_10936,N_10939);
xnor U11287 (N_11287,N_11053,N_10749);
nor U11288 (N_11288,N_10729,N_10519);
and U11289 (N_11289,N_11209,N_10774);
nand U11290 (N_11290,N_10742,N_10617);
xnor U11291 (N_11291,N_10835,N_10960);
nor U11292 (N_11292,N_10591,N_10544);
and U11293 (N_11293,N_10785,N_10612);
nor U11294 (N_11294,N_10534,N_11083);
nand U11295 (N_11295,N_10561,N_10751);
nand U11296 (N_11296,N_11150,N_10648);
or U11297 (N_11297,N_10636,N_10821);
or U11298 (N_11298,N_11190,N_11071);
or U11299 (N_11299,N_11245,N_11137);
or U11300 (N_11300,N_10856,N_10540);
xnor U11301 (N_11301,N_10815,N_10737);
and U11302 (N_11302,N_11124,N_11087);
and U11303 (N_11303,N_10752,N_10747);
xnor U11304 (N_11304,N_11122,N_10997);
nor U11305 (N_11305,N_11184,N_10641);
and U11306 (N_11306,N_10686,N_10644);
nor U11307 (N_11307,N_10924,N_10607);
nand U11308 (N_11308,N_11248,N_11179);
nor U11309 (N_11309,N_10590,N_10780);
nor U11310 (N_11310,N_10643,N_11154);
and U11311 (N_11311,N_10870,N_10721);
nand U11312 (N_11312,N_10977,N_11215);
or U11313 (N_11313,N_10839,N_11157);
and U11314 (N_11314,N_10842,N_10825);
nand U11315 (N_11315,N_10670,N_10706);
or U11316 (N_11316,N_10954,N_11066);
and U11317 (N_11317,N_11226,N_10831);
xnor U11318 (N_11318,N_10989,N_10871);
nor U11319 (N_11319,N_10868,N_10802);
and U11320 (N_11320,N_10570,N_11081);
or U11321 (N_11321,N_11140,N_11188);
nand U11322 (N_11322,N_10862,N_10609);
or U11323 (N_11323,N_10857,N_10589);
nor U11324 (N_11324,N_11173,N_10613);
nor U11325 (N_11325,N_10504,N_11094);
nor U11326 (N_11326,N_11048,N_11149);
nand U11327 (N_11327,N_10773,N_10698);
or U11328 (N_11328,N_10704,N_11146);
and U11329 (N_11329,N_10677,N_10808);
nand U11330 (N_11330,N_10959,N_11067);
and U11331 (N_11331,N_10853,N_10517);
and U11332 (N_11332,N_10801,N_10552);
nor U11333 (N_11333,N_10642,N_10674);
xnor U11334 (N_11334,N_10770,N_10678);
nor U11335 (N_11335,N_10880,N_10716);
or U11336 (N_11336,N_10820,N_10837);
or U11337 (N_11337,N_11040,N_10524);
and U11338 (N_11338,N_11131,N_10750);
and U11339 (N_11339,N_10503,N_10757);
nand U11340 (N_11340,N_10788,N_11194);
and U11341 (N_11341,N_10685,N_10592);
or U11342 (N_11342,N_10941,N_11107);
nand U11343 (N_11343,N_10818,N_10882);
nand U11344 (N_11344,N_10762,N_11203);
nand U11345 (N_11345,N_10881,N_10703);
nor U11346 (N_11346,N_10823,N_10624);
nand U11347 (N_11347,N_10666,N_11023);
and U11348 (N_11348,N_11235,N_10824);
or U11349 (N_11349,N_11180,N_11161);
xor U11350 (N_11350,N_10659,N_11085);
nand U11351 (N_11351,N_11207,N_11043);
nand U11352 (N_11352,N_10580,N_10611);
or U11353 (N_11353,N_10877,N_10778);
and U11354 (N_11354,N_10845,N_10994);
and U11355 (N_11355,N_11114,N_10861);
nand U11356 (N_11356,N_10556,N_10826);
nand U11357 (N_11357,N_10731,N_10595);
and U11358 (N_11358,N_10707,N_10947);
nand U11359 (N_11359,N_10664,N_11042);
nor U11360 (N_11360,N_10964,N_10967);
xnor U11361 (N_11361,N_10972,N_10799);
nor U11362 (N_11362,N_11202,N_10629);
nand U11363 (N_11363,N_10653,N_11090);
nor U11364 (N_11364,N_10657,N_10724);
nand U11365 (N_11365,N_11055,N_10650);
nor U11366 (N_11366,N_11063,N_10649);
or U11367 (N_11367,N_10593,N_10579);
or U11368 (N_11368,N_10847,N_11132);
and U11369 (N_11369,N_10658,N_11151);
nand U11370 (N_11370,N_11001,N_11177);
or U11371 (N_11371,N_10614,N_10511);
nand U11372 (N_11372,N_10569,N_10610);
and U11373 (N_11373,N_11125,N_10771);
nand U11374 (N_11374,N_10879,N_10776);
and U11375 (N_11375,N_10509,N_10973);
nor U11376 (N_11376,N_10542,N_10985);
nor U11377 (N_11377,N_10702,N_11162);
nand U11378 (N_11378,N_10891,N_11035);
or U11379 (N_11379,N_11110,N_10833);
and U11380 (N_11380,N_10661,N_11045);
nor U11381 (N_11381,N_11232,N_10797);
nor U11382 (N_11382,N_11115,N_10623);
nor U11383 (N_11383,N_11121,N_10622);
or U11384 (N_11384,N_11096,N_10740);
or U11385 (N_11385,N_10836,N_10547);
nor U11386 (N_11386,N_10598,N_10726);
nand U11387 (N_11387,N_11089,N_11017);
or U11388 (N_11388,N_11126,N_10537);
nand U11389 (N_11389,N_10638,N_10691);
and U11390 (N_11390,N_10717,N_11139);
nor U11391 (N_11391,N_10838,N_11156);
and U11392 (N_11392,N_11210,N_10874);
nand U11393 (N_11393,N_11214,N_10738);
and U11394 (N_11394,N_10912,N_10683);
nand U11395 (N_11395,N_11223,N_10849);
and U11396 (N_11396,N_10654,N_11093);
or U11397 (N_11397,N_10766,N_11116);
nand U11398 (N_11398,N_11075,N_10974);
nor U11399 (N_11399,N_10523,N_11022);
and U11400 (N_11400,N_10907,N_11041);
nand U11401 (N_11401,N_11051,N_10535);
xor U11402 (N_11402,N_11238,N_11174);
xnor U11403 (N_11403,N_11204,N_10712);
and U11404 (N_11404,N_10530,N_10777);
and U11405 (N_11405,N_11020,N_10890);
nand U11406 (N_11406,N_10633,N_11144);
and U11407 (N_11407,N_10886,N_10574);
or U11408 (N_11408,N_10969,N_10745);
or U11409 (N_11409,N_11185,N_10730);
nor U11410 (N_11410,N_10564,N_10898);
and U11411 (N_11411,N_10996,N_10507);
nand U11412 (N_11412,N_10631,N_11097);
or U11413 (N_11413,N_10988,N_11218);
nor U11414 (N_11414,N_10525,N_10562);
xor U11415 (N_11415,N_11102,N_10804);
and U11416 (N_11416,N_10915,N_11008);
and U11417 (N_11417,N_10667,N_11155);
or U11418 (N_11418,N_10896,N_11120);
or U11419 (N_11419,N_10656,N_11021);
xnor U11420 (N_11420,N_10950,N_11246);
nor U11421 (N_11421,N_10735,N_10560);
xnor U11422 (N_11422,N_10787,N_11148);
and U11423 (N_11423,N_11061,N_10546);
or U11424 (N_11424,N_10652,N_10758);
or U11425 (N_11425,N_10998,N_10906);
and U11426 (N_11426,N_10734,N_10908);
or U11427 (N_11427,N_10965,N_11182);
nand U11428 (N_11428,N_10987,N_11079);
nand U11429 (N_11429,N_11052,N_11072);
nor U11430 (N_11430,N_10575,N_10710);
nand U11431 (N_11431,N_11231,N_10596);
and U11432 (N_11432,N_10571,N_10536);
nor U11433 (N_11433,N_10621,N_10970);
or U11434 (N_11434,N_10810,N_11228);
nor U11435 (N_11435,N_10672,N_10584);
or U11436 (N_11436,N_10978,N_10843);
nand U11437 (N_11437,N_10655,N_10508);
xor U11438 (N_11438,N_10984,N_11211);
xor U11439 (N_11439,N_11069,N_10863);
nand U11440 (N_11440,N_10768,N_11046);
and U11441 (N_11441,N_11220,N_11086);
and U11442 (N_11442,N_11187,N_10714);
nand U11443 (N_11443,N_11186,N_10505);
or U11444 (N_11444,N_10700,N_11059);
or U11445 (N_11445,N_10789,N_11239);
and U11446 (N_11446,N_10705,N_10563);
or U11447 (N_11447,N_11175,N_10963);
and U11448 (N_11448,N_10919,N_10951);
nor U11449 (N_11449,N_11153,N_10899);
or U11450 (N_11450,N_10733,N_11205);
nor U11451 (N_11451,N_10743,N_10521);
or U11452 (N_11452,N_10781,N_10813);
nor U11453 (N_11453,N_10627,N_10551);
and U11454 (N_11454,N_11012,N_11171);
and U11455 (N_11455,N_10581,N_10688);
and U11456 (N_11456,N_11044,N_11176);
or U11457 (N_11457,N_11025,N_10764);
and U11458 (N_11458,N_11033,N_10516);
nand U11459 (N_11459,N_11159,N_10501);
and U11460 (N_11460,N_10859,N_11129);
and U11461 (N_11461,N_10500,N_11074);
or U11462 (N_11462,N_10888,N_10604);
nor U11463 (N_11463,N_11249,N_10746);
or U11464 (N_11464,N_10754,N_10981);
nor U11465 (N_11465,N_10566,N_10628);
nor U11466 (N_11466,N_10531,N_10690);
nand U11467 (N_11467,N_10952,N_10946);
nor U11468 (N_11468,N_10526,N_11172);
nand U11469 (N_11469,N_11244,N_11112);
and U11470 (N_11470,N_11101,N_10594);
nor U11471 (N_11471,N_10533,N_10933);
nor U11472 (N_11472,N_11130,N_10720);
nor U11473 (N_11473,N_10792,N_10701);
or U11474 (N_11474,N_10958,N_10761);
nand U11475 (N_11475,N_10605,N_10510);
nor U11476 (N_11476,N_10640,N_10548);
and U11477 (N_11477,N_11241,N_10852);
xor U11478 (N_11478,N_10512,N_10817);
nand U11479 (N_11479,N_10732,N_10962);
nor U11480 (N_11480,N_11004,N_10851);
nor U11481 (N_11481,N_10728,N_10669);
nand U11482 (N_11482,N_10841,N_11024);
and U11483 (N_11483,N_10634,N_10558);
nand U11484 (N_11484,N_11108,N_10518);
nor U11485 (N_11485,N_10736,N_10860);
nor U11486 (N_11486,N_10929,N_10884);
or U11487 (N_11487,N_10559,N_11167);
and U11488 (N_11488,N_10602,N_10827);
nor U11489 (N_11489,N_10942,N_10744);
nand U11490 (N_11490,N_11236,N_11018);
nor U11491 (N_11491,N_11217,N_11077);
nor U11492 (N_11492,N_10943,N_10795);
or U11493 (N_11493,N_10887,N_11031);
nor U11494 (N_11494,N_10840,N_10759);
or U11495 (N_11495,N_10798,N_10681);
and U11496 (N_11496,N_10549,N_10673);
and U11497 (N_11497,N_10539,N_10920);
nor U11498 (N_11498,N_10786,N_10976);
xnor U11499 (N_11499,N_10926,N_11163);
nor U11500 (N_11500,N_11208,N_10708);
nor U11501 (N_11501,N_10872,N_11147);
nor U11502 (N_11502,N_10979,N_10572);
nor U11503 (N_11503,N_10875,N_10600);
and U11504 (N_11504,N_10692,N_10680);
nand U11505 (N_11505,N_10883,N_11113);
nand U11506 (N_11506,N_10968,N_11111);
or U11507 (N_11507,N_11160,N_10922);
nor U11508 (N_11508,N_11135,N_10923);
nor U11509 (N_11509,N_10993,N_10567);
or U11510 (N_11510,N_10588,N_10980);
nor U11511 (N_11511,N_11091,N_10846);
and U11512 (N_11512,N_10910,N_10991);
or U11513 (N_11513,N_11060,N_11143);
xor U11514 (N_11514,N_10671,N_10858);
nor U11515 (N_11515,N_10927,N_10930);
nor U11516 (N_11516,N_10889,N_11193);
nand U11517 (N_11517,N_11065,N_11237);
nand U11518 (N_11518,N_11158,N_10695);
xor U11519 (N_11519,N_10934,N_10830);
and U11520 (N_11520,N_10645,N_11106);
nor U11521 (N_11521,N_10662,N_10739);
nor U11522 (N_11522,N_11028,N_11233);
nor U11523 (N_11523,N_10615,N_10725);
nor U11524 (N_11524,N_10576,N_11240);
nand U11525 (N_11525,N_10864,N_11078);
or U11526 (N_11526,N_10793,N_10921);
and U11527 (N_11527,N_11103,N_10687);
nand U11528 (N_11528,N_11219,N_11029);
and U11529 (N_11529,N_10618,N_10582);
and U11530 (N_11530,N_10783,N_11007);
and U11531 (N_11531,N_10646,N_10900);
or U11532 (N_11532,N_10866,N_10506);
and U11533 (N_11533,N_10573,N_10557);
xor U11534 (N_11534,N_11058,N_11222);
and U11535 (N_11535,N_11196,N_10513);
nor U11536 (N_11536,N_10855,N_11127);
and U11537 (N_11537,N_11198,N_10639);
and U11538 (N_11538,N_11064,N_10814);
nand U11539 (N_11539,N_11216,N_10948);
xor U11540 (N_11540,N_10800,N_11039);
nor U11541 (N_11541,N_10937,N_10945);
xor U11542 (N_11542,N_10971,N_11006);
nand U11543 (N_11543,N_10844,N_11056);
nor U11544 (N_11544,N_11243,N_11032);
and U11545 (N_11545,N_10719,N_10953);
nand U11546 (N_11546,N_11234,N_11178);
or U11547 (N_11547,N_10713,N_10597);
nor U11548 (N_11548,N_10723,N_10543);
and U11549 (N_11549,N_10782,N_10599);
or U11550 (N_11550,N_10925,N_10794);
and U11551 (N_11551,N_10616,N_10741);
or U11552 (N_11552,N_11027,N_11104);
nand U11553 (N_11553,N_11084,N_10715);
nand U11554 (N_11554,N_11229,N_11092);
or U11555 (N_11555,N_11009,N_10917);
or U11556 (N_11556,N_10502,N_10532);
and U11557 (N_11557,N_10928,N_10903);
nand U11558 (N_11558,N_11076,N_11181);
nor U11559 (N_11559,N_10755,N_11183);
xor U11560 (N_11560,N_10772,N_10709);
nor U11561 (N_11561,N_11095,N_11099);
or U11562 (N_11562,N_11168,N_10676);
and U11563 (N_11563,N_10834,N_11057);
xnor U11564 (N_11564,N_10679,N_11034);
nor U11565 (N_11565,N_11128,N_10515);
nor U11566 (N_11566,N_11197,N_10983);
nand U11567 (N_11567,N_11118,N_10663);
and U11568 (N_11568,N_10816,N_11142);
nand U11569 (N_11569,N_10990,N_11050);
nand U11570 (N_11570,N_10869,N_10606);
and U11571 (N_11571,N_10854,N_10932);
nor U11572 (N_11572,N_10885,N_10756);
and U11573 (N_11573,N_11105,N_10697);
and U11574 (N_11574,N_10819,N_10748);
nor U11575 (N_11575,N_10545,N_11062);
nor U11576 (N_11576,N_11098,N_10722);
and U11577 (N_11577,N_10619,N_11195);
and U11578 (N_11578,N_10760,N_10632);
nand U11579 (N_11579,N_11014,N_11049);
or U11580 (N_11580,N_11100,N_10541);
and U11581 (N_11581,N_11133,N_10694);
or U11582 (N_11582,N_10585,N_10651);
or U11583 (N_11583,N_10822,N_11003);
nor U11584 (N_11584,N_10828,N_10909);
or U11585 (N_11585,N_10918,N_10949);
or U11586 (N_11586,N_10902,N_10911);
nand U11587 (N_11587,N_11073,N_11026);
or U11588 (N_11588,N_11136,N_10966);
nand U11589 (N_11589,N_10769,N_10565);
nand U11590 (N_11590,N_10803,N_11206);
or U11591 (N_11591,N_10775,N_10865);
and U11592 (N_11592,N_11037,N_10796);
xor U11593 (N_11593,N_11070,N_10753);
or U11594 (N_11594,N_10601,N_10807);
and U11595 (N_11595,N_11224,N_10805);
nand U11596 (N_11596,N_10527,N_10696);
and U11597 (N_11597,N_11117,N_10935);
and U11598 (N_11598,N_11191,N_10811);
nor U11599 (N_11599,N_10938,N_10897);
nand U11600 (N_11600,N_10529,N_11119);
nor U11601 (N_11601,N_11123,N_11047);
or U11602 (N_11602,N_11189,N_10992);
and U11603 (N_11603,N_10784,N_10982);
and U11604 (N_11604,N_10913,N_10587);
nand U11605 (N_11605,N_10578,N_10873);
and U11606 (N_11606,N_11164,N_10901);
nand U11607 (N_11607,N_11200,N_10538);
nor U11608 (N_11608,N_10940,N_10608);
nor U11609 (N_11609,N_11152,N_10693);
nand U11610 (N_11610,N_10999,N_11015);
nand U11611 (N_11611,N_10895,N_11038);
or U11612 (N_11612,N_10829,N_10894);
and U11613 (N_11613,N_10568,N_10878);
nand U11614 (N_11614,N_10832,N_11169);
nand U11615 (N_11615,N_10763,N_10520);
nor U11616 (N_11616,N_10555,N_11088);
nor U11617 (N_11617,N_11068,N_11010);
nand U11618 (N_11618,N_11011,N_11002);
nand U11619 (N_11619,N_11000,N_10848);
and U11620 (N_11620,N_10675,N_10790);
or U11621 (N_11621,N_10791,N_10637);
nor U11622 (N_11622,N_11005,N_10986);
or U11623 (N_11623,N_10554,N_10975);
nor U11624 (N_11624,N_10635,N_10514);
xnor U11625 (N_11625,N_10750,N_10783);
nor U11626 (N_11626,N_10670,N_10702);
and U11627 (N_11627,N_10837,N_10917);
nand U11628 (N_11628,N_10940,N_11057);
and U11629 (N_11629,N_10687,N_11187);
or U11630 (N_11630,N_10853,N_10860);
and U11631 (N_11631,N_11134,N_11236);
nor U11632 (N_11632,N_10734,N_10882);
nor U11633 (N_11633,N_11192,N_10911);
xor U11634 (N_11634,N_10684,N_10872);
nor U11635 (N_11635,N_11209,N_10671);
nor U11636 (N_11636,N_10835,N_10563);
nor U11637 (N_11637,N_10752,N_10662);
nor U11638 (N_11638,N_10563,N_10965);
and U11639 (N_11639,N_11231,N_11197);
or U11640 (N_11640,N_10596,N_10951);
nand U11641 (N_11641,N_11229,N_11118);
nor U11642 (N_11642,N_10648,N_11111);
or U11643 (N_11643,N_10947,N_10875);
nor U11644 (N_11644,N_10685,N_11248);
and U11645 (N_11645,N_11102,N_10994);
or U11646 (N_11646,N_10883,N_10507);
and U11647 (N_11647,N_10516,N_11228);
and U11648 (N_11648,N_10861,N_10615);
nor U11649 (N_11649,N_11159,N_11066);
xor U11650 (N_11650,N_11080,N_10597);
nor U11651 (N_11651,N_10997,N_10723);
or U11652 (N_11652,N_10506,N_11069);
xnor U11653 (N_11653,N_10515,N_11142);
nor U11654 (N_11654,N_10882,N_10968);
or U11655 (N_11655,N_10973,N_10743);
or U11656 (N_11656,N_10746,N_10571);
and U11657 (N_11657,N_11027,N_10608);
and U11658 (N_11658,N_11202,N_11047);
nor U11659 (N_11659,N_10505,N_11045);
nor U11660 (N_11660,N_10790,N_11055);
and U11661 (N_11661,N_10857,N_10923);
xnor U11662 (N_11662,N_11111,N_10979);
nor U11663 (N_11663,N_10992,N_10705);
nor U11664 (N_11664,N_10864,N_11170);
and U11665 (N_11665,N_11150,N_11242);
nand U11666 (N_11666,N_10853,N_10861);
or U11667 (N_11667,N_10732,N_10855);
nor U11668 (N_11668,N_10821,N_10993);
or U11669 (N_11669,N_11053,N_10971);
and U11670 (N_11670,N_10848,N_11100);
xnor U11671 (N_11671,N_10940,N_11147);
xnor U11672 (N_11672,N_10928,N_10995);
and U11673 (N_11673,N_10870,N_10633);
and U11674 (N_11674,N_10608,N_10663);
nor U11675 (N_11675,N_10504,N_11081);
or U11676 (N_11676,N_10512,N_11175);
and U11677 (N_11677,N_10929,N_11153);
xnor U11678 (N_11678,N_10941,N_10926);
or U11679 (N_11679,N_10881,N_10747);
nand U11680 (N_11680,N_11078,N_10991);
and U11681 (N_11681,N_11006,N_11114);
xor U11682 (N_11682,N_10739,N_11201);
nor U11683 (N_11683,N_11068,N_10827);
nand U11684 (N_11684,N_11182,N_10974);
and U11685 (N_11685,N_10933,N_11123);
or U11686 (N_11686,N_10505,N_10545);
nand U11687 (N_11687,N_10742,N_11083);
and U11688 (N_11688,N_10902,N_10667);
or U11689 (N_11689,N_10598,N_10900);
and U11690 (N_11690,N_10717,N_10568);
or U11691 (N_11691,N_10829,N_10844);
nand U11692 (N_11692,N_10838,N_10957);
xnor U11693 (N_11693,N_11023,N_10780);
xor U11694 (N_11694,N_10559,N_10618);
or U11695 (N_11695,N_10569,N_10876);
nor U11696 (N_11696,N_11075,N_11049);
and U11697 (N_11697,N_11084,N_10501);
or U11698 (N_11698,N_10628,N_11041);
or U11699 (N_11699,N_10609,N_10635);
nor U11700 (N_11700,N_10538,N_10875);
and U11701 (N_11701,N_10639,N_10768);
nor U11702 (N_11702,N_10973,N_10596);
nor U11703 (N_11703,N_11095,N_11211);
and U11704 (N_11704,N_11033,N_10710);
nor U11705 (N_11705,N_10949,N_10990);
and U11706 (N_11706,N_10997,N_10972);
nor U11707 (N_11707,N_11006,N_11179);
xor U11708 (N_11708,N_10552,N_10708);
xnor U11709 (N_11709,N_10563,N_10519);
or U11710 (N_11710,N_10619,N_10880);
and U11711 (N_11711,N_10998,N_10612);
nand U11712 (N_11712,N_10976,N_11237);
xor U11713 (N_11713,N_11140,N_10914);
xor U11714 (N_11714,N_11007,N_11073);
nor U11715 (N_11715,N_10983,N_10679);
xor U11716 (N_11716,N_10866,N_10653);
xnor U11717 (N_11717,N_11017,N_10540);
nand U11718 (N_11718,N_10715,N_10573);
and U11719 (N_11719,N_10646,N_11035);
nor U11720 (N_11720,N_11110,N_11208);
nand U11721 (N_11721,N_11205,N_11106);
nand U11722 (N_11722,N_10586,N_10719);
or U11723 (N_11723,N_10849,N_10891);
nor U11724 (N_11724,N_11163,N_10557);
or U11725 (N_11725,N_10573,N_10925);
nor U11726 (N_11726,N_10701,N_10537);
xor U11727 (N_11727,N_10587,N_11126);
or U11728 (N_11728,N_10711,N_10859);
or U11729 (N_11729,N_10787,N_10736);
nor U11730 (N_11730,N_10701,N_10536);
nand U11731 (N_11731,N_10815,N_10819);
or U11732 (N_11732,N_10946,N_10660);
xnor U11733 (N_11733,N_10527,N_10991);
and U11734 (N_11734,N_10894,N_11050);
nor U11735 (N_11735,N_10534,N_11223);
or U11736 (N_11736,N_10524,N_10966);
nor U11737 (N_11737,N_10808,N_11187);
and U11738 (N_11738,N_10614,N_11201);
nand U11739 (N_11739,N_10990,N_10758);
and U11740 (N_11740,N_10734,N_11034);
nor U11741 (N_11741,N_10993,N_10696);
or U11742 (N_11742,N_11027,N_11220);
or U11743 (N_11743,N_11236,N_10781);
or U11744 (N_11744,N_11027,N_10769);
nand U11745 (N_11745,N_10677,N_11154);
or U11746 (N_11746,N_11186,N_10809);
or U11747 (N_11747,N_10907,N_10830);
or U11748 (N_11748,N_10564,N_10891);
nand U11749 (N_11749,N_10670,N_11030);
or U11750 (N_11750,N_11015,N_10995);
nand U11751 (N_11751,N_10652,N_10869);
or U11752 (N_11752,N_11128,N_10581);
nand U11753 (N_11753,N_10658,N_10609);
or U11754 (N_11754,N_10608,N_10595);
nor U11755 (N_11755,N_10537,N_10859);
xnor U11756 (N_11756,N_10536,N_10932);
and U11757 (N_11757,N_10561,N_10674);
nand U11758 (N_11758,N_11235,N_11028);
or U11759 (N_11759,N_10897,N_10842);
nor U11760 (N_11760,N_11148,N_11083);
or U11761 (N_11761,N_10730,N_11229);
or U11762 (N_11762,N_11168,N_10898);
or U11763 (N_11763,N_10899,N_10831);
and U11764 (N_11764,N_10751,N_10892);
nor U11765 (N_11765,N_11091,N_10733);
xor U11766 (N_11766,N_10530,N_10651);
xor U11767 (N_11767,N_11209,N_11229);
xor U11768 (N_11768,N_10631,N_10595);
or U11769 (N_11769,N_10857,N_10619);
nand U11770 (N_11770,N_11202,N_10583);
nor U11771 (N_11771,N_10919,N_11196);
nor U11772 (N_11772,N_10985,N_11037);
nor U11773 (N_11773,N_11231,N_11166);
nor U11774 (N_11774,N_11065,N_10680);
and U11775 (N_11775,N_10561,N_10544);
or U11776 (N_11776,N_10606,N_11128);
nand U11777 (N_11777,N_10939,N_10630);
xnor U11778 (N_11778,N_10789,N_10678);
nor U11779 (N_11779,N_10933,N_10882);
nand U11780 (N_11780,N_10583,N_10888);
or U11781 (N_11781,N_10965,N_10906);
nand U11782 (N_11782,N_11074,N_11029);
or U11783 (N_11783,N_10653,N_10536);
nand U11784 (N_11784,N_11214,N_10543);
or U11785 (N_11785,N_11027,N_11003);
or U11786 (N_11786,N_10693,N_10771);
nor U11787 (N_11787,N_10777,N_10916);
nand U11788 (N_11788,N_10674,N_11247);
and U11789 (N_11789,N_11004,N_11160);
nor U11790 (N_11790,N_11026,N_10572);
and U11791 (N_11791,N_10881,N_10929);
or U11792 (N_11792,N_10651,N_10928);
nand U11793 (N_11793,N_10574,N_10751);
nand U11794 (N_11794,N_10816,N_11117);
nor U11795 (N_11795,N_10528,N_11141);
and U11796 (N_11796,N_10769,N_10766);
nor U11797 (N_11797,N_10738,N_11201);
nand U11798 (N_11798,N_10870,N_11076);
nor U11799 (N_11799,N_10520,N_10594);
or U11800 (N_11800,N_10937,N_10652);
or U11801 (N_11801,N_10888,N_11174);
nand U11802 (N_11802,N_11077,N_10512);
nand U11803 (N_11803,N_10615,N_11084);
or U11804 (N_11804,N_10986,N_11024);
nor U11805 (N_11805,N_10505,N_10958);
nand U11806 (N_11806,N_10590,N_10911);
nor U11807 (N_11807,N_11081,N_10824);
and U11808 (N_11808,N_10630,N_10783);
and U11809 (N_11809,N_10862,N_10531);
xor U11810 (N_11810,N_10672,N_10698);
xnor U11811 (N_11811,N_11136,N_11008);
nor U11812 (N_11812,N_10982,N_10720);
and U11813 (N_11813,N_10986,N_11132);
nor U11814 (N_11814,N_11034,N_11097);
and U11815 (N_11815,N_10608,N_10702);
and U11816 (N_11816,N_11231,N_11249);
xor U11817 (N_11817,N_10685,N_10773);
or U11818 (N_11818,N_11021,N_10733);
and U11819 (N_11819,N_10981,N_10890);
nand U11820 (N_11820,N_10770,N_11047);
xnor U11821 (N_11821,N_10675,N_11081);
or U11822 (N_11822,N_10668,N_10735);
and U11823 (N_11823,N_11063,N_11214);
xor U11824 (N_11824,N_11210,N_11142);
or U11825 (N_11825,N_11093,N_10625);
nor U11826 (N_11826,N_10937,N_10952);
nand U11827 (N_11827,N_10679,N_10863);
and U11828 (N_11828,N_10942,N_10843);
xnor U11829 (N_11829,N_10627,N_10509);
and U11830 (N_11830,N_10790,N_10928);
or U11831 (N_11831,N_10505,N_10957);
or U11832 (N_11832,N_10917,N_11185);
nand U11833 (N_11833,N_10879,N_10621);
and U11834 (N_11834,N_10915,N_10785);
nand U11835 (N_11835,N_10900,N_10783);
nand U11836 (N_11836,N_11036,N_10508);
and U11837 (N_11837,N_10689,N_10895);
or U11838 (N_11838,N_10951,N_10837);
nor U11839 (N_11839,N_10737,N_10792);
or U11840 (N_11840,N_11062,N_11194);
nand U11841 (N_11841,N_10968,N_10562);
nor U11842 (N_11842,N_10856,N_10824);
or U11843 (N_11843,N_10737,N_11132);
and U11844 (N_11844,N_10748,N_10803);
or U11845 (N_11845,N_10567,N_10962);
nand U11846 (N_11846,N_10756,N_10801);
or U11847 (N_11847,N_10830,N_10856);
nor U11848 (N_11848,N_10883,N_11057);
nand U11849 (N_11849,N_10927,N_10777);
nor U11850 (N_11850,N_10891,N_10614);
nand U11851 (N_11851,N_10720,N_10837);
or U11852 (N_11852,N_10870,N_10523);
or U11853 (N_11853,N_11229,N_10676);
nor U11854 (N_11854,N_11084,N_10695);
and U11855 (N_11855,N_10742,N_11195);
or U11856 (N_11856,N_10735,N_10608);
xnor U11857 (N_11857,N_11029,N_11062);
nand U11858 (N_11858,N_11113,N_10762);
nor U11859 (N_11859,N_10796,N_10789);
or U11860 (N_11860,N_11218,N_10691);
nand U11861 (N_11861,N_10634,N_10924);
nor U11862 (N_11862,N_10940,N_10972);
nand U11863 (N_11863,N_11137,N_10972);
xnor U11864 (N_11864,N_11133,N_11151);
nor U11865 (N_11865,N_10543,N_11174);
or U11866 (N_11866,N_10949,N_11086);
nand U11867 (N_11867,N_10683,N_10705);
or U11868 (N_11868,N_11114,N_10749);
or U11869 (N_11869,N_10626,N_10933);
and U11870 (N_11870,N_10991,N_11022);
xnor U11871 (N_11871,N_10778,N_10757);
or U11872 (N_11872,N_11036,N_10965);
and U11873 (N_11873,N_11173,N_10979);
xor U11874 (N_11874,N_10600,N_11090);
nor U11875 (N_11875,N_10855,N_11164);
nand U11876 (N_11876,N_10919,N_11084);
or U11877 (N_11877,N_10878,N_11211);
nand U11878 (N_11878,N_10964,N_11232);
and U11879 (N_11879,N_10812,N_10740);
nor U11880 (N_11880,N_10938,N_10774);
or U11881 (N_11881,N_10547,N_10651);
nand U11882 (N_11882,N_11179,N_10661);
and U11883 (N_11883,N_10714,N_11000);
and U11884 (N_11884,N_10917,N_10929);
and U11885 (N_11885,N_11093,N_10864);
and U11886 (N_11886,N_10709,N_10972);
nor U11887 (N_11887,N_10602,N_10707);
nor U11888 (N_11888,N_10904,N_10931);
and U11889 (N_11889,N_11196,N_10636);
nor U11890 (N_11890,N_10637,N_10548);
or U11891 (N_11891,N_10824,N_10922);
and U11892 (N_11892,N_10543,N_10797);
nand U11893 (N_11893,N_10840,N_10995);
or U11894 (N_11894,N_10999,N_11138);
nand U11895 (N_11895,N_11042,N_11083);
nor U11896 (N_11896,N_10552,N_10980);
and U11897 (N_11897,N_11072,N_10673);
and U11898 (N_11898,N_10508,N_10969);
or U11899 (N_11899,N_10797,N_11019);
nor U11900 (N_11900,N_10635,N_10584);
xor U11901 (N_11901,N_10580,N_10882);
or U11902 (N_11902,N_10773,N_10985);
and U11903 (N_11903,N_11037,N_10780);
or U11904 (N_11904,N_10592,N_10599);
and U11905 (N_11905,N_10782,N_10867);
nor U11906 (N_11906,N_11144,N_10845);
and U11907 (N_11907,N_10932,N_10804);
nor U11908 (N_11908,N_10538,N_11011);
or U11909 (N_11909,N_10903,N_10891);
and U11910 (N_11910,N_10568,N_10686);
nor U11911 (N_11911,N_10682,N_10881);
nor U11912 (N_11912,N_11206,N_10981);
and U11913 (N_11913,N_10788,N_10906);
xor U11914 (N_11914,N_10710,N_10843);
xor U11915 (N_11915,N_10555,N_10584);
nand U11916 (N_11916,N_11240,N_10844);
or U11917 (N_11917,N_10584,N_10519);
or U11918 (N_11918,N_10859,N_10727);
nor U11919 (N_11919,N_10661,N_11085);
nor U11920 (N_11920,N_10831,N_11127);
nor U11921 (N_11921,N_11217,N_10906);
and U11922 (N_11922,N_10662,N_10780);
nand U11923 (N_11923,N_10806,N_11007);
nand U11924 (N_11924,N_10961,N_11060);
nand U11925 (N_11925,N_10912,N_11024);
nor U11926 (N_11926,N_11032,N_10960);
nand U11927 (N_11927,N_10543,N_10595);
nand U11928 (N_11928,N_10611,N_11172);
and U11929 (N_11929,N_10890,N_11013);
nor U11930 (N_11930,N_11061,N_10711);
nand U11931 (N_11931,N_10918,N_10970);
xor U11932 (N_11932,N_10796,N_10937);
and U11933 (N_11933,N_10561,N_10821);
nor U11934 (N_11934,N_10620,N_10997);
and U11935 (N_11935,N_11147,N_11091);
or U11936 (N_11936,N_10689,N_11218);
nand U11937 (N_11937,N_10668,N_10718);
nand U11938 (N_11938,N_10704,N_10699);
and U11939 (N_11939,N_11075,N_11018);
nor U11940 (N_11940,N_10641,N_10512);
xnor U11941 (N_11941,N_11103,N_10900);
and U11942 (N_11942,N_10544,N_11139);
nand U11943 (N_11943,N_10716,N_10894);
nand U11944 (N_11944,N_10618,N_10739);
nand U11945 (N_11945,N_11243,N_11027);
and U11946 (N_11946,N_11021,N_10841);
xnor U11947 (N_11947,N_11009,N_10794);
nor U11948 (N_11948,N_10578,N_11035);
nand U11949 (N_11949,N_10698,N_11234);
or U11950 (N_11950,N_11078,N_10556);
nor U11951 (N_11951,N_10986,N_11042);
nand U11952 (N_11952,N_10758,N_10639);
xor U11953 (N_11953,N_11182,N_10642);
xnor U11954 (N_11954,N_10818,N_11237);
and U11955 (N_11955,N_11031,N_10900);
nand U11956 (N_11956,N_11249,N_10723);
or U11957 (N_11957,N_11178,N_10883);
or U11958 (N_11958,N_10724,N_11141);
xnor U11959 (N_11959,N_11023,N_10646);
or U11960 (N_11960,N_10644,N_10805);
and U11961 (N_11961,N_10654,N_11191);
or U11962 (N_11962,N_10532,N_10600);
or U11963 (N_11963,N_11040,N_10912);
nand U11964 (N_11964,N_10559,N_10647);
nor U11965 (N_11965,N_10827,N_10563);
or U11966 (N_11966,N_11205,N_11177);
or U11967 (N_11967,N_11108,N_11133);
or U11968 (N_11968,N_10849,N_10664);
or U11969 (N_11969,N_10729,N_11238);
and U11970 (N_11970,N_10980,N_11216);
nor U11971 (N_11971,N_11019,N_10828);
or U11972 (N_11972,N_10835,N_10661);
and U11973 (N_11973,N_10820,N_11078);
nor U11974 (N_11974,N_11199,N_10688);
and U11975 (N_11975,N_11133,N_10917);
or U11976 (N_11976,N_10622,N_10840);
and U11977 (N_11977,N_10570,N_10932);
nor U11978 (N_11978,N_10903,N_10999);
nand U11979 (N_11979,N_10632,N_10576);
nand U11980 (N_11980,N_10699,N_10751);
and U11981 (N_11981,N_10723,N_10900);
xor U11982 (N_11982,N_11020,N_10506);
or U11983 (N_11983,N_11215,N_10930);
nor U11984 (N_11984,N_11136,N_10506);
nor U11985 (N_11985,N_10767,N_10941);
nor U11986 (N_11986,N_11151,N_10757);
and U11987 (N_11987,N_10613,N_11062);
and U11988 (N_11988,N_11135,N_10523);
nor U11989 (N_11989,N_11143,N_11064);
nand U11990 (N_11990,N_10673,N_10601);
nand U11991 (N_11991,N_10500,N_10888);
and U11992 (N_11992,N_10892,N_10956);
xor U11993 (N_11993,N_10688,N_10882);
nor U11994 (N_11994,N_10917,N_11244);
and U11995 (N_11995,N_11149,N_10934);
xnor U11996 (N_11996,N_11118,N_11014);
xor U11997 (N_11997,N_10764,N_11141);
nand U11998 (N_11998,N_10552,N_10998);
and U11999 (N_11999,N_11021,N_10768);
or U12000 (N_12000,N_11844,N_11362);
xnor U12001 (N_12001,N_11736,N_11607);
nor U12002 (N_12002,N_11419,N_11831);
nor U12003 (N_12003,N_11320,N_11905);
nand U12004 (N_12004,N_11542,N_11481);
nand U12005 (N_12005,N_11696,N_11325);
xnor U12006 (N_12006,N_11346,N_11726);
nor U12007 (N_12007,N_11490,N_11958);
or U12008 (N_12008,N_11530,N_11763);
nor U12009 (N_12009,N_11775,N_11523);
nand U12010 (N_12010,N_11665,N_11977);
nor U12011 (N_12011,N_11917,N_11838);
nand U12012 (N_12012,N_11491,N_11280);
or U12013 (N_12013,N_11779,N_11326);
and U12014 (N_12014,N_11305,N_11798);
or U12015 (N_12015,N_11477,N_11940);
xor U12016 (N_12016,N_11332,N_11376);
or U12017 (N_12017,N_11906,N_11423);
xnor U12018 (N_12018,N_11276,N_11399);
or U12019 (N_12019,N_11316,N_11283);
nand U12020 (N_12020,N_11790,N_11270);
nand U12021 (N_12021,N_11581,N_11650);
nor U12022 (N_12022,N_11662,N_11427);
and U12023 (N_12023,N_11816,N_11635);
nand U12024 (N_12024,N_11558,N_11680);
or U12025 (N_12025,N_11928,N_11502);
xor U12026 (N_12026,N_11646,N_11686);
nor U12027 (N_12027,N_11911,N_11337);
or U12028 (N_12028,N_11832,N_11625);
and U12029 (N_12029,N_11478,N_11438);
xnor U12030 (N_12030,N_11408,N_11693);
xnor U12031 (N_12031,N_11651,N_11367);
nand U12032 (N_12032,N_11666,N_11366);
or U12033 (N_12033,N_11683,N_11489);
nor U12034 (N_12034,N_11347,N_11770);
or U12035 (N_12035,N_11596,N_11772);
or U12036 (N_12036,N_11406,N_11484);
nand U12037 (N_12037,N_11468,N_11973);
nand U12038 (N_12038,N_11262,N_11654);
or U12039 (N_12039,N_11519,N_11479);
and U12040 (N_12040,N_11791,N_11513);
xor U12041 (N_12041,N_11488,N_11821);
nand U12042 (N_12042,N_11543,N_11339);
nor U12043 (N_12043,N_11372,N_11254);
and U12044 (N_12044,N_11876,N_11774);
or U12045 (N_12045,N_11360,N_11971);
or U12046 (N_12046,N_11585,N_11766);
nor U12047 (N_12047,N_11375,N_11935);
nand U12048 (N_12048,N_11507,N_11556);
or U12049 (N_12049,N_11279,N_11559);
and U12050 (N_12050,N_11861,N_11573);
nand U12051 (N_12051,N_11512,N_11572);
xnor U12052 (N_12052,N_11994,N_11350);
nor U12053 (N_12053,N_11398,N_11595);
xnor U12054 (N_12054,N_11801,N_11975);
and U12055 (N_12055,N_11892,N_11609);
or U12056 (N_12056,N_11717,N_11296);
nor U12057 (N_12057,N_11890,N_11273);
and U12058 (N_12058,N_11674,N_11638);
or U12059 (N_12059,N_11454,N_11834);
nor U12060 (N_12060,N_11628,N_11447);
nor U12061 (N_12061,N_11370,N_11867);
nand U12062 (N_12062,N_11714,N_11528);
nand U12063 (N_12063,N_11443,N_11255);
nand U12064 (N_12064,N_11846,N_11944);
xor U12065 (N_12065,N_11794,N_11516);
and U12066 (N_12066,N_11531,N_11286);
and U12067 (N_12067,N_11356,N_11985);
nor U12068 (N_12068,N_11250,N_11970);
nand U12069 (N_12069,N_11950,N_11411);
and U12070 (N_12070,N_11744,N_11587);
and U12071 (N_12071,N_11565,N_11421);
nand U12072 (N_12072,N_11632,N_11263);
or U12073 (N_12073,N_11862,N_11592);
nor U12074 (N_12074,N_11453,N_11505);
nor U12075 (N_12075,N_11451,N_11997);
xor U12076 (N_12076,N_11742,N_11939);
and U12077 (N_12077,N_11681,N_11333);
and U12078 (N_12078,N_11534,N_11981);
nand U12079 (N_12079,N_11999,N_11599);
or U12080 (N_12080,N_11449,N_11749);
or U12081 (N_12081,N_11752,N_11377);
nand U12082 (N_12082,N_11723,N_11336);
or U12083 (N_12083,N_11335,N_11793);
and U12084 (N_12084,N_11927,N_11498);
nand U12085 (N_12085,N_11967,N_11682);
or U12086 (N_12086,N_11466,N_11327);
nor U12087 (N_12087,N_11987,N_11968);
and U12088 (N_12088,N_11315,N_11483);
or U12089 (N_12089,N_11877,N_11746);
or U12090 (N_12090,N_11261,N_11989);
or U12091 (N_12091,N_11792,N_11643);
nand U12092 (N_12092,N_11458,N_11824);
and U12093 (N_12093,N_11393,N_11597);
nand U12094 (N_12094,N_11750,N_11331);
nand U12095 (N_12095,N_11946,N_11422);
or U12096 (N_12096,N_11503,N_11308);
or U12097 (N_12097,N_11402,N_11610);
nor U12098 (N_12098,N_11341,N_11990);
nand U12099 (N_12099,N_11330,N_11323);
xor U12100 (N_12100,N_11358,N_11383);
and U12101 (N_12101,N_11252,N_11656);
and U12102 (N_12102,N_11904,N_11839);
nor U12103 (N_12103,N_11873,N_11539);
nand U12104 (N_12104,N_11567,N_11678);
and U12105 (N_12105,N_11521,N_11941);
and U12106 (N_12106,N_11591,N_11836);
nor U12107 (N_12107,N_11340,N_11663);
or U12108 (N_12108,N_11475,N_11322);
or U12109 (N_12109,N_11524,N_11275);
and U12110 (N_12110,N_11430,N_11590);
or U12111 (N_12111,N_11274,N_11753);
nand U12112 (N_12112,N_11795,N_11948);
nand U12113 (N_12113,N_11444,N_11329);
or U12114 (N_12114,N_11933,N_11776);
or U12115 (N_12115,N_11389,N_11511);
or U12116 (N_12116,N_11708,N_11704);
and U12117 (N_12117,N_11781,N_11299);
nand U12118 (N_12118,N_11853,N_11504);
and U12119 (N_12119,N_11517,N_11961);
or U12120 (N_12120,N_11756,N_11380);
and U12121 (N_12121,N_11334,N_11854);
or U12122 (N_12122,N_11442,N_11537);
nor U12123 (N_12123,N_11536,N_11768);
or U12124 (N_12124,N_11583,N_11538);
nand U12125 (N_12125,N_11891,N_11864);
nand U12126 (N_12126,N_11314,N_11762);
and U12127 (N_12127,N_11922,N_11745);
or U12128 (N_12128,N_11979,N_11709);
or U12129 (N_12129,N_11829,N_11951);
and U12130 (N_12130,N_11574,N_11550);
and U12131 (N_12131,N_11555,N_11761);
nand U12132 (N_12132,N_11920,N_11472);
and U12133 (N_12133,N_11306,N_11827);
xnor U12134 (N_12134,N_11957,N_11807);
nand U12135 (N_12135,N_11445,N_11557);
and U12136 (N_12136,N_11668,N_11553);
nand U12137 (N_12137,N_11469,N_11353);
xnor U12138 (N_12138,N_11301,N_11623);
or U12139 (N_12139,N_11485,N_11740);
nand U12140 (N_12140,N_11780,N_11812);
nand U12141 (N_12141,N_11374,N_11461);
or U12142 (N_12142,N_11570,N_11782);
nand U12143 (N_12143,N_11634,N_11527);
nor U12144 (N_12144,N_11936,N_11272);
nand U12145 (N_12145,N_11738,N_11494);
or U12146 (N_12146,N_11788,N_11344);
nand U12147 (N_12147,N_11799,N_11382);
xnor U12148 (N_12148,N_11568,N_11850);
nand U12149 (N_12149,N_11878,N_11866);
and U12150 (N_12150,N_11577,N_11998);
nand U12151 (N_12151,N_11966,N_11437);
nor U12152 (N_12152,N_11995,N_11817);
nor U12153 (N_12153,N_11857,N_11787);
or U12154 (N_12154,N_11943,N_11264);
or U12155 (N_12155,N_11338,N_11659);
or U12156 (N_12156,N_11364,N_11289);
or U12157 (N_12157,N_11849,N_11614);
xnor U12158 (N_12158,N_11390,N_11830);
nor U12159 (N_12159,N_11303,N_11368);
or U12160 (N_12160,N_11391,N_11582);
nand U12161 (N_12161,N_11518,N_11897);
nand U12162 (N_12162,N_11992,N_11884);
and U12163 (N_12163,N_11835,N_11395);
nor U12164 (N_12164,N_11433,N_11624);
nor U12165 (N_12165,N_11352,N_11739);
and U12166 (N_12166,N_11667,N_11520);
and U12167 (N_12167,N_11741,N_11881);
nor U12168 (N_12168,N_11983,N_11673);
and U12169 (N_12169,N_11809,N_11621);
xor U12170 (N_12170,N_11471,N_11713);
nand U12171 (N_12171,N_11616,N_11578);
or U12172 (N_12172,N_11729,N_11868);
and U12173 (N_12173,N_11914,N_11622);
xor U12174 (N_12174,N_11688,N_11655);
and U12175 (N_12175,N_11955,N_11769);
xnor U12176 (N_12176,N_11435,N_11647);
nand U12177 (N_12177,N_11953,N_11889);
xor U12178 (N_12178,N_11942,N_11594);
nand U12179 (N_12179,N_11978,N_11473);
and U12180 (N_12180,N_11893,N_11566);
or U12181 (N_12181,N_11754,N_11584);
and U12182 (N_12182,N_11586,N_11425);
nor U12183 (N_12183,N_11912,N_11418);
nor U12184 (N_12184,N_11748,N_11480);
and U12185 (N_12185,N_11560,N_11938);
nor U12186 (N_12186,N_11661,N_11563);
or U12187 (N_12187,N_11349,N_11710);
and U12188 (N_12188,N_11860,N_11436);
and U12189 (N_12189,N_11548,N_11545);
nor U12190 (N_12190,N_11764,N_11400);
or U12191 (N_12191,N_11902,N_11260);
nand U12192 (N_12192,N_11253,N_11923);
and U12193 (N_12193,N_11732,N_11734);
nor U12194 (N_12194,N_11387,N_11900);
nor U12195 (N_12195,N_11915,N_11882);
or U12196 (N_12196,N_11974,N_11903);
or U12197 (N_12197,N_11986,N_11354);
nor U12198 (N_12198,N_11388,N_11644);
nand U12199 (N_12199,N_11298,N_11404);
and U12200 (N_12200,N_11464,N_11934);
nor U12201 (N_12201,N_11956,N_11608);
and U12202 (N_12202,N_11820,N_11533);
and U12203 (N_12203,N_11277,N_11886);
nor U12204 (N_12204,N_11965,N_11588);
nand U12205 (N_12205,N_11291,N_11639);
nand U12206 (N_12206,N_11465,N_11345);
nor U12207 (N_12207,N_11258,N_11660);
or U12208 (N_12208,N_11653,N_11712);
nand U12209 (N_12209,N_11589,N_11724);
nor U12210 (N_12210,N_11493,N_11302);
xnor U12211 (N_12211,N_11879,N_11514);
nor U12212 (N_12212,N_11649,N_11629);
nor U12213 (N_12213,N_11806,N_11721);
nor U12214 (N_12214,N_11615,N_11529);
and U12215 (N_12215,N_11924,N_11424);
nand U12216 (N_12216,N_11962,N_11960);
and U12217 (N_12217,N_11672,N_11727);
nor U12218 (N_12218,N_11805,N_11869);
or U12219 (N_12219,N_11932,N_11313);
or U12220 (N_12220,N_11909,N_11417);
or U12221 (N_12221,N_11281,N_11571);
and U12222 (N_12222,N_11880,N_11486);
xor U12223 (N_12223,N_11618,N_11474);
nand U12224 (N_12224,N_11642,N_11637);
nand U12225 (N_12225,N_11718,N_11626);
or U12226 (N_12226,N_11457,N_11716);
and U12227 (N_12227,N_11728,N_11747);
nor U12228 (N_12228,N_11684,N_11532);
nor U12229 (N_12229,N_11949,N_11848);
nor U12230 (N_12230,N_11546,N_11870);
nand U12231 (N_12231,N_11972,N_11993);
or U12232 (N_12232,N_11707,N_11725);
and U12233 (N_12233,N_11899,N_11640);
or U12234 (N_12234,N_11365,N_11575);
and U12235 (N_12235,N_11720,N_11508);
and U12236 (N_12236,N_11845,N_11602);
nor U12237 (N_12237,N_11251,N_11913);
nor U12238 (N_12238,N_11910,N_11414);
and U12239 (N_12239,N_11434,N_11576);
nor U12240 (N_12240,N_11361,N_11819);
nand U12241 (N_12241,N_11669,N_11373);
nor U12242 (N_12242,N_11648,N_11540);
nor U12243 (N_12243,N_11996,N_11369);
nor U12244 (N_12244,N_11658,N_11657);
nand U12245 (N_12245,N_11789,N_11432);
and U12246 (N_12246,N_11883,N_11701);
or U12247 (N_12247,N_11705,N_11357);
or U12248 (N_12248,N_11319,N_11679);
xnor U12249 (N_12249,N_11561,N_11901);
nor U12250 (N_12250,N_11413,N_11363);
nor U12251 (N_12251,N_11378,N_11440);
and U12252 (N_12252,N_11875,N_11429);
or U12253 (N_12253,N_11737,N_11271);
and U12254 (N_12254,N_11784,N_11722);
nand U12255 (N_12255,N_11921,N_11492);
nand U12256 (N_12256,N_11702,N_11814);
or U12257 (N_12257,N_11612,N_11982);
and U12258 (N_12258,N_11605,N_11929);
nand U12259 (N_12259,N_11297,N_11525);
and U12260 (N_12260,N_11535,N_11952);
nor U12261 (N_12261,N_11415,N_11448);
nand U12262 (N_12262,N_11851,N_11888);
or U12263 (N_12263,N_11268,N_11343);
nand U12264 (N_12264,N_11825,N_11569);
and U12265 (N_12265,N_11863,N_11822);
nand U12266 (N_12266,N_11828,N_11630);
or U12267 (N_12267,N_11412,N_11731);
or U12268 (N_12268,N_11783,N_11501);
nor U12269 (N_12269,N_11416,N_11476);
nor U12270 (N_12270,N_11773,N_11617);
or U12271 (N_12271,N_11470,N_11266);
xnor U12272 (N_12272,N_11606,N_11410);
or U12273 (N_12273,N_11833,N_11930);
nor U12274 (N_12274,N_11664,N_11976);
nor U12275 (N_12275,N_11459,N_11947);
nand U12276 (N_12276,N_11706,N_11631);
nor U12277 (N_12277,N_11500,N_11856);
and U12278 (N_12278,N_11991,N_11452);
nor U12279 (N_12279,N_11311,N_11964);
or U12280 (N_12280,N_11564,N_11499);
nand U12281 (N_12281,N_11495,N_11269);
or U12282 (N_12282,N_11694,N_11758);
or U12283 (N_12283,N_11670,N_11645);
xor U12284 (N_12284,N_11348,N_11916);
nor U12285 (N_12285,N_11677,N_11907);
nand U12286 (N_12286,N_11619,N_11858);
or U12287 (N_12287,N_11671,N_11803);
nand U12288 (N_12288,N_11580,N_11441);
or U12289 (N_12289,N_11810,N_11379);
nor U12290 (N_12290,N_11818,N_11321);
nand U12291 (N_12291,N_11431,N_11926);
nand U12292 (N_12292,N_11307,N_11755);
and U12293 (N_12293,N_11735,N_11759);
nor U12294 (N_12294,N_11874,N_11808);
and U12295 (N_12295,N_11652,N_11603);
xnor U12296 (N_12296,N_11796,N_11446);
and U12297 (N_12297,N_11551,N_11401);
nand U12298 (N_12298,N_11439,N_11544);
nor U12299 (N_12299,N_11837,N_11403);
and U12300 (N_12300,N_11386,N_11777);
or U12301 (N_12301,N_11547,N_11522);
nand U12302 (N_12302,N_11611,N_11815);
nand U12303 (N_12303,N_11697,N_11450);
or U12304 (N_12304,N_11895,N_11259);
or U12305 (N_12305,N_11381,N_11842);
xor U12306 (N_12306,N_11785,N_11823);
and U12307 (N_12307,N_11887,N_11385);
nand U12308 (N_12308,N_11872,N_11420);
or U12309 (N_12309,N_11552,N_11885);
nor U12310 (N_12310,N_11925,N_11797);
xnor U12311 (N_12311,N_11937,N_11394);
and U12312 (N_12312,N_11549,N_11257);
and U12313 (N_12313,N_11562,N_11765);
xnor U12314 (N_12314,N_11287,N_11526);
or U12315 (N_12315,N_11865,N_11278);
nor U12316 (N_12316,N_11730,N_11692);
or U12317 (N_12317,N_11898,N_11908);
xnor U12318 (N_12318,N_11392,N_11675);
xor U12319 (N_12319,N_11715,N_11288);
nand U12320 (N_12320,N_11641,N_11963);
and U12321 (N_12321,N_11317,N_11691);
nor U12322 (N_12322,N_11351,N_11598);
nand U12323 (N_12323,N_11371,N_11554);
and U12324 (N_12324,N_11256,N_11871);
or U12325 (N_12325,N_11919,N_11984);
nand U12326 (N_12326,N_11859,N_11328);
nand U12327 (N_12327,N_11396,N_11676);
and U12328 (N_12328,N_11294,N_11342);
nand U12329 (N_12329,N_11760,N_11355);
nand U12330 (N_12330,N_11309,N_11988);
nor U12331 (N_12331,N_11843,N_11959);
or U12332 (N_12332,N_11267,N_11409);
nor U12333 (N_12333,N_11292,N_11600);
and U12334 (N_12334,N_11304,N_11636);
or U12335 (N_12335,N_11295,N_11620);
nor U12336 (N_12336,N_11397,N_11767);
nor U12337 (N_12337,N_11931,N_11751);
or U12338 (N_12338,N_11800,N_11462);
or U12339 (N_12339,N_11690,N_11506);
nor U12340 (N_12340,N_11407,N_11593);
or U12341 (N_12341,N_11687,N_11685);
nand U12342 (N_12342,N_11384,N_11633);
nor U12343 (N_12343,N_11711,N_11487);
and U12344 (N_12344,N_11310,N_11743);
xor U12345 (N_12345,N_11852,N_11456);
nand U12346 (N_12346,N_11778,N_11613);
and U12347 (N_12347,N_11733,N_11579);
or U12348 (N_12348,N_11282,N_11509);
or U12349 (N_12349,N_11698,N_11945);
and U12350 (N_12350,N_11463,N_11695);
or U12351 (N_12351,N_11467,N_11954);
and U12352 (N_12352,N_11840,N_11757);
nand U12353 (N_12353,N_11426,N_11719);
nand U12354 (N_12354,N_11359,N_11405);
and U12355 (N_12355,N_11300,N_11703);
and U12356 (N_12356,N_11896,N_11510);
and U12357 (N_12357,N_11541,N_11699);
or U12358 (N_12358,N_11700,N_11813);
and U12359 (N_12359,N_11293,N_11771);
nand U12360 (N_12360,N_11689,N_11627);
xnor U12361 (N_12361,N_11515,N_11601);
nor U12362 (N_12362,N_11980,N_11811);
and U12363 (N_12363,N_11497,N_11802);
nor U12364 (N_12364,N_11312,N_11786);
and U12365 (N_12365,N_11284,N_11455);
nor U12366 (N_12366,N_11290,N_11804);
or U12367 (N_12367,N_11496,N_11482);
nand U12368 (N_12368,N_11918,N_11855);
and U12369 (N_12369,N_11826,N_11604);
nor U12370 (N_12370,N_11460,N_11841);
nor U12371 (N_12371,N_11285,N_11428);
nor U12372 (N_12372,N_11265,N_11847);
or U12373 (N_12373,N_11318,N_11969);
or U12374 (N_12374,N_11894,N_11324);
and U12375 (N_12375,N_11745,N_11514);
nand U12376 (N_12376,N_11256,N_11806);
nor U12377 (N_12377,N_11754,N_11399);
nand U12378 (N_12378,N_11337,N_11643);
and U12379 (N_12379,N_11389,N_11282);
or U12380 (N_12380,N_11953,N_11502);
nand U12381 (N_12381,N_11676,N_11717);
nand U12382 (N_12382,N_11956,N_11978);
or U12383 (N_12383,N_11563,N_11810);
and U12384 (N_12384,N_11410,N_11926);
nand U12385 (N_12385,N_11429,N_11766);
or U12386 (N_12386,N_11502,N_11555);
xnor U12387 (N_12387,N_11872,N_11833);
or U12388 (N_12388,N_11736,N_11654);
nor U12389 (N_12389,N_11333,N_11486);
nor U12390 (N_12390,N_11726,N_11814);
and U12391 (N_12391,N_11899,N_11761);
nor U12392 (N_12392,N_11584,N_11866);
and U12393 (N_12393,N_11639,N_11511);
or U12394 (N_12394,N_11878,N_11812);
nand U12395 (N_12395,N_11432,N_11679);
and U12396 (N_12396,N_11832,N_11537);
or U12397 (N_12397,N_11545,N_11367);
and U12398 (N_12398,N_11888,N_11280);
or U12399 (N_12399,N_11272,N_11782);
nand U12400 (N_12400,N_11816,N_11600);
and U12401 (N_12401,N_11566,N_11558);
nand U12402 (N_12402,N_11460,N_11944);
xor U12403 (N_12403,N_11821,N_11359);
nand U12404 (N_12404,N_11815,N_11527);
nor U12405 (N_12405,N_11819,N_11334);
or U12406 (N_12406,N_11692,N_11973);
nand U12407 (N_12407,N_11321,N_11883);
and U12408 (N_12408,N_11250,N_11452);
or U12409 (N_12409,N_11897,N_11928);
nand U12410 (N_12410,N_11284,N_11555);
xor U12411 (N_12411,N_11615,N_11689);
or U12412 (N_12412,N_11941,N_11774);
nand U12413 (N_12413,N_11390,N_11571);
nand U12414 (N_12414,N_11744,N_11356);
and U12415 (N_12415,N_11569,N_11706);
xnor U12416 (N_12416,N_11770,N_11530);
nand U12417 (N_12417,N_11801,N_11346);
and U12418 (N_12418,N_11999,N_11331);
xnor U12419 (N_12419,N_11667,N_11524);
nor U12420 (N_12420,N_11762,N_11896);
and U12421 (N_12421,N_11477,N_11906);
nand U12422 (N_12422,N_11656,N_11324);
nor U12423 (N_12423,N_11707,N_11759);
nand U12424 (N_12424,N_11759,N_11494);
and U12425 (N_12425,N_11997,N_11279);
and U12426 (N_12426,N_11886,N_11803);
nor U12427 (N_12427,N_11391,N_11848);
and U12428 (N_12428,N_11537,N_11937);
and U12429 (N_12429,N_11516,N_11577);
nand U12430 (N_12430,N_11270,N_11948);
or U12431 (N_12431,N_11875,N_11665);
xor U12432 (N_12432,N_11638,N_11469);
and U12433 (N_12433,N_11874,N_11958);
nand U12434 (N_12434,N_11264,N_11406);
and U12435 (N_12435,N_11598,N_11985);
xor U12436 (N_12436,N_11403,N_11542);
nor U12437 (N_12437,N_11389,N_11961);
or U12438 (N_12438,N_11786,N_11918);
xnor U12439 (N_12439,N_11823,N_11257);
or U12440 (N_12440,N_11879,N_11652);
nand U12441 (N_12441,N_11997,N_11407);
and U12442 (N_12442,N_11797,N_11470);
and U12443 (N_12443,N_11541,N_11556);
nand U12444 (N_12444,N_11826,N_11273);
nand U12445 (N_12445,N_11391,N_11804);
xor U12446 (N_12446,N_11577,N_11649);
and U12447 (N_12447,N_11833,N_11477);
nor U12448 (N_12448,N_11484,N_11275);
and U12449 (N_12449,N_11653,N_11436);
xor U12450 (N_12450,N_11663,N_11474);
and U12451 (N_12451,N_11537,N_11391);
nor U12452 (N_12452,N_11592,N_11411);
and U12453 (N_12453,N_11259,N_11700);
and U12454 (N_12454,N_11976,N_11464);
nor U12455 (N_12455,N_11281,N_11999);
nor U12456 (N_12456,N_11599,N_11413);
xor U12457 (N_12457,N_11636,N_11286);
or U12458 (N_12458,N_11798,N_11849);
and U12459 (N_12459,N_11955,N_11482);
xnor U12460 (N_12460,N_11955,N_11481);
nand U12461 (N_12461,N_11940,N_11414);
nand U12462 (N_12462,N_11851,N_11643);
or U12463 (N_12463,N_11320,N_11626);
or U12464 (N_12464,N_11261,N_11927);
and U12465 (N_12465,N_11894,N_11429);
or U12466 (N_12466,N_11754,N_11327);
nand U12467 (N_12467,N_11562,N_11812);
nor U12468 (N_12468,N_11445,N_11635);
nor U12469 (N_12469,N_11867,N_11472);
and U12470 (N_12470,N_11592,N_11301);
or U12471 (N_12471,N_11252,N_11423);
nor U12472 (N_12472,N_11549,N_11607);
nor U12473 (N_12473,N_11775,N_11472);
and U12474 (N_12474,N_11471,N_11715);
and U12475 (N_12475,N_11694,N_11327);
nor U12476 (N_12476,N_11836,N_11991);
nand U12477 (N_12477,N_11350,N_11739);
or U12478 (N_12478,N_11350,N_11728);
nor U12479 (N_12479,N_11937,N_11501);
nor U12480 (N_12480,N_11533,N_11933);
nand U12481 (N_12481,N_11776,N_11542);
and U12482 (N_12482,N_11738,N_11769);
nor U12483 (N_12483,N_11830,N_11255);
or U12484 (N_12484,N_11557,N_11779);
and U12485 (N_12485,N_11887,N_11759);
nand U12486 (N_12486,N_11544,N_11492);
xnor U12487 (N_12487,N_11959,N_11859);
or U12488 (N_12488,N_11523,N_11346);
xor U12489 (N_12489,N_11865,N_11545);
or U12490 (N_12490,N_11642,N_11351);
or U12491 (N_12491,N_11337,N_11956);
and U12492 (N_12492,N_11688,N_11854);
xor U12493 (N_12493,N_11814,N_11600);
or U12494 (N_12494,N_11660,N_11954);
and U12495 (N_12495,N_11469,N_11333);
and U12496 (N_12496,N_11398,N_11453);
nand U12497 (N_12497,N_11887,N_11769);
and U12498 (N_12498,N_11455,N_11936);
or U12499 (N_12499,N_11988,N_11467);
and U12500 (N_12500,N_11674,N_11582);
or U12501 (N_12501,N_11438,N_11439);
or U12502 (N_12502,N_11907,N_11956);
or U12503 (N_12503,N_11806,N_11595);
and U12504 (N_12504,N_11359,N_11836);
nand U12505 (N_12505,N_11314,N_11666);
and U12506 (N_12506,N_11742,N_11706);
or U12507 (N_12507,N_11910,N_11881);
nand U12508 (N_12508,N_11888,N_11277);
nor U12509 (N_12509,N_11488,N_11458);
and U12510 (N_12510,N_11984,N_11321);
nor U12511 (N_12511,N_11933,N_11775);
and U12512 (N_12512,N_11426,N_11481);
nor U12513 (N_12513,N_11850,N_11317);
and U12514 (N_12514,N_11962,N_11922);
and U12515 (N_12515,N_11778,N_11984);
or U12516 (N_12516,N_11471,N_11509);
nor U12517 (N_12517,N_11522,N_11690);
or U12518 (N_12518,N_11278,N_11404);
or U12519 (N_12519,N_11695,N_11827);
nor U12520 (N_12520,N_11342,N_11590);
or U12521 (N_12521,N_11915,N_11560);
nor U12522 (N_12522,N_11724,N_11555);
nand U12523 (N_12523,N_11372,N_11891);
or U12524 (N_12524,N_11329,N_11758);
nand U12525 (N_12525,N_11331,N_11304);
or U12526 (N_12526,N_11488,N_11757);
and U12527 (N_12527,N_11893,N_11804);
and U12528 (N_12528,N_11743,N_11516);
nand U12529 (N_12529,N_11727,N_11426);
nor U12530 (N_12530,N_11713,N_11907);
or U12531 (N_12531,N_11710,N_11331);
or U12532 (N_12532,N_11630,N_11399);
nor U12533 (N_12533,N_11854,N_11783);
or U12534 (N_12534,N_11269,N_11446);
xnor U12535 (N_12535,N_11958,N_11262);
xor U12536 (N_12536,N_11961,N_11412);
xor U12537 (N_12537,N_11889,N_11378);
nand U12538 (N_12538,N_11704,N_11325);
and U12539 (N_12539,N_11851,N_11615);
nand U12540 (N_12540,N_11715,N_11545);
nand U12541 (N_12541,N_11939,N_11518);
or U12542 (N_12542,N_11566,N_11284);
xor U12543 (N_12543,N_11562,N_11513);
nor U12544 (N_12544,N_11932,N_11848);
nand U12545 (N_12545,N_11808,N_11774);
and U12546 (N_12546,N_11394,N_11541);
xnor U12547 (N_12547,N_11994,N_11711);
nand U12548 (N_12548,N_11557,N_11768);
xor U12549 (N_12549,N_11795,N_11815);
xnor U12550 (N_12550,N_11294,N_11768);
nand U12551 (N_12551,N_11854,N_11793);
or U12552 (N_12552,N_11506,N_11983);
or U12553 (N_12553,N_11272,N_11430);
nand U12554 (N_12554,N_11420,N_11936);
or U12555 (N_12555,N_11268,N_11594);
nor U12556 (N_12556,N_11280,N_11752);
and U12557 (N_12557,N_11758,N_11845);
and U12558 (N_12558,N_11540,N_11405);
nor U12559 (N_12559,N_11884,N_11876);
nor U12560 (N_12560,N_11907,N_11941);
nand U12561 (N_12561,N_11554,N_11835);
or U12562 (N_12562,N_11473,N_11260);
nand U12563 (N_12563,N_11530,N_11872);
nand U12564 (N_12564,N_11542,N_11308);
nand U12565 (N_12565,N_11815,N_11464);
nor U12566 (N_12566,N_11922,N_11874);
and U12567 (N_12567,N_11484,N_11678);
and U12568 (N_12568,N_11934,N_11263);
nand U12569 (N_12569,N_11966,N_11417);
nand U12570 (N_12570,N_11898,N_11799);
nand U12571 (N_12571,N_11439,N_11433);
or U12572 (N_12572,N_11771,N_11902);
or U12573 (N_12573,N_11455,N_11371);
nor U12574 (N_12574,N_11663,N_11768);
or U12575 (N_12575,N_11582,N_11727);
xnor U12576 (N_12576,N_11698,N_11378);
xnor U12577 (N_12577,N_11726,N_11423);
and U12578 (N_12578,N_11598,N_11624);
nor U12579 (N_12579,N_11533,N_11275);
nand U12580 (N_12580,N_11250,N_11274);
nor U12581 (N_12581,N_11847,N_11445);
nand U12582 (N_12582,N_11737,N_11276);
and U12583 (N_12583,N_11860,N_11772);
nand U12584 (N_12584,N_11744,N_11658);
or U12585 (N_12585,N_11496,N_11253);
nor U12586 (N_12586,N_11862,N_11855);
or U12587 (N_12587,N_11739,N_11661);
nor U12588 (N_12588,N_11777,N_11441);
nor U12589 (N_12589,N_11362,N_11939);
nand U12590 (N_12590,N_11324,N_11968);
nand U12591 (N_12591,N_11639,N_11760);
nor U12592 (N_12592,N_11399,N_11855);
or U12593 (N_12593,N_11321,N_11370);
or U12594 (N_12594,N_11831,N_11683);
nor U12595 (N_12595,N_11900,N_11313);
nor U12596 (N_12596,N_11551,N_11459);
and U12597 (N_12597,N_11996,N_11773);
nor U12598 (N_12598,N_11759,N_11904);
nand U12599 (N_12599,N_11570,N_11746);
and U12600 (N_12600,N_11565,N_11489);
nand U12601 (N_12601,N_11705,N_11772);
nor U12602 (N_12602,N_11785,N_11532);
xor U12603 (N_12603,N_11803,N_11702);
nand U12604 (N_12604,N_11528,N_11462);
nand U12605 (N_12605,N_11952,N_11450);
nor U12606 (N_12606,N_11349,N_11762);
or U12607 (N_12607,N_11408,N_11672);
or U12608 (N_12608,N_11802,N_11872);
xor U12609 (N_12609,N_11353,N_11905);
nor U12610 (N_12610,N_11913,N_11442);
nand U12611 (N_12611,N_11317,N_11916);
nand U12612 (N_12612,N_11482,N_11329);
nand U12613 (N_12613,N_11388,N_11342);
and U12614 (N_12614,N_11968,N_11274);
and U12615 (N_12615,N_11605,N_11494);
and U12616 (N_12616,N_11546,N_11410);
nor U12617 (N_12617,N_11663,N_11469);
nand U12618 (N_12618,N_11334,N_11647);
or U12619 (N_12619,N_11393,N_11321);
and U12620 (N_12620,N_11798,N_11579);
and U12621 (N_12621,N_11692,N_11769);
nor U12622 (N_12622,N_11428,N_11328);
or U12623 (N_12623,N_11922,N_11319);
or U12624 (N_12624,N_11841,N_11291);
and U12625 (N_12625,N_11521,N_11545);
nand U12626 (N_12626,N_11567,N_11921);
xor U12627 (N_12627,N_11419,N_11472);
nor U12628 (N_12628,N_11481,N_11504);
nand U12629 (N_12629,N_11600,N_11406);
and U12630 (N_12630,N_11514,N_11650);
nor U12631 (N_12631,N_11374,N_11369);
and U12632 (N_12632,N_11759,N_11938);
nand U12633 (N_12633,N_11976,N_11458);
and U12634 (N_12634,N_11297,N_11592);
xor U12635 (N_12635,N_11297,N_11418);
or U12636 (N_12636,N_11499,N_11632);
nor U12637 (N_12637,N_11414,N_11534);
nand U12638 (N_12638,N_11657,N_11282);
or U12639 (N_12639,N_11357,N_11827);
nand U12640 (N_12640,N_11507,N_11823);
and U12641 (N_12641,N_11777,N_11944);
and U12642 (N_12642,N_11942,N_11556);
and U12643 (N_12643,N_11277,N_11948);
or U12644 (N_12644,N_11773,N_11554);
nand U12645 (N_12645,N_11688,N_11394);
nor U12646 (N_12646,N_11449,N_11310);
nand U12647 (N_12647,N_11826,N_11421);
xnor U12648 (N_12648,N_11895,N_11402);
nor U12649 (N_12649,N_11750,N_11899);
nor U12650 (N_12650,N_11389,N_11832);
nor U12651 (N_12651,N_11402,N_11430);
xnor U12652 (N_12652,N_11655,N_11347);
nand U12653 (N_12653,N_11887,N_11909);
nand U12654 (N_12654,N_11538,N_11980);
nand U12655 (N_12655,N_11878,N_11493);
nand U12656 (N_12656,N_11391,N_11842);
or U12657 (N_12657,N_11617,N_11942);
nand U12658 (N_12658,N_11815,N_11433);
nand U12659 (N_12659,N_11767,N_11654);
and U12660 (N_12660,N_11765,N_11385);
and U12661 (N_12661,N_11976,N_11865);
nand U12662 (N_12662,N_11821,N_11355);
nor U12663 (N_12663,N_11256,N_11359);
and U12664 (N_12664,N_11336,N_11888);
or U12665 (N_12665,N_11621,N_11548);
and U12666 (N_12666,N_11961,N_11879);
and U12667 (N_12667,N_11729,N_11801);
xor U12668 (N_12668,N_11855,N_11539);
nand U12669 (N_12669,N_11904,N_11764);
and U12670 (N_12670,N_11422,N_11652);
nor U12671 (N_12671,N_11700,N_11419);
xor U12672 (N_12672,N_11571,N_11380);
or U12673 (N_12673,N_11765,N_11324);
nor U12674 (N_12674,N_11797,N_11724);
and U12675 (N_12675,N_11871,N_11923);
and U12676 (N_12676,N_11642,N_11279);
or U12677 (N_12677,N_11905,N_11574);
nor U12678 (N_12678,N_11723,N_11842);
and U12679 (N_12679,N_11410,N_11918);
nor U12680 (N_12680,N_11839,N_11607);
nor U12681 (N_12681,N_11370,N_11803);
xor U12682 (N_12682,N_11646,N_11422);
or U12683 (N_12683,N_11730,N_11257);
nand U12684 (N_12684,N_11502,N_11889);
nand U12685 (N_12685,N_11729,N_11537);
nor U12686 (N_12686,N_11267,N_11920);
nor U12687 (N_12687,N_11678,N_11413);
nand U12688 (N_12688,N_11579,N_11819);
nor U12689 (N_12689,N_11931,N_11622);
nor U12690 (N_12690,N_11989,N_11948);
nand U12691 (N_12691,N_11786,N_11277);
and U12692 (N_12692,N_11410,N_11738);
nor U12693 (N_12693,N_11910,N_11269);
or U12694 (N_12694,N_11945,N_11857);
and U12695 (N_12695,N_11435,N_11538);
nor U12696 (N_12696,N_11843,N_11421);
or U12697 (N_12697,N_11395,N_11468);
nor U12698 (N_12698,N_11771,N_11273);
or U12699 (N_12699,N_11876,N_11359);
nand U12700 (N_12700,N_11500,N_11713);
and U12701 (N_12701,N_11540,N_11682);
nor U12702 (N_12702,N_11398,N_11290);
or U12703 (N_12703,N_11439,N_11376);
or U12704 (N_12704,N_11729,N_11547);
and U12705 (N_12705,N_11462,N_11365);
or U12706 (N_12706,N_11612,N_11866);
and U12707 (N_12707,N_11266,N_11690);
or U12708 (N_12708,N_11582,N_11657);
or U12709 (N_12709,N_11508,N_11411);
nand U12710 (N_12710,N_11887,N_11471);
nand U12711 (N_12711,N_11778,N_11597);
nor U12712 (N_12712,N_11784,N_11802);
or U12713 (N_12713,N_11482,N_11679);
nor U12714 (N_12714,N_11854,N_11498);
nand U12715 (N_12715,N_11513,N_11664);
or U12716 (N_12716,N_11613,N_11653);
and U12717 (N_12717,N_11871,N_11483);
nor U12718 (N_12718,N_11518,N_11413);
or U12719 (N_12719,N_11797,N_11363);
xnor U12720 (N_12720,N_11683,N_11305);
or U12721 (N_12721,N_11850,N_11684);
nand U12722 (N_12722,N_11668,N_11696);
or U12723 (N_12723,N_11657,N_11277);
xor U12724 (N_12724,N_11606,N_11735);
nand U12725 (N_12725,N_11256,N_11267);
nor U12726 (N_12726,N_11797,N_11542);
nand U12727 (N_12727,N_11449,N_11461);
and U12728 (N_12728,N_11475,N_11765);
xnor U12729 (N_12729,N_11408,N_11603);
and U12730 (N_12730,N_11660,N_11944);
nand U12731 (N_12731,N_11465,N_11993);
xnor U12732 (N_12732,N_11447,N_11493);
and U12733 (N_12733,N_11835,N_11253);
or U12734 (N_12734,N_11830,N_11893);
nand U12735 (N_12735,N_11250,N_11304);
nor U12736 (N_12736,N_11606,N_11403);
and U12737 (N_12737,N_11930,N_11805);
nor U12738 (N_12738,N_11915,N_11266);
xor U12739 (N_12739,N_11553,N_11558);
nand U12740 (N_12740,N_11446,N_11829);
nor U12741 (N_12741,N_11549,N_11421);
nand U12742 (N_12742,N_11278,N_11627);
and U12743 (N_12743,N_11671,N_11485);
xor U12744 (N_12744,N_11874,N_11349);
nand U12745 (N_12745,N_11955,N_11992);
or U12746 (N_12746,N_11892,N_11371);
nor U12747 (N_12747,N_11517,N_11514);
or U12748 (N_12748,N_11558,N_11377);
or U12749 (N_12749,N_11571,N_11711);
or U12750 (N_12750,N_12182,N_12693);
or U12751 (N_12751,N_12365,N_12039);
or U12752 (N_12752,N_12421,N_12580);
nand U12753 (N_12753,N_12400,N_12438);
and U12754 (N_12754,N_12196,N_12246);
and U12755 (N_12755,N_12640,N_12709);
nor U12756 (N_12756,N_12096,N_12689);
nor U12757 (N_12757,N_12407,N_12243);
nor U12758 (N_12758,N_12467,N_12167);
nor U12759 (N_12759,N_12489,N_12075);
and U12760 (N_12760,N_12569,N_12229);
or U12761 (N_12761,N_12054,N_12221);
or U12762 (N_12762,N_12244,N_12117);
nand U12763 (N_12763,N_12644,N_12639);
nor U12764 (N_12764,N_12195,N_12727);
xnor U12765 (N_12765,N_12710,N_12017);
or U12766 (N_12766,N_12323,N_12216);
or U12767 (N_12767,N_12366,N_12690);
or U12768 (N_12768,N_12070,N_12735);
and U12769 (N_12769,N_12386,N_12086);
or U12770 (N_12770,N_12416,N_12642);
nand U12771 (N_12771,N_12480,N_12240);
nand U12772 (N_12772,N_12695,N_12312);
xor U12773 (N_12773,N_12171,N_12277);
nand U12774 (N_12774,N_12413,N_12140);
and U12775 (N_12775,N_12013,N_12372);
xnor U12776 (N_12776,N_12295,N_12543);
nand U12777 (N_12777,N_12576,N_12278);
nor U12778 (N_12778,N_12652,N_12211);
nand U12779 (N_12779,N_12354,N_12322);
and U12780 (N_12780,N_12739,N_12414);
nor U12781 (N_12781,N_12577,N_12311);
or U12782 (N_12782,N_12090,N_12380);
or U12783 (N_12783,N_12687,N_12160);
and U12784 (N_12784,N_12135,N_12628);
nand U12785 (N_12785,N_12335,N_12749);
and U12786 (N_12786,N_12499,N_12383);
nand U12787 (N_12787,N_12236,N_12044);
or U12788 (N_12788,N_12494,N_12447);
nor U12789 (N_12789,N_12694,N_12194);
or U12790 (N_12790,N_12597,N_12052);
or U12791 (N_12791,N_12342,N_12641);
nand U12792 (N_12792,N_12152,N_12225);
nand U12793 (N_12793,N_12622,N_12495);
or U12794 (N_12794,N_12223,N_12742);
nor U12795 (N_12795,N_12179,N_12053);
nand U12796 (N_12796,N_12371,N_12344);
nor U12797 (N_12797,N_12014,N_12566);
and U12798 (N_12798,N_12638,N_12536);
or U12799 (N_12799,N_12190,N_12439);
or U12800 (N_12800,N_12479,N_12591);
nand U12801 (N_12801,N_12363,N_12408);
nand U12802 (N_12802,N_12058,N_12581);
and U12803 (N_12803,N_12381,N_12219);
and U12804 (N_12804,N_12538,N_12614);
and U12805 (N_12805,N_12074,N_12304);
nor U12806 (N_12806,N_12141,N_12517);
or U12807 (N_12807,N_12247,N_12401);
nor U12808 (N_12808,N_12301,N_12481);
nand U12809 (N_12809,N_12071,N_12012);
xor U12810 (N_12810,N_12526,N_12426);
nand U12811 (N_12811,N_12588,N_12065);
nand U12812 (N_12812,N_12136,N_12392);
or U12813 (N_12813,N_12422,N_12567);
nor U12814 (N_12814,N_12001,N_12706);
or U12815 (N_12815,N_12209,N_12121);
nor U12816 (N_12816,N_12298,N_12393);
or U12817 (N_12817,N_12450,N_12748);
xnor U12818 (N_12818,N_12570,N_12395);
nand U12819 (N_12819,N_12181,N_12037);
nor U12820 (N_12820,N_12169,N_12154);
and U12821 (N_12821,N_12064,N_12230);
nor U12822 (N_12822,N_12725,N_12453);
and U12823 (N_12823,N_12271,N_12255);
or U12824 (N_12824,N_12305,N_12189);
nor U12825 (N_12825,N_12003,N_12329);
and U12826 (N_12826,N_12726,N_12267);
and U12827 (N_12827,N_12069,N_12505);
nand U12828 (N_12828,N_12470,N_12062);
or U12829 (N_12829,N_12680,N_12732);
or U12830 (N_12830,N_12532,N_12704);
nand U12831 (N_12831,N_12529,N_12143);
nor U12832 (N_12832,N_12620,N_12006);
or U12833 (N_12833,N_12463,N_12523);
nand U12834 (N_12834,N_12343,N_12428);
nor U12835 (N_12835,N_12712,N_12441);
xor U12836 (N_12836,N_12516,N_12242);
xnor U12837 (N_12837,N_12585,N_12681);
xor U12838 (N_12838,N_12034,N_12382);
and U12839 (N_12839,N_12207,N_12296);
or U12840 (N_12840,N_12430,N_12351);
xnor U12841 (N_12841,N_12515,N_12276);
nand U12842 (N_12842,N_12369,N_12410);
and U12843 (N_12843,N_12418,N_12518);
nand U12844 (N_12844,N_12352,N_12485);
nor U12845 (N_12845,N_12056,N_12741);
xnor U12846 (N_12846,N_12434,N_12227);
nor U12847 (N_12847,N_12707,N_12708);
and U12848 (N_12848,N_12718,N_12653);
xor U12849 (N_12849,N_12320,N_12579);
and U12850 (N_12850,N_12294,N_12367);
and U12851 (N_12851,N_12153,N_12284);
and U12852 (N_12852,N_12405,N_12126);
or U12853 (N_12853,N_12389,N_12297);
xor U12854 (N_12854,N_12613,N_12004);
nand U12855 (N_12855,N_12107,N_12457);
xnor U12856 (N_12856,N_12192,N_12662);
nor U12857 (N_12857,N_12593,N_12101);
and U12858 (N_12858,N_12250,N_12161);
and U12859 (N_12859,N_12024,N_12714);
and U12860 (N_12860,N_12604,N_12539);
or U12861 (N_12861,N_12172,N_12345);
nor U12862 (N_12862,N_12292,N_12321);
nor U12863 (N_12863,N_12643,N_12509);
or U12864 (N_12864,N_12645,N_12347);
or U12865 (N_12865,N_12715,N_12258);
and U12866 (N_12866,N_12130,N_12289);
and U12867 (N_12867,N_12089,N_12477);
nor U12868 (N_12868,N_12719,N_12656);
nor U12869 (N_12869,N_12688,N_12098);
nor U12870 (N_12870,N_12226,N_12487);
xnor U12871 (N_12871,N_12616,N_12631);
and U12872 (N_12872,N_12233,N_12370);
and U12873 (N_12873,N_12600,N_12299);
xor U12874 (N_12874,N_12185,N_12562);
and U12875 (N_12875,N_12699,N_12376);
xnor U12876 (N_12876,N_12568,N_12711);
and U12877 (N_12877,N_12474,N_12429);
and U12878 (N_12878,N_12455,N_12435);
xnor U12879 (N_12879,N_12549,N_12164);
xor U12880 (N_12880,N_12578,N_12647);
nand U12881 (N_12881,N_12602,N_12026);
xor U12882 (N_12882,N_12397,N_12286);
and U12883 (N_12883,N_12498,N_12103);
nand U12884 (N_12884,N_12125,N_12235);
or U12885 (N_12885,N_12419,N_12521);
or U12886 (N_12886,N_12609,N_12355);
xnor U12887 (N_12887,N_12059,N_12658);
or U12888 (N_12888,N_12083,N_12184);
or U12889 (N_12889,N_12358,N_12350);
and U12890 (N_12890,N_12346,N_12599);
nor U12891 (N_12891,N_12624,N_12092);
nor U12892 (N_12892,N_12050,N_12134);
and U12893 (N_12893,N_12519,N_12049);
or U12894 (N_12894,N_12073,N_12348);
nor U12895 (N_12895,N_12398,N_12374);
nor U12896 (N_12896,N_12176,N_12402);
or U12897 (N_12897,N_12565,N_12678);
and U12898 (N_12898,N_12551,N_12700);
and U12899 (N_12899,N_12334,N_12068);
and U12900 (N_12900,N_12105,N_12476);
and U12901 (N_12901,N_12210,N_12066);
and U12902 (N_12902,N_12032,N_12239);
or U12903 (N_12903,N_12091,N_12657);
or U12904 (N_12904,N_12087,N_12492);
nor U12905 (N_12905,N_12288,N_12061);
nor U12906 (N_12906,N_12603,N_12731);
and U12907 (N_12907,N_12046,N_12208);
or U12908 (N_12908,N_12723,N_12260);
and U12909 (N_12909,N_12610,N_12635);
nand U12910 (N_12910,N_12452,N_12472);
nor U12911 (N_12911,N_12559,N_12215);
and U12912 (N_12912,N_12633,N_12282);
nand U12913 (N_12913,N_12275,N_12461);
xnor U12914 (N_12914,N_12145,N_12333);
and U12915 (N_12915,N_12630,N_12033);
nor U12916 (N_12916,N_12387,N_12394);
nor U12917 (N_12917,N_12595,N_12510);
nor U12918 (N_12918,N_12142,N_12571);
and U12919 (N_12919,N_12331,N_12500);
nor U12920 (N_12920,N_12019,N_12200);
or U12921 (N_12921,N_12637,N_12425);
and U12922 (N_12922,N_12078,N_12448);
and U12923 (N_12923,N_12212,N_12406);
xnor U12924 (N_12924,N_12738,N_12676);
nand U12925 (N_12925,N_12608,N_12665);
or U12926 (N_12926,N_12253,N_12116);
nor U12927 (N_12927,N_12632,N_12097);
nor U12928 (N_12928,N_12390,N_12100);
and U12929 (N_12929,N_12546,N_12507);
xor U12930 (N_12930,N_12224,N_12303);
nor U12931 (N_12931,N_12378,N_12466);
xor U12932 (N_12932,N_12646,N_12651);
and U12933 (N_12933,N_12339,N_12318);
or U12934 (N_12934,N_12490,N_12206);
or U12935 (N_12935,N_12664,N_12133);
and U12936 (N_12936,N_12486,N_12512);
and U12937 (N_12937,N_12548,N_12468);
xnor U12938 (N_12938,N_12677,N_12259);
nand U12939 (N_12939,N_12205,N_12005);
or U12940 (N_12940,N_12057,N_12574);
and U12941 (N_12941,N_12533,N_12237);
and U12942 (N_12942,N_12084,N_12621);
or U12943 (N_12943,N_12491,N_12550);
nor U12944 (N_12944,N_12541,N_12668);
xnor U12945 (N_12945,N_12148,N_12112);
or U12946 (N_12946,N_12745,N_12048);
nor U12947 (N_12947,N_12252,N_12018);
and U12948 (N_12948,N_12552,N_12248);
nor U12949 (N_12949,N_12021,N_12131);
nand U12950 (N_12950,N_12332,N_12445);
nor U12951 (N_12951,N_12623,N_12409);
and U12952 (N_12952,N_12129,N_12627);
nor U12953 (N_12953,N_12040,N_12330);
xor U12954 (N_12954,N_12222,N_12666);
nand U12955 (N_12955,N_12138,N_12349);
xor U12956 (N_12956,N_12264,N_12340);
or U12957 (N_12957,N_12634,N_12009);
nand U12958 (N_12958,N_12093,N_12031);
and U12959 (N_12959,N_12488,N_12612);
nand U12960 (N_12960,N_12188,N_12478);
nor U12961 (N_12961,N_12314,N_12213);
and U12962 (N_12962,N_12482,N_12473);
xor U12963 (N_12963,N_12572,N_12307);
xnor U12964 (N_12964,N_12177,N_12265);
or U12965 (N_12965,N_12669,N_12234);
nor U12966 (N_12966,N_12217,N_12263);
nor U12967 (N_12967,N_12460,N_12442);
nand U12968 (N_12968,N_12674,N_12396);
nor U12969 (N_12969,N_12325,N_12415);
and U12970 (N_12970,N_12615,N_12589);
nor U12971 (N_12971,N_12673,N_12175);
and U12972 (N_12972,N_12022,N_12611);
nor U12973 (N_12973,N_12557,N_12186);
nor U12974 (N_12974,N_12016,N_12156);
nor U12975 (N_12975,N_12436,N_12456);
or U12976 (N_12976,N_12251,N_12683);
or U12977 (N_12977,N_12734,N_12684);
nor U12978 (N_12978,N_12041,N_12283);
nand U12979 (N_12979,N_12232,N_12147);
and U12980 (N_12980,N_12051,N_12081);
nand U12981 (N_12981,N_12174,N_12535);
nand U12982 (N_12982,N_12015,N_12508);
nor U12983 (N_12983,N_12137,N_12203);
and U12984 (N_12984,N_12660,N_12261);
nor U12985 (N_12985,N_12537,N_12170);
and U12986 (N_12986,N_12679,N_12705);
nand U12987 (N_12987,N_12183,N_12391);
nor U12988 (N_12988,N_12558,N_12420);
and U12989 (N_12989,N_12564,N_12357);
nor U12990 (N_12990,N_12454,N_12178);
and U12991 (N_12991,N_12113,N_12173);
nand U12992 (N_12992,N_12446,N_12555);
nand U12993 (N_12993,N_12360,N_12262);
or U12994 (N_12994,N_12290,N_12404);
nand U12995 (N_12995,N_12029,N_12379);
nor U12996 (N_12996,N_12440,N_12055);
nor U12997 (N_12997,N_12503,N_12327);
nand U12998 (N_12998,N_12035,N_12661);
and U12999 (N_12999,N_12109,N_12736);
or U13000 (N_13000,N_12522,N_12010);
or U13001 (N_13001,N_12285,N_12554);
and U13002 (N_13002,N_12682,N_12531);
and U13003 (N_13003,N_12636,N_12513);
nor U13004 (N_13004,N_12716,N_12095);
or U13005 (N_13005,N_12218,N_12431);
or U13006 (N_13006,N_12118,N_12204);
nor U13007 (N_13007,N_12724,N_12362);
and U13008 (N_13008,N_12659,N_12165);
and U13009 (N_13009,N_12520,N_12123);
xnor U13010 (N_13010,N_12654,N_12493);
and U13011 (N_13011,N_12746,N_12269);
nor U13012 (N_13012,N_12341,N_12720);
and U13013 (N_13013,N_12146,N_12228);
or U13014 (N_13014,N_12128,N_12080);
or U13015 (N_13015,N_12692,N_12459);
nor U13016 (N_13016,N_12256,N_12155);
and U13017 (N_13017,N_12427,N_12601);
nor U13018 (N_13018,N_12308,N_12249);
nand U13019 (N_13019,N_12702,N_12036);
xnor U13020 (N_13020,N_12592,N_12563);
nor U13021 (N_13021,N_12721,N_12011);
and U13022 (N_13022,N_12002,N_12686);
or U13023 (N_13023,N_12744,N_12245);
xor U13024 (N_13024,N_12045,N_12309);
xnor U13025 (N_13025,N_12497,N_12703);
and U13026 (N_13026,N_12027,N_12675);
and U13027 (N_13027,N_12619,N_12424);
nand U13028 (N_13028,N_12663,N_12443);
or U13029 (N_13029,N_12545,N_12586);
nand U13030 (N_13030,N_12149,N_12291);
or U13031 (N_13031,N_12399,N_12617);
and U13032 (N_13032,N_12279,N_12085);
and U13033 (N_13033,N_12475,N_12544);
or U13034 (N_13034,N_12698,N_12444);
nor U13035 (N_13035,N_12079,N_12722);
nand U13036 (N_13036,N_12368,N_12671);
or U13037 (N_13037,N_12582,N_12302);
and U13038 (N_13038,N_12306,N_12655);
and U13039 (N_13039,N_12484,N_12587);
nand U13040 (N_13040,N_12697,N_12102);
nand U13041 (N_13041,N_12583,N_12496);
and U13042 (N_13042,N_12120,N_12238);
or U13043 (N_13043,N_12534,N_12626);
nor U13044 (N_13044,N_12462,N_12573);
and U13045 (N_13045,N_12038,N_12605);
xnor U13046 (N_13046,N_12257,N_12127);
or U13047 (N_13047,N_12353,N_12685);
or U13048 (N_13048,N_12596,N_12007);
nor U13049 (N_13049,N_12575,N_12028);
nand U13050 (N_13050,N_12122,N_12187);
or U13051 (N_13051,N_12649,N_12606);
or U13052 (N_13052,N_12733,N_12648);
nand U13053 (N_13053,N_12144,N_12412);
and U13054 (N_13054,N_12319,N_12110);
nand U13055 (N_13055,N_12514,N_12124);
or U13056 (N_13056,N_12008,N_12088);
nand U13057 (N_13057,N_12502,N_12168);
nor U13058 (N_13058,N_12730,N_12743);
or U13059 (N_13059,N_12701,N_12139);
and U13060 (N_13060,N_12525,N_12072);
nand U13061 (N_13061,N_12315,N_12272);
and U13062 (N_13062,N_12670,N_12471);
and U13063 (N_13063,N_12300,N_12202);
and U13064 (N_13064,N_12157,N_12162);
nand U13065 (N_13065,N_12199,N_12584);
or U13066 (N_13066,N_12530,N_12191);
or U13067 (N_13067,N_12667,N_12728);
nor U13068 (N_13068,N_12464,N_12293);
and U13069 (N_13069,N_12449,N_12197);
nor U13070 (N_13070,N_12458,N_12553);
nor U13071 (N_13071,N_12099,N_12151);
nand U13072 (N_13072,N_12326,N_12384);
and U13073 (N_13073,N_12163,N_12273);
and U13074 (N_13074,N_12629,N_12220);
or U13075 (N_13075,N_12524,N_12119);
nand U13076 (N_13076,N_12506,N_12542);
nor U13077 (N_13077,N_12356,N_12511);
or U13078 (N_13078,N_12063,N_12403);
nor U13079 (N_13079,N_12737,N_12433);
xor U13080 (N_13080,N_12231,N_12483);
and U13081 (N_13081,N_12316,N_12310);
and U13082 (N_13082,N_12077,N_12313);
and U13083 (N_13083,N_12594,N_12336);
and U13084 (N_13084,N_12067,N_12159);
or U13085 (N_13085,N_12469,N_12625);
or U13086 (N_13086,N_12411,N_12451);
nand U13087 (N_13087,N_12740,N_12437);
or U13088 (N_13088,N_12254,N_12560);
or U13089 (N_13089,N_12025,N_12023);
and U13090 (N_13090,N_12432,N_12020);
nand U13091 (N_13091,N_12747,N_12556);
and U13092 (N_13092,N_12043,N_12047);
xnor U13093 (N_13093,N_12270,N_12359);
nand U13094 (N_13094,N_12000,N_12180);
or U13095 (N_13095,N_12590,N_12287);
nand U13096 (N_13096,N_12377,N_12650);
and U13097 (N_13097,N_12696,N_12198);
or U13098 (N_13098,N_12501,N_12373);
nor U13099 (N_13099,N_12528,N_12201);
xor U13100 (N_13100,N_12672,N_12104);
nand U13101 (N_13101,N_12423,N_12150);
xnor U13102 (N_13102,N_12076,N_12281);
nand U13103 (N_13103,N_12691,N_12193);
or U13104 (N_13104,N_12042,N_12111);
and U13105 (N_13105,N_12717,N_12375);
or U13106 (N_13106,N_12527,N_12166);
and U13107 (N_13107,N_12094,N_12266);
nor U13108 (N_13108,N_12328,N_12274);
nor U13109 (N_13109,N_12132,N_12317);
and U13110 (N_13110,N_12338,N_12280);
nand U13111 (N_13111,N_12115,N_12547);
nor U13112 (N_13112,N_12618,N_12060);
and U13113 (N_13113,N_12214,N_12114);
nor U13114 (N_13114,N_12337,N_12268);
nor U13115 (N_13115,N_12729,N_12713);
nand U13116 (N_13116,N_12607,N_12417);
nand U13117 (N_13117,N_12108,N_12158);
xor U13118 (N_13118,N_12385,N_12361);
nor U13119 (N_13119,N_12540,N_12082);
nand U13120 (N_13120,N_12030,N_12504);
nand U13121 (N_13121,N_12598,N_12364);
and U13122 (N_13122,N_12388,N_12106);
or U13123 (N_13123,N_12324,N_12561);
or U13124 (N_13124,N_12465,N_12241);
or U13125 (N_13125,N_12336,N_12574);
xor U13126 (N_13126,N_12595,N_12622);
and U13127 (N_13127,N_12236,N_12350);
or U13128 (N_13128,N_12096,N_12410);
or U13129 (N_13129,N_12330,N_12675);
or U13130 (N_13130,N_12514,N_12380);
nand U13131 (N_13131,N_12181,N_12640);
nand U13132 (N_13132,N_12736,N_12127);
and U13133 (N_13133,N_12576,N_12388);
nand U13134 (N_13134,N_12651,N_12396);
and U13135 (N_13135,N_12345,N_12524);
and U13136 (N_13136,N_12207,N_12056);
or U13137 (N_13137,N_12196,N_12685);
nand U13138 (N_13138,N_12623,N_12702);
nor U13139 (N_13139,N_12332,N_12319);
nand U13140 (N_13140,N_12172,N_12590);
or U13141 (N_13141,N_12571,N_12044);
or U13142 (N_13142,N_12315,N_12745);
nor U13143 (N_13143,N_12692,N_12223);
nand U13144 (N_13144,N_12045,N_12158);
and U13145 (N_13145,N_12619,N_12202);
and U13146 (N_13146,N_12012,N_12395);
and U13147 (N_13147,N_12278,N_12234);
nor U13148 (N_13148,N_12127,N_12600);
nor U13149 (N_13149,N_12711,N_12606);
nor U13150 (N_13150,N_12034,N_12217);
nand U13151 (N_13151,N_12008,N_12310);
or U13152 (N_13152,N_12592,N_12703);
xor U13153 (N_13153,N_12404,N_12302);
nor U13154 (N_13154,N_12319,N_12517);
or U13155 (N_13155,N_12648,N_12689);
nor U13156 (N_13156,N_12254,N_12630);
and U13157 (N_13157,N_12396,N_12548);
xnor U13158 (N_13158,N_12087,N_12514);
or U13159 (N_13159,N_12131,N_12626);
or U13160 (N_13160,N_12740,N_12115);
and U13161 (N_13161,N_12355,N_12157);
nand U13162 (N_13162,N_12450,N_12205);
and U13163 (N_13163,N_12063,N_12072);
or U13164 (N_13164,N_12685,N_12410);
nor U13165 (N_13165,N_12391,N_12659);
nand U13166 (N_13166,N_12311,N_12729);
or U13167 (N_13167,N_12347,N_12275);
or U13168 (N_13168,N_12202,N_12555);
nand U13169 (N_13169,N_12253,N_12221);
or U13170 (N_13170,N_12155,N_12393);
xnor U13171 (N_13171,N_12289,N_12406);
nand U13172 (N_13172,N_12010,N_12217);
nand U13173 (N_13173,N_12345,N_12349);
xor U13174 (N_13174,N_12064,N_12706);
nor U13175 (N_13175,N_12085,N_12368);
and U13176 (N_13176,N_12647,N_12386);
or U13177 (N_13177,N_12448,N_12483);
nand U13178 (N_13178,N_12034,N_12397);
xnor U13179 (N_13179,N_12658,N_12097);
and U13180 (N_13180,N_12250,N_12739);
nand U13181 (N_13181,N_12710,N_12486);
xnor U13182 (N_13182,N_12159,N_12174);
nor U13183 (N_13183,N_12702,N_12723);
nand U13184 (N_13184,N_12501,N_12208);
xor U13185 (N_13185,N_12379,N_12339);
and U13186 (N_13186,N_12024,N_12296);
or U13187 (N_13187,N_12238,N_12009);
and U13188 (N_13188,N_12220,N_12699);
nor U13189 (N_13189,N_12364,N_12551);
or U13190 (N_13190,N_12294,N_12050);
or U13191 (N_13191,N_12055,N_12066);
or U13192 (N_13192,N_12694,N_12490);
and U13193 (N_13193,N_12348,N_12660);
and U13194 (N_13194,N_12379,N_12745);
nor U13195 (N_13195,N_12256,N_12341);
xor U13196 (N_13196,N_12347,N_12284);
nor U13197 (N_13197,N_12209,N_12746);
xnor U13198 (N_13198,N_12319,N_12445);
nand U13199 (N_13199,N_12637,N_12096);
and U13200 (N_13200,N_12300,N_12494);
nor U13201 (N_13201,N_12711,N_12331);
or U13202 (N_13202,N_12662,N_12421);
nand U13203 (N_13203,N_12081,N_12517);
nand U13204 (N_13204,N_12161,N_12579);
and U13205 (N_13205,N_12502,N_12547);
and U13206 (N_13206,N_12196,N_12330);
and U13207 (N_13207,N_12629,N_12090);
xor U13208 (N_13208,N_12665,N_12288);
nand U13209 (N_13209,N_12276,N_12091);
nor U13210 (N_13210,N_12201,N_12352);
or U13211 (N_13211,N_12190,N_12666);
nor U13212 (N_13212,N_12652,N_12184);
and U13213 (N_13213,N_12140,N_12280);
and U13214 (N_13214,N_12638,N_12220);
nand U13215 (N_13215,N_12509,N_12676);
nor U13216 (N_13216,N_12181,N_12584);
xor U13217 (N_13217,N_12230,N_12380);
nand U13218 (N_13218,N_12618,N_12276);
or U13219 (N_13219,N_12263,N_12570);
or U13220 (N_13220,N_12153,N_12081);
or U13221 (N_13221,N_12079,N_12684);
nand U13222 (N_13222,N_12418,N_12721);
or U13223 (N_13223,N_12067,N_12086);
nand U13224 (N_13224,N_12439,N_12531);
nor U13225 (N_13225,N_12103,N_12479);
or U13226 (N_13226,N_12381,N_12530);
nand U13227 (N_13227,N_12011,N_12467);
xnor U13228 (N_13228,N_12006,N_12749);
nand U13229 (N_13229,N_12675,N_12404);
nand U13230 (N_13230,N_12502,N_12222);
and U13231 (N_13231,N_12642,N_12187);
and U13232 (N_13232,N_12372,N_12665);
and U13233 (N_13233,N_12124,N_12328);
and U13234 (N_13234,N_12409,N_12691);
or U13235 (N_13235,N_12559,N_12599);
nor U13236 (N_13236,N_12679,N_12521);
nor U13237 (N_13237,N_12528,N_12352);
nand U13238 (N_13238,N_12144,N_12679);
or U13239 (N_13239,N_12589,N_12602);
and U13240 (N_13240,N_12130,N_12576);
nor U13241 (N_13241,N_12666,N_12329);
or U13242 (N_13242,N_12042,N_12035);
nand U13243 (N_13243,N_12351,N_12632);
or U13244 (N_13244,N_12184,N_12206);
or U13245 (N_13245,N_12530,N_12379);
nand U13246 (N_13246,N_12363,N_12264);
and U13247 (N_13247,N_12210,N_12549);
nor U13248 (N_13248,N_12371,N_12461);
nor U13249 (N_13249,N_12098,N_12531);
nor U13250 (N_13250,N_12715,N_12349);
nand U13251 (N_13251,N_12214,N_12217);
and U13252 (N_13252,N_12527,N_12105);
and U13253 (N_13253,N_12428,N_12515);
nand U13254 (N_13254,N_12443,N_12020);
and U13255 (N_13255,N_12734,N_12203);
nand U13256 (N_13256,N_12071,N_12346);
nor U13257 (N_13257,N_12290,N_12610);
and U13258 (N_13258,N_12624,N_12189);
nor U13259 (N_13259,N_12626,N_12650);
nand U13260 (N_13260,N_12139,N_12697);
or U13261 (N_13261,N_12273,N_12324);
nand U13262 (N_13262,N_12204,N_12688);
nand U13263 (N_13263,N_12549,N_12204);
or U13264 (N_13264,N_12066,N_12257);
or U13265 (N_13265,N_12597,N_12313);
nand U13266 (N_13266,N_12519,N_12243);
nand U13267 (N_13267,N_12177,N_12433);
nor U13268 (N_13268,N_12521,N_12208);
xor U13269 (N_13269,N_12356,N_12361);
and U13270 (N_13270,N_12398,N_12313);
nand U13271 (N_13271,N_12097,N_12328);
nor U13272 (N_13272,N_12058,N_12273);
nor U13273 (N_13273,N_12667,N_12445);
nor U13274 (N_13274,N_12318,N_12043);
and U13275 (N_13275,N_12360,N_12400);
or U13276 (N_13276,N_12134,N_12186);
and U13277 (N_13277,N_12079,N_12336);
or U13278 (N_13278,N_12345,N_12738);
or U13279 (N_13279,N_12180,N_12616);
and U13280 (N_13280,N_12625,N_12647);
and U13281 (N_13281,N_12269,N_12614);
nand U13282 (N_13282,N_12684,N_12477);
or U13283 (N_13283,N_12346,N_12341);
nor U13284 (N_13284,N_12454,N_12290);
and U13285 (N_13285,N_12597,N_12582);
and U13286 (N_13286,N_12486,N_12378);
xor U13287 (N_13287,N_12333,N_12403);
nor U13288 (N_13288,N_12154,N_12629);
nand U13289 (N_13289,N_12470,N_12566);
and U13290 (N_13290,N_12241,N_12014);
nor U13291 (N_13291,N_12506,N_12122);
or U13292 (N_13292,N_12278,N_12381);
nor U13293 (N_13293,N_12632,N_12270);
nor U13294 (N_13294,N_12695,N_12047);
nand U13295 (N_13295,N_12379,N_12239);
and U13296 (N_13296,N_12086,N_12644);
nand U13297 (N_13297,N_12384,N_12450);
nand U13298 (N_13298,N_12147,N_12296);
nor U13299 (N_13299,N_12255,N_12188);
nor U13300 (N_13300,N_12662,N_12055);
or U13301 (N_13301,N_12179,N_12455);
or U13302 (N_13302,N_12528,N_12510);
or U13303 (N_13303,N_12138,N_12325);
xnor U13304 (N_13304,N_12108,N_12554);
and U13305 (N_13305,N_12216,N_12196);
or U13306 (N_13306,N_12084,N_12241);
xor U13307 (N_13307,N_12211,N_12424);
nand U13308 (N_13308,N_12100,N_12076);
nand U13309 (N_13309,N_12394,N_12130);
nor U13310 (N_13310,N_12691,N_12449);
nor U13311 (N_13311,N_12221,N_12370);
or U13312 (N_13312,N_12114,N_12082);
or U13313 (N_13313,N_12110,N_12464);
xor U13314 (N_13314,N_12442,N_12049);
and U13315 (N_13315,N_12608,N_12430);
nor U13316 (N_13316,N_12446,N_12666);
nor U13317 (N_13317,N_12198,N_12018);
nor U13318 (N_13318,N_12119,N_12614);
nor U13319 (N_13319,N_12077,N_12641);
or U13320 (N_13320,N_12537,N_12021);
nor U13321 (N_13321,N_12478,N_12245);
nand U13322 (N_13322,N_12429,N_12171);
nor U13323 (N_13323,N_12189,N_12298);
xor U13324 (N_13324,N_12710,N_12618);
and U13325 (N_13325,N_12052,N_12236);
and U13326 (N_13326,N_12447,N_12680);
nand U13327 (N_13327,N_12472,N_12481);
and U13328 (N_13328,N_12642,N_12600);
and U13329 (N_13329,N_12498,N_12311);
and U13330 (N_13330,N_12033,N_12456);
xnor U13331 (N_13331,N_12522,N_12382);
nand U13332 (N_13332,N_12748,N_12516);
nor U13333 (N_13333,N_12584,N_12299);
nor U13334 (N_13334,N_12605,N_12016);
nand U13335 (N_13335,N_12251,N_12258);
nor U13336 (N_13336,N_12515,N_12203);
or U13337 (N_13337,N_12312,N_12346);
and U13338 (N_13338,N_12063,N_12021);
nand U13339 (N_13339,N_12393,N_12580);
or U13340 (N_13340,N_12463,N_12396);
nor U13341 (N_13341,N_12645,N_12285);
and U13342 (N_13342,N_12441,N_12247);
or U13343 (N_13343,N_12520,N_12393);
and U13344 (N_13344,N_12566,N_12747);
and U13345 (N_13345,N_12192,N_12340);
nor U13346 (N_13346,N_12014,N_12094);
nor U13347 (N_13347,N_12093,N_12739);
and U13348 (N_13348,N_12564,N_12005);
and U13349 (N_13349,N_12722,N_12162);
nor U13350 (N_13350,N_12703,N_12269);
nor U13351 (N_13351,N_12142,N_12186);
and U13352 (N_13352,N_12166,N_12062);
nand U13353 (N_13353,N_12204,N_12221);
nand U13354 (N_13354,N_12176,N_12151);
and U13355 (N_13355,N_12482,N_12713);
or U13356 (N_13356,N_12506,N_12462);
nand U13357 (N_13357,N_12478,N_12581);
and U13358 (N_13358,N_12338,N_12079);
and U13359 (N_13359,N_12303,N_12051);
nand U13360 (N_13360,N_12014,N_12654);
nand U13361 (N_13361,N_12596,N_12453);
and U13362 (N_13362,N_12287,N_12274);
and U13363 (N_13363,N_12083,N_12141);
and U13364 (N_13364,N_12721,N_12395);
nor U13365 (N_13365,N_12359,N_12382);
and U13366 (N_13366,N_12689,N_12327);
or U13367 (N_13367,N_12063,N_12035);
and U13368 (N_13368,N_12669,N_12224);
xor U13369 (N_13369,N_12635,N_12202);
nand U13370 (N_13370,N_12259,N_12612);
xor U13371 (N_13371,N_12220,N_12286);
and U13372 (N_13372,N_12588,N_12510);
and U13373 (N_13373,N_12652,N_12064);
and U13374 (N_13374,N_12639,N_12080);
nor U13375 (N_13375,N_12330,N_12579);
and U13376 (N_13376,N_12150,N_12133);
or U13377 (N_13377,N_12748,N_12597);
nor U13378 (N_13378,N_12598,N_12442);
nor U13379 (N_13379,N_12662,N_12634);
nor U13380 (N_13380,N_12624,N_12184);
nand U13381 (N_13381,N_12366,N_12224);
nand U13382 (N_13382,N_12472,N_12213);
xor U13383 (N_13383,N_12638,N_12071);
nor U13384 (N_13384,N_12297,N_12487);
nand U13385 (N_13385,N_12004,N_12697);
nand U13386 (N_13386,N_12456,N_12463);
or U13387 (N_13387,N_12720,N_12562);
and U13388 (N_13388,N_12571,N_12168);
nand U13389 (N_13389,N_12238,N_12588);
nor U13390 (N_13390,N_12648,N_12281);
nand U13391 (N_13391,N_12099,N_12372);
or U13392 (N_13392,N_12611,N_12387);
xor U13393 (N_13393,N_12213,N_12616);
nand U13394 (N_13394,N_12084,N_12419);
and U13395 (N_13395,N_12267,N_12398);
and U13396 (N_13396,N_12456,N_12137);
nand U13397 (N_13397,N_12456,N_12424);
nor U13398 (N_13398,N_12344,N_12571);
or U13399 (N_13399,N_12732,N_12010);
nand U13400 (N_13400,N_12076,N_12503);
or U13401 (N_13401,N_12702,N_12440);
and U13402 (N_13402,N_12261,N_12148);
nor U13403 (N_13403,N_12327,N_12607);
and U13404 (N_13404,N_12022,N_12741);
nor U13405 (N_13405,N_12193,N_12651);
and U13406 (N_13406,N_12491,N_12563);
nand U13407 (N_13407,N_12585,N_12102);
nand U13408 (N_13408,N_12477,N_12722);
nor U13409 (N_13409,N_12442,N_12372);
or U13410 (N_13410,N_12739,N_12698);
or U13411 (N_13411,N_12356,N_12670);
and U13412 (N_13412,N_12310,N_12301);
nor U13413 (N_13413,N_12086,N_12280);
nand U13414 (N_13414,N_12654,N_12425);
or U13415 (N_13415,N_12352,N_12652);
or U13416 (N_13416,N_12041,N_12355);
nor U13417 (N_13417,N_12450,N_12536);
or U13418 (N_13418,N_12513,N_12031);
nand U13419 (N_13419,N_12353,N_12700);
nand U13420 (N_13420,N_12099,N_12736);
nand U13421 (N_13421,N_12014,N_12316);
and U13422 (N_13422,N_12337,N_12219);
nor U13423 (N_13423,N_12308,N_12329);
nand U13424 (N_13424,N_12490,N_12652);
nand U13425 (N_13425,N_12593,N_12011);
nand U13426 (N_13426,N_12035,N_12455);
or U13427 (N_13427,N_12501,N_12500);
nand U13428 (N_13428,N_12316,N_12407);
or U13429 (N_13429,N_12383,N_12433);
nor U13430 (N_13430,N_12093,N_12388);
and U13431 (N_13431,N_12344,N_12055);
and U13432 (N_13432,N_12430,N_12714);
or U13433 (N_13433,N_12625,N_12206);
xor U13434 (N_13434,N_12434,N_12258);
or U13435 (N_13435,N_12744,N_12023);
and U13436 (N_13436,N_12274,N_12651);
and U13437 (N_13437,N_12428,N_12288);
nor U13438 (N_13438,N_12358,N_12406);
or U13439 (N_13439,N_12662,N_12457);
and U13440 (N_13440,N_12719,N_12422);
and U13441 (N_13441,N_12260,N_12215);
and U13442 (N_13442,N_12116,N_12465);
nand U13443 (N_13443,N_12046,N_12265);
xor U13444 (N_13444,N_12145,N_12148);
or U13445 (N_13445,N_12482,N_12636);
and U13446 (N_13446,N_12474,N_12354);
nand U13447 (N_13447,N_12432,N_12328);
nand U13448 (N_13448,N_12139,N_12532);
xnor U13449 (N_13449,N_12136,N_12459);
or U13450 (N_13450,N_12396,N_12334);
nand U13451 (N_13451,N_12094,N_12049);
nor U13452 (N_13452,N_12065,N_12654);
nand U13453 (N_13453,N_12574,N_12666);
and U13454 (N_13454,N_12741,N_12211);
nand U13455 (N_13455,N_12586,N_12279);
and U13456 (N_13456,N_12485,N_12730);
nand U13457 (N_13457,N_12310,N_12637);
xnor U13458 (N_13458,N_12341,N_12312);
nand U13459 (N_13459,N_12310,N_12608);
or U13460 (N_13460,N_12468,N_12545);
or U13461 (N_13461,N_12348,N_12658);
and U13462 (N_13462,N_12514,N_12235);
and U13463 (N_13463,N_12332,N_12146);
nor U13464 (N_13464,N_12427,N_12694);
nor U13465 (N_13465,N_12582,N_12031);
or U13466 (N_13466,N_12065,N_12163);
and U13467 (N_13467,N_12281,N_12530);
and U13468 (N_13468,N_12455,N_12668);
or U13469 (N_13469,N_12523,N_12242);
nor U13470 (N_13470,N_12230,N_12142);
and U13471 (N_13471,N_12244,N_12037);
nand U13472 (N_13472,N_12388,N_12134);
nor U13473 (N_13473,N_12716,N_12645);
and U13474 (N_13474,N_12298,N_12161);
nand U13475 (N_13475,N_12081,N_12210);
nor U13476 (N_13476,N_12088,N_12093);
nor U13477 (N_13477,N_12283,N_12604);
or U13478 (N_13478,N_12415,N_12520);
or U13479 (N_13479,N_12063,N_12553);
or U13480 (N_13480,N_12032,N_12140);
or U13481 (N_13481,N_12708,N_12394);
or U13482 (N_13482,N_12346,N_12579);
nand U13483 (N_13483,N_12389,N_12527);
and U13484 (N_13484,N_12082,N_12453);
xor U13485 (N_13485,N_12075,N_12173);
nand U13486 (N_13486,N_12291,N_12634);
nor U13487 (N_13487,N_12026,N_12146);
and U13488 (N_13488,N_12393,N_12646);
nor U13489 (N_13489,N_12566,N_12224);
and U13490 (N_13490,N_12383,N_12547);
nor U13491 (N_13491,N_12334,N_12126);
nor U13492 (N_13492,N_12213,N_12051);
nand U13493 (N_13493,N_12228,N_12137);
nor U13494 (N_13494,N_12283,N_12719);
nand U13495 (N_13495,N_12699,N_12498);
nor U13496 (N_13496,N_12231,N_12342);
or U13497 (N_13497,N_12383,N_12429);
nand U13498 (N_13498,N_12654,N_12063);
nor U13499 (N_13499,N_12206,N_12311);
or U13500 (N_13500,N_13308,N_13402);
and U13501 (N_13501,N_12829,N_13020);
xor U13502 (N_13502,N_13255,N_13215);
and U13503 (N_13503,N_12982,N_13167);
nor U13504 (N_13504,N_13250,N_13471);
nor U13505 (N_13505,N_13490,N_12959);
nor U13506 (N_13506,N_13370,N_12825);
and U13507 (N_13507,N_13364,N_12776);
or U13508 (N_13508,N_12951,N_13210);
nor U13509 (N_13509,N_13314,N_13484);
nand U13510 (N_13510,N_12901,N_13428);
nand U13511 (N_13511,N_13104,N_13351);
or U13512 (N_13512,N_12865,N_13360);
nor U13513 (N_13513,N_13257,N_12996);
or U13514 (N_13514,N_13294,N_12957);
nand U13515 (N_13515,N_13131,N_13328);
nand U13516 (N_13516,N_12758,N_12930);
nor U13517 (N_13517,N_12977,N_13405);
and U13518 (N_13518,N_13253,N_13404);
and U13519 (N_13519,N_12874,N_13208);
nor U13520 (N_13520,N_13482,N_13305);
nor U13521 (N_13521,N_13320,N_13176);
or U13522 (N_13522,N_13162,N_12782);
or U13523 (N_13523,N_13281,N_13128);
nor U13524 (N_13524,N_13237,N_13437);
and U13525 (N_13525,N_13019,N_13129);
and U13526 (N_13526,N_13075,N_12859);
xor U13527 (N_13527,N_13262,N_13054);
nand U13528 (N_13528,N_12904,N_13443);
and U13529 (N_13529,N_12897,N_12999);
or U13530 (N_13530,N_12946,N_13301);
nor U13531 (N_13531,N_13093,N_12841);
and U13532 (N_13532,N_12845,N_12954);
xor U13533 (N_13533,N_13122,N_13171);
or U13534 (N_13534,N_13359,N_13053);
or U13535 (N_13535,N_12953,N_13102);
nand U13536 (N_13536,N_13483,N_13426);
or U13537 (N_13537,N_13466,N_12933);
nor U13538 (N_13538,N_12932,N_13442);
nor U13539 (N_13539,N_13086,N_13295);
nand U13540 (N_13540,N_13392,N_13383);
or U13541 (N_13541,N_12773,N_13284);
nand U13542 (N_13542,N_13292,N_13347);
nand U13543 (N_13543,N_13217,N_12971);
or U13544 (N_13544,N_13307,N_13407);
nand U13545 (N_13545,N_12763,N_13494);
nor U13546 (N_13546,N_12820,N_13472);
nor U13547 (N_13547,N_12936,N_12772);
and U13548 (N_13548,N_13495,N_13225);
and U13549 (N_13549,N_13356,N_13423);
or U13550 (N_13550,N_12849,N_13000);
xnor U13551 (N_13551,N_13350,N_12784);
nand U13552 (N_13552,N_12764,N_13487);
and U13553 (N_13553,N_13398,N_13087);
nand U13554 (N_13554,N_13427,N_13012);
or U13555 (N_13555,N_13143,N_13375);
xor U13556 (N_13556,N_13189,N_13488);
nor U13557 (N_13557,N_13203,N_12760);
xnor U13558 (N_13558,N_13408,N_13411);
or U13559 (N_13559,N_13455,N_13485);
nand U13560 (N_13560,N_13146,N_13017);
and U13561 (N_13561,N_13151,N_13373);
nor U13562 (N_13562,N_12805,N_13417);
nor U13563 (N_13563,N_13154,N_13254);
nand U13564 (N_13564,N_13174,N_12872);
xnor U13565 (N_13565,N_12927,N_13070);
nor U13566 (N_13566,N_13333,N_13479);
xor U13567 (N_13567,N_12816,N_13361);
or U13568 (N_13568,N_13365,N_12903);
nand U13569 (N_13569,N_13452,N_13195);
or U13570 (N_13570,N_13298,N_13246);
nand U13571 (N_13571,N_13186,N_13352);
nand U13572 (N_13572,N_13394,N_12912);
or U13573 (N_13573,N_12910,N_12774);
and U13574 (N_13574,N_12900,N_13205);
and U13575 (N_13575,N_13409,N_13214);
xor U13576 (N_13576,N_13011,N_12920);
and U13577 (N_13577,N_13429,N_13192);
and U13578 (N_13578,N_12831,N_13156);
nand U13579 (N_13579,N_13457,N_13413);
or U13580 (N_13580,N_13449,N_13163);
nand U13581 (N_13581,N_12828,N_13458);
nand U13582 (N_13582,N_13387,N_13088);
or U13583 (N_13583,N_12935,N_13311);
and U13584 (N_13584,N_13058,N_13029);
nand U13585 (N_13585,N_13296,N_12992);
nand U13586 (N_13586,N_12949,N_13172);
nand U13587 (N_13587,N_12755,N_13376);
nor U13588 (N_13588,N_13273,N_13468);
or U13589 (N_13589,N_13021,N_12907);
nor U13590 (N_13590,N_13047,N_13321);
nand U13591 (N_13591,N_13346,N_13132);
or U13592 (N_13592,N_13285,N_12973);
nor U13593 (N_13593,N_12810,N_13362);
and U13594 (N_13594,N_13059,N_12881);
nand U13595 (N_13595,N_13043,N_13282);
nor U13596 (N_13596,N_12842,N_12843);
nor U13597 (N_13597,N_12906,N_13196);
and U13598 (N_13598,N_12824,N_13152);
and U13599 (N_13599,N_12861,N_12998);
and U13600 (N_13600,N_12750,N_12937);
or U13601 (N_13601,N_13177,N_12846);
xor U13602 (N_13602,N_12968,N_12924);
or U13603 (N_13603,N_12974,N_13006);
nor U13604 (N_13604,N_12873,N_13231);
nor U13605 (N_13605,N_13459,N_12783);
and U13606 (N_13606,N_13139,N_13319);
or U13607 (N_13607,N_12812,N_13261);
nor U13608 (N_13608,N_13233,N_12798);
nor U13609 (N_13609,N_13276,N_13473);
nor U13610 (N_13610,N_13015,N_13467);
and U13611 (N_13611,N_12925,N_13022);
nand U13612 (N_13612,N_13100,N_13330);
nand U13613 (N_13613,N_13068,N_12787);
nand U13614 (N_13614,N_13126,N_12852);
and U13615 (N_13615,N_13289,N_13393);
xor U13616 (N_13616,N_13209,N_12970);
nor U13617 (N_13617,N_13341,N_13031);
xnor U13618 (N_13618,N_12860,N_12980);
nand U13619 (N_13619,N_13050,N_13226);
and U13620 (N_13620,N_13194,N_13439);
or U13621 (N_13621,N_13046,N_13310);
or U13622 (N_13622,N_12839,N_12766);
nor U13623 (N_13623,N_13300,N_13099);
nor U13624 (N_13624,N_13158,N_13110);
xnor U13625 (N_13625,N_12791,N_13096);
or U13626 (N_13626,N_12891,N_13182);
nor U13627 (N_13627,N_13366,N_13159);
nor U13628 (N_13628,N_13180,N_13188);
nand U13629 (N_13629,N_12942,N_13083);
nor U13630 (N_13630,N_13041,N_13441);
nor U13631 (N_13631,N_12851,N_12975);
nand U13632 (N_13632,N_13090,N_12794);
or U13633 (N_13633,N_13169,N_13232);
nor U13634 (N_13634,N_12837,N_12768);
nor U13635 (N_13635,N_13291,N_13322);
nand U13636 (N_13636,N_13092,N_12834);
or U13637 (N_13637,N_12887,N_13389);
nor U13638 (N_13638,N_13496,N_13016);
and U13639 (N_13639,N_13200,N_12853);
nand U13640 (N_13640,N_13134,N_12754);
nor U13641 (N_13641,N_12803,N_13007);
or U13642 (N_13642,N_13034,N_13297);
xnor U13643 (N_13643,N_12960,N_13249);
or U13644 (N_13644,N_12862,N_13438);
and U13645 (N_13645,N_12938,N_13363);
or U13646 (N_13646,N_13002,N_13142);
and U13647 (N_13647,N_13185,N_13386);
or U13648 (N_13648,N_13299,N_13368);
or U13649 (N_13649,N_13127,N_13241);
or U13650 (N_13650,N_13206,N_12940);
nand U13651 (N_13651,N_13238,N_13306);
nand U13652 (N_13652,N_13211,N_13014);
nor U13653 (N_13653,N_12969,N_13179);
nor U13654 (N_13654,N_13181,N_13095);
nand U13655 (N_13655,N_12921,N_12955);
and U13656 (N_13656,N_13332,N_13312);
or U13657 (N_13657,N_12914,N_13039);
nand U13658 (N_13658,N_12775,N_13260);
or U13659 (N_13659,N_13227,N_13009);
or U13660 (N_13660,N_13304,N_13097);
or U13661 (N_13661,N_13435,N_13028);
or U13662 (N_13662,N_13042,N_13130);
or U13663 (N_13663,N_13264,N_13349);
or U13664 (N_13664,N_13178,N_12789);
nor U13665 (N_13665,N_13219,N_13119);
and U13666 (N_13666,N_13372,N_13265);
or U13667 (N_13667,N_13339,N_12950);
nor U13668 (N_13668,N_12945,N_13414);
nor U13669 (N_13669,N_12847,N_13266);
nand U13670 (N_13670,N_13344,N_13433);
nand U13671 (N_13671,N_13116,N_12922);
nand U13672 (N_13672,N_12818,N_13140);
or U13673 (N_13673,N_12870,N_13108);
xor U13674 (N_13674,N_12815,N_13069);
or U13675 (N_13675,N_13161,N_12780);
and U13676 (N_13676,N_13079,N_13412);
nor U13677 (N_13677,N_13474,N_13157);
nor U13678 (N_13678,N_13138,N_12855);
or U13679 (N_13679,N_12896,N_13044);
nor U13680 (N_13680,N_13168,N_13406);
nand U13681 (N_13681,N_13460,N_13248);
xnor U13682 (N_13682,N_13327,N_13036);
and U13683 (N_13683,N_13230,N_12895);
nand U13684 (N_13684,N_13037,N_12918);
nand U13685 (N_13685,N_13074,N_13144);
nand U13686 (N_13686,N_12993,N_13049);
and U13687 (N_13687,N_13018,N_12928);
nand U13688 (N_13688,N_12813,N_12757);
and U13689 (N_13689,N_13170,N_12885);
xor U13690 (N_13690,N_13223,N_12804);
and U13691 (N_13691,N_13493,N_13397);
and U13692 (N_13692,N_13424,N_12826);
nand U13693 (N_13693,N_12868,N_13064);
xor U13694 (N_13694,N_12788,N_13173);
or U13695 (N_13695,N_12759,N_13183);
xnor U13696 (N_13696,N_13288,N_13057);
or U13697 (N_13697,N_13084,N_13160);
or U13698 (N_13698,N_13354,N_13481);
and U13699 (N_13699,N_13107,N_13316);
nor U13700 (N_13700,N_13270,N_12795);
nor U13701 (N_13701,N_13447,N_13245);
nor U13702 (N_13702,N_13274,N_12879);
xor U13703 (N_13703,N_13147,N_13150);
nand U13704 (N_13704,N_13491,N_13032);
nor U13705 (N_13705,N_13343,N_13335);
and U13706 (N_13706,N_13420,N_13089);
nor U13707 (N_13707,N_13071,N_12835);
or U13708 (N_13708,N_12817,N_13111);
nand U13709 (N_13709,N_13415,N_13198);
nand U13710 (N_13710,N_13045,N_13113);
nor U13711 (N_13711,N_13052,N_13303);
nand U13712 (N_13712,N_12800,N_13348);
nor U13713 (N_13713,N_12844,N_12854);
or U13714 (N_13714,N_13085,N_13061);
and U13715 (N_13715,N_13212,N_12871);
and U13716 (N_13716,N_13388,N_13023);
and U13717 (N_13717,N_13258,N_12943);
nor U13718 (N_13718,N_13358,N_12913);
and U13719 (N_13719,N_12858,N_13486);
or U13720 (N_13720,N_13165,N_12893);
nor U13721 (N_13721,N_13451,N_13027);
nor U13722 (N_13722,N_13117,N_13199);
and U13723 (N_13723,N_13272,N_12911);
nor U13724 (N_13724,N_12939,N_13367);
xor U13725 (N_13725,N_13422,N_13076);
nand U13726 (N_13726,N_12988,N_13229);
nor U13727 (N_13727,N_13425,N_12880);
and U13728 (N_13728,N_13381,N_13244);
nand U13729 (N_13729,N_13379,N_13242);
nand U13730 (N_13730,N_13003,N_13155);
and U13731 (N_13731,N_12948,N_13164);
or U13732 (N_13732,N_13463,N_13324);
nand U13733 (N_13733,N_13399,N_13419);
nand U13734 (N_13734,N_13004,N_13030);
nand U13735 (N_13735,N_13240,N_13499);
or U13736 (N_13736,N_13072,N_13228);
and U13737 (N_13737,N_13166,N_12876);
and U13738 (N_13738,N_13317,N_13213);
and U13739 (N_13739,N_13302,N_13187);
nor U13740 (N_13740,N_13446,N_13444);
and U13741 (N_13741,N_13202,N_13063);
and U13742 (N_13742,N_12864,N_13337);
or U13743 (N_13743,N_13403,N_12827);
or U13744 (N_13744,N_12899,N_13410);
nor U13745 (N_13745,N_13338,N_13251);
and U13746 (N_13746,N_13184,N_13325);
and U13747 (N_13747,N_12963,N_13135);
or U13748 (N_13748,N_12956,N_12850);
nor U13749 (N_13749,N_12807,N_13440);
nand U13750 (N_13750,N_13461,N_12799);
and U13751 (N_13751,N_12909,N_13293);
nand U13752 (N_13752,N_12984,N_12833);
nor U13753 (N_13753,N_13033,N_13121);
nor U13754 (N_13754,N_12765,N_13222);
and U13755 (N_13755,N_12994,N_13390);
or U13756 (N_13756,N_13465,N_13277);
and U13757 (N_13757,N_13066,N_13118);
nor U13758 (N_13758,N_13476,N_13077);
nor U13759 (N_13759,N_12915,N_13224);
nor U13760 (N_13760,N_13120,N_13220);
nand U13761 (N_13761,N_13469,N_12785);
nand U13762 (N_13762,N_12867,N_13124);
nor U13763 (N_13763,N_13286,N_12808);
xnor U13764 (N_13764,N_12769,N_13005);
nand U13765 (N_13765,N_13374,N_13221);
and U13766 (N_13766,N_12814,N_13342);
or U13767 (N_13767,N_12964,N_13326);
nor U13768 (N_13768,N_13141,N_13263);
and U13769 (N_13769,N_13355,N_13283);
and U13770 (N_13770,N_13051,N_13391);
nor U13771 (N_13771,N_12989,N_12756);
and U13772 (N_13772,N_13329,N_12877);
xor U13773 (N_13773,N_13204,N_12806);
and U13774 (N_13774,N_12886,N_13137);
nand U13775 (N_13775,N_13048,N_13145);
nor U13776 (N_13776,N_13498,N_13353);
xnor U13777 (N_13777,N_13218,N_13136);
nor U13778 (N_13778,N_13256,N_12952);
or U13779 (N_13779,N_12823,N_13243);
nand U13780 (N_13780,N_13401,N_13497);
or U13781 (N_13781,N_13094,N_13456);
and U13782 (N_13782,N_13269,N_13489);
and U13783 (N_13783,N_13318,N_13025);
or U13784 (N_13784,N_13436,N_12781);
xnor U13785 (N_13785,N_13336,N_13013);
or U13786 (N_13786,N_13331,N_13287);
nor U13787 (N_13787,N_12875,N_13271);
and U13788 (N_13788,N_12836,N_13395);
nor U13789 (N_13789,N_12819,N_13323);
nor U13790 (N_13790,N_12767,N_13421);
nand U13791 (N_13791,N_13026,N_13385);
nor U13792 (N_13792,N_13216,N_13475);
or U13793 (N_13793,N_13035,N_12884);
and U13794 (N_13794,N_13056,N_12838);
nor U13795 (N_13795,N_12917,N_13252);
nand U13796 (N_13796,N_13345,N_12797);
nor U13797 (N_13797,N_13448,N_12902);
and U13798 (N_13798,N_13492,N_12995);
nor U13799 (N_13799,N_12779,N_12986);
nand U13800 (N_13800,N_13236,N_13462);
xor U13801 (N_13801,N_13091,N_13073);
and U13802 (N_13802,N_13081,N_12863);
nand U13803 (N_13803,N_12792,N_12972);
nor U13804 (N_13804,N_12809,N_13377);
and U13805 (N_13805,N_12923,N_13430);
or U13806 (N_13806,N_12856,N_13259);
and U13807 (N_13807,N_12753,N_13434);
and U13808 (N_13808,N_13478,N_12979);
nor U13809 (N_13809,N_13247,N_12944);
nor U13810 (N_13810,N_12941,N_12905);
or U13811 (N_13811,N_13123,N_12889);
or U13812 (N_13812,N_12934,N_12857);
and U13813 (N_13813,N_12976,N_13278);
and U13814 (N_13814,N_13290,N_12991);
or U13815 (N_13815,N_12796,N_12840);
nor U13816 (N_13816,N_13101,N_12966);
and U13817 (N_13817,N_13065,N_13105);
or U13818 (N_13818,N_13432,N_13445);
and U13819 (N_13819,N_13114,N_12892);
nand U13820 (N_13820,N_13280,N_13470);
and U13821 (N_13821,N_13149,N_13010);
nand U13822 (N_13822,N_13418,N_12822);
nand U13823 (N_13823,N_12790,N_13098);
or U13824 (N_13824,N_13477,N_12961);
or U13825 (N_13825,N_12965,N_12882);
and U13826 (N_13826,N_12752,N_13201);
and U13827 (N_13827,N_13024,N_12978);
xor U13828 (N_13828,N_13190,N_13380);
nand U13829 (N_13829,N_13334,N_13384);
and U13830 (N_13830,N_13340,N_12777);
nand U13831 (N_13831,N_13382,N_13400);
or U13832 (N_13832,N_12751,N_12926);
and U13833 (N_13833,N_13431,N_13133);
or U13834 (N_13834,N_13040,N_13067);
or U13835 (N_13835,N_13112,N_13235);
or U13836 (N_13836,N_13109,N_13239);
xor U13837 (N_13837,N_13309,N_13008);
nor U13838 (N_13838,N_12981,N_12821);
nor U13839 (N_13839,N_12987,N_13313);
or U13840 (N_13840,N_12997,N_12786);
and U13841 (N_13841,N_13115,N_12983);
or U13842 (N_13842,N_12811,N_12848);
or U13843 (N_13843,N_12778,N_13315);
nand U13844 (N_13844,N_12947,N_12890);
nor U13845 (N_13845,N_13378,N_12919);
or U13846 (N_13846,N_12883,N_13197);
and U13847 (N_13847,N_13454,N_12898);
nor U13848 (N_13848,N_13191,N_13396);
or U13849 (N_13849,N_13453,N_13038);
nand U13850 (N_13850,N_12916,N_12869);
nand U13851 (N_13851,N_12990,N_13480);
or U13852 (N_13852,N_13080,N_13062);
or U13853 (N_13853,N_13106,N_12832);
or U13854 (N_13854,N_13078,N_13369);
nor U13855 (N_13855,N_12962,N_12908);
nand U13856 (N_13856,N_12967,N_12888);
and U13857 (N_13857,N_12762,N_13207);
xnor U13858 (N_13858,N_13153,N_13234);
nor U13859 (N_13859,N_12929,N_13055);
or U13860 (N_13860,N_12878,N_13450);
xor U13861 (N_13861,N_13193,N_13275);
nor U13862 (N_13862,N_12771,N_13268);
and U13863 (N_13863,N_12985,N_12958);
or U13864 (N_13864,N_13371,N_13103);
and U13865 (N_13865,N_13060,N_12801);
nand U13866 (N_13866,N_13279,N_12866);
and U13867 (N_13867,N_13148,N_12761);
nor U13868 (N_13868,N_13357,N_12770);
nand U13869 (N_13869,N_13175,N_12894);
or U13870 (N_13870,N_13001,N_12830);
and U13871 (N_13871,N_13464,N_12802);
nand U13872 (N_13872,N_13267,N_13082);
nor U13873 (N_13873,N_13125,N_12931);
or U13874 (N_13874,N_12793,N_13416);
nor U13875 (N_13875,N_13223,N_12852);
nor U13876 (N_13876,N_13000,N_13008);
xor U13877 (N_13877,N_12786,N_12976);
or U13878 (N_13878,N_13114,N_12828);
nor U13879 (N_13879,N_12850,N_13045);
and U13880 (N_13880,N_13100,N_12854);
xnor U13881 (N_13881,N_13466,N_13498);
and U13882 (N_13882,N_13092,N_12976);
xnor U13883 (N_13883,N_12761,N_12926);
nor U13884 (N_13884,N_13417,N_12765);
nand U13885 (N_13885,N_12790,N_13211);
nor U13886 (N_13886,N_13272,N_13188);
nand U13887 (N_13887,N_13089,N_13348);
nor U13888 (N_13888,N_12952,N_13264);
nand U13889 (N_13889,N_13154,N_12761);
and U13890 (N_13890,N_13128,N_12840);
nand U13891 (N_13891,N_12908,N_13156);
xor U13892 (N_13892,N_13480,N_12780);
or U13893 (N_13893,N_13273,N_13322);
and U13894 (N_13894,N_13395,N_13115);
and U13895 (N_13895,N_12835,N_12988);
or U13896 (N_13896,N_12753,N_13251);
xnor U13897 (N_13897,N_13150,N_13141);
nor U13898 (N_13898,N_13043,N_13066);
nor U13899 (N_13899,N_13156,N_13056);
nand U13900 (N_13900,N_12985,N_13271);
and U13901 (N_13901,N_13487,N_13389);
nand U13902 (N_13902,N_13371,N_13453);
nor U13903 (N_13903,N_12873,N_12750);
nand U13904 (N_13904,N_13299,N_13270);
or U13905 (N_13905,N_13083,N_12974);
and U13906 (N_13906,N_13476,N_12878);
nor U13907 (N_13907,N_12986,N_12947);
nand U13908 (N_13908,N_13439,N_13352);
nor U13909 (N_13909,N_13092,N_13481);
and U13910 (N_13910,N_13305,N_12817);
and U13911 (N_13911,N_13230,N_13380);
and U13912 (N_13912,N_12893,N_13239);
and U13913 (N_13913,N_12908,N_13387);
nand U13914 (N_13914,N_12783,N_13431);
and U13915 (N_13915,N_13195,N_12814);
nand U13916 (N_13916,N_12899,N_12818);
or U13917 (N_13917,N_13062,N_13078);
nand U13918 (N_13918,N_13376,N_13053);
nand U13919 (N_13919,N_13032,N_13314);
and U13920 (N_13920,N_13170,N_12886);
nor U13921 (N_13921,N_13325,N_12932);
nor U13922 (N_13922,N_12830,N_13425);
nor U13923 (N_13923,N_12759,N_12854);
nor U13924 (N_13924,N_12943,N_13481);
nor U13925 (N_13925,N_13405,N_13480);
or U13926 (N_13926,N_13089,N_13243);
or U13927 (N_13927,N_12777,N_12832);
and U13928 (N_13928,N_13100,N_13267);
or U13929 (N_13929,N_13108,N_12973);
nor U13930 (N_13930,N_13346,N_13265);
nand U13931 (N_13931,N_13337,N_12894);
nand U13932 (N_13932,N_12949,N_13202);
xor U13933 (N_13933,N_12869,N_13366);
and U13934 (N_13934,N_13243,N_13465);
and U13935 (N_13935,N_13450,N_12925);
nor U13936 (N_13936,N_12833,N_13090);
xor U13937 (N_13937,N_13434,N_13309);
xnor U13938 (N_13938,N_13103,N_13262);
nor U13939 (N_13939,N_13308,N_13036);
or U13940 (N_13940,N_12958,N_13138);
nand U13941 (N_13941,N_13473,N_13184);
nand U13942 (N_13942,N_13092,N_13251);
nor U13943 (N_13943,N_13224,N_12972);
xor U13944 (N_13944,N_12867,N_13270);
nor U13945 (N_13945,N_12973,N_12934);
nor U13946 (N_13946,N_13189,N_13380);
nor U13947 (N_13947,N_12878,N_13487);
xor U13948 (N_13948,N_13241,N_12802);
and U13949 (N_13949,N_13242,N_13071);
or U13950 (N_13950,N_13160,N_13048);
or U13951 (N_13951,N_13313,N_13082);
and U13952 (N_13952,N_13314,N_12785);
nand U13953 (N_13953,N_13068,N_12940);
and U13954 (N_13954,N_12787,N_13254);
or U13955 (N_13955,N_12827,N_13246);
nand U13956 (N_13956,N_12755,N_12877);
nand U13957 (N_13957,N_13252,N_13448);
or U13958 (N_13958,N_13054,N_13393);
nand U13959 (N_13959,N_12980,N_12891);
and U13960 (N_13960,N_13083,N_12822);
and U13961 (N_13961,N_13154,N_13427);
or U13962 (N_13962,N_12825,N_13082);
or U13963 (N_13963,N_13121,N_12844);
or U13964 (N_13964,N_13233,N_13061);
xnor U13965 (N_13965,N_12764,N_12875);
or U13966 (N_13966,N_13299,N_13473);
and U13967 (N_13967,N_12793,N_12953);
or U13968 (N_13968,N_12777,N_12892);
nand U13969 (N_13969,N_12882,N_13069);
or U13970 (N_13970,N_12832,N_12884);
nor U13971 (N_13971,N_13099,N_12829);
nand U13972 (N_13972,N_13366,N_13060);
and U13973 (N_13973,N_13460,N_13174);
or U13974 (N_13974,N_13410,N_13437);
or U13975 (N_13975,N_13266,N_13260);
xnor U13976 (N_13976,N_13320,N_13220);
and U13977 (N_13977,N_13435,N_13295);
xor U13978 (N_13978,N_13258,N_12923);
nand U13979 (N_13979,N_12903,N_12761);
or U13980 (N_13980,N_13242,N_13016);
nand U13981 (N_13981,N_13431,N_13394);
nand U13982 (N_13982,N_13409,N_13322);
and U13983 (N_13983,N_12868,N_12942);
nor U13984 (N_13984,N_13367,N_13292);
and U13985 (N_13985,N_12984,N_13373);
or U13986 (N_13986,N_12778,N_12804);
nor U13987 (N_13987,N_12788,N_13074);
nand U13988 (N_13988,N_13274,N_13138);
xor U13989 (N_13989,N_13494,N_13451);
or U13990 (N_13990,N_13212,N_13035);
nand U13991 (N_13991,N_12807,N_12906);
and U13992 (N_13992,N_13220,N_12898);
nand U13993 (N_13993,N_12842,N_13053);
nor U13994 (N_13994,N_12826,N_13390);
and U13995 (N_13995,N_13206,N_13414);
or U13996 (N_13996,N_13463,N_12875);
nor U13997 (N_13997,N_13054,N_13068);
or U13998 (N_13998,N_13468,N_13112);
nor U13999 (N_13999,N_13399,N_13388);
nand U14000 (N_14000,N_12752,N_13023);
and U14001 (N_14001,N_13252,N_13440);
nor U14002 (N_14002,N_12864,N_12970);
xnor U14003 (N_14003,N_13250,N_13375);
and U14004 (N_14004,N_13481,N_13056);
or U14005 (N_14005,N_12757,N_13042);
nor U14006 (N_14006,N_13041,N_12961);
and U14007 (N_14007,N_13226,N_13380);
and U14008 (N_14008,N_13052,N_12809);
nand U14009 (N_14009,N_12810,N_13482);
nand U14010 (N_14010,N_13379,N_12945);
and U14011 (N_14011,N_12879,N_13356);
nor U14012 (N_14012,N_13430,N_13002);
nor U14013 (N_14013,N_13284,N_13121);
xnor U14014 (N_14014,N_12877,N_13176);
nor U14015 (N_14015,N_13205,N_13475);
nand U14016 (N_14016,N_12792,N_12874);
and U14017 (N_14017,N_13270,N_12942);
nand U14018 (N_14018,N_13243,N_13118);
and U14019 (N_14019,N_12877,N_12888);
and U14020 (N_14020,N_13198,N_12953);
and U14021 (N_14021,N_12885,N_13048);
and U14022 (N_14022,N_13071,N_12841);
nand U14023 (N_14023,N_13205,N_13462);
nor U14024 (N_14024,N_12818,N_12822);
or U14025 (N_14025,N_13315,N_12753);
nor U14026 (N_14026,N_12813,N_12851);
xnor U14027 (N_14027,N_13198,N_12764);
and U14028 (N_14028,N_12956,N_12859);
nor U14029 (N_14029,N_12767,N_13238);
or U14030 (N_14030,N_13344,N_13438);
and U14031 (N_14031,N_13055,N_13260);
and U14032 (N_14032,N_13005,N_13106);
nor U14033 (N_14033,N_12980,N_13492);
nor U14034 (N_14034,N_13411,N_13211);
xnor U14035 (N_14035,N_13005,N_12874);
or U14036 (N_14036,N_12753,N_13428);
nor U14037 (N_14037,N_13075,N_13470);
nor U14038 (N_14038,N_13478,N_13443);
nand U14039 (N_14039,N_13026,N_13154);
nor U14040 (N_14040,N_13379,N_12949);
xnor U14041 (N_14041,N_12803,N_13423);
or U14042 (N_14042,N_13293,N_13051);
and U14043 (N_14043,N_12940,N_12796);
or U14044 (N_14044,N_12907,N_13244);
nor U14045 (N_14045,N_13124,N_13339);
or U14046 (N_14046,N_13323,N_12777);
nor U14047 (N_14047,N_13348,N_13168);
or U14048 (N_14048,N_13262,N_13459);
and U14049 (N_14049,N_13190,N_13412);
nand U14050 (N_14050,N_13147,N_12820);
nor U14051 (N_14051,N_13471,N_13251);
nand U14052 (N_14052,N_12875,N_13221);
or U14053 (N_14053,N_13299,N_13411);
or U14054 (N_14054,N_13426,N_12786);
and U14055 (N_14055,N_12960,N_12908);
or U14056 (N_14056,N_13355,N_13258);
or U14057 (N_14057,N_13477,N_12765);
or U14058 (N_14058,N_12753,N_13466);
and U14059 (N_14059,N_13246,N_12870);
or U14060 (N_14060,N_12802,N_13060);
xnor U14061 (N_14061,N_12786,N_13064);
nor U14062 (N_14062,N_12875,N_13111);
or U14063 (N_14063,N_12961,N_12959);
nor U14064 (N_14064,N_12928,N_13459);
nand U14065 (N_14065,N_13240,N_13012);
nand U14066 (N_14066,N_13426,N_13150);
nor U14067 (N_14067,N_12936,N_13165);
xnor U14068 (N_14068,N_13329,N_13362);
or U14069 (N_14069,N_13012,N_13215);
and U14070 (N_14070,N_12855,N_13229);
nand U14071 (N_14071,N_13466,N_13252);
and U14072 (N_14072,N_13364,N_12794);
or U14073 (N_14073,N_12806,N_13068);
or U14074 (N_14074,N_12967,N_12832);
and U14075 (N_14075,N_12750,N_12851);
nand U14076 (N_14076,N_13138,N_13310);
nor U14077 (N_14077,N_12794,N_13188);
xnor U14078 (N_14078,N_13220,N_13110);
or U14079 (N_14079,N_12985,N_13499);
nor U14080 (N_14080,N_13475,N_13496);
and U14081 (N_14081,N_13410,N_12963);
or U14082 (N_14082,N_13292,N_12854);
nand U14083 (N_14083,N_13406,N_13183);
and U14084 (N_14084,N_13110,N_13355);
and U14085 (N_14085,N_13235,N_13123);
nor U14086 (N_14086,N_13270,N_13127);
or U14087 (N_14087,N_12932,N_13223);
nand U14088 (N_14088,N_13048,N_12984);
nand U14089 (N_14089,N_13340,N_13038);
and U14090 (N_14090,N_13055,N_13056);
and U14091 (N_14091,N_13286,N_13239);
or U14092 (N_14092,N_12819,N_13158);
nand U14093 (N_14093,N_13464,N_12848);
and U14094 (N_14094,N_13321,N_13074);
nand U14095 (N_14095,N_13487,N_13064);
xor U14096 (N_14096,N_13312,N_13198);
or U14097 (N_14097,N_12936,N_13229);
nand U14098 (N_14098,N_13400,N_13076);
or U14099 (N_14099,N_13118,N_13115);
nand U14100 (N_14100,N_13213,N_13401);
nor U14101 (N_14101,N_13063,N_13307);
or U14102 (N_14102,N_12833,N_13461);
nor U14103 (N_14103,N_13057,N_12879);
nor U14104 (N_14104,N_13202,N_12845);
nor U14105 (N_14105,N_12767,N_13153);
and U14106 (N_14106,N_12893,N_13064);
nor U14107 (N_14107,N_13281,N_12955);
nor U14108 (N_14108,N_13205,N_12881);
and U14109 (N_14109,N_12772,N_13163);
and U14110 (N_14110,N_13405,N_12852);
and U14111 (N_14111,N_12769,N_12993);
or U14112 (N_14112,N_13119,N_13060);
nor U14113 (N_14113,N_13162,N_13119);
nor U14114 (N_14114,N_13457,N_13017);
and U14115 (N_14115,N_13408,N_13499);
or U14116 (N_14116,N_13253,N_12936);
xor U14117 (N_14117,N_13470,N_12890);
nor U14118 (N_14118,N_13294,N_13206);
nor U14119 (N_14119,N_13037,N_13022);
nor U14120 (N_14120,N_13215,N_12997);
xor U14121 (N_14121,N_13398,N_12797);
nand U14122 (N_14122,N_13314,N_12787);
or U14123 (N_14123,N_13074,N_12783);
or U14124 (N_14124,N_13343,N_13319);
nor U14125 (N_14125,N_13261,N_12892);
nor U14126 (N_14126,N_13214,N_12939);
nor U14127 (N_14127,N_12759,N_13353);
nor U14128 (N_14128,N_13043,N_13341);
nor U14129 (N_14129,N_13319,N_12984);
xnor U14130 (N_14130,N_13077,N_12911);
or U14131 (N_14131,N_12782,N_13098);
or U14132 (N_14132,N_12973,N_13355);
and U14133 (N_14133,N_13315,N_12970);
and U14134 (N_14134,N_13450,N_13262);
nor U14135 (N_14135,N_13176,N_13453);
nor U14136 (N_14136,N_12930,N_13340);
or U14137 (N_14137,N_13315,N_12866);
and U14138 (N_14138,N_12774,N_13246);
and U14139 (N_14139,N_12945,N_13098);
or U14140 (N_14140,N_13383,N_12931);
nand U14141 (N_14141,N_13324,N_12800);
nand U14142 (N_14142,N_13128,N_12991);
and U14143 (N_14143,N_12944,N_13257);
nand U14144 (N_14144,N_13070,N_13185);
xor U14145 (N_14145,N_13147,N_13045);
and U14146 (N_14146,N_12804,N_12918);
or U14147 (N_14147,N_13022,N_12799);
nand U14148 (N_14148,N_12815,N_13021);
or U14149 (N_14149,N_13109,N_13381);
and U14150 (N_14150,N_13195,N_12765);
or U14151 (N_14151,N_13139,N_13165);
nor U14152 (N_14152,N_13070,N_13377);
nor U14153 (N_14153,N_13446,N_12862);
or U14154 (N_14154,N_13276,N_12961);
and U14155 (N_14155,N_13279,N_13091);
nor U14156 (N_14156,N_13215,N_13051);
nor U14157 (N_14157,N_12849,N_13053);
nand U14158 (N_14158,N_13308,N_13386);
nor U14159 (N_14159,N_13301,N_13127);
and U14160 (N_14160,N_13220,N_13200);
or U14161 (N_14161,N_12825,N_13141);
or U14162 (N_14162,N_12839,N_13274);
or U14163 (N_14163,N_13242,N_13496);
or U14164 (N_14164,N_13166,N_12967);
and U14165 (N_14165,N_13162,N_13300);
nor U14166 (N_14166,N_13076,N_13379);
or U14167 (N_14167,N_12984,N_13015);
or U14168 (N_14168,N_12873,N_12811);
and U14169 (N_14169,N_13126,N_13495);
or U14170 (N_14170,N_13475,N_12841);
or U14171 (N_14171,N_12797,N_12919);
or U14172 (N_14172,N_13172,N_13468);
nor U14173 (N_14173,N_13442,N_13257);
or U14174 (N_14174,N_12986,N_12751);
or U14175 (N_14175,N_13312,N_13047);
nor U14176 (N_14176,N_13188,N_12786);
and U14177 (N_14177,N_12955,N_13049);
xor U14178 (N_14178,N_12792,N_13301);
nor U14179 (N_14179,N_13075,N_13303);
nor U14180 (N_14180,N_12849,N_13344);
xor U14181 (N_14181,N_13320,N_13159);
and U14182 (N_14182,N_13174,N_12785);
nor U14183 (N_14183,N_12753,N_13250);
nor U14184 (N_14184,N_13029,N_12762);
or U14185 (N_14185,N_12947,N_12895);
nor U14186 (N_14186,N_12830,N_13329);
nor U14187 (N_14187,N_13025,N_13341);
and U14188 (N_14188,N_13060,N_13436);
nand U14189 (N_14189,N_13375,N_13413);
or U14190 (N_14190,N_12811,N_12874);
or U14191 (N_14191,N_13316,N_13295);
or U14192 (N_14192,N_12981,N_12768);
nand U14193 (N_14193,N_12981,N_12894);
nand U14194 (N_14194,N_13377,N_12781);
or U14195 (N_14195,N_13031,N_12859);
or U14196 (N_14196,N_13299,N_12924);
and U14197 (N_14197,N_13254,N_13260);
and U14198 (N_14198,N_12968,N_13014);
nor U14199 (N_14199,N_12964,N_13208);
or U14200 (N_14200,N_13388,N_12990);
nand U14201 (N_14201,N_13076,N_13185);
and U14202 (N_14202,N_13332,N_13465);
or U14203 (N_14203,N_12865,N_13026);
nor U14204 (N_14204,N_12817,N_13361);
xnor U14205 (N_14205,N_12998,N_13397);
or U14206 (N_14206,N_13252,N_13353);
nor U14207 (N_14207,N_13357,N_12752);
nor U14208 (N_14208,N_13433,N_12968);
nand U14209 (N_14209,N_13007,N_13158);
nor U14210 (N_14210,N_13199,N_13449);
or U14211 (N_14211,N_12936,N_13124);
or U14212 (N_14212,N_13148,N_12867);
xnor U14213 (N_14213,N_12978,N_13131);
or U14214 (N_14214,N_13184,N_13365);
and U14215 (N_14215,N_13385,N_12781);
or U14216 (N_14216,N_12907,N_13197);
nor U14217 (N_14217,N_12879,N_13430);
nor U14218 (N_14218,N_13264,N_13429);
nand U14219 (N_14219,N_13308,N_12767);
nor U14220 (N_14220,N_13169,N_13203);
and U14221 (N_14221,N_13337,N_13333);
and U14222 (N_14222,N_12758,N_13144);
xnor U14223 (N_14223,N_13332,N_13338);
and U14224 (N_14224,N_13112,N_13414);
and U14225 (N_14225,N_12975,N_13115);
nand U14226 (N_14226,N_13157,N_13111);
nor U14227 (N_14227,N_13024,N_13314);
nand U14228 (N_14228,N_12932,N_13143);
and U14229 (N_14229,N_12968,N_13168);
and U14230 (N_14230,N_13104,N_12863);
and U14231 (N_14231,N_13047,N_12891);
or U14232 (N_14232,N_12928,N_13150);
or U14233 (N_14233,N_13391,N_13393);
and U14234 (N_14234,N_13113,N_13310);
nor U14235 (N_14235,N_13387,N_13079);
and U14236 (N_14236,N_13233,N_13238);
nor U14237 (N_14237,N_13044,N_13010);
or U14238 (N_14238,N_13157,N_13278);
nor U14239 (N_14239,N_13050,N_12826);
nand U14240 (N_14240,N_12811,N_13368);
nor U14241 (N_14241,N_13401,N_12817);
nand U14242 (N_14242,N_13479,N_12997);
and U14243 (N_14243,N_13405,N_13100);
nand U14244 (N_14244,N_13470,N_13131);
nand U14245 (N_14245,N_13365,N_13009);
xnor U14246 (N_14246,N_13297,N_12850);
nor U14247 (N_14247,N_12843,N_13238);
or U14248 (N_14248,N_12772,N_13278);
or U14249 (N_14249,N_13441,N_13047);
and U14250 (N_14250,N_14189,N_13529);
nor U14251 (N_14251,N_13848,N_13669);
nand U14252 (N_14252,N_14084,N_14022);
nor U14253 (N_14253,N_13824,N_14014);
and U14254 (N_14254,N_13999,N_13524);
nor U14255 (N_14255,N_13715,N_13511);
and U14256 (N_14256,N_14168,N_13677);
and U14257 (N_14257,N_13589,N_13724);
or U14258 (N_14258,N_13618,N_13569);
nand U14259 (N_14259,N_14034,N_13615);
xor U14260 (N_14260,N_13915,N_13776);
or U14261 (N_14261,N_13813,N_13705);
nor U14262 (N_14262,N_13782,N_13796);
nor U14263 (N_14263,N_13559,N_13988);
nand U14264 (N_14264,N_14248,N_13532);
xor U14265 (N_14265,N_14123,N_14030);
nor U14266 (N_14266,N_14057,N_13706);
xor U14267 (N_14267,N_14135,N_14134);
and U14268 (N_14268,N_14213,N_13568);
nand U14269 (N_14269,N_14040,N_13594);
and U14270 (N_14270,N_13979,N_13579);
and U14271 (N_14271,N_14182,N_13621);
or U14272 (N_14272,N_13780,N_13993);
or U14273 (N_14273,N_14092,N_14199);
and U14274 (N_14274,N_13968,N_14105);
nand U14275 (N_14275,N_13881,N_13897);
and U14276 (N_14276,N_13907,N_14138);
nor U14277 (N_14277,N_13743,N_13974);
and U14278 (N_14278,N_13631,N_14107);
and U14279 (N_14279,N_14028,N_13673);
or U14280 (N_14280,N_13707,N_14001);
or U14281 (N_14281,N_13711,N_13967);
nor U14282 (N_14282,N_14020,N_13903);
nor U14283 (N_14283,N_13650,N_13938);
or U14284 (N_14284,N_13850,N_14125);
or U14285 (N_14285,N_13630,N_14231);
nor U14286 (N_14286,N_13871,N_13522);
nor U14287 (N_14287,N_13771,N_13633);
and U14288 (N_14288,N_13998,N_13525);
nor U14289 (N_14289,N_14216,N_14017);
and U14290 (N_14290,N_14065,N_14212);
or U14291 (N_14291,N_13550,N_13504);
nand U14292 (N_14292,N_13545,N_13858);
xor U14293 (N_14293,N_13681,N_13508);
nand U14294 (N_14294,N_14095,N_13582);
or U14295 (N_14295,N_14140,N_13767);
nand U14296 (N_14296,N_13657,N_13847);
nor U14297 (N_14297,N_13624,N_13756);
or U14298 (N_14298,N_14176,N_13639);
nor U14299 (N_14299,N_14245,N_14188);
or U14300 (N_14300,N_13626,N_13870);
nand U14301 (N_14301,N_13797,N_13562);
nand U14302 (N_14302,N_14163,N_13928);
and U14303 (N_14303,N_14037,N_13539);
or U14304 (N_14304,N_13766,N_13893);
nor U14305 (N_14305,N_13917,N_13619);
and U14306 (N_14306,N_14166,N_13695);
nor U14307 (N_14307,N_13795,N_13890);
nor U14308 (N_14308,N_13640,N_14081);
or U14309 (N_14309,N_13959,N_14136);
xor U14310 (N_14310,N_14099,N_14012);
or U14311 (N_14311,N_13859,N_13831);
nand U14312 (N_14312,N_14227,N_13609);
nand U14313 (N_14313,N_13679,N_13612);
and U14314 (N_14314,N_13670,N_14104);
and U14315 (N_14315,N_13973,N_13722);
nand U14316 (N_14316,N_13977,N_14002);
nor U14317 (N_14317,N_13586,N_13906);
nor U14318 (N_14318,N_14165,N_13622);
and U14319 (N_14319,N_13882,N_13838);
nor U14320 (N_14320,N_14101,N_14203);
nand U14321 (N_14321,N_14169,N_13734);
nand U14322 (N_14322,N_14214,N_14187);
xnor U14323 (N_14323,N_13865,N_14208);
nor U14324 (N_14324,N_14246,N_14023);
nor U14325 (N_14325,N_14016,N_13638);
xnor U14326 (N_14326,N_13606,N_13512);
nor U14327 (N_14327,N_13720,N_14031);
and U14328 (N_14328,N_13943,N_13623);
or U14329 (N_14329,N_13814,N_14019);
and U14330 (N_14330,N_13526,N_13717);
or U14331 (N_14331,N_14149,N_13970);
or U14332 (N_14332,N_13656,N_13768);
nor U14333 (N_14333,N_13965,N_13904);
or U14334 (N_14334,N_14050,N_13598);
nand U14335 (N_14335,N_13761,N_13517);
or U14336 (N_14336,N_13674,N_14229);
or U14337 (N_14337,N_13936,N_14180);
nand U14338 (N_14338,N_13520,N_13625);
and U14339 (N_14339,N_13689,N_14052);
nor U14340 (N_14340,N_14064,N_14085);
xnor U14341 (N_14341,N_14077,N_14209);
and U14342 (N_14342,N_13763,N_14228);
nand U14343 (N_14343,N_13949,N_13688);
or U14344 (N_14344,N_13690,N_13827);
or U14345 (N_14345,N_13610,N_13672);
or U14346 (N_14346,N_13651,N_13918);
or U14347 (N_14347,N_13649,N_14011);
nor U14348 (N_14348,N_13701,N_14058);
or U14349 (N_14349,N_13889,N_13564);
and U14350 (N_14350,N_13509,N_13742);
nor U14351 (N_14351,N_13770,N_14167);
nor U14352 (N_14352,N_13913,N_14106);
or U14353 (N_14353,N_14056,N_14151);
nor U14354 (N_14354,N_13960,N_14021);
nand U14355 (N_14355,N_13927,N_13527);
or U14356 (N_14356,N_13851,N_14003);
or U14357 (N_14357,N_14100,N_14075);
or U14358 (N_14358,N_13931,N_13984);
nand U14359 (N_14359,N_14154,N_13678);
nor U14360 (N_14360,N_13544,N_14000);
nand U14361 (N_14361,N_13832,N_13935);
nand U14362 (N_14362,N_13671,N_13788);
nor U14363 (N_14363,N_13641,N_13985);
nand U14364 (N_14364,N_13945,N_13876);
nand U14365 (N_14365,N_13798,N_13593);
nor U14366 (N_14366,N_13694,N_13596);
and U14367 (N_14367,N_13933,N_14211);
or U14368 (N_14368,N_13801,N_13737);
nand U14369 (N_14369,N_13953,N_13987);
nor U14370 (N_14370,N_13940,N_14029);
nand U14371 (N_14371,N_14087,N_13833);
or U14372 (N_14372,N_14156,N_13994);
or U14373 (N_14373,N_14171,N_14150);
nand U14374 (N_14374,N_13786,N_14072);
and U14375 (N_14375,N_14082,N_13822);
nor U14376 (N_14376,N_13930,N_13874);
and U14377 (N_14377,N_13732,N_13958);
or U14378 (N_14378,N_13744,N_13546);
or U14379 (N_14379,N_13675,N_14242);
nand U14380 (N_14380,N_13686,N_13789);
or U14381 (N_14381,N_13759,N_14131);
nor U14382 (N_14382,N_14184,N_14226);
nor U14383 (N_14383,N_13603,N_13941);
nor U14384 (N_14384,N_13912,N_13629);
nor U14385 (N_14385,N_13805,N_14179);
nand U14386 (N_14386,N_13607,N_13978);
nor U14387 (N_14387,N_14009,N_13836);
and U14388 (N_14388,N_13964,N_14066);
and U14389 (N_14389,N_14088,N_14132);
and U14390 (N_14390,N_13852,N_13567);
and U14391 (N_14391,N_14083,N_13839);
and U14392 (N_14392,N_14111,N_13667);
nand U14393 (N_14393,N_14054,N_13557);
xor U14394 (N_14394,N_14233,N_13575);
or U14395 (N_14395,N_14006,N_13572);
xnor U14396 (N_14396,N_13856,N_13862);
nor U14397 (N_14397,N_13902,N_13723);
nor U14398 (N_14398,N_13661,N_13793);
or U14399 (N_14399,N_13600,N_13540);
nand U14400 (N_14400,N_14224,N_13773);
nand U14401 (N_14401,N_13548,N_13692);
nand U14402 (N_14402,N_14121,N_14210);
or U14403 (N_14403,N_13595,N_13729);
or U14404 (N_14404,N_14235,N_13659);
xor U14405 (N_14405,N_14005,N_13652);
or U14406 (N_14406,N_13986,N_13749);
nor U14407 (N_14407,N_13887,N_13829);
xor U14408 (N_14408,N_13861,N_14115);
and U14409 (N_14409,N_13516,N_13841);
nand U14410 (N_14410,N_13542,N_13844);
nand U14411 (N_14411,N_13704,N_14007);
nor U14412 (N_14412,N_13635,N_13911);
and U14413 (N_14413,N_14128,N_13591);
nand U14414 (N_14414,N_13541,N_13860);
or U14415 (N_14415,N_13510,N_13716);
or U14416 (N_14416,N_13885,N_14061);
or U14417 (N_14417,N_14080,N_14147);
xor U14418 (N_14418,N_13736,N_13983);
xor U14419 (N_14419,N_13642,N_14143);
and U14420 (N_14420,N_14234,N_14076);
or U14421 (N_14421,N_14157,N_13685);
xnor U14422 (N_14422,N_13730,N_13519);
or U14423 (N_14423,N_13721,N_13563);
and U14424 (N_14424,N_13819,N_13817);
or U14425 (N_14425,N_13785,N_13555);
or U14426 (N_14426,N_13739,N_14183);
nor U14427 (N_14427,N_13894,N_13561);
or U14428 (N_14428,N_13895,N_13997);
nand U14429 (N_14429,N_14198,N_13901);
nor U14430 (N_14430,N_13571,N_13605);
and U14431 (N_14431,N_13834,N_14027);
and U14432 (N_14432,N_13845,N_14159);
nor U14433 (N_14433,N_13864,N_14238);
or U14434 (N_14434,N_13758,N_13614);
nor U14435 (N_14435,N_13896,N_13696);
nor U14436 (N_14436,N_13608,N_13923);
nor U14437 (N_14437,N_13627,N_13857);
and U14438 (N_14438,N_13764,N_14139);
nor U14439 (N_14439,N_13731,N_13753);
nor U14440 (N_14440,N_14215,N_13637);
nand U14441 (N_14441,N_13728,N_13570);
nand U14442 (N_14442,N_13636,N_14113);
nand U14443 (N_14443,N_13663,N_13698);
or U14444 (N_14444,N_13939,N_14118);
nor U14445 (N_14445,N_14218,N_13826);
xnor U14446 (N_14446,N_13925,N_13735);
nor U14447 (N_14447,N_13837,N_13573);
and U14448 (N_14448,N_14059,N_14127);
or U14449 (N_14449,N_14243,N_13556);
nand U14450 (N_14450,N_14200,N_13765);
or U14451 (N_14451,N_14133,N_14232);
xor U14452 (N_14452,N_14053,N_14186);
nor U14453 (N_14453,N_13937,N_13791);
or U14454 (N_14454,N_13799,N_13809);
nor U14455 (N_14455,N_14222,N_13942);
and U14456 (N_14456,N_13719,N_13760);
nor U14457 (N_14457,N_14196,N_13956);
nor U14458 (N_14458,N_13872,N_13910);
or U14459 (N_14459,N_13762,N_13566);
or U14460 (N_14460,N_14114,N_14221);
nor U14461 (N_14461,N_14249,N_13613);
nand U14462 (N_14462,N_14201,N_13971);
or U14463 (N_14463,N_14060,N_13835);
nand U14464 (N_14464,N_13533,N_13883);
nand U14465 (N_14465,N_13617,N_13703);
nor U14466 (N_14466,N_13855,N_14062);
xnor U14467 (N_14467,N_13687,N_13750);
and U14468 (N_14468,N_14145,N_13995);
xnor U14469 (N_14469,N_13957,N_14108);
and U14470 (N_14470,N_13553,N_13807);
and U14471 (N_14471,N_13843,N_13769);
or U14472 (N_14472,N_13554,N_13628);
and U14473 (N_14473,N_13891,N_13697);
nand U14474 (N_14474,N_14074,N_13513);
and U14475 (N_14475,N_13547,N_14070);
xnor U14476 (N_14476,N_13585,N_13952);
nor U14477 (N_14477,N_14142,N_13515);
and U14478 (N_14478,N_13800,N_13849);
and U14479 (N_14479,N_13867,N_13774);
and U14480 (N_14480,N_13576,N_13950);
nand U14481 (N_14481,N_13592,N_14191);
and U14482 (N_14482,N_13726,N_13501);
nor U14483 (N_14483,N_13514,N_13989);
or U14484 (N_14484,N_13620,N_13955);
and U14485 (N_14485,N_13751,N_13682);
nor U14486 (N_14486,N_13846,N_14045);
nand U14487 (N_14487,N_14116,N_13934);
nor U14488 (N_14488,N_13951,N_13745);
or U14489 (N_14489,N_14130,N_14090);
or U14490 (N_14490,N_14086,N_14117);
nand U14491 (N_14491,N_13748,N_13602);
nand U14492 (N_14492,N_13693,N_13565);
xnor U14493 (N_14493,N_14144,N_13787);
nor U14494 (N_14494,N_13772,N_13803);
xnor U14495 (N_14495,N_13944,N_13683);
nand U14496 (N_14496,N_13991,N_13919);
or U14497 (N_14497,N_14096,N_13990);
nand U14498 (N_14498,N_14041,N_13712);
and U14499 (N_14499,N_14068,N_13583);
xnor U14500 (N_14500,N_13752,N_13665);
nand U14501 (N_14501,N_13812,N_14119);
or U14502 (N_14502,N_13543,N_13574);
and U14503 (N_14503,N_13815,N_13905);
or U14504 (N_14504,N_13821,N_14036);
and U14505 (N_14505,N_13794,N_13924);
nand U14506 (N_14506,N_14071,N_13727);
nand U14507 (N_14507,N_14110,N_14120);
nand U14508 (N_14508,N_13975,N_13863);
and U14509 (N_14509,N_13899,N_13962);
or U14510 (N_14510,N_13804,N_13502);
xor U14511 (N_14511,N_13653,N_14236);
or U14512 (N_14512,N_13580,N_14069);
and U14513 (N_14513,N_14089,N_13680);
nand U14514 (N_14514,N_13708,N_14044);
and U14515 (N_14515,N_13714,N_14164);
or U14516 (N_14516,N_13811,N_14109);
or U14517 (N_14517,N_14170,N_14073);
or U14518 (N_14518,N_14042,N_13668);
nor U14519 (N_14519,N_13777,N_13892);
xor U14520 (N_14520,N_13741,N_13664);
or U14521 (N_14521,N_14103,N_14004);
and U14522 (N_14522,N_13818,N_13718);
nand U14523 (N_14523,N_13992,N_14207);
and U14524 (N_14524,N_13597,N_13733);
nand U14525 (N_14525,N_13710,N_14102);
nor U14526 (N_14526,N_14097,N_13880);
nor U14527 (N_14527,N_14174,N_14008);
nor U14528 (N_14528,N_13725,N_14204);
nor U14529 (N_14529,N_13521,N_13775);
nor U14530 (N_14530,N_13662,N_14172);
and U14531 (N_14531,N_13535,N_13888);
or U14532 (N_14532,N_13587,N_14032);
nor U14533 (N_14533,N_14197,N_13868);
nand U14534 (N_14534,N_14223,N_13947);
and U14535 (N_14535,N_14033,N_13781);
nand U14536 (N_14536,N_14155,N_14146);
nor U14537 (N_14537,N_13816,N_13961);
nor U14538 (N_14538,N_14112,N_13792);
nor U14539 (N_14539,N_14239,N_13740);
nor U14540 (N_14540,N_14173,N_13560);
nand U14541 (N_14541,N_14202,N_14177);
and U14542 (N_14542,N_13702,N_13932);
and U14543 (N_14543,N_14047,N_14094);
nor U14544 (N_14544,N_13972,N_13981);
or U14545 (N_14545,N_14241,N_14230);
or U14546 (N_14546,N_13842,N_13666);
nor U14547 (N_14547,N_14079,N_13898);
nand U14548 (N_14548,N_13581,N_14193);
nor U14549 (N_14549,N_14039,N_14217);
or U14550 (N_14550,N_13783,N_14126);
nor U14551 (N_14551,N_13660,N_13537);
nand U14552 (N_14552,N_14158,N_13963);
nand U14553 (N_14553,N_14122,N_14205);
nand U14554 (N_14554,N_14192,N_13503);
xnor U14555 (N_14555,N_13996,N_13507);
and U14556 (N_14556,N_13590,N_13634);
or U14557 (N_14557,N_13908,N_13806);
or U14558 (N_14558,N_14148,N_14048);
and U14559 (N_14559,N_14046,N_14067);
nor U14560 (N_14560,N_14162,N_13921);
and U14561 (N_14561,N_13577,N_14181);
nor U14562 (N_14562,N_13578,N_13909);
or U14563 (N_14563,N_13518,N_14078);
nor U14564 (N_14564,N_14018,N_13601);
nor U14565 (N_14565,N_13875,N_14237);
nand U14566 (N_14566,N_14244,N_14190);
and U14567 (N_14567,N_14063,N_13810);
xor U14568 (N_14568,N_13691,N_13922);
or U14569 (N_14569,N_14038,N_13500);
nand U14570 (N_14570,N_14093,N_13920);
xnor U14571 (N_14571,N_14043,N_14195);
nand U14572 (N_14572,N_14049,N_14013);
and U14573 (N_14573,N_13825,N_13709);
or U14574 (N_14574,N_13877,N_13643);
or U14575 (N_14575,N_14025,N_13530);
or U14576 (N_14576,N_13878,N_13754);
nor U14577 (N_14577,N_13755,N_14153);
nor U14578 (N_14578,N_13523,N_13549);
nand U14579 (N_14579,N_14024,N_13886);
xor U14580 (N_14580,N_13757,N_13611);
xor U14581 (N_14581,N_13853,N_14247);
and U14582 (N_14582,N_13528,N_14137);
nand U14583 (N_14583,N_13969,N_13599);
or U14584 (N_14584,N_13632,N_13820);
and U14585 (N_14585,N_13790,N_13648);
nand U14586 (N_14586,N_13976,N_13802);
and U14587 (N_14587,N_13713,N_13746);
or U14588 (N_14588,N_13840,N_14010);
or U14589 (N_14589,N_14160,N_14185);
and U14590 (N_14590,N_14152,N_13866);
nand U14591 (N_14591,N_13531,N_13929);
and U14592 (N_14592,N_14026,N_13616);
nor U14593 (N_14593,N_13946,N_14141);
nor U14594 (N_14594,N_13884,N_14240);
nand U14595 (N_14595,N_13699,N_13954);
xor U14596 (N_14596,N_13552,N_14098);
and U14597 (N_14597,N_14220,N_13700);
nand U14598 (N_14598,N_13646,N_13966);
and U14599 (N_14599,N_13823,N_13879);
nand U14600 (N_14600,N_14055,N_13980);
and U14601 (N_14601,N_13505,N_13684);
nand U14602 (N_14602,N_14161,N_14124);
and U14603 (N_14603,N_13645,N_13779);
nand U14604 (N_14604,N_13854,N_13982);
nor U14605 (N_14605,N_14015,N_13551);
and U14606 (N_14606,N_13914,N_14178);
nand U14607 (N_14607,N_13584,N_14219);
and U14608 (N_14608,N_14129,N_14206);
and U14609 (N_14609,N_14091,N_13869);
nor U14610 (N_14610,N_13604,N_13558);
and U14611 (N_14611,N_13784,N_13948);
nand U14612 (N_14612,N_14035,N_13873);
and U14613 (N_14613,N_13654,N_13828);
nor U14614 (N_14614,N_13644,N_14225);
nor U14615 (N_14615,N_13538,N_13808);
or U14616 (N_14616,N_13536,N_13738);
nor U14617 (N_14617,N_13647,N_13676);
nor U14618 (N_14618,N_13534,N_13588);
and U14619 (N_14619,N_13830,N_13916);
and U14620 (N_14620,N_13900,N_14194);
or U14621 (N_14621,N_13926,N_13778);
and U14622 (N_14622,N_14051,N_13658);
and U14623 (N_14623,N_13747,N_14175);
and U14624 (N_14624,N_13655,N_13506);
nor U14625 (N_14625,N_14208,N_13814);
or U14626 (N_14626,N_13728,N_14134);
nand U14627 (N_14627,N_13673,N_13808);
nor U14628 (N_14628,N_14095,N_13659);
and U14629 (N_14629,N_13751,N_13506);
or U14630 (N_14630,N_13934,N_14086);
nor U14631 (N_14631,N_14242,N_14147);
and U14632 (N_14632,N_14019,N_14098);
xnor U14633 (N_14633,N_13510,N_13999);
nand U14634 (N_14634,N_13677,N_13799);
nand U14635 (N_14635,N_13916,N_13977);
or U14636 (N_14636,N_14165,N_13555);
or U14637 (N_14637,N_14024,N_13640);
and U14638 (N_14638,N_13615,N_14058);
nand U14639 (N_14639,N_14047,N_14089);
and U14640 (N_14640,N_13959,N_14111);
or U14641 (N_14641,N_14094,N_14088);
and U14642 (N_14642,N_13982,N_13521);
and U14643 (N_14643,N_13924,N_13915);
and U14644 (N_14644,N_14183,N_13611);
xor U14645 (N_14645,N_14056,N_14068);
and U14646 (N_14646,N_14009,N_13701);
and U14647 (N_14647,N_14130,N_13721);
xor U14648 (N_14648,N_13660,N_13671);
nor U14649 (N_14649,N_13681,N_13808);
or U14650 (N_14650,N_14019,N_14023);
nor U14651 (N_14651,N_13753,N_13709);
and U14652 (N_14652,N_14199,N_13820);
and U14653 (N_14653,N_14157,N_14079);
nor U14654 (N_14654,N_13586,N_14236);
nand U14655 (N_14655,N_13602,N_14090);
nor U14656 (N_14656,N_13677,N_13998);
and U14657 (N_14657,N_14174,N_13521);
nand U14658 (N_14658,N_13860,N_13730);
and U14659 (N_14659,N_13538,N_13876);
and U14660 (N_14660,N_13795,N_13998);
nor U14661 (N_14661,N_13555,N_14031);
nor U14662 (N_14662,N_14073,N_13796);
nand U14663 (N_14663,N_13592,N_14195);
and U14664 (N_14664,N_13977,N_13784);
nand U14665 (N_14665,N_13752,N_13554);
and U14666 (N_14666,N_14215,N_14244);
xor U14667 (N_14667,N_13961,N_14101);
and U14668 (N_14668,N_14248,N_14210);
or U14669 (N_14669,N_13832,N_14246);
nor U14670 (N_14670,N_14067,N_13735);
and U14671 (N_14671,N_14149,N_13871);
nor U14672 (N_14672,N_13684,N_13525);
nand U14673 (N_14673,N_13504,N_13831);
nand U14674 (N_14674,N_14179,N_14190);
nor U14675 (N_14675,N_13952,N_14063);
and U14676 (N_14676,N_13918,N_13921);
nor U14677 (N_14677,N_13812,N_13579);
nand U14678 (N_14678,N_14037,N_14154);
nand U14679 (N_14679,N_13911,N_13982);
xnor U14680 (N_14680,N_13652,N_13539);
nor U14681 (N_14681,N_14002,N_13937);
nand U14682 (N_14682,N_13530,N_13904);
or U14683 (N_14683,N_14106,N_13960);
nor U14684 (N_14684,N_13764,N_14223);
nand U14685 (N_14685,N_13810,N_14138);
nor U14686 (N_14686,N_13646,N_13755);
or U14687 (N_14687,N_13948,N_13563);
nor U14688 (N_14688,N_13517,N_13845);
xnor U14689 (N_14689,N_14074,N_13615);
xnor U14690 (N_14690,N_14121,N_14224);
or U14691 (N_14691,N_13570,N_14121);
and U14692 (N_14692,N_13699,N_13521);
or U14693 (N_14693,N_13580,N_14012);
or U14694 (N_14694,N_13707,N_14022);
and U14695 (N_14695,N_13714,N_13875);
or U14696 (N_14696,N_13582,N_14139);
and U14697 (N_14697,N_13915,N_13760);
nand U14698 (N_14698,N_13729,N_14124);
nand U14699 (N_14699,N_13789,N_13951);
nor U14700 (N_14700,N_13867,N_14152);
nor U14701 (N_14701,N_13957,N_13996);
or U14702 (N_14702,N_14243,N_13824);
nand U14703 (N_14703,N_14088,N_14195);
or U14704 (N_14704,N_13831,N_13759);
or U14705 (N_14705,N_13553,N_13702);
or U14706 (N_14706,N_13772,N_13688);
and U14707 (N_14707,N_14119,N_13680);
nor U14708 (N_14708,N_13852,N_13775);
or U14709 (N_14709,N_13780,N_13976);
nand U14710 (N_14710,N_13768,N_13930);
nor U14711 (N_14711,N_13518,N_14032);
nor U14712 (N_14712,N_13765,N_14246);
and U14713 (N_14713,N_13900,N_13691);
nand U14714 (N_14714,N_14025,N_13510);
nand U14715 (N_14715,N_14218,N_14151);
and U14716 (N_14716,N_13514,N_14225);
or U14717 (N_14717,N_13574,N_13784);
and U14718 (N_14718,N_13619,N_13527);
nor U14719 (N_14719,N_13690,N_13997);
nor U14720 (N_14720,N_14179,N_13883);
nor U14721 (N_14721,N_13511,N_14066);
nor U14722 (N_14722,N_13661,N_14009);
nand U14723 (N_14723,N_13688,N_13719);
nand U14724 (N_14724,N_13965,N_13609);
and U14725 (N_14725,N_13970,N_13591);
and U14726 (N_14726,N_13546,N_14207);
or U14727 (N_14727,N_13849,N_14197);
nand U14728 (N_14728,N_14106,N_13720);
and U14729 (N_14729,N_14197,N_13502);
and U14730 (N_14730,N_14159,N_13524);
and U14731 (N_14731,N_13587,N_14231);
and U14732 (N_14732,N_14121,N_13732);
and U14733 (N_14733,N_13727,N_14157);
nand U14734 (N_14734,N_13743,N_13754);
nor U14735 (N_14735,N_13905,N_13819);
and U14736 (N_14736,N_13509,N_13854);
nor U14737 (N_14737,N_14212,N_14042);
nor U14738 (N_14738,N_13676,N_14026);
xnor U14739 (N_14739,N_13558,N_13960);
nor U14740 (N_14740,N_13878,N_13987);
or U14741 (N_14741,N_13820,N_14138);
and U14742 (N_14742,N_13546,N_14056);
nand U14743 (N_14743,N_14129,N_14233);
and U14744 (N_14744,N_14099,N_13576);
and U14745 (N_14745,N_14247,N_14014);
xor U14746 (N_14746,N_14108,N_13710);
xor U14747 (N_14747,N_14200,N_14131);
and U14748 (N_14748,N_13928,N_13815);
and U14749 (N_14749,N_14120,N_13530);
or U14750 (N_14750,N_13831,N_14196);
or U14751 (N_14751,N_13845,N_13740);
or U14752 (N_14752,N_13596,N_14074);
nor U14753 (N_14753,N_14178,N_13785);
or U14754 (N_14754,N_14054,N_14061);
nor U14755 (N_14755,N_13975,N_13970);
and U14756 (N_14756,N_14042,N_13753);
nand U14757 (N_14757,N_13828,N_13582);
xor U14758 (N_14758,N_14026,N_13937);
nand U14759 (N_14759,N_14140,N_13659);
or U14760 (N_14760,N_13609,N_14105);
nand U14761 (N_14761,N_13958,N_13810);
and U14762 (N_14762,N_14244,N_13834);
and U14763 (N_14763,N_13736,N_13797);
xor U14764 (N_14764,N_14204,N_13508);
and U14765 (N_14765,N_13820,N_13526);
nor U14766 (N_14766,N_13531,N_13935);
nor U14767 (N_14767,N_14052,N_13973);
and U14768 (N_14768,N_14055,N_14056);
nor U14769 (N_14769,N_13718,N_13927);
nand U14770 (N_14770,N_14010,N_13508);
and U14771 (N_14771,N_13637,N_14010);
nor U14772 (N_14772,N_13697,N_14054);
nor U14773 (N_14773,N_14133,N_13738);
nor U14774 (N_14774,N_13962,N_13741);
and U14775 (N_14775,N_13868,N_13875);
nand U14776 (N_14776,N_14209,N_13802);
or U14777 (N_14777,N_14084,N_14236);
or U14778 (N_14778,N_13521,N_14123);
nor U14779 (N_14779,N_13733,N_14125);
nor U14780 (N_14780,N_14212,N_13878);
nor U14781 (N_14781,N_14018,N_14134);
or U14782 (N_14782,N_14057,N_13933);
or U14783 (N_14783,N_13600,N_14102);
nand U14784 (N_14784,N_13910,N_13537);
xor U14785 (N_14785,N_13963,N_13654);
or U14786 (N_14786,N_13918,N_13512);
nor U14787 (N_14787,N_13917,N_13790);
nand U14788 (N_14788,N_13517,N_13838);
nand U14789 (N_14789,N_13582,N_14101);
xor U14790 (N_14790,N_13816,N_13552);
nor U14791 (N_14791,N_14133,N_13708);
nor U14792 (N_14792,N_13607,N_13603);
or U14793 (N_14793,N_14177,N_13840);
nand U14794 (N_14794,N_13978,N_13670);
nor U14795 (N_14795,N_14076,N_13785);
nand U14796 (N_14796,N_13656,N_14212);
xor U14797 (N_14797,N_13752,N_14103);
nor U14798 (N_14798,N_13725,N_14208);
or U14799 (N_14799,N_13874,N_13590);
or U14800 (N_14800,N_13965,N_13783);
nand U14801 (N_14801,N_13753,N_14009);
and U14802 (N_14802,N_13665,N_14156);
nand U14803 (N_14803,N_13757,N_13944);
nand U14804 (N_14804,N_13968,N_13999);
or U14805 (N_14805,N_14187,N_14096);
nand U14806 (N_14806,N_13602,N_13719);
xnor U14807 (N_14807,N_13582,N_14208);
nand U14808 (N_14808,N_13860,N_14069);
nand U14809 (N_14809,N_14156,N_13980);
nand U14810 (N_14810,N_14235,N_13893);
and U14811 (N_14811,N_13925,N_14210);
nor U14812 (N_14812,N_13512,N_13669);
and U14813 (N_14813,N_13585,N_14041);
xor U14814 (N_14814,N_14244,N_13773);
nand U14815 (N_14815,N_13866,N_13978);
xnor U14816 (N_14816,N_13829,N_13511);
nor U14817 (N_14817,N_14068,N_14176);
or U14818 (N_14818,N_13833,N_14128);
or U14819 (N_14819,N_13969,N_14129);
or U14820 (N_14820,N_13565,N_13680);
and U14821 (N_14821,N_13929,N_13546);
and U14822 (N_14822,N_14218,N_13942);
nand U14823 (N_14823,N_13856,N_13811);
nor U14824 (N_14824,N_14017,N_13518);
nor U14825 (N_14825,N_13608,N_13815);
nor U14826 (N_14826,N_13602,N_14029);
nor U14827 (N_14827,N_13654,N_14035);
or U14828 (N_14828,N_13925,N_14240);
nand U14829 (N_14829,N_13727,N_14049);
or U14830 (N_14830,N_13588,N_13571);
and U14831 (N_14831,N_13544,N_14063);
and U14832 (N_14832,N_14016,N_14001);
nand U14833 (N_14833,N_14079,N_13643);
and U14834 (N_14834,N_13552,N_14022);
nor U14835 (N_14835,N_13925,N_13978);
nand U14836 (N_14836,N_13886,N_14150);
nand U14837 (N_14837,N_14215,N_14205);
and U14838 (N_14838,N_13920,N_13996);
nor U14839 (N_14839,N_14118,N_13700);
xnor U14840 (N_14840,N_13625,N_13940);
nand U14841 (N_14841,N_13775,N_13841);
and U14842 (N_14842,N_14086,N_13830);
nand U14843 (N_14843,N_14011,N_13686);
nor U14844 (N_14844,N_13951,N_13843);
nand U14845 (N_14845,N_14168,N_13988);
nand U14846 (N_14846,N_13696,N_13913);
nand U14847 (N_14847,N_13587,N_13867);
xnor U14848 (N_14848,N_13593,N_14094);
nor U14849 (N_14849,N_13643,N_13645);
and U14850 (N_14850,N_13970,N_13733);
nor U14851 (N_14851,N_13716,N_13806);
nand U14852 (N_14852,N_13878,N_13659);
or U14853 (N_14853,N_14154,N_13952);
nand U14854 (N_14854,N_13831,N_13895);
and U14855 (N_14855,N_13766,N_13510);
nand U14856 (N_14856,N_14040,N_13862);
or U14857 (N_14857,N_13749,N_14033);
or U14858 (N_14858,N_13820,N_13541);
and U14859 (N_14859,N_14243,N_13833);
nand U14860 (N_14860,N_13988,N_13888);
or U14861 (N_14861,N_13749,N_13512);
nor U14862 (N_14862,N_13588,N_14197);
nand U14863 (N_14863,N_14003,N_14221);
nand U14864 (N_14864,N_14046,N_13588);
xor U14865 (N_14865,N_13722,N_14215);
and U14866 (N_14866,N_13922,N_13759);
nor U14867 (N_14867,N_13595,N_13984);
nor U14868 (N_14868,N_14189,N_14054);
or U14869 (N_14869,N_14087,N_13506);
nand U14870 (N_14870,N_13885,N_13830);
or U14871 (N_14871,N_13731,N_14239);
nand U14872 (N_14872,N_14027,N_13840);
or U14873 (N_14873,N_13521,N_14243);
or U14874 (N_14874,N_13609,N_13904);
and U14875 (N_14875,N_14192,N_13928);
nand U14876 (N_14876,N_14000,N_13756);
xnor U14877 (N_14877,N_13691,N_13832);
or U14878 (N_14878,N_14129,N_13635);
and U14879 (N_14879,N_13881,N_13924);
nor U14880 (N_14880,N_14142,N_13550);
or U14881 (N_14881,N_13633,N_13529);
nand U14882 (N_14882,N_13665,N_13824);
nand U14883 (N_14883,N_14105,N_13881);
or U14884 (N_14884,N_14041,N_14176);
nand U14885 (N_14885,N_14105,N_13543);
nand U14886 (N_14886,N_13765,N_13866);
nor U14887 (N_14887,N_14002,N_13545);
and U14888 (N_14888,N_13524,N_14229);
nor U14889 (N_14889,N_14008,N_13804);
nand U14890 (N_14890,N_13956,N_13913);
or U14891 (N_14891,N_13535,N_13579);
or U14892 (N_14892,N_13965,N_13786);
nor U14893 (N_14893,N_14132,N_14017);
or U14894 (N_14894,N_13848,N_13599);
xnor U14895 (N_14895,N_13517,N_14125);
nand U14896 (N_14896,N_13704,N_13682);
or U14897 (N_14897,N_14039,N_13717);
nand U14898 (N_14898,N_13820,N_14129);
nand U14899 (N_14899,N_13933,N_14007);
nor U14900 (N_14900,N_13671,N_14004);
or U14901 (N_14901,N_13902,N_13858);
xor U14902 (N_14902,N_13737,N_14097);
xnor U14903 (N_14903,N_14078,N_13851);
nand U14904 (N_14904,N_13693,N_14083);
nand U14905 (N_14905,N_13544,N_13506);
nand U14906 (N_14906,N_13525,N_14058);
nor U14907 (N_14907,N_14028,N_13566);
nor U14908 (N_14908,N_13775,N_13580);
or U14909 (N_14909,N_13790,N_14141);
or U14910 (N_14910,N_14011,N_14202);
and U14911 (N_14911,N_14244,N_14248);
nor U14912 (N_14912,N_13564,N_14160);
nand U14913 (N_14913,N_14002,N_13915);
nand U14914 (N_14914,N_14096,N_13526);
or U14915 (N_14915,N_13745,N_13539);
nand U14916 (N_14916,N_14107,N_14231);
nor U14917 (N_14917,N_13558,N_14105);
or U14918 (N_14918,N_14092,N_13536);
or U14919 (N_14919,N_13878,N_14042);
nand U14920 (N_14920,N_13874,N_13746);
nor U14921 (N_14921,N_13791,N_14130);
and U14922 (N_14922,N_13926,N_14068);
nor U14923 (N_14923,N_13808,N_14073);
nor U14924 (N_14924,N_13538,N_13690);
nor U14925 (N_14925,N_13694,N_13756);
and U14926 (N_14926,N_13684,N_13622);
or U14927 (N_14927,N_14148,N_13932);
and U14928 (N_14928,N_14073,N_13924);
nand U14929 (N_14929,N_13957,N_14087);
nor U14930 (N_14930,N_14188,N_14216);
or U14931 (N_14931,N_13747,N_13889);
nand U14932 (N_14932,N_14187,N_13843);
nand U14933 (N_14933,N_13852,N_13636);
or U14934 (N_14934,N_13573,N_13779);
xnor U14935 (N_14935,N_13503,N_13877);
nand U14936 (N_14936,N_13980,N_13870);
nand U14937 (N_14937,N_14022,N_13826);
nor U14938 (N_14938,N_14162,N_14229);
or U14939 (N_14939,N_13693,N_14141);
or U14940 (N_14940,N_13580,N_13897);
nand U14941 (N_14941,N_13541,N_14168);
or U14942 (N_14942,N_14127,N_13629);
nor U14943 (N_14943,N_13548,N_14057);
nand U14944 (N_14944,N_13673,N_13736);
and U14945 (N_14945,N_13920,N_13536);
xnor U14946 (N_14946,N_13598,N_14151);
nor U14947 (N_14947,N_14164,N_13827);
or U14948 (N_14948,N_13708,N_13792);
or U14949 (N_14949,N_13939,N_13963);
or U14950 (N_14950,N_13505,N_14222);
nand U14951 (N_14951,N_13834,N_13580);
xor U14952 (N_14952,N_14202,N_13929);
and U14953 (N_14953,N_13621,N_13974);
nand U14954 (N_14954,N_13548,N_13641);
nor U14955 (N_14955,N_14168,N_13504);
xnor U14956 (N_14956,N_13503,N_13595);
and U14957 (N_14957,N_13853,N_14072);
nor U14958 (N_14958,N_14100,N_13718);
nand U14959 (N_14959,N_13665,N_14119);
and U14960 (N_14960,N_13662,N_14132);
nand U14961 (N_14961,N_13876,N_13527);
nor U14962 (N_14962,N_13829,N_13578);
and U14963 (N_14963,N_14238,N_14060);
or U14964 (N_14964,N_13850,N_13764);
nand U14965 (N_14965,N_14177,N_13891);
or U14966 (N_14966,N_13683,N_14150);
nor U14967 (N_14967,N_13960,N_13510);
xnor U14968 (N_14968,N_13762,N_13701);
or U14969 (N_14969,N_13554,N_13822);
nand U14970 (N_14970,N_14069,N_13981);
and U14971 (N_14971,N_13979,N_13690);
and U14972 (N_14972,N_13930,N_13752);
and U14973 (N_14973,N_13881,N_14207);
nor U14974 (N_14974,N_13967,N_14102);
or U14975 (N_14975,N_13510,N_13728);
nand U14976 (N_14976,N_14011,N_14141);
or U14977 (N_14977,N_13691,N_13833);
and U14978 (N_14978,N_14185,N_13520);
nand U14979 (N_14979,N_14064,N_14002);
nand U14980 (N_14980,N_14120,N_14094);
nor U14981 (N_14981,N_13973,N_13936);
nand U14982 (N_14982,N_14164,N_13823);
and U14983 (N_14983,N_13805,N_13877);
or U14984 (N_14984,N_14013,N_13927);
nor U14985 (N_14985,N_13519,N_13785);
nand U14986 (N_14986,N_13747,N_13546);
and U14987 (N_14987,N_14060,N_14180);
nor U14988 (N_14988,N_14069,N_14210);
nand U14989 (N_14989,N_14197,N_13967);
nor U14990 (N_14990,N_13723,N_13536);
or U14991 (N_14991,N_13780,N_13846);
or U14992 (N_14992,N_13804,N_13551);
xor U14993 (N_14993,N_14187,N_13864);
or U14994 (N_14994,N_13691,N_13751);
nor U14995 (N_14995,N_13512,N_13863);
nor U14996 (N_14996,N_13777,N_14076);
and U14997 (N_14997,N_13757,N_14118);
xor U14998 (N_14998,N_13759,N_13619);
nand U14999 (N_14999,N_14189,N_14022);
or UO_0 (O_0,N_14267,N_14469);
and UO_1 (O_1,N_14991,N_14681);
or UO_2 (O_2,N_14397,N_14440);
and UO_3 (O_3,N_14865,N_14254);
and UO_4 (O_4,N_14492,N_14750);
nor UO_5 (O_5,N_14886,N_14639);
nor UO_6 (O_6,N_14498,N_14420);
or UO_7 (O_7,N_14474,N_14996);
nor UO_8 (O_8,N_14418,N_14411);
or UO_9 (O_9,N_14346,N_14501);
nor UO_10 (O_10,N_14803,N_14818);
xor UO_11 (O_11,N_14392,N_14867);
and UO_12 (O_12,N_14964,N_14793);
or UO_13 (O_13,N_14298,N_14527);
nor UO_14 (O_14,N_14836,N_14443);
and UO_15 (O_15,N_14723,N_14599);
or UO_16 (O_16,N_14568,N_14591);
nor UO_17 (O_17,N_14938,N_14871);
nand UO_18 (O_18,N_14559,N_14995);
and UO_19 (O_19,N_14481,N_14905);
nand UO_20 (O_20,N_14330,N_14837);
nand UO_21 (O_21,N_14699,N_14708);
nor UO_22 (O_22,N_14783,N_14388);
xnor UO_23 (O_23,N_14590,N_14302);
and UO_24 (O_24,N_14777,N_14584);
and UO_25 (O_25,N_14759,N_14490);
nor UO_26 (O_26,N_14265,N_14484);
xnor UO_27 (O_27,N_14778,N_14744);
nor UO_28 (O_28,N_14850,N_14251);
nand UO_29 (O_29,N_14350,N_14339);
nor UO_30 (O_30,N_14911,N_14847);
nand UO_31 (O_31,N_14977,N_14518);
and UO_32 (O_32,N_14948,N_14696);
or UO_33 (O_33,N_14770,N_14712);
and UO_34 (O_34,N_14672,N_14675);
xnor UO_35 (O_35,N_14534,N_14371);
nor UO_36 (O_36,N_14937,N_14961);
and UO_37 (O_37,N_14337,N_14835);
nor UO_38 (O_38,N_14451,N_14382);
xor UO_39 (O_39,N_14665,N_14300);
nor UO_40 (O_40,N_14407,N_14378);
nand UO_41 (O_41,N_14351,N_14494);
and UO_42 (O_42,N_14507,N_14500);
and UO_43 (O_43,N_14406,N_14508);
nor UO_44 (O_44,N_14612,N_14873);
nor UO_45 (O_45,N_14656,N_14756);
or UO_46 (O_46,N_14523,N_14618);
and UO_47 (O_47,N_14611,N_14806);
or UO_48 (O_48,N_14594,N_14506);
and UO_49 (O_49,N_14972,N_14983);
and UO_50 (O_50,N_14684,N_14697);
and UO_51 (O_51,N_14277,N_14547);
nand UO_52 (O_52,N_14914,N_14532);
or UO_53 (O_53,N_14817,N_14496);
nand UO_54 (O_54,N_14540,N_14487);
and UO_55 (O_55,N_14311,N_14811);
xnor UO_56 (O_56,N_14260,N_14321);
nand UO_57 (O_57,N_14864,N_14673);
nor UO_58 (O_58,N_14557,N_14910);
xor UO_59 (O_59,N_14934,N_14965);
nand UO_60 (O_60,N_14586,N_14688);
or UO_61 (O_61,N_14472,N_14638);
and UO_62 (O_62,N_14709,N_14876);
and UO_63 (O_63,N_14585,N_14990);
or UO_64 (O_64,N_14630,N_14784);
or UO_65 (O_65,N_14762,N_14671);
nor UO_66 (O_66,N_14366,N_14257);
or UO_67 (O_67,N_14979,N_14434);
or UO_68 (O_68,N_14644,N_14537);
nor UO_69 (O_69,N_14936,N_14520);
nand UO_70 (O_70,N_14450,N_14291);
and UO_71 (O_71,N_14881,N_14926);
nor UO_72 (O_72,N_14308,N_14413);
nor UO_73 (O_73,N_14619,N_14389);
nor UO_74 (O_74,N_14652,N_14600);
nor UO_75 (O_75,N_14538,N_14323);
xnor UO_76 (O_76,N_14814,N_14651);
and UO_77 (O_77,N_14399,N_14355);
nand UO_78 (O_78,N_14356,N_14909);
xnor UO_79 (O_79,N_14889,N_14766);
and UO_80 (O_80,N_14788,N_14272);
and UO_81 (O_81,N_14931,N_14274);
nor UO_82 (O_82,N_14479,N_14952);
nand UO_83 (O_83,N_14513,N_14657);
nand UO_84 (O_84,N_14482,N_14779);
or UO_85 (O_85,N_14276,N_14561);
or UO_86 (O_86,N_14641,N_14872);
or UO_87 (O_87,N_14264,N_14765);
nand UO_88 (O_88,N_14893,N_14429);
nor UO_89 (O_89,N_14691,N_14349);
nand UO_90 (O_90,N_14383,N_14604);
and UO_91 (O_91,N_14992,N_14963);
nand UO_92 (O_92,N_14796,N_14632);
or UO_93 (O_93,N_14425,N_14376);
nand UO_94 (O_94,N_14592,N_14751);
nand UO_95 (O_95,N_14564,N_14296);
and UO_96 (O_96,N_14860,N_14928);
nand UO_97 (O_97,N_14757,N_14966);
and UO_98 (O_98,N_14567,N_14623);
nand UO_99 (O_99,N_14859,N_14993);
or UO_100 (O_100,N_14858,N_14405);
xor UO_101 (O_101,N_14918,N_14721);
xor UO_102 (O_102,N_14637,N_14791);
or UO_103 (O_103,N_14259,N_14728);
nor UO_104 (O_104,N_14875,N_14477);
or UO_105 (O_105,N_14398,N_14700);
or UO_106 (O_106,N_14813,N_14908);
xnor UO_107 (O_107,N_14312,N_14581);
or UO_108 (O_108,N_14655,N_14566);
xor UO_109 (O_109,N_14999,N_14364);
or UO_110 (O_110,N_14774,N_14271);
nor UO_111 (O_111,N_14760,N_14576);
or UO_112 (O_112,N_14845,N_14896);
nor UO_113 (O_113,N_14338,N_14299);
and UO_114 (O_114,N_14678,N_14569);
nand UO_115 (O_115,N_14748,N_14325);
nand UO_116 (O_116,N_14278,N_14828);
xor UO_117 (O_117,N_14769,N_14446);
and UO_118 (O_118,N_14431,N_14626);
and UO_119 (O_119,N_14548,N_14714);
nand UO_120 (O_120,N_14862,N_14840);
nor UO_121 (O_121,N_14453,N_14797);
and UO_122 (O_122,N_14949,N_14415);
or UO_123 (O_123,N_14461,N_14578);
xor UO_124 (O_124,N_14821,N_14574);
and UO_125 (O_125,N_14807,N_14973);
and UO_126 (O_126,N_14336,N_14679);
or UO_127 (O_127,N_14725,N_14776);
or UO_128 (O_128,N_14854,N_14416);
nor UO_129 (O_129,N_14307,N_14556);
nand UO_130 (O_130,N_14393,N_14802);
nor UO_131 (O_131,N_14322,N_14826);
nor UO_132 (O_132,N_14648,N_14629);
or UO_133 (O_133,N_14795,N_14794);
nor UO_134 (O_134,N_14386,N_14633);
and UO_135 (O_135,N_14452,N_14605);
and UO_136 (O_136,N_14941,N_14674);
and UO_137 (O_137,N_14654,N_14717);
or UO_138 (O_138,N_14823,N_14250);
nor UO_139 (O_139,N_14782,N_14562);
or UO_140 (O_140,N_14362,N_14888);
or UO_141 (O_141,N_14516,N_14704);
or UO_142 (O_142,N_14841,N_14852);
and UO_143 (O_143,N_14683,N_14305);
nand UO_144 (O_144,N_14292,N_14583);
or UO_145 (O_145,N_14402,N_14953);
nand UO_146 (O_146,N_14607,N_14763);
nand UO_147 (O_147,N_14460,N_14805);
xor UO_148 (O_148,N_14912,N_14543);
or UO_149 (O_149,N_14514,N_14846);
nand UO_150 (O_150,N_14622,N_14660);
nand UO_151 (O_151,N_14891,N_14359);
xor UO_152 (O_152,N_14377,N_14409);
or UO_153 (O_153,N_14832,N_14736);
xnor UO_154 (O_154,N_14447,N_14943);
nor UO_155 (O_155,N_14869,N_14384);
or UO_156 (O_156,N_14334,N_14710);
and UO_157 (O_157,N_14772,N_14601);
and UO_158 (O_158,N_14758,N_14617);
nand UO_159 (O_159,N_14404,N_14502);
xor UO_160 (O_160,N_14809,N_14635);
nor UO_161 (O_161,N_14539,N_14801);
nor UO_162 (O_162,N_14468,N_14255);
or UO_163 (O_163,N_14764,N_14668);
and UO_164 (O_164,N_14531,N_14987);
nor UO_165 (O_165,N_14483,N_14331);
or UO_166 (O_166,N_14974,N_14833);
nand UO_167 (O_167,N_14844,N_14722);
or UO_168 (O_168,N_14454,N_14658);
and UO_169 (O_169,N_14902,N_14642);
and UO_170 (O_170,N_14495,N_14473);
nand UO_171 (O_171,N_14917,N_14438);
and UO_172 (O_172,N_14609,N_14874);
nor UO_173 (O_173,N_14640,N_14853);
or UO_174 (O_174,N_14426,N_14649);
nand UO_175 (O_175,N_14470,N_14895);
or UO_176 (O_176,N_14742,N_14326);
nor UO_177 (O_177,N_14503,N_14324);
xnor UO_178 (O_178,N_14646,N_14436);
or UO_179 (O_179,N_14702,N_14295);
xnor UO_180 (O_180,N_14551,N_14706);
or UO_181 (O_181,N_14462,N_14690);
nor UO_182 (O_182,N_14478,N_14439);
and UO_183 (O_183,N_14923,N_14903);
nand UO_184 (O_184,N_14560,N_14713);
or UO_185 (O_185,N_14631,N_14705);
nand UO_186 (O_186,N_14512,N_14947);
nand UO_187 (O_187,N_14410,N_14373);
and UO_188 (O_188,N_14353,N_14283);
nand UO_189 (O_189,N_14830,N_14951);
nand UO_190 (O_190,N_14768,N_14374);
nand UO_191 (O_191,N_14510,N_14269);
or UO_192 (O_192,N_14703,N_14724);
nand UO_193 (O_193,N_14975,N_14345);
xnor UO_194 (O_194,N_14739,N_14491);
nor UO_195 (O_195,N_14505,N_14417);
or UO_196 (O_196,N_14695,N_14301);
or UO_197 (O_197,N_14882,N_14341);
or UO_198 (O_198,N_14414,N_14587);
nand UO_199 (O_199,N_14885,N_14541);
or UO_200 (O_200,N_14395,N_14958);
or UO_201 (O_201,N_14616,N_14843);
nand UO_202 (O_202,N_14615,N_14314);
nor UO_203 (O_203,N_14666,N_14424);
and UO_204 (O_204,N_14980,N_14734);
or UO_205 (O_205,N_14596,N_14927);
nand UO_206 (O_206,N_14771,N_14819);
nand UO_207 (O_207,N_14489,N_14754);
nand UO_208 (O_208,N_14707,N_14579);
nand UO_209 (O_209,N_14627,N_14729);
or UO_210 (O_210,N_14313,N_14998);
xor UO_211 (O_211,N_14986,N_14432);
xor UO_212 (O_212,N_14281,N_14730);
nand UO_213 (O_213,N_14342,N_14575);
nor UO_214 (O_214,N_14266,N_14892);
nor UO_215 (O_215,N_14863,N_14256);
nand UO_216 (O_216,N_14643,N_14954);
nor UO_217 (O_217,N_14361,N_14368);
or UO_218 (O_218,N_14906,N_14303);
and UO_219 (O_219,N_14284,N_14970);
and UO_220 (O_220,N_14775,N_14645);
or UO_221 (O_221,N_14682,N_14433);
nand UO_222 (O_222,N_14509,N_14767);
or UO_223 (O_223,N_14427,N_14925);
or UO_224 (O_224,N_14464,N_14667);
xnor UO_225 (O_225,N_14499,N_14827);
nor UO_226 (O_226,N_14270,N_14554);
or UO_227 (O_227,N_14456,N_14620);
or UO_228 (O_228,N_14316,N_14394);
or UO_229 (O_229,N_14780,N_14856);
nand UO_230 (O_230,N_14476,N_14812);
xor UO_231 (O_231,N_14825,N_14530);
or UO_232 (O_232,N_14711,N_14329);
and UO_233 (O_233,N_14957,N_14955);
or UO_234 (O_234,N_14577,N_14380);
and UO_235 (O_235,N_14969,N_14422);
or UO_236 (O_236,N_14465,N_14851);
nor UO_237 (O_237,N_14752,N_14360);
or UO_238 (O_238,N_14740,N_14304);
xnor UO_239 (O_239,N_14610,N_14890);
and UO_240 (O_240,N_14428,N_14718);
and UO_241 (O_241,N_14982,N_14838);
nand UO_242 (O_242,N_14449,N_14275);
and UO_243 (O_243,N_14379,N_14899);
nor UO_244 (O_244,N_14262,N_14933);
and UO_245 (O_245,N_14400,N_14787);
nor UO_246 (O_246,N_14920,N_14458);
or UO_247 (O_247,N_14781,N_14820);
and UO_248 (O_248,N_14901,N_14968);
nand UO_249 (O_249,N_14582,N_14686);
xor UO_250 (O_250,N_14897,N_14363);
nor UO_251 (O_251,N_14997,N_14870);
nor UO_252 (O_252,N_14287,N_14603);
or UO_253 (O_253,N_14286,N_14661);
or UO_254 (O_254,N_14375,N_14685);
nor UO_255 (O_255,N_14544,N_14401);
nor UO_256 (O_256,N_14533,N_14810);
and UO_257 (O_257,N_14753,N_14877);
nor UO_258 (O_258,N_14921,N_14340);
xnor UO_259 (O_259,N_14261,N_14290);
nand UO_260 (O_260,N_14868,N_14799);
and UO_261 (O_261,N_14677,N_14521);
xor UO_262 (O_262,N_14597,N_14546);
nor UO_263 (O_263,N_14669,N_14466);
nand UO_264 (O_264,N_14732,N_14297);
or UO_265 (O_265,N_14459,N_14317);
nand UO_266 (O_266,N_14790,N_14515);
and UO_267 (O_267,N_14357,N_14430);
or UO_268 (O_268,N_14919,N_14602);
nand UO_269 (O_269,N_14369,N_14745);
xor UO_270 (O_270,N_14288,N_14621);
nor UO_271 (O_271,N_14391,N_14913);
nor UO_272 (O_272,N_14589,N_14894);
nor UO_273 (O_273,N_14989,N_14735);
and UO_274 (O_274,N_14967,N_14659);
and UO_275 (O_275,N_14976,N_14940);
nand UO_276 (O_276,N_14570,N_14370);
xnor UO_277 (O_277,N_14984,N_14580);
nand UO_278 (O_278,N_14485,N_14692);
and UO_279 (O_279,N_14552,N_14822);
xnor UO_280 (O_280,N_14831,N_14628);
or UO_281 (O_281,N_14253,N_14800);
nand UO_282 (O_282,N_14842,N_14526);
and UO_283 (O_283,N_14444,N_14318);
nor UO_284 (O_284,N_14571,N_14358);
or UO_285 (O_285,N_14731,N_14932);
or UO_286 (O_286,N_14785,N_14593);
nand UO_287 (O_287,N_14613,N_14789);
xnor UO_288 (O_288,N_14493,N_14598);
nand UO_289 (O_289,N_14719,N_14344);
xnor UO_290 (O_290,N_14252,N_14985);
and UO_291 (O_291,N_14857,N_14480);
nand UO_292 (O_292,N_14348,N_14504);
nand UO_293 (O_293,N_14445,N_14285);
or UO_294 (O_294,N_14848,N_14647);
nor UO_295 (O_295,N_14282,N_14588);
nor UO_296 (O_296,N_14606,N_14834);
and UO_297 (O_297,N_14550,N_14878);
and UO_298 (O_298,N_14945,N_14457);
or UO_299 (O_299,N_14555,N_14372);
nor UO_300 (O_300,N_14930,N_14309);
xnor UO_301 (O_301,N_14693,N_14536);
or UO_302 (O_302,N_14390,N_14475);
nor UO_303 (O_303,N_14978,N_14517);
xnor UO_304 (O_304,N_14944,N_14524);
nor UO_305 (O_305,N_14535,N_14663);
or UO_306 (O_306,N_14289,N_14935);
nor UO_307 (O_307,N_14467,N_14916);
or UO_308 (O_308,N_14542,N_14808);
nor UO_309 (O_309,N_14887,N_14367);
nor UO_310 (O_310,N_14545,N_14662);
nand UO_311 (O_311,N_14981,N_14804);
nand UO_312 (O_312,N_14866,N_14761);
xnor UO_313 (O_313,N_14907,N_14924);
xor UO_314 (O_314,N_14319,N_14962);
or UO_315 (O_315,N_14563,N_14347);
nand UO_316 (O_316,N_14939,N_14861);
or UO_317 (O_317,N_14898,N_14488);
nand UO_318 (O_318,N_14694,N_14403);
or UO_319 (O_319,N_14792,N_14273);
or UO_320 (O_320,N_14883,N_14595);
or UO_321 (O_321,N_14497,N_14994);
nor UO_322 (O_322,N_14715,N_14636);
or UO_323 (O_323,N_14798,N_14315);
and UO_324 (O_324,N_14396,N_14293);
nor UO_325 (O_325,N_14650,N_14354);
nor UO_326 (O_326,N_14884,N_14716);
nand UO_327 (O_327,N_14511,N_14471);
xor UO_328 (O_328,N_14689,N_14855);
and UO_329 (O_329,N_14519,N_14676);
nand UO_330 (O_330,N_14327,N_14333);
nand UO_331 (O_331,N_14335,N_14558);
nand UO_332 (O_332,N_14528,N_14608);
nor UO_333 (O_333,N_14815,N_14687);
nor UO_334 (O_334,N_14680,N_14988);
or UO_335 (O_335,N_14701,N_14922);
xor UO_336 (O_336,N_14829,N_14614);
or UO_337 (O_337,N_14786,N_14448);
and UO_338 (O_338,N_14653,N_14343);
nor UO_339 (O_339,N_14741,N_14733);
and UO_340 (O_340,N_14381,N_14279);
nor UO_341 (O_341,N_14565,N_14720);
and UO_342 (O_342,N_14900,N_14320);
and UO_343 (O_343,N_14306,N_14971);
xnor UO_344 (O_344,N_14664,N_14572);
xor UO_345 (O_345,N_14956,N_14352);
nor UO_346 (O_346,N_14332,N_14950);
and UO_347 (O_347,N_14435,N_14929);
nand UO_348 (O_348,N_14423,N_14529);
or UO_349 (O_349,N_14749,N_14387);
xnor UO_350 (O_350,N_14737,N_14522);
nand UO_351 (O_351,N_14573,N_14879);
nand UO_352 (O_352,N_14904,N_14746);
and UO_353 (O_353,N_14960,N_14942);
nand UO_354 (O_354,N_14412,N_14421);
nor UO_355 (O_355,N_14280,N_14310);
nor UO_356 (O_356,N_14839,N_14553);
and UO_357 (O_357,N_14743,N_14268);
xnor UO_358 (O_358,N_14915,N_14747);
nand UO_359 (O_359,N_14437,N_14263);
nor UO_360 (O_360,N_14625,N_14549);
nor UO_361 (O_361,N_14365,N_14880);
or UO_362 (O_362,N_14442,N_14773);
or UO_363 (O_363,N_14441,N_14634);
nor UO_364 (O_364,N_14738,N_14824);
and UO_365 (O_365,N_14408,N_14755);
or UO_366 (O_366,N_14385,N_14726);
nand UO_367 (O_367,N_14455,N_14486);
nand UO_368 (O_368,N_14727,N_14419);
or UO_369 (O_369,N_14463,N_14670);
nor UO_370 (O_370,N_14959,N_14698);
nor UO_371 (O_371,N_14946,N_14624);
xor UO_372 (O_372,N_14328,N_14258);
or UO_373 (O_373,N_14816,N_14849);
xor UO_374 (O_374,N_14294,N_14525);
nand UO_375 (O_375,N_14777,N_14965);
nand UO_376 (O_376,N_14959,N_14888);
nor UO_377 (O_377,N_14765,N_14513);
or UO_378 (O_378,N_14550,N_14739);
and UO_379 (O_379,N_14555,N_14303);
nor UO_380 (O_380,N_14749,N_14815);
nand UO_381 (O_381,N_14980,N_14943);
nor UO_382 (O_382,N_14404,N_14920);
nor UO_383 (O_383,N_14966,N_14545);
and UO_384 (O_384,N_14744,N_14583);
xnor UO_385 (O_385,N_14577,N_14724);
nor UO_386 (O_386,N_14277,N_14757);
nand UO_387 (O_387,N_14465,N_14423);
nor UO_388 (O_388,N_14939,N_14744);
xnor UO_389 (O_389,N_14431,N_14962);
nand UO_390 (O_390,N_14447,N_14997);
or UO_391 (O_391,N_14561,N_14848);
and UO_392 (O_392,N_14838,N_14662);
xor UO_393 (O_393,N_14746,N_14938);
nand UO_394 (O_394,N_14379,N_14528);
and UO_395 (O_395,N_14572,N_14268);
nor UO_396 (O_396,N_14705,N_14647);
and UO_397 (O_397,N_14835,N_14291);
and UO_398 (O_398,N_14418,N_14665);
and UO_399 (O_399,N_14841,N_14483);
and UO_400 (O_400,N_14555,N_14487);
and UO_401 (O_401,N_14301,N_14374);
and UO_402 (O_402,N_14251,N_14983);
or UO_403 (O_403,N_14841,N_14468);
and UO_404 (O_404,N_14667,N_14849);
and UO_405 (O_405,N_14334,N_14609);
nor UO_406 (O_406,N_14518,N_14494);
nand UO_407 (O_407,N_14714,N_14784);
or UO_408 (O_408,N_14373,N_14381);
nand UO_409 (O_409,N_14767,N_14948);
and UO_410 (O_410,N_14315,N_14503);
nor UO_411 (O_411,N_14626,N_14898);
or UO_412 (O_412,N_14480,N_14754);
nand UO_413 (O_413,N_14302,N_14593);
and UO_414 (O_414,N_14543,N_14428);
or UO_415 (O_415,N_14934,N_14836);
nand UO_416 (O_416,N_14317,N_14280);
nor UO_417 (O_417,N_14449,N_14709);
and UO_418 (O_418,N_14793,N_14845);
nand UO_419 (O_419,N_14797,N_14892);
and UO_420 (O_420,N_14399,N_14691);
nand UO_421 (O_421,N_14890,N_14651);
nand UO_422 (O_422,N_14787,N_14624);
nand UO_423 (O_423,N_14370,N_14485);
xor UO_424 (O_424,N_14883,N_14932);
nand UO_425 (O_425,N_14561,N_14804);
or UO_426 (O_426,N_14946,N_14328);
nor UO_427 (O_427,N_14662,N_14303);
nand UO_428 (O_428,N_14607,N_14327);
and UO_429 (O_429,N_14312,N_14926);
and UO_430 (O_430,N_14492,N_14998);
nand UO_431 (O_431,N_14993,N_14280);
xor UO_432 (O_432,N_14307,N_14792);
nand UO_433 (O_433,N_14612,N_14324);
or UO_434 (O_434,N_14265,N_14649);
nor UO_435 (O_435,N_14818,N_14748);
nor UO_436 (O_436,N_14721,N_14650);
xnor UO_437 (O_437,N_14450,N_14453);
nand UO_438 (O_438,N_14881,N_14942);
or UO_439 (O_439,N_14563,N_14362);
or UO_440 (O_440,N_14279,N_14317);
or UO_441 (O_441,N_14270,N_14297);
or UO_442 (O_442,N_14259,N_14927);
nor UO_443 (O_443,N_14526,N_14415);
nor UO_444 (O_444,N_14848,N_14927);
and UO_445 (O_445,N_14399,N_14440);
and UO_446 (O_446,N_14756,N_14762);
or UO_447 (O_447,N_14621,N_14457);
or UO_448 (O_448,N_14309,N_14881);
nand UO_449 (O_449,N_14581,N_14939);
nor UO_450 (O_450,N_14758,N_14379);
nor UO_451 (O_451,N_14370,N_14860);
or UO_452 (O_452,N_14914,N_14390);
and UO_453 (O_453,N_14792,N_14672);
and UO_454 (O_454,N_14691,N_14505);
and UO_455 (O_455,N_14928,N_14287);
or UO_456 (O_456,N_14253,N_14947);
nor UO_457 (O_457,N_14628,N_14816);
and UO_458 (O_458,N_14948,N_14601);
xor UO_459 (O_459,N_14915,N_14668);
xnor UO_460 (O_460,N_14678,N_14991);
nand UO_461 (O_461,N_14920,N_14836);
and UO_462 (O_462,N_14841,N_14860);
or UO_463 (O_463,N_14334,N_14425);
or UO_464 (O_464,N_14868,N_14714);
nand UO_465 (O_465,N_14291,N_14278);
xor UO_466 (O_466,N_14364,N_14840);
nand UO_467 (O_467,N_14422,N_14944);
nor UO_468 (O_468,N_14651,N_14401);
xnor UO_469 (O_469,N_14548,N_14795);
nor UO_470 (O_470,N_14266,N_14782);
or UO_471 (O_471,N_14735,N_14854);
and UO_472 (O_472,N_14288,N_14410);
and UO_473 (O_473,N_14293,N_14295);
nand UO_474 (O_474,N_14434,N_14344);
and UO_475 (O_475,N_14332,N_14679);
and UO_476 (O_476,N_14521,N_14290);
and UO_477 (O_477,N_14927,N_14802);
nand UO_478 (O_478,N_14747,N_14971);
nor UO_479 (O_479,N_14672,N_14690);
or UO_480 (O_480,N_14895,N_14298);
or UO_481 (O_481,N_14355,N_14713);
and UO_482 (O_482,N_14631,N_14693);
or UO_483 (O_483,N_14788,N_14290);
or UO_484 (O_484,N_14497,N_14409);
or UO_485 (O_485,N_14798,N_14465);
and UO_486 (O_486,N_14675,N_14277);
nand UO_487 (O_487,N_14719,N_14771);
or UO_488 (O_488,N_14914,N_14768);
and UO_489 (O_489,N_14613,N_14679);
xor UO_490 (O_490,N_14488,N_14422);
xor UO_491 (O_491,N_14291,N_14708);
nand UO_492 (O_492,N_14394,N_14670);
nor UO_493 (O_493,N_14328,N_14302);
or UO_494 (O_494,N_14780,N_14629);
nor UO_495 (O_495,N_14570,N_14486);
and UO_496 (O_496,N_14705,N_14383);
nand UO_497 (O_497,N_14972,N_14800);
or UO_498 (O_498,N_14745,N_14417);
or UO_499 (O_499,N_14846,N_14900);
and UO_500 (O_500,N_14791,N_14510);
nor UO_501 (O_501,N_14488,N_14809);
nand UO_502 (O_502,N_14541,N_14940);
nand UO_503 (O_503,N_14826,N_14837);
nor UO_504 (O_504,N_14741,N_14381);
or UO_505 (O_505,N_14876,N_14805);
or UO_506 (O_506,N_14307,N_14911);
and UO_507 (O_507,N_14848,N_14420);
nor UO_508 (O_508,N_14645,N_14963);
nand UO_509 (O_509,N_14724,N_14314);
or UO_510 (O_510,N_14470,N_14667);
xor UO_511 (O_511,N_14383,N_14670);
and UO_512 (O_512,N_14927,N_14477);
nand UO_513 (O_513,N_14288,N_14942);
and UO_514 (O_514,N_14347,N_14969);
xnor UO_515 (O_515,N_14766,N_14470);
or UO_516 (O_516,N_14342,N_14444);
or UO_517 (O_517,N_14841,N_14983);
nor UO_518 (O_518,N_14788,N_14280);
or UO_519 (O_519,N_14357,N_14992);
nand UO_520 (O_520,N_14354,N_14702);
nand UO_521 (O_521,N_14775,N_14688);
and UO_522 (O_522,N_14908,N_14616);
or UO_523 (O_523,N_14540,N_14475);
or UO_524 (O_524,N_14316,N_14975);
nor UO_525 (O_525,N_14645,N_14525);
and UO_526 (O_526,N_14400,N_14709);
or UO_527 (O_527,N_14909,N_14438);
nor UO_528 (O_528,N_14328,N_14772);
and UO_529 (O_529,N_14614,N_14280);
or UO_530 (O_530,N_14622,N_14546);
nand UO_531 (O_531,N_14427,N_14836);
nand UO_532 (O_532,N_14580,N_14594);
and UO_533 (O_533,N_14621,N_14653);
and UO_534 (O_534,N_14598,N_14930);
nor UO_535 (O_535,N_14437,N_14733);
nand UO_536 (O_536,N_14332,N_14915);
xnor UO_537 (O_537,N_14436,N_14566);
xor UO_538 (O_538,N_14661,N_14930);
and UO_539 (O_539,N_14279,N_14868);
xnor UO_540 (O_540,N_14569,N_14493);
nand UO_541 (O_541,N_14646,N_14731);
or UO_542 (O_542,N_14478,N_14972);
nor UO_543 (O_543,N_14731,N_14694);
nand UO_544 (O_544,N_14638,N_14367);
nor UO_545 (O_545,N_14767,N_14724);
nor UO_546 (O_546,N_14875,N_14804);
nand UO_547 (O_547,N_14251,N_14545);
nand UO_548 (O_548,N_14739,N_14263);
and UO_549 (O_549,N_14884,N_14450);
xnor UO_550 (O_550,N_14764,N_14648);
or UO_551 (O_551,N_14731,N_14262);
nand UO_552 (O_552,N_14466,N_14674);
and UO_553 (O_553,N_14692,N_14527);
nand UO_554 (O_554,N_14994,N_14626);
or UO_555 (O_555,N_14711,N_14362);
and UO_556 (O_556,N_14274,N_14458);
xnor UO_557 (O_557,N_14466,N_14860);
xnor UO_558 (O_558,N_14374,N_14367);
and UO_559 (O_559,N_14354,N_14911);
or UO_560 (O_560,N_14806,N_14841);
nor UO_561 (O_561,N_14397,N_14340);
nor UO_562 (O_562,N_14840,N_14469);
nor UO_563 (O_563,N_14330,N_14555);
nor UO_564 (O_564,N_14414,N_14626);
and UO_565 (O_565,N_14435,N_14972);
nand UO_566 (O_566,N_14604,N_14842);
xnor UO_567 (O_567,N_14514,N_14864);
or UO_568 (O_568,N_14349,N_14443);
nand UO_569 (O_569,N_14736,N_14746);
and UO_570 (O_570,N_14385,N_14597);
or UO_571 (O_571,N_14632,N_14473);
nand UO_572 (O_572,N_14759,N_14670);
and UO_573 (O_573,N_14522,N_14777);
and UO_574 (O_574,N_14923,N_14317);
nor UO_575 (O_575,N_14268,N_14300);
and UO_576 (O_576,N_14604,N_14576);
and UO_577 (O_577,N_14267,N_14312);
nor UO_578 (O_578,N_14608,N_14562);
nand UO_579 (O_579,N_14650,N_14641);
nor UO_580 (O_580,N_14793,N_14902);
nor UO_581 (O_581,N_14663,N_14760);
and UO_582 (O_582,N_14640,N_14540);
xnor UO_583 (O_583,N_14715,N_14873);
and UO_584 (O_584,N_14553,N_14517);
and UO_585 (O_585,N_14281,N_14392);
and UO_586 (O_586,N_14826,N_14378);
xor UO_587 (O_587,N_14429,N_14607);
or UO_588 (O_588,N_14737,N_14266);
and UO_589 (O_589,N_14377,N_14790);
or UO_590 (O_590,N_14948,N_14748);
or UO_591 (O_591,N_14250,N_14576);
or UO_592 (O_592,N_14539,N_14654);
nor UO_593 (O_593,N_14914,N_14907);
or UO_594 (O_594,N_14712,N_14844);
nand UO_595 (O_595,N_14486,N_14481);
or UO_596 (O_596,N_14723,N_14707);
nand UO_597 (O_597,N_14761,N_14806);
or UO_598 (O_598,N_14995,N_14369);
nand UO_599 (O_599,N_14475,N_14794);
xor UO_600 (O_600,N_14466,N_14901);
or UO_601 (O_601,N_14999,N_14486);
or UO_602 (O_602,N_14866,N_14890);
xnor UO_603 (O_603,N_14440,N_14675);
and UO_604 (O_604,N_14839,N_14654);
nor UO_605 (O_605,N_14971,N_14446);
nor UO_606 (O_606,N_14829,N_14366);
nor UO_607 (O_607,N_14278,N_14614);
or UO_608 (O_608,N_14926,N_14797);
or UO_609 (O_609,N_14905,N_14537);
and UO_610 (O_610,N_14261,N_14884);
or UO_611 (O_611,N_14969,N_14818);
or UO_612 (O_612,N_14476,N_14416);
nand UO_613 (O_613,N_14821,N_14829);
and UO_614 (O_614,N_14789,N_14616);
or UO_615 (O_615,N_14740,N_14345);
nand UO_616 (O_616,N_14263,N_14910);
and UO_617 (O_617,N_14454,N_14366);
or UO_618 (O_618,N_14308,N_14625);
and UO_619 (O_619,N_14274,N_14477);
or UO_620 (O_620,N_14618,N_14782);
xnor UO_621 (O_621,N_14409,N_14327);
nor UO_622 (O_622,N_14892,N_14844);
or UO_623 (O_623,N_14313,N_14912);
and UO_624 (O_624,N_14367,N_14425);
or UO_625 (O_625,N_14898,N_14684);
nor UO_626 (O_626,N_14435,N_14586);
or UO_627 (O_627,N_14471,N_14465);
and UO_628 (O_628,N_14779,N_14658);
nand UO_629 (O_629,N_14842,N_14780);
and UO_630 (O_630,N_14845,N_14952);
nor UO_631 (O_631,N_14908,N_14606);
or UO_632 (O_632,N_14580,N_14414);
nor UO_633 (O_633,N_14830,N_14884);
nor UO_634 (O_634,N_14896,N_14867);
nand UO_635 (O_635,N_14926,N_14822);
and UO_636 (O_636,N_14921,N_14717);
nor UO_637 (O_637,N_14871,N_14497);
or UO_638 (O_638,N_14604,N_14837);
nor UO_639 (O_639,N_14306,N_14524);
nand UO_640 (O_640,N_14435,N_14861);
or UO_641 (O_641,N_14400,N_14951);
and UO_642 (O_642,N_14359,N_14820);
nor UO_643 (O_643,N_14677,N_14673);
and UO_644 (O_644,N_14535,N_14962);
or UO_645 (O_645,N_14554,N_14751);
xor UO_646 (O_646,N_14446,N_14779);
nor UO_647 (O_647,N_14789,N_14637);
nand UO_648 (O_648,N_14532,N_14406);
and UO_649 (O_649,N_14861,N_14357);
and UO_650 (O_650,N_14485,N_14556);
nand UO_651 (O_651,N_14908,N_14507);
nor UO_652 (O_652,N_14422,N_14782);
or UO_653 (O_653,N_14514,N_14998);
nand UO_654 (O_654,N_14538,N_14551);
nand UO_655 (O_655,N_14296,N_14319);
nor UO_656 (O_656,N_14709,N_14631);
nand UO_657 (O_657,N_14613,N_14300);
nor UO_658 (O_658,N_14495,N_14667);
nand UO_659 (O_659,N_14951,N_14818);
nand UO_660 (O_660,N_14590,N_14997);
or UO_661 (O_661,N_14538,N_14739);
or UO_662 (O_662,N_14365,N_14567);
nand UO_663 (O_663,N_14778,N_14494);
and UO_664 (O_664,N_14804,N_14701);
nand UO_665 (O_665,N_14509,N_14891);
nor UO_666 (O_666,N_14673,N_14981);
nand UO_667 (O_667,N_14840,N_14441);
nor UO_668 (O_668,N_14502,N_14532);
or UO_669 (O_669,N_14864,N_14411);
or UO_670 (O_670,N_14699,N_14278);
nand UO_671 (O_671,N_14675,N_14505);
nor UO_672 (O_672,N_14448,N_14971);
nor UO_673 (O_673,N_14894,N_14869);
nand UO_674 (O_674,N_14273,N_14550);
and UO_675 (O_675,N_14616,N_14947);
nor UO_676 (O_676,N_14995,N_14806);
nand UO_677 (O_677,N_14754,N_14774);
and UO_678 (O_678,N_14973,N_14785);
and UO_679 (O_679,N_14262,N_14948);
and UO_680 (O_680,N_14479,N_14887);
nor UO_681 (O_681,N_14869,N_14682);
nand UO_682 (O_682,N_14941,N_14987);
or UO_683 (O_683,N_14704,N_14348);
nor UO_684 (O_684,N_14898,N_14908);
and UO_685 (O_685,N_14669,N_14592);
or UO_686 (O_686,N_14446,N_14529);
or UO_687 (O_687,N_14346,N_14446);
nand UO_688 (O_688,N_14999,N_14670);
or UO_689 (O_689,N_14446,N_14308);
nor UO_690 (O_690,N_14653,N_14784);
or UO_691 (O_691,N_14356,N_14893);
or UO_692 (O_692,N_14779,N_14478);
nor UO_693 (O_693,N_14537,N_14821);
nand UO_694 (O_694,N_14650,N_14760);
and UO_695 (O_695,N_14766,N_14392);
xnor UO_696 (O_696,N_14250,N_14666);
and UO_697 (O_697,N_14833,N_14363);
or UO_698 (O_698,N_14485,N_14891);
and UO_699 (O_699,N_14661,N_14537);
nor UO_700 (O_700,N_14457,N_14729);
xnor UO_701 (O_701,N_14874,N_14999);
nand UO_702 (O_702,N_14963,N_14631);
or UO_703 (O_703,N_14265,N_14600);
xnor UO_704 (O_704,N_14572,N_14285);
and UO_705 (O_705,N_14675,N_14413);
nor UO_706 (O_706,N_14995,N_14735);
and UO_707 (O_707,N_14453,N_14692);
and UO_708 (O_708,N_14363,N_14740);
and UO_709 (O_709,N_14754,N_14923);
and UO_710 (O_710,N_14705,N_14274);
or UO_711 (O_711,N_14667,N_14480);
or UO_712 (O_712,N_14599,N_14677);
and UO_713 (O_713,N_14544,N_14699);
nor UO_714 (O_714,N_14484,N_14731);
or UO_715 (O_715,N_14471,N_14713);
nand UO_716 (O_716,N_14885,N_14722);
xnor UO_717 (O_717,N_14356,N_14791);
nand UO_718 (O_718,N_14740,N_14959);
nor UO_719 (O_719,N_14766,N_14377);
and UO_720 (O_720,N_14505,N_14276);
nand UO_721 (O_721,N_14965,N_14588);
xnor UO_722 (O_722,N_14785,N_14451);
or UO_723 (O_723,N_14532,N_14665);
nor UO_724 (O_724,N_14683,N_14295);
nand UO_725 (O_725,N_14400,N_14827);
and UO_726 (O_726,N_14451,N_14606);
xnor UO_727 (O_727,N_14861,N_14672);
and UO_728 (O_728,N_14954,N_14606);
and UO_729 (O_729,N_14856,N_14881);
and UO_730 (O_730,N_14669,N_14363);
or UO_731 (O_731,N_14572,N_14928);
or UO_732 (O_732,N_14432,N_14444);
nand UO_733 (O_733,N_14613,N_14948);
nor UO_734 (O_734,N_14539,N_14787);
and UO_735 (O_735,N_14470,N_14567);
xor UO_736 (O_736,N_14857,N_14885);
nor UO_737 (O_737,N_14767,N_14961);
or UO_738 (O_738,N_14276,N_14288);
xnor UO_739 (O_739,N_14888,N_14780);
and UO_740 (O_740,N_14513,N_14746);
nor UO_741 (O_741,N_14516,N_14958);
nand UO_742 (O_742,N_14625,N_14724);
and UO_743 (O_743,N_14703,N_14709);
or UO_744 (O_744,N_14303,N_14549);
nor UO_745 (O_745,N_14864,N_14725);
nor UO_746 (O_746,N_14528,N_14672);
nor UO_747 (O_747,N_14857,N_14350);
and UO_748 (O_748,N_14917,N_14856);
nor UO_749 (O_749,N_14881,N_14920);
xor UO_750 (O_750,N_14483,N_14621);
nand UO_751 (O_751,N_14674,N_14757);
or UO_752 (O_752,N_14858,N_14580);
nor UO_753 (O_753,N_14381,N_14802);
xor UO_754 (O_754,N_14539,N_14805);
or UO_755 (O_755,N_14334,N_14931);
nand UO_756 (O_756,N_14443,N_14755);
and UO_757 (O_757,N_14918,N_14930);
nor UO_758 (O_758,N_14268,N_14505);
and UO_759 (O_759,N_14869,N_14964);
and UO_760 (O_760,N_14328,N_14964);
nor UO_761 (O_761,N_14849,N_14544);
and UO_762 (O_762,N_14323,N_14725);
or UO_763 (O_763,N_14913,N_14579);
nor UO_764 (O_764,N_14928,N_14680);
nor UO_765 (O_765,N_14466,N_14386);
or UO_766 (O_766,N_14719,N_14889);
and UO_767 (O_767,N_14890,N_14589);
xor UO_768 (O_768,N_14787,N_14362);
nor UO_769 (O_769,N_14664,N_14920);
nand UO_770 (O_770,N_14380,N_14533);
nor UO_771 (O_771,N_14618,N_14921);
and UO_772 (O_772,N_14832,N_14702);
xnor UO_773 (O_773,N_14839,N_14683);
nand UO_774 (O_774,N_14788,N_14824);
or UO_775 (O_775,N_14655,N_14719);
or UO_776 (O_776,N_14569,N_14289);
and UO_777 (O_777,N_14499,N_14348);
and UO_778 (O_778,N_14448,N_14444);
nor UO_779 (O_779,N_14570,N_14504);
and UO_780 (O_780,N_14657,N_14875);
nand UO_781 (O_781,N_14570,N_14719);
or UO_782 (O_782,N_14383,N_14710);
nor UO_783 (O_783,N_14431,N_14631);
xnor UO_784 (O_784,N_14688,N_14426);
nor UO_785 (O_785,N_14590,N_14433);
nor UO_786 (O_786,N_14306,N_14762);
nand UO_787 (O_787,N_14602,N_14583);
nor UO_788 (O_788,N_14790,N_14588);
nor UO_789 (O_789,N_14946,N_14725);
and UO_790 (O_790,N_14654,N_14871);
nor UO_791 (O_791,N_14566,N_14439);
or UO_792 (O_792,N_14976,N_14845);
nand UO_793 (O_793,N_14299,N_14809);
nand UO_794 (O_794,N_14861,N_14392);
nor UO_795 (O_795,N_14945,N_14563);
xnor UO_796 (O_796,N_14442,N_14546);
nor UO_797 (O_797,N_14432,N_14485);
or UO_798 (O_798,N_14924,N_14426);
and UO_799 (O_799,N_14604,N_14925);
xnor UO_800 (O_800,N_14995,N_14751);
and UO_801 (O_801,N_14380,N_14667);
nor UO_802 (O_802,N_14408,N_14837);
and UO_803 (O_803,N_14584,N_14910);
or UO_804 (O_804,N_14378,N_14667);
or UO_805 (O_805,N_14479,N_14957);
nand UO_806 (O_806,N_14685,N_14739);
and UO_807 (O_807,N_14823,N_14819);
nor UO_808 (O_808,N_14719,N_14419);
and UO_809 (O_809,N_14422,N_14612);
nand UO_810 (O_810,N_14292,N_14657);
and UO_811 (O_811,N_14539,N_14362);
xnor UO_812 (O_812,N_14448,N_14771);
and UO_813 (O_813,N_14547,N_14296);
nor UO_814 (O_814,N_14701,N_14359);
nor UO_815 (O_815,N_14999,N_14645);
xnor UO_816 (O_816,N_14386,N_14786);
nor UO_817 (O_817,N_14975,N_14733);
xnor UO_818 (O_818,N_14759,N_14629);
nand UO_819 (O_819,N_14562,N_14502);
nand UO_820 (O_820,N_14549,N_14265);
nand UO_821 (O_821,N_14346,N_14355);
or UO_822 (O_822,N_14565,N_14742);
xor UO_823 (O_823,N_14710,N_14793);
nor UO_824 (O_824,N_14367,N_14866);
and UO_825 (O_825,N_14474,N_14363);
nor UO_826 (O_826,N_14779,N_14486);
nor UO_827 (O_827,N_14773,N_14684);
nor UO_828 (O_828,N_14478,N_14255);
xnor UO_829 (O_829,N_14923,N_14811);
nand UO_830 (O_830,N_14761,N_14764);
nand UO_831 (O_831,N_14741,N_14490);
nand UO_832 (O_832,N_14644,N_14865);
and UO_833 (O_833,N_14446,N_14949);
nor UO_834 (O_834,N_14670,N_14572);
nor UO_835 (O_835,N_14369,N_14908);
or UO_836 (O_836,N_14514,N_14883);
and UO_837 (O_837,N_14789,N_14728);
or UO_838 (O_838,N_14430,N_14942);
or UO_839 (O_839,N_14252,N_14296);
and UO_840 (O_840,N_14693,N_14278);
nand UO_841 (O_841,N_14596,N_14661);
nand UO_842 (O_842,N_14922,N_14923);
or UO_843 (O_843,N_14723,N_14738);
nand UO_844 (O_844,N_14959,N_14467);
xnor UO_845 (O_845,N_14301,N_14441);
nand UO_846 (O_846,N_14730,N_14964);
nor UO_847 (O_847,N_14511,N_14740);
nand UO_848 (O_848,N_14922,N_14900);
and UO_849 (O_849,N_14401,N_14612);
or UO_850 (O_850,N_14752,N_14539);
nand UO_851 (O_851,N_14279,N_14853);
nand UO_852 (O_852,N_14589,N_14854);
nand UO_853 (O_853,N_14354,N_14850);
or UO_854 (O_854,N_14924,N_14958);
or UO_855 (O_855,N_14288,N_14323);
and UO_856 (O_856,N_14316,N_14675);
or UO_857 (O_857,N_14902,N_14570);
nand UO_858 (O_858,N_14569,N_14367);
xor UO_859 (O_859,N_14578,N_14703);
nor UO_860 (O_860,N_14943,N_14818);
nor UO_861 (O_861,N_14924,N_14748);
xnor UO_862 (O_862,N_14456,N_14749);
xor UO_863 (O_863,N_14886,N_14531);
and UO_864 (O_864,N_14325,N_14397);
nand UO_865 (O_865,N_14482,N_14309);
nor UO_866 (O_866,N_14974,N_14595);
nor UO_867 (O_867,N_14260,N_14972);
nor UO_868 (O_868,N_14586,N_14821);
or UO_869 (O_869,N_14513,N_14903);
or UO_870 (O_870,N_14297,N_14641);
nand UO_871 (O_871,N_14618,N_14544);
nor UO_872 (O_872,N_14615,N_14830);
or UO_873 (O_873,N_14695,N_14931);
nor UO_874 (O_874,N_14625,N_14707);
or UO_875 (O_875,N_14675,N_14366);
nand UO_876 (O_876,N_14752,N_14939);
and UO_877 (O_877,N_14545,N_14482);
nand UO_878 (O_878,N_14946,N_14650);
or UO_879 (O_879,N_14522,N_14975);
or UO_880 (O_880,N_14814,N_14751);
nor UO_881 (O_881,N_14313,N_14757);
nor UO_882 (O_882,N_14342,N_14981);
nor UO_883 (O_883,N_14682,N_14332);
xnor UO_884 (O_884,N_14594,N_14443);
xor UO_885 (O_885,N_14682,N_14286);
nor UO_886 (O_886,N_14471,N_14598);
nor UO_887 (O_887,N_14496,N_14684);
nor UO_888 (O_888,N_14875,N_14771);
and UO_889 (O_889,N_14820,N_14835);
and UO_890 (O_890,N_14859,N_14945);
nand UO_891 (O_891,N_14259,N_14354);
nand UO_892 (O_892,N_14465,N_14972);
nor UO_893 (O_893,N_14276,N_14997);
and UO_894 (O_894,N_14615,N_14763);
or UO_895 (O_895,N_14264,N_14388);
or UO_896 (O_896,N_14410,N_14937);
nand UO_897 (O_897,N_14921,N_14927);
or UO_898 (O_898,N_14801,N_14757);
xnor UO_899 (O_899,N_14860,N_14914);
nor UO_900 (O_900,N_14774,N_14411);
or UO_901 (O_901,N_14687,N_14873);
xnor UO_902 (O_902,N_14452,N_14714);
nor UO_903 (O_903,N_14624,N_14961);
nor UO_904 (O_904,N_14475,N_14413);
nand UO_905 (O_905,N_14918,N_14841);
and UO_906 (O_906,N_14450,N_14789);
and UO_907 (O_907,N_14520,N_14642);
xnor UO_908 (O_908,N_14399,N_14362);
or UO_909 (O_909,N_14906,N_14386);
or UO_910 (O_910,N_14699,N_14656);
or UO_911 (O_911,N_14469,N_14585);
nor UO_912 (O_912,N_14383,N_14578);
xor UO_913 (O_913,N_14519,N_14982);
and UO_914 (O_914,N_14617,N_14744);
or UO_915 (O_915,N_14333,N_14288);
and UO_916 (O_916,N_14638,N_14690);
and UO_917 (O_917,N_14886,N_14274);
nor UO_918 (O_918,N_14948,N_14355);
nor UO_919 (O_919,N_14290,N_14468);
nand UO_920 (O_920,N_14292,N_14367);
or UO_921 (O_921,N_14673,N_14966);
and UO_922 (O_922,N_14389,N_14556);
xor UO_923 (O_923,N_14463,N_14285);
and UO_924 (O_924,N_14281,N_14261);
or UO_925 (O_925,N_14302,N_14300);
and UO_926 (O_926,N_14726,N_14560);
or UO_927 (O_927,N_14774,N_14348);
and UO_928 (O_928,N_14630,N_14976);
nand UO_929 (O_929,N_14512,N_14372);
nor UO_930 (O_930,N_14697,N_14450);
xnor UO_931 (O_931,N_14939,N_14395);
nand UO_932 (O_932,N_14548,N_14524);
nand UO_933 (O_933,N_14600,N_14583);
xnor UO_934 (O_934,N_14742,N_14842);
nor UO_935 (O_935,N_14991,N_14422);
nor UO_936 (O_936,N_14365,N_14872);
nand UO_937 (O_937,N_14278,N_14675);
or UO_938 (O_938,N_14342,N_14617);
and UO_939 (O_939,N_14618,N_14364);
and UO_940 (O_940,N_14484,N_14684);
nor UO_941 (O_941,N_14954,N_14847);
nor UO_942 (O_942,N_14679,N_14282);
nor UO_943 (O_943,N_14689,N_14717);
nor UO_944 (O_944,N_14455,N_14369);
and UO_945 (O_945,N_14577,N_14268);
nand UO_946 (O_946,N_14385,N_14757);
nor UO_947 (O_947,N_14519,N_14744);
xnor UO_948 (O_948,N_14770,N_14645);
nor UO_949 (O_949,N_14571,N_14572);
nand UO_950 (O_950,N_14878,N_14438);
nor UO_951 (O_951,N_14589,N_14865);
nor UO_952 (O_952,N_14500,N_14406);
xnor UO_953 (O_953,N_14258,N_14453);
xor UO_954 (O_954,N_14350,N_14567);
nand UO_955 (O_955,N_14558,N_14607);
nor UO_956 (O_956,N_14738,N_14947);
nand UO_957 (O_957,N_14470,N_14367);
or UO_958 (O_958,N_14639,N_14674);
nand UO_959 (O_959,N_14408,N_14945);
nor UO_960 (O_960,N_14451,N_14622);
nand UO_961 (O_961,N_14731,N_14777);
or UO_962 (O_962,N_14948,N_14303);
nand UO_963 (O_963,N_14317,N_14281);
and UO_964 (O_964,N_14257,N_14824);
and UO_965 (O_965,N_14913,N_14819);
or UO_966 (O_966,N_14509,N_14920);
or UO_967 (O_967,N_14296,N_14630);
or UO_968 (O_968,N_14583,N_14522);
or UO_969 (O_969,N_14302,N_14348);
nand UO_970 (O_970,N_14332,N_14883);
nor UO_971 (O_971,N_14335,N_14354);
and UO_972 (O_972,N_14759,N_14919);
nor UO_973 (O_973,N_14259,N_14832);
or UO_974 (O_974,N_14579,N_14706);
nand UO_975 (O_975,N_14706,N_14716);
nand UO_976 (O_976,N_14420,N_14859);
or UO_977 (O_977,N_14827,N_14929);
or UO_978 (O_978,N_14270,N_14490);
nand UO_979 (O_979,N_14601,N_14616);
nand UO_980 (O_980,N_14517,N_14557);
and UO_981 (O_981,N_14893,N_14602);
and UO_982 (O_982,N_14620,N_14528);
nor UO_983 (O_983,N_14435,N_14261);
nor UO_984 (O_984,N_14816,N_14754);
nand UO_985 (O_985,N_14882,N_14597);
nand UO_986 (O_986,N_14769,N_14616);
and UO_987 (O_987,N_14623,N_14553);
nor UO_988 (O_988,N_14492,N_14994);
nand UO_989 (O_989,N_14580,N_14394);
nand UO_990 (O_990,N_14608,N_14632);
and UO_991 (O_991,N_14670,N_14460);
nand UO_992 (O_992,N_14811,N_14908);
or UO_993 (O_993,N_14328,N_14443);
or UO_994 (O_994,N_14491,N_14407);
or UO_995 (O_995,N_14361,N_14568);
nor UO_996 (O_996,N_14989,N_14667);
nor UO_997 (O_997,N_14634,N_14802);
nand UO_998 (O_998,N_14381,N_14738);
or UO_999 (O_999,N_14839,N_14443);
nor UO_1000 (O_1000,N_14512,N_14783);
and UO_1001 (O_1001,N_14525,N_14684);
and UO_1002 (O_1002,N_14576,N_14406);
or UO_1003 (O_1003,N_14892,N_14992);
or UO_1004 (O_1004,N_14454,N_14730);
or UO_1005 (O_1005,N_14728,N_14753);
nor UO_1006 (O_1006,N_14880,N_14997);
and UO_1007 (O_1007,N_14523,N_14694);
and UO_1008 (O_1008,N_14900,N_14262);
nand UO_1009 (O_1009,N_14747,N_14804);
or UO_1010 (O_1010,N_14502,N_14756);
nor UO_1011 (O_1011,N_14838,N_14454);
and UO_1012 (O_1012,N_14599,N_14977);
nand UO_1013 (O_1013,N_14790,N_14312);
or UO_1014 (O_1014,N_14691,N_14357);
and UO_1015 (O_1015,N_14641,N_14439);
and UO_1016 (O_1016,N_14636,N_14946);
nor UO_1017 (O_1017,N_14754,N_14334);
nand UO_1018 (O_1018,N_14694,N_14384);
and UO_1019 (O_1019,N_14711,N_14987);
xor UO_1020 (O_1020,N_14970,N_14494);
or UO_1021 (O_1021,N_14526,N_14485);
or UO_1022 (O_1022,N_14583,N_14694);
nand UO_1023 (O_1023,N_14538,N_14507);
nor UO_1024 (O_1024,N_14848,N_14754);
nand UO_1025 (O_1025,N_14360,N_14374);
and UO_1026 (O_1026,N_14523,N_14614);
xor UO_1027 (O_1027,N_14671,N_14498);
xor UO_1028 (O_1028,N_14361,N_14535);
and UO_1029 (O_1029,N_14491,N_14384);
and UO_1030 (O_1030,N_14591,N_14579);
and UO_1031 (O_1031,N_14740,N_14844);
nor UO_1032 (O_1032,N_14447,N_14987);
and UO_1033 (O_1033,N_14312,N_14966);
nor UO_1034 (O_1034,N_14391,N_14326);
or UO_1035 (O_1035,N_14913,N_14733);
or UO_1036 (O_1036,N_14567,N_14726);
or UO_1037 (O_1037,N_14408,N_14911);
or UO_1038 (O_1038,N_14957,N_14471);
or UO_1039 (O_1039,N_14465,N_14748);
xnor UO_1040 (O_1040,N_14769,N_14783);
nand UO_1041 (O_1041,N_14819,N_14972);
or UO_1042 (O_1042,N_14802,N_14403);
and UO_1043 (O_1043,N_14694,N_14357);
nor UO_1044 (O_1044,N_14830,N_14806);
and UO_1045 (O_1045,N_14875,N_14573);
nor UO_1046 (O_1046,N_14746,N_14667);
nor UO_1047 (O_1047,N_14989,N_14404);
or UO_1048 (O_1048,N_14526,N_14383);
nand UO_1049 (O_1049,N_14678,N_14327);
nand UO_1050 (O_1050,N_14378,N_14483);
xor UO_1051 (O_1051,N_14538,N_14893);
nand UO_1052 (O_1052,N_14315,N_14443);
nor UO_1053 (O_1053,N_14964,N_14633);
or UO_1054 (O_1054,N_14833,N_14614);
nor UO_1055 (O_1055,N_14590,N_14684);
and UO_1056 (O_1056,N_14990,N_14335);
or UO_1057 (O_1057,N_14316,N_14758);
nor UO_1058 (O_1058,N_14632,N_14788);
nand UO_1059 (O_1059,N_14614,N_14967);
nand UO_1060 (O_1060,N_14727,N_14483);
nand UO_1061 (O_1061,N_14925,N_14257);
nor UO_1062 (O_1062,N_14671,N_14615);
nand UO_1063 (O_1063,N_14656,N_14960);
and UO_1064 (O_1064,N_14627,N_14429);
xor UO_1065 (O_1065,N_14449,N_14476);
and UO_1066 (O_1066,N_14284,N_14434);
or UO_1067 (O_1067,N_14284,N_14343);
nor UO_1068 (O_1068,N_14381,N_14362);
nor UO_1069 (O_1069,N_14994,N_14822);
nor UO_1070 (O_1070,N_14608,N_14385);
or UO_1071 (O_1071,N_14841,N_14309);
nand UO_1072 (O_1072,N_14853,N_14560);
and UO_1073 (O_1073,N_14814,N_14266);
or UO_1074 (O_1074,N_14274,N_14334);
or UO_1075 (O_1075,N_14612,N_14431);
or UO_1076 (O_1076,N_14941,N_14755);
or UO_1077 (O_1077,N_14490,N_14977);
or UO_1078 (O_1078,N_14901,N_14348);
nand UO_1079 (O_1079,N_14894,N_14282);
nand UO_1080 (O_1080,N_14743,N_14755);
nand UO_1081 (O_1081,N_14895,N_14280);
nand UO_1082 (O_1082,N_14268,N_14993);
xnor UO_1083 (O_1083,N_14260,N_14375);
nand UO_1084 (O_1084,N_14541,N_14683);
or UO_1085 (O_1085,N_14901,N_14470);
nand UO_1086 (O_1086,N_14362,N_14869);
nor UO_1087 (O_1087,N_14616,N_14608);
nor UO_1088 (O_1088,N_14800,N_14470);
or UO_1089 (O_1089,N_14531,N_14796);
and UO_1090 (O_1090,N_14799,N_14705);
nand UO_1091 (O_1091,N_14278,N_14473);
or UO_1092 (O_1092,N_14879,N_14873);
or UO_1093 (O_1093,N_14760,N_14453);
nand UO_1094 (O_1094,N_14289,N_14797);
nand UO_1095 (O_1095,N_14275,N_14946);
nand UO_1096 (O_1096,N_14798,N_14932);
or UO_1097 (O_1097,N_14761,N_14338);
or UO_1098 (O_1098,N_14644,N_14532);
or UO_1099 (O_1099,N_14753,N_14371);
xor UO_1100 (O_1100,N_14869,N_14913);
and UO_1101 (O_1101,N_14869,N_14441);
xor UO_1102 (O_1102,N_14949,N_14596);
nand UO_1103 (O_1103,N_14350,N_14783);
and UO_1104 (O_1104,N_14891,N_14360);
nor UO_1105 (O_1105,N_14647,N_14494);
nor UO_1106 (O_1106,N_14547,N_14758);
nand UO_1107 (O_1107,N_14818,N_14382);
or UO_1108 (O_1108,N_14495,N_14915);
nor UO_1109 (O_1109,N_14414,N_14757);
xnor UO_1110 (O_1110,N_14306,N_14820);
nand UO_1111 (O_1111,N_14860,N_14440);
and UO_1112 (O_1112,N_14271,N_14672);
nand UO_1113 (O_1113,N_14422,N_14703);
nand UO_1114 (O_1114,N_14865,N_14928);
or UO_1115 (O_1115,N_14895,N_14908);
nand UO_1116 (O_1116,N_14275,N_14871);
nand UO_1117 (O_1117,N_14701,N_14941);
xnor UO_1118 (O_1118,N_14990,N_14297);
and UO_1119 (O_1119,N_14695,N_14838);
nor UO_1120 (O_1120,N_14414,N_14471);
and UO_1121 (O_1121,N_14472,N_14749);
and UO_1122 (O_1122,N_14651,N_14372);
nand UO_1123 (O_1123,N_14530,N_14789);
and UO_1124 (O_1124,N_14434,N_14982);
or UO_1125 (O_1125,N_14467,N_14724);
and UO_1126 (O_1126,N_14336,N_14650);
nand UO_1127 (O_1127,N_14739,N_14912);
or UO_1128 (O_1128,N_14792,N_14952);
nor UO_1129 (O_1129,N_14315,N_14652);
nor UO_1130 (O_1130,N_14558,N_14434);
and UO_1131 (O_1131,N_14833,N_14391);
or UO_1132 (O_1132,N_14793,N_14614);
or UO_1133 (O_1133,N_14682,N_14522);
nand UO_1134 (O_1134,N_14364,N_14474);
nand UO_1135 (O_1135,N_14610,N_14762);
or UO_1136 (O_1136,N_14524,N_14663);
or UO_1137 (O_1137,N_14610,N_14412);
nand UO_1138 (O_1138,N_14574,N_14601);
nand UO_1139 (O_1139,N_14642,N_14463);
xnor UO_1140 (O_1140,N_14516,N_14757);
xnor UO_1141 (O_1141,N_14497,N_14976);
nand UO_1142 (O_1142,N_14737,N_14598);
and UO_1143 (O_1143,N_14823,N_14383);
nand UO_1144 (O_1144,N_14464,N_14783);
nand UO_1145 (O_1145,N_14842,N_14750);
nand UO_1146 (O_1146,N_14305,N_14587);
nor UO_1147 (O_1147,N_14845,N_14883);
nor UO_1148 (O_1148,N_14733,N_14471);
and UO_1149 (O_1149,N_14727,N_14663);
nand UO_1150 (O_1150,N_14886,N_14991);
xor UO_1151 (O_1151,N_14767,N_14982);
nor UO_1152 (O_1152,N_14470,N_14278);
or UO_1153 (O_1153,N_14990,N_14808);
xor UO_1154 (O_1154,N_14309,N_14483);
and UO_1155 (O_1155,N_14294,N_14978);
xnor UO_1156 (O_1156,N_14837,N_14481);
nor UO_1157 (O_1157,N_14601,N_14476);
xor UO_1158 (O_1158,N_14714,N_14480);
xor UO_1159 (O_1159,N_14816,N_14773);
and UO_1160 (O_1160,N_14710,N_14409);
or UO_1161 (O_1161,N_14844,N_14475);
or UO_1162 (O_1162,N_14717,N_14901);
nor UO_1163 (O_1163,N_14521,N_14863);
and UO_1164 (O_1164,N_14999,N_14416);
nor UO_1165 (O_1165,N_14937,N_14849);
nor UO_1166 (O_1166,N_14942,N_14320);
nand UO_1167 (O_1167,N_14639,N_14344);
and UO_1168 (O_1168,N_14290,N_14754);
nand UO_1169 (O_1169,N_14913,N_14887);
xnor UO_1170 (O_1170,N_14749,N_14604);
nor UO_1171 (O_1171,N_14467,N_14289);
or UO_1172 (O_1172,N_14485,N_14351);
nor UO_1173 (O_1173,N_14298,N_14995);
nor UO_1174 (O_1174,N_14782,N_14453);
nand UO_1175 (O_1175,N_14821,N_14666);
xor UO_1176 (O_1176,N_14694,N_14567);
or UO_1177 (O_1177,N_14360,N_14772);
xor UO_1178 (O_1178,N_14746,N_14711);
or UO_1179 (O_1179,N_14806,N_14893);
nor UO_1180 (O_1180,N_14414,N_14449);
nand UO_1181 (O_1181,N_14746,N_14985);
or UO_1182 (O_1182,N_14997,N_14913);
nor UO_1183 (O_1183,N_14762,N_14909);
or UO_1184 (O_1184,N_14297,N_14903);
nand UO_1185 (O_1185,N_14659,N_14638);
and UO_1186 (O_1186,N_14509,N_14517);
and UO_1187 (O_1187,N_14310,N_14416);
nor UO_1188 (O_1188,N_14836,N_14732);
or UO_1189 (O_1189,N_14721,N_14538);
or UO_1190 (O_1190,N_14558,N_14609);
nor UO_1191 (O_1191,N_14612,N_14645);
nand UO_1192 (O_1192,N_14965,N_14583);
nor UO_1193 (O_1193,N_14412,N_14775);
and UO_1194 (O_1194,N_14298,N_14628);
nand UO_1195 (O_1195,N_14501,N_14603);
nand UO_1196 (O_1196,N_14492,N_14253);
or UO_1197 (O_1197,N_14584,N_14530);
nand UO_1198 (O_1198,N_14968,N_14750);
nor UO_1199 (O_1199,N_14532,N_14571);
nand UO_1200 (O_1200,N_14761,N_14843);
or UO_1201 (O_1201,N_14796,N_14279);
or UO_1202 (O_1202,N_14400,N_14336);
or UO_1203 (O_1203,N_14448,N_14936);
or UO_1204 (O_1204,N_14471,N_14544);
nor UO_1205 (O_1205,N_14351,N_14894);
nand UO_1206 (O_1206,N_14380,N_14783);
and UO_1207 (O_1207,N_14659,N_14936);
and UO_1208 (O_1208,N_14993,N_14844);
or UO_1209 (O_1209,N_14912,N_14374);
nand UO_1210 (O_1210,N_14823,N_14930);
or UO_1211 (O_1211,N_14575,N_14615);
and UO_1212 (O_1212,N_14554,N_14884);
nor UO_1213 (O_1213,N_14881,N_14894);
nand UO_1214 (O_1214,N_14376,N_14561);
or UO_1215 (O_1215,N_14833,N_14688);
or UO_1216 (O_1216,N_14968,N_14638);
or UO_1217 (O_1217,N_14440,N_14327);
nand UO_1218 (O_1218,N_14611,N_14578);
nor UO_1219 (O_1219,N_14542,N_14615);
nand UO_1220 (O_1220,N_14961,N_14597);
nor UO_1221 (O_1221,N_14662,N_14678);
nor UO_1222 (O_1222,N_14310,N_14592);
xor UO_1223 (O_1223,N_14594,N_14884);
nor UO_1224 (O_1224,N_14540,N_14920);
nand UO_1225 (O_1225,N_14429,N_14808);
and UO_1226 (O_1226,N_14631,N_14622);
nor UO_1227 (O_1227,N_14831,N_14483);
and UO_1228 (O_1228,N_14338,N_14559);
and UO_1229 (O_1229,N_14776,N_14485);
nand UO_1230 (O_1230,N_14345,N_14286);
nor UO_1231 (O_1231,N_14642,N_14779);
nand UO_1232 (O_1232,N_14619,N_14928);
nand UO_1233 (O_1233,N_14574,N_14516);
nand UO_1234 (O_1234,N_14603,N_14423);
and UO_1235 (O_1235,N_14572,N_14927);
or UO_1236 (O_1236,N_14288,N_14781);
nor UO_1237 (O_1237,N_14628,N_14413);
and UO_1238 (O_1238,N_14266,N_14368);
or UO_1239 (O_1239,N_14862,N_14642);
and UO_1240 (O_1240,N_14732,N_14537);
and UO_1241 (O_1241,N_14882,N_14916);
and UO_1242 (O_1242,N_14457,N_14438);
nand UO_1243 (O_1243,N_14521,N_14629);
and UO_1244 (O_1244,N_14887,N_14606);
or UO_1245 (O_1245,N_14319,N_14884);
and UO_1246 (O_1246,N_14512,N_14812);
or UO_1247 (O_1247,N_14657,N_14554);
or UO_1248 (O_1248,N_14629,N_14978);
nand UO_1249 (O_1249,N_14504,N_14252);
nor UO_1250 (O_1250,N_14600,N_14530);
and UO_1251 (O_1251,N_14313,N_14848);
nand UO_1252 (O_1252,N_14910,N_14499);
nand UO_1253 (O_1253,N_14433,N_14722);
or UO_1254 (O_1254,N_14706,N_14959);
nor UO_1255 (O_1255,N_14680,N_14285);
nor UO_1256 (O_1256,N_14768,N_14907);
nor UO_1257 (O_1257,N_14561,N_14515);
or UO_1258 (O_1258,N_14538,N_14289);
xnor UO_1259 (O_1259,N_14305,N_14596);
or UO_1260 (O_1260,N_14454,N_14777);
and UO_1261 (O_1261,N_14498,N_14915);
and UO_1262 (O_1262,N_14326,N_14732);
nand UO_1263 (O_1263,N_14816,N_14882);
or UO_1264 (O_1264,N_14842,N_14878);
nand UO_1265 (O_1265,N_14864,N_14450);
or UO_1266 (O_1266,N_14549,N_14748);
xor UO_1267 (O_1267,N_14562,N_14526);
nand UO_1268 (O_1268,N_14646,N_14550);
and UO_1269 (O_1269,N_14690,N_14990);
and UO_1270 (O_1270,N_14260,N_14507);
nand UO_1271 (O_1271,N_14529,N_14923);
nand UO_1272 (O_1272,N_14534,N_14699);
nand UO_1273 (O_1273,N_14460,N_14401);
and UO_1274 (O_1274,N_14583,N_14924);
and UO_1275 (O_1275,N_14964,N_14500);
xnor UO_1276 (O_1276,N_14558,N_14782);
or UO_1277 (O_1277,N_14699,N_14602);
and UO_1278 (O_1278,N_14990,N_14975);
and UO_1279 (O_1279,N_14629,N_14859);
or UO_1280 (O_1280,N_14255,N_14469);
xor UO_1281 (O_1281,N_14817,N_14869);
nand UO_1282 (O_1282,N_14915,N_14997);
nor UO_1283 (O_1283,N_14556,N_14759);
and UO_1284 (O_1284,N_14650,N_14860);
or UO_1285 (O_1285,N_14545,N_14825);
and UO_1286 (O_1286,N_14876,N_14979);
nand UO_1287 (O_1287,N_14338,N_14893);
nor UO_1288 (O_1288,N_14865,N_14378);
nand UO_1289 (O_1289,N_14357,N_14576);
nand UO_1290 (O_1290,N_14298,N_14789);
and UO_1291 (O_1291,N_14447,N_14731);
xor UO_1292 (O_1292,N_14988,N_14484);
or UO_1293 (O_1293,N_14668,N_14552);
or UO_1294 (O_1294,N_14599,N_14992);
and UO_1295 (O_1295,N_14459,N_14993);
or UO_1296 (O_1296,N_14954,N_14700);
nand UO_1297 (O_1297,N_14748,N_14537);
nand UO_1298 (O_1298,N_14743,N_14413);
nor UO_1299 (O_1299,N_14937,N_14689);
or UO_1300 (O_1300,N_14846,N_14427);
and UO_1301 (O_1301,N_14326,N_14500);
and UO_1302 (O_1302,N_14787,N_14434);
or UO_1303 (O_1303,N_14821,N_14335);
nor UO_1304 (O_1304,N_14377,N_14361);
xor UO_1305 (O_1305,N_14481,N_14445);
and UO_1306 (O_1306,N_14734,N_14407);
nor UO_1307 (O_1307,N_14316,N_14593);
nand UO_1308 (O_1308,N_14399,N_14531);
nor UO_1309 (O_1309,N_14539,N_14547);
or UO_1310 (O_1310,N_14676,N_14709);
and UO_1311 (O_1311,N_14756,N_14536);
and UO_1312 (O_1312,N_14513,N_14421);
and UO_1313 (O_1313,N_14378,N_14733);
or UO_1314 (O_1314,N_14315,N_14758);
and UO_1315 (O_1315,N_14851,N_14322);
nor UO_1316 (O_1316,N_14344,N_14869);
or UO_1317 (O_1317,N_14276,N_14702);
nand UO_1318 (O_1318,N_14963,N_14842);
xor UO_1319 (O_1319,N_14728,N_14423);
xnor UO_1320 (O_1320,N_14899,N_14717);
nand UO_1321 (O_1321,N_14605,N_14923);
and UO_1322 (O_1322,N_14854,N_14660);
nand UO_1323 (O_1323,N_14311,N_14760);
nor UO_1324 (O_1324,N_14598,N_14799);
nand UO_1325 (O_1325,N_14405,N_14370);
nor UO_1326 (O_1326,N_14596,N_14381);
or UO_1327 (O_1327,N_14678,N_14799);
nand UO_1328 (O_1328,N_14577,N_14360);
nor UO_1329 (O_1329,N_14703,N_14442);
and UO_1330 (O_1330,N_14508,N_14874);
xor UO_1331 (O_1331,N_14393,N_14966);
nand UO_1332 (O_1332,N_14479,N_14276);
or UO_1333 (O_1333,N_14991,N_14603);
nand UO_1334 (O_1334,N_14420,N_14870);
nor UO_1335 (O_1335,N_14689,N_14646);
and UO_1336 (O_1336,N_14809,N_14978);
nand UO_1337 (O_1337,N_14476,N_14619);
xnor UO_1338 (O_1338,N_14803,N_14611);
nand UO_1339 (O_1339,N_14446,N_14590);
and UO_1340 (O_1340,N_14478,N_14592);
and UO_1341 (O_1341,N_14315,N_14662);
or UO_1342 (O_1342,N_14606,N_14257);
and UO_1343 (O_1343,N_14301,N_14457);
xnor UO_1344 (O_1344,N_14860,N_14522);
nand UO_1345 (O_1345,N_14548,N_14448);
and UO_1346 (O_1346,N_14539,N_14681);
nand UO_1347 (O_1347,N_14880,N_14281);
nand UO_1348 (O_1348,N_14666,N_14732);
or UO_1349 (O_1349,N_14863,N_14983);
nand UO_1350 (O_1350,N_14465,N_14650);
or UO_1351 (O_1351,N_14993,N_14541);
xor UO_1352 (O_1352,N_14354,N_14893);
and UO_1353 (O_1353,N_14729,N_14511);
xor UO_1354 (O_1354,N_14550,N_14698);
and UO_1355 (O_1355,N_14356,N_14921);
and UO_1356 (O_1356,N_14283,N_14503);
or UO_1357 (O_1357,N_14590,N_14652);
nand UO_1358 (O_1358,N_14639,N_14955);
or UO_1359 (O_1359,N_14442,N_14523);
xor UO_1360 (O_1360,N_14761,N_14756);
nor UO_1361 (O_1361,N_14303,N_14413);
and UO_1362 (O_1362,N_14991,N_14755);
nand UO_1363 (O_1363,N_14560,N_14743);
nor UO_1364 (O_1364,N_14746,N_14597);
nor UO_1365 (O_1365,N_14354,N_14898);
nor UO_1366 (O_1366,N_14803,N_14739);
nor UO_1367 (O_1367,N_14586,N_14809);
and UO_1368 (O_1368,N_14266,N_14722);
and UO_1369 (O_1369,N_14433,N_14766);
nor UO_1370 (O_1370,N_14650,N_14909);
and UO_1371 (O_1371,N_14701,N_14801);
xor UO_1372 (O_1372,N_14665,N_14380);
and UO_1373 (O_1373,N_14594,N_14670);
nand UO_1374 (O_1374,N_14415,N_14732);
nand UO_1375 (O_1375,N_14252,N_14478);
nand UO_1376 (O_1376,N_14692,N_14693);
nor UO_1377 (O_1377,N_14861,N_14976);
or UO_1378 (O_1378,N_14594,N_14808);
or UO_1379 (O_1379,N_14908,N_14495);
or UO_1380 (O_1380,N_14949,N_14250);
nor UO_1381 (O_1381,N_14443,N_14946);
or UO_1382 (O_1382,N_14553,N_14611);
and UO_1383 (O_1383,N_14281,N_14255);
or UO_1384 (O_1384,N_14523,N_14877);
and UO_1385 (O_1385,N_14878,N_14341);
nand UO_1386 (O_1386,N_14840,N_14634);
nand UO_1387 (O_1387,N_14340,N_14639);
nand UO_1388 (O_1388,N_14662,N_14390);
nor UO_1389 (O_1389,N_14880,N_14827);
or UO_1390 (O_1390,N_14774,N_14378);
nand UO_1391 (O_1391,N_14888,N_14949);
nand UO_1392 (O_1392,N_14558,N_14665);
nand UO_1393 (O_1393,N_14936,N_14886);
or UO_1394 (O_1394,N_14343,N_14517);
or UO_1395 (O_1395,N_14385,N_14453);
nor UO_1396 (O_1396,N_14601,N_14991);
nand UO_1397 (O_1397,N_14906,N_14535);
nor UO_1398 (O_1398,N_14616,N_14527);
or UO_1399 (O_1399,N_14608,N_14705);
nor UO_1400 (O_1400,N_14770,N_14290);
or UO_1401 (O_1401,N_14697,N_14886);
nor UO_1402 (O_1402,N_14945,N_14739);
nor UO_1403 (O_1403,N_14367,N_14780);
and UO_1404 (O_1404,N_14740,N_14746);
or UO_1405 (O_1405,N_14391,N_14265);
or UO_1406 (O_1406,N_14571,N_14325);
nor UO_1407 (O_1407,N_14293,N_14732);
nor UO_1408 (O_1408,N_14490,N_14880);
xor UO_1409 (O_1409,N_14721,N_14568);
nor UO_1410 (O_1410,N_14937,N_14866);
or UO_1411 (O_1411,N_14384,N_14732);
xor UO_1412 (O_1412,N_14390,N_14997);
or UO_1413 (O_1413,N_14662,N_14487);
and UO_1414 (O_1414,N_14800,N_14671);
nand UO_1415 (O_1415,N_14363,N_14348);
or UO_1416 (O_1416,N_14626,N_14756);
and UO_1417 (O_1417,N_14618,N_14585);
and UO_1418 (O_1418,N_14857,N_14326);
or UO_1419 (O_1419,N_14705,N_14515);
nand UO_1420 (O_1420,N_14969,N_14713);
or UO_1421 (O_1421,N_14955,N_14737);
or UO_1422 (O_1422,N_14721,N_14556);
and UO_1423 (O_1423,N_14574,N_14702);
nand UO_1424 (O_1424,N_14837,N_14319);
nand UO_1425 (O_1425,N_14503,N_14929);
or UO_1426 (O_1426,N_14255,N_14972);
and UO_1427 (O_1427,N_14413,N_14793);
nor UO_1428 (O_1428,N_14281,N_14513);
or UO_1429 (O_1429,N_14904,N_14536);
nand UO_1430 (O_1430,N_14370,N_14730);
nand UO_1431 (O_1431,N_14322,N_14423);
or UO_1432 (O_1432,N_14825,N_14863);
and UO_1433 (O_1433,N_14404,N_14547);
or UO_1434 (O_1434,N_14863,N_14472);
or UO_1435 (O_1435,N_14411,N_14512);
nand UO_1436 (O_1436,N_14742,N_14628);
xnor UO_1437 (O_1437,N_14837,N_14514);
xnor UO_1438 (O_1438,N_14470,N_14397);
nor UO_1439 (O_1439,N_14295,N_14617);
or UO_1440 (O_1440,N_14402,N_14308);
and UO_1441 (O_1441,N_14874,N_14431);
nor UO_1442 (O_1442,N_14877,N_14502);
nor UO_1443 (O_1443,N_14462,N_14864);
nand UO_1444 (O_1444,N_14719,N_14453);
nand UO_1445 (O_1445,N_14865,N_14590);
nand UO_1446 (O_1446,N_14758,N_14727);
and UO_1447 (O_1447,N_14878,N_14405);
xnor UO_1448 (O_1448,N_14994,N_14868);
and UO_1449 (O_1449,N_14994,N_14913);
xnor UO_1450 (O_1450,N_14744,N_14640);
and UO_1451 (O_1451,N_14587,N_14391);
nand UO_1452 (O_1452,N_14602,N_14483);
nand UO_1453 (O_1453,N_14864,N_14317);
or UO_1454 (O_1454,N_14764,N_14563);
nand UO_1455 (O_1455,N_14587,N_14315);
nor UO_1456 (O_1456,N_14343,N_14738);
or UO_1457 (O_1457,N_14928,N_14977);
or UO_1458 (O_1458,N_14431,N_14940);
nor UO_1459 (O_1459,N_14431,N_14664);
nor UO_1460 (O_1460,N_14507,N_14727);
nand UO_1461 (O_1461,N_14423,N_14300);
nand UO_1462 (O_1462,N_14651,N_14784);
xnor UO_1463 (O_1463,N_14597,N_14888);
xnor UO_1464 (O_1464,N_14945,N_14970);
xor UO_1465 (O_1465,N_14288,N_14543);
nor UO_1466 (O_1466,N_14632,N_14570);
nor UO_1467 (O_1467,N_14661,N_14938);
and UO_1468 (O_1468,N_14774,N_14819);
or UO_1469 (O_1469,N_14315,N_14440);
and UO_1470 (O_1470,N_14464,N_14574);
nand UO_1471 (O_1471,N_14799,N_14927);
nor UO_1472 (O_1472,N_14325,N_14718);
and UO_1473 (O_1473,N_14644,N_14312);
or UO_1474 (O_1474,N_14257,N_14407);
nand UO_1475 (O_1475,N_14388,N_14343);
nor UO_1476 (O_1476,N_14753,N_14378);
and UO_1477 (O_1477,N_14611,N_14743);
nor UO_1478 (O_1478,N_14655,N_14876);
and UO_1479 (O_1479,N_14580,N_14450);
or UO_1480 (O_1480,N_14432,N_14583);
and UO_1481 (O_1481,N_14822,N_14804);
nor UO_1482 (O_1482,N_14325,N_14704);
nor UO_1483 (O_1483,N_14508,N_14781);
or UO_1484 (O_1484,N_14640,N_14687);
nand UO_1485 (O_1485,N_14998,N_14519);
or UO_1486 (O_1486,N_14505,N_14999);
nand UO_1487 (O_1487,N_14939,N_14285);
and UO_1488 (O_1488,N_14821,N_14861);
or UO_1489 (O_1489,N_14686,N_14884);
nor UO_1490 (O_1490,N_14458,N_14687);
and UO_1491 (O_1491,N_14794,N_14405);
and UO_1492 (O_1492,N_14873,N_14971);
and UO_1493 (O_1493,N_14744,N_14672);
nor UO_1494 (O_1494,N_14669,N_14314);
nand UO_1495 (O_1495,N_14484,N_14870);
nand UO_1496 (O_1496,N_14721,N_14879);
or UO_1497 (O_1497,N_14534,N_14709);
or UO_1498 (O_1498,N_14372,N_14350);
or UO_1499 (O_1499,N_14779,N_14255);
nand UO_1500 (O_1500,N_14657,N_14668);
xnor UO_1501 (O_1501,N_14324,N_14790);
nand UO_1502 (O_1502,N_14904,N_14976);
and UO_1503 (O_1503,N_14255,N_14481);
or UO_1504 (O_1504,N_14318,N_14445);
nand UO_1505 (O_1505,N_14941,N_14943);
or UO_1506 (O_1506,N_14304,N_14616);
nor UO_1507 (O_1507,N_14345,N_14868);
nand UO_1508 (O_1508,N_14333,N_14317);
nor UO_1509 (O_1509,N_14481,N_14561);
nor UO_1510 (O_1510,N_14680,N_14376);
nor UO_1511 (O_1511,N_14316,N_14835);
nor UO_1512 (O_1512,N_14344,N_14660);
and UO_1513 (O_1513,N_14976,N_14688);
or UO_1514 (O_1514,N_14398,N_14424);
and UO_1515 (O_1515,N_14387,N_14395);
or UO_1516 (O_1516,N_14570,N_14361);
or UO_1517 (O_1517,N_14286,N_14383);
nor UO_1518 (O_1518,N_14318,N_14848);
and UO_1519 (O_1519,N_14615,N_14376);
nor UO_1520 (O_1520,N_14560,N_14372);
or UO_1521 (O_1521,N_14676,N_14566);
nand UO_1522 (O_1522,N_14682,N_14703);
nand UO_1523 (O_1523,N_14251,N_14320);
nor UO_1524 (O_1524,N_14356,N_14430);
nor UO_1525 (O_1525,N_14317,N_14663);
xor UO_1526 (O_1526,N_14915,N_14912);
nand UO_1527 (O_1527,N_14757,N_14917);
or UO_1528 (O_1528,N_14352,N_14863);
and UO_1529 (O_1529,N_14340,N_14428);
nor UO_1530 (O_1530,N_14767,N_14725);
xor UO_1531 (O_1531,N_14460,N_14339);
nor UO_1532 (O_1532,N_14489,N_14727);
or UO_1533 (O_1533,N_14381,N_14429);
nor UO_1534 (O_1534,N_14312,N_14799);
xor UO_1535 (O_1535,N_14987,N_14295);
nor UO_1536 (O_1536,N_14311,N_14635);
or UO_1537 (O_1537,N_14347,N_14678);
nor UO_1538 (O_1538,N_14931,N_14678);
nand UO_1539 (O_1539,N_14675,N_14649);
nor UO_1540 (O_1540,N_14872,N_14602);
or UO_1541 (O_1541,N_14340,N_14400);
or UO_1542 (O_1542,N_14492,N_14785);
and UO_1543 (O_1543,N_14955,N_14393);
nand UO_1544 (O_1544,N_14905,N_14913);
and UO_1545 (O_1545,N_14620,N_14981);
and UO_1546 (O_1546,N_14331,N_14697);
nand UO_1547 (O_1547,N_14705,N_14930);
nand UO_1548 (O_1548,N_14340,N_14265);
xnor UO_1549 (O_1549,N_14468,N_14291);
nor UO_1550 (O_1550,N_14901,N_14528);
or UO_1551 (O_1551,N_14744,N_14993);
nor UO_1552 (O_1552,N_14265,N_14342);
nor UO_1553 (O_1553,N_14802,N_14646);
nor UO_1554 (O_1554,N_14903,N_14420);
nand UO_1555 (O_1555,N_14687,N_14301);
and UO_1556 (O_1556,N_14960,N_14955);
nor UO_1557 (O_1557,N_14682,N_14289);
and UO_1558 (O_1558,N_14430,N_14300);
or UO_1559 (O_1559,N_14824,N_14999);
nor UO_1560 (O_1560,N_14395,N_14342);
nand UO_1561 (O_1561,N_14842,N_14771);
nand UO_1562 (O_1562,N_14857,N_14340);
nor UO_1563 (O_1563,N_14618,N_14659);
nand UO_1564 (O_1564,N_14621,N_14430);
nand UO_1565 (O_1565,N_14625,N_14948);
nor UO_1566 (O_1566,N_14822,N_14739);
nor UO_1567 (O_1567,N_14723,N_14257);
or UO_1568 (O_1568,N_14286,N_14923);
and UO_1569 (O_1569,N_14343,N_14593);
nand UO_1570 (O_1570,N_14998,N_14696);
nand UO_1571 (O_1571,N_14704,N_14448);
or UO_1572 (O_1572,N_14921,N_14823);
and UO_1573 (O_1573,N_14671,N_14643);
and UO_1574 (O_1574,N_14461,N_14789);
nand UO_1575 (O_1575,N_14935,N_14355);
xor UO_1576 (O_1576,N_14616,N_14889);
nand UO_1577 (O_1577,N_14348,N_14486);
nor UO_1578 (O_1578,N_14516,N_14412);
nand UO_1579 (O_1579,N_14361,N_14265);
nand UO_1580 (O_1580,N_14603,N_14357);
and UO_1581 (O_1581,N_14710,N_14538);
and UO_1582 (O_1582,N_14359,N_14512);
nor UO_1583 (O_1583,N_14777,N_14443);
nor UO_1584 (O_1584,N_14644,N_14561);
nor UO_1585 (O_1585,N_14716,N_14628);
nand UO_1586 (O_1586,N_14939,N_14909);
or UO_1587 (O_1587,N_14407,N_14394);
nor UO_1588 (O_1588,N_14505,N_14934);
and UO_1589 (O_1589,N_14790,N_14314);
nand UO_1590 (O_1590,N_14839,N_14835);
and UO_1591 (O_1591,N_14253,N_14839);
xnor UO_1592 (O_1592,N_14654,N_14404);
nor UO_1593 (O_1593,N_14814,N_14446);
nand UO_1594 (O_1594,N_14657,N_14807);
or UO_1595 (O_1595,N_14593,N_14980);
nor UO_1596 (O_1596,N_14517,N_14560);
or UO_1597 (O_1597,N_14928,N_14653);
or UO_1598 (O_1598,N_14625,N_14845);
nand UO_1599 (O_1599,N_14900,N_14896);
nor UO_1600 (O_1600,N_14483,N_14917);
or UO_1601 (O_1601,N_14838,N_14554);
or UO_1602 (O_1602,N_14311,N_14432);
and UO_1603 (O_1603,N_14847,N_14668);
or UO_1604 (O_1604,N_14819,N_14805);
nand UO_1605 (O_1605,N_14323,N_14548);
nand UO_1606 (O_1606,N_14800,N_14547);
xor UO_1607 (O_1607,N_14316,N_14614);
xnor UO_1608 (O_1608,N_14489,N_14548);
and UO_1609 (O_1609,N_14590,N_14911);
or UO_1610 (O_1610,N_14912,N_14529);
nor UO_1611 (O_1611,N_14903,N_14983);
and UO_1612 (O_1612,N_14807,N_14460);
nor UO_1613 (O_1613,N_14702,N_14892);
nor UO_1614 (O_1614,N_14425,N_14918);
nand UO_1615 (O_1615,N_14790,N_14547);
and UO_1616 (O_1616,N_14988,N_14374);
xor UO_1617 (O_1617,N_14989,N_14414);
xnor UO_1618 (O_1618,N_14722,N_14750);
or UO_1619 (O_1619,N_14734,N_14510);
nand UO_1620 (O_1620,N_14818,N_14957);
and UO_1621 (O_1621,N_14379,N_14787);
nand UO_1622 (O_1622,N_14798,N_14675);
or UO_1623 (O_1623,N_14922,N_14876);
nor UO_1624 (O_1624,N_14523,N_14275);
xor UO_1625 (O_1625,N_14894,N_14556);
or UO_1626 (O_1626,N_14774,N_14956);
and UO_1627 (O_1627,N_14724,N_14489);
xnor UO_1628 (O_1628,N_14881,N_14362);
nand UO_1629 (O_1629,N_14582,N_14577);
nand UO_1630 (O_1630,N_14605,N_14802);
xnor UO_1631 (O_1631,N_14573,N_14961);
nor UO_1632 (O_1632,N_14499,N_14540);
xnor UO_1633 (O_1633,N_14269,N_14782);
or UO_1634 (O_1634,N_14700,N_14301);
or UO_1635 (O_1635,N_14843,N_14308);
or UO_1636 (O_1636,N_14303,N_14867);
nand UO_1637 (O_1637,N_14689,N_14653);
nand UO_1638 (O_1638,N_14475,N_14836);
and UO_1639 (O_1639,N_14428,N_14969);
or UO_1640 (O_1640,N_14901,N_14908);
or UO_1641 (O_1641,N_14316,N_14550);
and UO_1642 (O_1642,N_14802,N_14678);
xor UO_1643 (O_1643,N_14363,N_14265);
and UO_1644 (O_1644,N_14891,N_14675);
nor UO_1645 (O_1645,N_14381,N_14256);
or UO_1646 (O_1646,N_14403,N_14895);
nand UO_1647 (O_1647,N_14733,N_14773);
xor UO_1648 (O_1648,N_14671,N_14631);
or UO_1649 (O_1649,N_14397,N_14316);
nor UO_1650 (O_1650,N_14598,N_14263);
and UO_1651 (O_1651,N_14672,N_14964);
and UO_1652 (O_1652,N_14950,N_14304);
or UO_1653 (O_1653,N_14683,N_14330);
and UO_1654 (O_1654,N_14994,N_14701);
and UO_1655 (O_1655,N_14863,N_14940);
and UO_1656 (O_1656,N_14651,N_14710);
nand UO_1657 (O_1657,N_14261,N_14877);
and UO_1658 (O_1658,N_14997,N_14745);
nor UO_1659 (O_1659,N_14615,N_14628);
nand UO_1660 (O_1660,N_14511,N_14571);
or UO_1661 (O_1661,N_14909,N_14497);
or UO_1662 (O_1662,N_14933,N_14649);
nand UO_1663 (O_1663,N_14893,N_14364);
and UO_1664 (O_1664,N_14800,N_14802);
and UO_1665 (O_1665,N_14595,N_14436);
or UO_1666 (O_1666,N_14372,N_14362);
nand UO_1667 (O_1667,N_14959,N_14519);
and UO_1668 (O_1668,N_14458,N_14366);
nand UO_1669 (O_1669,N_14773,N_14862);
or UO_1670 (O_1670,N_14627,N_14427);
nand UO_1671 (O_1671,N_14889,N_14733);
nand UO_1672 (O_1672,N_14582,N_14594);
nor UO_1673 (O_1673,N_14486,N_14391);
nor UO_1674 (O_1674,N_14762,N_14396);
or UO_1675 (O_1675,N_14497,N_14536);
or UO_1676 (O_1676,N_14639,N_14573);
and UO_1677 (O_1677,N_14530,N_14454);
nand UO_1678 (O_1678,N_14307,N_14475);
nor UO_1679 (O_1679,N_14887,N_14570);
nand UO_1680 (O_1680,N_14565,N_14375);
nand UO_1681 (O_1681,N_14376,N_14610);
nor UO_1682 (O_1682,N_14565,N_14598);
and UO_1683 (O_1683,N_14545,N_14370);
nor UO_1684 (O_1684,N_14946,N_14383);
or UO_1685 (O_1685,N_14658,N_14465);
or UO_1686 (O_1686,N_14615,N_14872);
or UO_1687 (O_1687,N_14604,N_14294);
or UO_1688 (O_1688,N_14348,N_14317);
nand UO_1689 (O_1689,N_14250,N_14699);
nor UO_1690 (O_1690,N_14785,N_14548);
or UO_1691 (O_1691,N_14322,N_14293);
nor UO_1692 (O_1692,N_14425,N_14502);
nand UO_1693 (O_1693,N_14740,N_14437);
nor UO_1694 (O_1694,N_14490,N_14293);
or UO_1695 (O_1695,N_14615,N_14853);
or UO_1696 (O_1696,N_14877,N_14994);
and UO_1697 (O_1697,N_14449,N_14816);
and UO_1698 (O_1698,N_14301,N_14872);
nor UO_1699 (O_1699,N_14739,N_14473);
xor UO_1700 (O_1700,N_14853,N_14583);
or UO_1701 (O_1701,N_14465,N_14488);
nand UO_1702 (O_1702,N_14675,N_14409);
nor UO_1703 (O_1703,N_14663,N_14597);
nand UO_1704 (O_1704,N_14386,N_14262);
nand UO_1705 (O_1705,N_14370,N_14666);
and UO_1706 (O_1706,N_14649,N_14262);
nand UO_1707 (O_1707,N_14895,N_14902);
or UO_1708 (O_1708,N_14419,N_14961);
nand UO_1709 (O_1709,N_14911,N_14594);
xnor UO_1710 (O_1710,N_14554,N_14632);
or UO_1711 (O_1711,N_14927,N_14587);
xnor UO_1712 (O_1712,N_14572,N_14849);
or UO_1713 (O_1713,N_14559,N_14945);
and UO_1714 (O_1714,N_14704,N_14734);
nor UO_1715 (O_1715,N_14401,N_14316);
or UO_1716 (O_1716,N_14445,N_14802);
nor UO_1717 (O_1717,N_14296,N_14479);
nor UO_1718 (O_1718,N_14507,N_14504);
nand UO_1719 (O_1719,N_14514,N_14774);
and UO_1720 (O_1720,N_14392,N_14933);
nor UO_1721 (O_1721,N_14353,N_14446);
nand UO_1722 (O_1722,N_14705,N_14888);
and UO_1723 (O_1723,N_14913,N_14460);
nor UO_1724 (O_1724,N_14419,N_14772);
nand UO_1725 (O_1725,N_14901,N_14784);
nand UO_1726 (O_1726,N_14445,N_14434);
nand UO_1727 (O_1727,N_14712,N_14891);
nor UO_1728 (O_1728,N_14914,N_14562);
nand UO_1729 (O_1729,N_14691,N_14474);
xor UO_1730 (O_1730,N_14786,N_14497);
nand UO_1731 (O_1731,N_14262,N_14657);
nand UO_1732 (O_1732,N_14561,N_14507);
xnor UO_1733 (O_1733,N_14581,N_14718);
and UO_1734 (O_1734,N_14379,N_14965);
or UO_1735 (O_1735,N_14263,N_14310);
or UO_1736 (O_1736,N_14551,N_14368);
or UO_1737 (O_1737,N_14366,N_14668);
nand UO_1738 (O_1738,N_14882,N_14747);
nor UO_1739 (O_1739,N_14759,N_14764);
or UO_1740 (O_1740,N_14339,N_14591);
or UO_1741 (O_1741,N_14729,N_14864);
or UO_1742 (O_1742,N_14250,N_14429);
or UO_1743 (O_1743,N_14866,N_14296);
xor UO_1744 (O_1744,N_14634,N_14422);
and UO_1745 (O_1745,N_14392,N_14725);
and UO_1746 (O_1746,N_14404,N_14816);
or UO_1747 (O_1747,N_14641,N_14706);
nor UO_1748 (O_1748,N_14290,N_14412);
xor UO_1749 (O_1749,N_14583,N_14667);
and UO_1750 (O_1750,N_14467,N_14965);
nand UO_1751 (O_1751,N_14742,N_14731);
nor UO_1752 (O_1752,N_14857,N_14924);
nand UO_1753 (O_1753,N_14797,N_14522);
or UO_1754 (O_1754,N_14434,N_14744);
or UO_1755 (O_1755,N_14868,N_14698);
nor UO_1756 (O_1756,N_14973,N_14333);
nand UO_1757 (O_1757,N_14688,N_14507);
nand UO_1758 (O_1758,N_14741,N_14965);
and UO_1759 (O_1759,N_14537,N_14612);
nand UO_1760 (O_1760,N_14376,N_14894);
or UO_1761 (O_1761,N_14416,N_14748);
and UO_1762 (O_1762,N_14674,N_14569);
nor UO_1763 (O_1763,N_14755,N_14520);
and UO_1764 (O_1764,N_14489,N_14529);
nor UO_1765 (O_1765,N_14660,N_14986);
and UO_1766 (O_1766,N_14378,N_14852);
nor UO_1767 (O_1767,N_14947,N_14605);
or UO_1768 (O_1768,N_14359,N_14965);
nor UO_1769 (O_1769,N_14624,N_14288);
nor UO_1770 (O_1770,N_14896,N_14880);
or UO_1771 (O_1771,N_14976,N_14291);
nor UO_1772 (O_1772,N_14523,N_14996);
xnor UO_1773 (O_1773,N_14622,N_14945);
and UO_1774 (O_1774,N_14506,N_14386);
nor UO_1775 (O_1775,N_14981,N_14594);
nand UO_1776 (O_1776,N_14798,N_14408);
nand UO_1777 (O_1777,N_14713,N_14700);
nand UO_1778 (O_1778,N_14528,N_14681);
xnor UO_1779 (O_1779,N_14584,N_14345);
nand UO_1780 (O_1780,N_14719,N_14816);
nand UO_1781 (O_1781,N_14936,N_14727);
nor UO_1782 (O_1782,N_14900,N_14441);
nor UO_1783 (O_1783,N_14498,N_14972);
nor UO_1784 (O_1784,N_14431,N_14502);
and UO_1785 (O_1785,N_14694,N_14818);
and UO_1786 (O_1786,N_14666,N_14633);
nand UO_1787 (O_1787,N_14340,N_14826);
or UO_1788 (O_1788,N_14824,N_14353);
nor UO_1789 (O_1789,N_14693,N_14420);
or UO_1790 (O_1790,N_14540,N_14357);
xnor UO_1791 (O_1791,N_14332,N_14409);
nor UO_1792 (O_1792,N_14297,N_14626);
or UO_1793 (O_1793,N_14572,N_14758);
xor UO_1794 (O_1794,N_14900,N_14309);
xor UO_1795 (O_1795,N_14251,N_14408);
nor UO_1796 (O_1796,N_14952,N_14322);
and UO_1797 (O_1797,N_14542,N_14503);
nand UO_1798 (O_1798,N_14674,N_14288);
and UO_1799 (O_1799,N_14634,N_14716);
or UO_1800 (O_1800,N_14364,N_14727);
nand UO_1801 (O_1801,N_14428,N_14750);
nor UO_1802 (O_1802,N_14828,N_14430);
nor UO_1803 (O_1803,N_14987,N_14642);
nand UO_1804 (O_1804,N_14592,N_14746);
nand UO_1805 (O_1805,N_14530,N_14988);
nand UO_1806 (O_1806,N_14762,N_14381);
nand UO_1807 (O_1807,N_14856,N_14365);
xnor UO_1808 (O_1808,N_14647,N_14257);
xnor UO_1809 (O_1809,N_14723,N_14812);
nand UO_1810 (O_1810,N_14952,N_14456);
xnor UO_1811 (O_1811,N_14353,N_14890);
and UO_1812 (O_1812,N_14423,N_14886);
xor UO_1813 (O_1813,N_14857,N_14834);
nor UO_1814 (O_1814,N_14906,N_14353);
nor UO_1815 (O_1815,N_14598,N_14942);
and UO_1816 (O_1816,N_14783,N_14612);
nand UO_1817 (O_1817,N_14371,N_14689);
or UO_1818 (O_1818,N_14434,N_14995);
nor UO_1819 (O_1819,N_14916,N_14493);
or UO_1820 (O_1820,N_14696,N_14547);
and UO_1821 (O_1821,N_14472,N_14573);
and UO_1822 (O_1822,N_14881,N_14553);
and UO_1823 (O_1823,N_14704,N_14639);
and UO_1824 (O_1824,N_14457,N_14929);
nor UO_1825 (O_1825,N_14749,N_14931);
nor UO_1826 (O_1826,N_14382,N_14932);
nor UO_1827 (O_1827,N_14610,N_14799);
and UO_1828 (O_1828,N_14377,N_14574);
xnor UO_1829 (O_1829,N_14935,N_14783);
nand UO_1830 (O_1830,N_14872,N_14966);
and UO_1831 (O_1831,N_14504,N_14544);
or UO_1832 (O_1832,N_14389,N_14764);
nand UO_1833 (O_1833,N_14548,N_14813);
or UO_1834 (O_1834,N_14996,N_14418);
xnor UO_1835 (O_1835,N_14492,N_14274);
nor UO_1836 (O_1836,N_14323,N_14280);
and UO_1837 (O_1837,N_14886,N_14299);
xnor UO_1838 (O_1838,N_14444,N_14781);
nand UO_1839 (O_1839,N_14998,N_14396);
and UO_1840 (O_1840,N_14287,N_14721);
or UO_1841 (O_1841,N_14884,N_14987);
or UO_1842 (O_1842,N_14686,N_14322);
nor UO_1843 (O_1843,N_14871,N_14605);
or UO_1844 (O_1844,N_14890,N_14781);
nor UO_1845 (O_1845,N_14354,N_14632);
nor UO_1846 (O_1846,N_14622,N_14808);
nor UO_1847 (O_1847,N_14970,N_14623);
nand UO_1848 (O_1848,N_14880,N_14753);
nand UO_1849 (O_1849,N_14650,N_14793);
nand UO_1850 (O_1850,N_14472,N_14262);
nor UO_1851 (O_1851,N_14671,N_14752);
or UO_1852 (O_1852,N_14695,N_14669);
nand UO_1853 (O_1853,N_14331,N_14978);
and UO_1854 (O_1854,N_14825,N_14884);
or UO_1855 (O_1855,N_14552,N_14279);
or UO_1856 (O_1856,N_14798,N_14657);
or UO_1857 (O_1857,N_14417,N_14817);
nand UO_1858 (O_1858,N_14255,N_14840);
and UO_1859 (O_1859,N_14796,N_14697);
and UO_1860 (O_1860,N_14481,N_14490);
or UO_1861 (O_1861,N_14451,N_14264);
or UO_1862 (O_1862,N_14774,N_14919);
and UO_1863 (O_1863,N_14871,N_14297);
and UO_1864 (O_1864,N_14803,N_14855);
nor UO_1865 (O_1865,N_14703,N_14603);
nor UO_1866 (O_1866,N_14873,N_14863);
nand UO_1867 (O_1867,N_14621,N_14393);
xnor UO_1868 (O_1868,N_14535,N_14799);
nor UO_1869 (O_1869,N_14591,N_14433);
nand UO_1870 (O_1870,N_14489,N_14362);
or UO_1871 (O_1871,N_14753,N_14474);
nor UO_1872 (O_1872,N_14781,N_14337);
or UO_1873 (O_1873,N_14310,N_14977);
xnor UO_1874 (O_1874,N_14463,N_14717);
or UO_1875 (O_1875,N_14383,N_14770);
and UO_1876 (O_1876,N_14320,N_14437);
xor UO_1877 (O_1877,N_14574,N_14781);
nand UO_1878 (O_1878,N_14412,N_14952);
nand UO_1879 (O_1879,N_14314,N_14824);
nor UO_1880 (O_1880,N_14710,N_14309);
nand UO_1881 (O_1881,N_14667,N_14638);
or UO_1882 (O_1882,N_14372,N_14487);
or UO_1883 (O_1883,N_14253,N_14391);
nor UO_1884 (O_1884,N_14468,N_14637);
nand UO_1885 (O_1885,N_14788,N_14263);
nand UO_1886 (O_1886,N_14699,N_14296);
nand UO_1887 (O_1887,N_14339,N_14483);
and UO_1888 (O_1888,N_14302,N_14815);
nand UO_1889 (O_1889,N_14463,N_14877);
or UO_1890 (O_1890,N_14405,N_14511);
or UO_1891 (O_1891,N_14842,N_14789);
or UO_1892 (O_1892,N_14984,N_14516);
and UO_1893 (O_1893,N_14709,N_14895);
xnor UO_1894 (O_1894,N_14877,N_14566);
or UO_1895 (O_1895,N_14996,N_14654);
xnor UO_1896 (O_1896,N_14447,N_14788);
nand UO_1897 (O_1897,N_14453,N_14715);
nor UO_1898 (O_1898,N_14304,N_14390);
and UO_1899 (O_1899,N_14950,N_14415);
xor UO_1900 (O_1900,N_14894,N_14752);
nand UO_1901 (O_1901,N_14914,N_14649);
and UO_1902 (O_1902,N_14351,N_14475);
nor UO_1903 (O_1903,N_14358,N_14397);
nor UO_1904 (O_1904,N_14433,N_14431);
and UO_1905 (O_1905,N_14560,N_14832);
nor UO_1906 (O_1906,N_14617,N_14640);
and UO_1907 (O_1907,N_14716,N_14485);
xor UO_1908 (O_1908,N_14406,N_14896);
nand UO_1909 (O_1909,N_14919,N_14599);
and UO_1910 (O_1910,N_14268,N_14784);
xnor UO_1911 (O_1911,N_14310,N_14306);
or UO_1912 (O_1912,N_14379,N_14773);
and UO_1913 (O_1913,N_14669,N_14693);
and UO_1914 (O_1914,N_14373,N_14938);
and UO_1915 (O_1915,N_14833,N_14619);
and UO_1916 (O_1916,N_14333,N_14826);
xor UO_1917 (O_1917,N_14893,N_14733);
nor UO_1918 (O_1918,N_14405,N_14993);
nand UO_1919 (O_1919,N_14354,N_14577);
nor UO_1920 (O_1920,N_14744,N_14881);
and UO_1921 (O_1921,N_14837,N_14477);
and UO_1922 (O_1922,N_14903,N_14609);
nor UO_1923 (O_1923,N_14917,N_14887);
or UO_1924 (O_1924,N_14951,N_14781);
nand UO_1925 (O_1925,N_14628,N_14984);
and UO_1926 (O_1926,N_14554,N_14307);
and UO_1927 (O_1927,N_14748,N_14467);
or UO_1928 (O_1928,N_14424,N_14878);
nand UO_1929 (O_1929,N_14800,N_14600);
and UO_1930 (O_1930,N_14838,N_14818);
or UO_1931 (O_1931,N_14368,N_14627);
and UO_1932 (O_1932,N_14964,N_14728);
nand UO_1933 (O_1933,N_14251,N_14785);
nor UO_1934 (O_1934,N_14858,N_14542);
and UO_1935 (O_1935,N_14629,N_14361);
and UO_1936 (O_1936,N_14338,N_14404);
or UO_1937 (O_1937,N_14721,N_14467);
nor UO_1938 (O_1938,N_14399,N_14477);
xor UO_1939 (O_1939,N_14968,N_14926);
or UO_1940 (O_1940,N_14334,N_14730);
nand UO_1941 (O_1941,N_14802,N_14355);
and UO_1942 (O_1942,N_14344,N_14990);
nand UO_1943 (O_1943,N_14607,N_14283);
and UO_1944 (O_1944,N_14305,N_14503);
nor UO_1945 (O_1945,N_14939,N_14486);
nand UO_1946 (O_1946,N_14980,N_14649);
xnor UO_1947 (O_1947,N_14989,N_14618);
or UO_1948 (O_1948,N_14537,N_14815);
and UO_1949 (O_1949,N_14835,N_14391);
or UO_1950 (O_1950,N_14413,N_14893);
nor UO_1951 (O_1951,N_14362,N_14364);
nand UO_1952 (O_1952,N_14785,N_14830);
nor UO_1953 (O_1953,N_14421,N_14976);
nor UO_1954 (O_1954,N_14376,N_14664);
nor UO_1955 (O_1955,N_14892,N_14852);
or UO_1956 (O_1956,N_14271,N_14408);
nand UO_1957 (O_1957,N_14736,N_14451);
nand UO_1958 (O_1958,N_14715,N_14993);
xnor UO_1959 (O_1959,N_14932,N_14936);
or UO_1960 (O_1960,N_14629,N_14569);
xor UO_1961 (O_1961,N_14579,N_14505);
or UO_1962 (O_1962,N_14361,N_14823);
nor UO_1963 (O_1963,N_14261,N_14584);
xnor UO_1964 (O_1964,N_14820,N_14467);
and UO_1965 (O_1965,N_14524,N_14278);
or UO_1966 (O_1966,N_14493,N_14520);
or UO_1967 (O_1967,N_14896,N_14876);
or UO_1968 (O_1968,N_14577,N_14541);
or UO_1969 (O_1969,N_14369,N_14533);
xor UO_1970 (O_1970,N_14518,N_14617);
xor UO_1971 (O_1971,N_14661,N_14511);
or UO_1972 (O_1972,N_14264,N_14586);
nor UO_1973 (O_1973,N_14624,N_14477);
or UO_1974 (O_1974,N_14667,N_14322);
or UO_1975 (O_1975,N_14471,N_14528);
xnor UO_1976 (O_1976,N_14849,N_14600);
or UO_1977 (O_1977,N_14685,N_14433);
nor UO_1978 (O_1978,N_14437,N_14859);
and UO_1979 (O_1979,N_14392,N_14439);
nand UO_1980 (O_1980,N_14852,N_14669);
nand UO_1981 (O_1981,N_14991,N_14972);
or UO_1982 (O_1982,N_14275,N_14888);
and UO_1983 (O_1983,N_14418,N_14991);
and UO_1984 (O_1984,N_14564,N_14918);
or UO_1985 (O_1985,N_14918,N_14781);
xnor UO_1986 (O_1986,N_14620,N_14344);
xnor UO_1987 (O_1987,N_14274,N_14778);
or UO_1988 (O_1988,N_14557,N_14555);
xor UO_1989 (O_1989,N_14756,N_14891);
nor UO_1990 (O_1990,N_14344,N_14485);
or UO_1991 (O_1991,N_14695,N_14589);
or UO_1992 (O_1992,N_14560,N_14599);
and UO_1993 (O_1993,N_14313,N_14276);
and UO_1994 (O_1994,N_14721,N_14781);
nand UO_1995 (O_1995,N_14840,N_14380);
nand UO_1996 (O_1996,N_14980,N_14689);
nand UO_1997 (O_1997,N_14551,N_14910);
and UO_1998 (O_1998,N_14628,N_14515);
or UO_1999 (O_1999,N_14570,N_14940);
endmodule