module basic_2000_20000_2500_80_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
or U0 (N_0,In_1181,In_1328);
nand U1 (N_1,In_1427,In_1190);
nor U2 (N_2,In_176,In_140);
or U3 (N_3,In_640,In_1914);
and U4 (N_4,In_1234,In_1399);
or U5 (N_5,In_851,In_1436);
xor U6 (N_6,In_1468,In_1969);
xnor U7 (N_7,In_701,In_1292);
nand U8 (N_8,In_62,In_213);
nand U9 (N_9,In_122,In_1522);
nor U10 (N_10,In_563,In_1432);
nor U11 (N_11,In_881,In_123);
and U12 (N_12,In_4,In_1222);
xor U13 (N_13,In_326,In_35);
and U14 (N_14,In_809,In_1070);
xor U15 (N_15,In_1995,In_22);
or U16 (N_16,In_559,In_312);
xnor U17 (N_17,In_1951,In_1441);
and U18 (N_18,In_1780,In_1838);
xor U19 (N_19,In_1183,In_166);
and U20 (N_20,In_2,In_369);
nand U21 (N_21,In_1697,In_1085);
xnor U22 (N_22,In_641,In_1918);
nor U23 (N_23,In_30,In_889);
nor U24 (N_24,In_1044,In_1011);
nand U25 (N_25,In_1477,In_1023);
xnor U26 (N_26,In_841,In_1345);
nor U27 (N_27,In_1628,In_1892);
xnor U28 (N_28,In_1739,In_224);
nand U29 (N_29,In_441,In_1776);
xnor U30 (N_30,In_1930,In_1316);
xor U31 (N_31,In_1157,In_277);
nor U32 (N_32,In_483,In_537);
nor U33 (N_33,In_446,In_1859);
xnor U34 (N_34,In_985,In_828);
nand U35 (N_35,In_207,In_34);
nand U36 (N_36,In_959,In_1241);
nand U37 (N_37,In_527,In_1252);
or U38 (N_38,In_908,In_1402);
nor U39 (N_39,In_1687,In_1799);
xnor U40 (N_40,In_1971,In_1643);
xnor U41 (N_41,In_87,In_576);
nor U42 (N_42,In_262,In_17);
xnor U43 (N_43,In_545,In_1945);
nor U44 (N_44,In_1510,In_1073);
xnor U45 (N_45,In_114,In_1996);
and U46 (N_46,In_967,In_625);
xor U47 (N_47,In_515,In_992);
and U48 (N_48,In_300,In_1863);
nand U49 (N_49,In_1661,In_109);
or U50 (N_50,In_448,In_907);
nand U51 (N_51,In_1396,In_105);
xnor U52 (N_52,In_665,In_84);
nand U53 (N_53,In_1123,In_1528);
nor U54 (N_54,In_204,In_539);
nor U55 (N_55,In_136,In_654);
and U56 (N_56,In_29,In_1054);
nand U57 (N_57,In_177,In_479);
or U58 (N_58,In_1832,In_1211);
nand U59 (N_59,In_264,In_1612);
nand U60 (N_60,In_139,In_577);
nor U61 (N_61,In_906,In_1437);
and U62 (N_62,In_1805,In_1609);
or U63 (N_63,In_1074,In_580);
and U64 (N_64,In_1923,In_647);
nand U65 (N_65,In_1052,In_533);
xor U66 (N_66,In_1125,In_606);
nor U67 (N_67,In_488,In_41);
nor U68 (N_68,In_1706,In_1281);
nor U69 (N_69,In_20,In_1658);
and U70 (N_70,In_952,In_1659);
nor U71 (N_71,In_1231,In_1501);
and U72 (N_72,In_116,In_1826);
nor U73 (N_73,In_411,In_940);
or U74 (N_74,In_484,In_591);
nor U75 (N_75,In_486,In_1188);
xor U76 (N_76,In_879,In_1931);
nor U77 (N_77,In_1048,In_1243);
nor U78 (N_78,In_356,In_953);
or U79 (N_79,In_248,In_226);
xnor U80 (N_80,In_1772,In_377);
or U81 (N_81,In_1937,In_816);
nor U82 (N_82,In_806,In_1414);
xnor U83 (N_83,In_1541,In_1709);
xnor U84 (N_84,In_541,In_694);
xor U85 (N_85,In_1299,In_1305);
nand U86 (N_86,In_1673,In_1089);
or U87 (N_87,In_1868,In_592);
xor U88 (N_88,In_666,In_547);
nor U89 (N_89,In_1081,In_958);
and U90 (N_90,In_1443,In_1888);
and U91 (N_91,In_535,In_1848);
or U92 (N_92,In_1444,In_1354);
xnor U93 (N_93,In_214,In_1397);
nand U94 (N_94,In_810,In_1341);
and U95 (N_95,In_987,In_1289);
and U96 (N_96,In_1994,In_876);
and U97 (N_97,In_1297,In_1733);
or U98 (N_98,In_1745,In_266);
nand U99 (N_99,In_936,In_511);
and U100 (N_100,In_236,In_1530);
and U101 (N_101,In_626,In_646);
nor U102 (N_102,In_10,In_1988);
nor U103 (N_103,In_587,In_1302);
and U104 (N_104,In_1214,In_1748);
nand U105 (N_105,In_1581,In_1910);
and U106 (N_106,In_1318,In_1600);
or U107 (N_107,In_517,In_822);
nand U108 (N_108,In_1703,In_423);
and U109 (N_109,In_943,In_1949);
xnor U110 (N_110,In_1864,In_241);
xnor U111 (N_111,In_1693,In_730);
or U112 (N_112,In_860,In_1880);
nand U113 (N_113,In_1166,In_426);
nor U114 (N_114,In_1415,In_279);
nor U115 (N_115,In_1456,In_1069);
nor U116 (N_116,In_400,In_282);
xnor U117 (N_117,In_83,In_930);
nor U118 (N_118,In_949,In_1891);
or U119 (N_119,In_614,In_1976);
xnor U120 (N_120,In_235,In_1831);
xor U121 (N_121,In_1948,In_74);
nand U122 (N_122,In_561,In_1090);
xnor U123 (N_123,In_1487,In_1425);
xor U124 (N_124,In_1632,In_751);
nor U125 (N_125,In_1224,In_181);
nor U126 (N_126,In_1010,In_1226);
and U127 (N_127,In_1064,In_1783);
nand U128 (N_128,In_399,In_1171);
nand U129 (N_129,In_501,In_970);
and U130 (N_130,In_685,In_320);
nor U131 (N_131,In_629,In_1865);
and U132 (N_132,In_595,In_314);
xnor U133 (N_133,In_897,In_565);
and U134 (N_134,In_47,In_842);
or U135 (N_135,In_1290,In_1607);
and U136 (N_136,In_219,In_1428);
or U137 (N_137,In_875,In_1883);
and U138 (N_138,In_1239,In_1959);
and U139 (N_139,In_1684,In_663);
and U140 (N_140,In_298,In_482);
or U141 (N_141,In_1964,In_289);
nand U142 (N_142,In_280,In_982);
or U143 (N_143,In_420,In_601);
nand U144 (N_144,In_508,In_604);
nand U145 (N_145,In_1887,In_1326);
xor U146 (N_146,In_459,In_364);
or U147 (N_147,In_336,In_1881);
or U148 (N_148,In_1018,In_1668);
or U149 (N_149,In_1087,In_684);
and U150 (N_150,In_630,In_243);
or U151 (N_151,In_832,In_821);
xor U152 (N_152,In_650,In_574);
and U153 (N_153,In_1932,In_1724);
or U154 (N_154,In_410,In_294);
or U155 (N_155,In_1198,In_1380);
or U156 (N_156,In_588,In_935);
nor U157 (N_157,In_1478,In_1989);
nor U158 (N_158,In_1814,In_598);
xor U159 (N_159,In_272,In_612);
and U160 (N_160,In_1068,In_1273);
nand U161 (N_161,In_119,In_994);
xor U162 (N_162,In_1306,In_1774);
nor U163 (N_163,In_1275,In_996);
nor U164 (N_164,In_424,In_709);
xor U165 (N_165,In_1473,In_1722);
xnor U166 (N_166,In_1347,In_600);
xnor U167 (N_167,In_569,In_1731);
or U168 (N_168,In_920,In_1531);
nor U169 (N_169,In_1463,In_164);
or U170 (N_170,In_1119,In_1498);
and U171 (N_171,In_1103,In_1768);
nor U172 (N_172,In_1764,In_1093);
and U173 (N_173,In_503,In_1182);
nand U174 (N_174,In_1288,In_1469);
nand U175 (N_175,In_288,In_1943);
xnor U176 (N_176,In_877,In_233);
nor U177 (N_177,In_444,In_807);
nand U178 (N_178,In_58,In_931);
and U179 (N_179,In_379,In_398);
xor U180 (N_180,In_1411,In_1741);
and U181 (N_181,In_1797,In_1997);
or U182 (N_182,In_1650,In_1586);
nor U183 (N_183,In_127,In_1867);
nor U184 (N_184,In_1955,In_658);
nand U185 (N_185,In_428,In_1927);
or U186 (N_186,In_975,In_826);
nand U187 (N_187,In_1192,In_1383);
xor U188 (N_188,In_137,In_1219);
or U189 (N_189,In_1815,In_361);
or U190 (N_190,In_1778,In_1409);
or U191 (N_191,In_597,In_1792);
or U192 (N_192,In_729,In_1453);
or U193 (N_193,In_1454,In_1141);
nand U194 (N_194,In_230,In_1912);
nor U195 (N_195,In_1753,In_1938);
nand U196 (N_196,In_1153,In_1533);
xor U197 (N_197,In_1941,In_357);
and U198 (N_198,In_1365,In_1816);
xor U199 (N_199,In_125,In_90);
xnor U200 (N_200,In_205,In_1156);
or U201 (N_201,In_330,In_1075);
and U202 (N_202,In_461,In_304);
nand U203 (N_203,In_1083,In_218);
xnor U204 (N_204,In_146,In_1806);
or U205 (N_205,In_1963,In_852);
nand U206 (N_206,In_1175,In_195);
xnor U207 (N_207,In_567,In_1337);
nand U208 (N_208,In_1670,In_1237);
nand U209 (N_209,In_1849,In_1269);
nand U210 (N_210,In_1015,In_1738);
xor U211 (N_211,In_391,In_1209);
xnor U212 (N_212,In_747,In_212);
nor U213 (N_213,In_182,In_396);
nand U214 (N_214,In_240,In_848);
nor U215 (N_215,In_1492,In_187);
nand U216 (N_216,In_1665,In_1150);
nand U217 (N_217,In_1187,In_458);
nor U218 (N_218,In_1812,In_494);
nor U219 (N_219,In_79,In_1755);
xnor U220 (N_220,In_1588,In_1489);
xnor U221 (N_221,In_937,In_815);
and U222 (N_222,In_750,In_939);
and U223 (N_223,In_575,In_1803);
and U224 (N_224,In_1475,In_1174);
xor U225 (N_225,In_1331,In_1715);
nand U226 (N_226,In_825,In_161);
nor U227 (N_227,In_1082,In_220);
nor U228 (N_228,In_291,In_1610);
nand U229 (N_229,In_1245,In_394);
xor U230 (N_230,In_1563,In_499);
and U231 (N_231,In_1340,In_788);
nor U232 (N_232,In_1556,In_476);
and U233 (N_233,In_775,In_1162);
nor U234 (N_234,In_1935,In_1524);
and U235 (N_235,In_259,In_664);
nand U236 (N_236,In_1363,In_1704);
xor U237 (N_237,In_104,In_234);
or U238 (N_238,In_733,In_111);
or U239 (N_239,In_28,In_523);
and U240 (N_240,In_753,In_301);
nand U241 (N_241,In_1749,In_573);
nor U242 (N_242,In_1681,In_305);
and U243 (N_243,In_892,In_1029);
nor U244 (N_244,In_1388,In_589);
and U245 (N_245,In_831,In_1372);
nor U246 (N_246,In_1841,In_1719);
nor U247 (N_247,In_429,In_1105);
nand U248 (N_248,In_1202,In_1993);
or U249 (N_249,In_874,In_1450);
nor U250 (N_250,In_667,N_89);
xnor U251 (N_251,N_150,In_638);
nand U252 (N_252,N_97,In_1484);
and U253 (N_253,In_926,In_71);
and U254 (N_254,In_1227,In_1303);
and U255 (N_255,In_752,In_705);
xnor U256 (N_256,In_1329,N_7);
xnor U257 (N_257,In_159,In_1424);
xnor U258 (N_258,N_100,In_1718);
xor U259 (N_259,N_49,In_1369);
xor U260 (N_260,In_1207,In_1856);
nand U261 (N_261,In_1506,In_1889);
nand U262 (N_262,N_87,In_1895);
and U263 (N_263,In_829,In_1493);
nand U264 (N_264,In_670,In_1904);
nor U265 (N_265,In_1500,In_986);
and U266 (N_266,In_925,N_24);
and U267 (N_267,N_223,In_325);
and U268 (N_268,In_1901,In_1);
or U269 (N_269,In_554,In_1407);
nor U270 (N_270,In_1417,In_38);
nand U271 (N_271,In_1961,In_1598);
and U272 (N_272,In_450,N_101);
or U273 (N_273,In_678,N_1);
nand U274 (N_274,In_862,In_55);
nand U275 (N_275,In_655,In_657);
nor U276 (N_276,In_171,In_1221);
and U277 (N_277,In_1319,In_169);
and U278 (N_278,In_491,In_308);
nor U279 (N_279,In_1132,In_342);
nand U280 (N_280,In_1977,In_106);
nand U281 (N_281,In_676,In_1565);
and U282 (N_282,In_228,In_1591);
and U283 (N_283,In_703,In_1053);
xnor U284 (N_284,N_169,In_1445);
and U285 (N_285,N_75,In_1108);
or U286 (N_286,In_1246,In_550);
and U287 (N_287,In_386,In_1128);
nand U288 (N_288,In_472,N_17);
xnor U289 (N_289,In_1678,In_487);
or U290 (N_290,In_1235,In_497);
and U291 (N_291,In_1804,In_1827);
nand U292 (N_292,N_76,In_1611);
xnor U293 (N_293,In_769,In_130);
nor U294 (N_294,In_1909,In_1457);
nor U295 (N_295,In_1946,In_1672);
and U296 (N_296,In_473,In_43);
nor U297 (N_297,In_1744,N_25);
nor U298 (N_298,In_888,N_72);
nand U299 (N_299,In_365,In_1301);
nor U300 (N_300,N_200,In_372);
nand U301 (N_301,In_1801,In_1197);
nor U302 (N_302,In_1377,In_1031);
or U303 (N_303,N_194,In_419);
or U304 (N_304,N_140,In_403);
and U305 (N_305,N_98,In_1555);
or U306 (N_306,In_37,N_171);
nand U307 (N_307,In_1462,N_113);
xnor U308 (N_308,In_1356,In_433);
and U309 (N_309,In_1152,In_1640);
xnor U310 (N_310,In_782,N_96);
xor U311 (N_311,In_303,In_1765);
and U312 (N_312,In_1422,In_1595);
or U313 (N_313,In_1271,In_93);
xnor U314 (N_314,In_1798,In_285);
nor U315 (N_315,N_173,N_27);
and U316 (N_316,N_67,In_1099);
nand U317 (N_317,In_1113,In_39);
and U318 (N_318,In_1335,In_763);
or U319 (N_319,In_1076,In_206);
nand U320 (N_320,In_1819,In_991);
and U321 (N_321,N_59,In_7);
xor U322 (N_322,In_244,In_1763);
nand U323 (N_323,In_1716,In_1720);
nor U324 (N_324,In_706,In_526);
nor U325 (N_325,In_295,In_1470);
and U326 (N_326,In_1272,N_30);
nand U327 (N_327,In_1728,In_1244);
or U328 (N_328,In_33,In_154);
nor U329 (N_329,In_1975,In_77);
and U330 (N_330,In_932,In_855);
xor U331 (N_331,In_1788,N_71);
nor U332 (N_332,In_864,In_964);
or U333 (N_333,N_230,In_452);
nor U334 (N_334,In_1857,In_1613);
nor U335 (N_335,In_898,In_1999);
nor U336 (N_336,In_1035,In_562);
nand U337 (N_337,In_468,In_1606);
or U338 (N_338,In_1717,In_1557);
and U339 (N_339,In_211,In_190);
nor U340 (N_340,In_1285,In_1526);
nor U341 (N_341,In_387,N_221);
nor U342 (N_342,N_26,In_1265);
and U343 (N_343,In_1519,In_714);
or U344 (N_344,In_1523,N_203);
or U345 (N_345,In_168,In_615);
or U346 (N_346,In_1042,In_680);
or U347 (N_347,In_1855,In_145);
nand U348 (N_348,N_185,In_1796);
or U349 (N_349,In_737,In_1117);
and U350 (N_350,In_1001,N_117);
nand U351 (N_351,In_422,In_675);
nand U352 (N_352,In_1810,In_1040);
nand U353 (N_353,In_1928,In_1858);
nand U354 (N_354,In_1727,In_1137);
xor U355 (N_355,In_689,In_1459);
or U356 (N_356,In_1631,In_1710);
and U357 (N_357,In_1974,In_1903);
and U358 (N_358,In_1133,N_186);
xor U359 (N_359,In_375,In_14);
and U360 (N_360,In_1616,In_1582);
or U361 (N_361,In_1594,In_500);
xnor U362 (N_362,In_1438,N_23);
nand U363 (N_363,In_794,In_972);
xnor U364 (N_364,In_229,In_984);
nor U365 (N_365,In_25,In_777);
nand U366 (N_366,In_734,N_79);
or U367 (N_367,In_103,In_844);
xor U368 (N_368,In_370,N_205);
nor U369 (N_369,In_337,In_1622);
nor U370 (N_370,In_1630,In_1638);
xnor U371 (N_371,In_120,In_89);
or U372 (N_372,In_275,In_699);
xor U373 (N_373,In_656,N_199);
nand U374 (N_374,In_1164,In_1713);
nand U375 (N_375,In_412,In_1078);
nor U376 (N_376,In_1100,In_1829);
xor U377 (N_377,In_1551,In_890);
and U378 (N_378,In_758,In_414);
or U379 (N_379,In_1061,In_1268);
xor U380 (N_380,In_922,In_1474);
nand U381 (N_381,In_948,In_1879);
nor U382 (N_382,N_19,N_122);
xnor U383 (N_383,In_586,In_1732);
nor U384 (N_384,In_1690,In_843);
nand U385 (N_385,In_1714,In_1548);
nand U386 (N_386,In_596,N_73);
nor U387 (N_387,In_965,In_389);
or U388 (N_388,N_246,N_170);
and U389 (N_389,In_69,In_1442);
nand U390 (N_390,In_724,In_552);
nor U391 (N_391,In_968,In_1247);
and U392 (N_392,In_409,In_695);
xor U393 (N_393,In_447,In_118);
and U394 (N_394,In_955,N_175);
or U395 (N_395,In_1106,In_1505);
and U396 (N_396,In_31,In_1692);
nor U397 (N_397,In_1159,In_327);
xnor U398 (N_398,N_161,N_92);
or U399 (N_399,In_969,In_1593);
nand U400 (N_400,In_915,In_1096);
or U401 (N_401,In_1917,In_1726);
nand U402 (N_402,N_245,N_183);
and U403 (N_403,In_649,In_196);
nand U404 (N_404,In_346,N_147);
or U405 (N_405,In_1036,In_349);
or U406 (N_406,In_49,In_530);
and U407 (N_407,In_184,N_120);
nor U408 (N_408,N_154,In_1038);
nor U409 (N_409,In_309,In_1885);
or U410 (N_410,In_1811,N_136);
or U411 (N_411,In_609,In_313);
nand U412 (N_412,N_177,In_302);
nor U413 (N_413,In_899,In_590);
nor U414 (N_414,In_1368,In_1680);
nand U415 (N_415,In_1566,N_115);
xor U416 (N_416,In_1458,In_253);
xnor U417 (N_417,In_923,In_696);
or U418 (N_418,In_1315,In_1908);
nand U419 (N_419,In_1338,In_1781);
or U420 (N_420,In_221,In_540);
nor U421 (N_421,N_209,In_1585);
and U422 (N_422,In_463,In_1967);
and U423 (N_423,In_12,In_1509);
or U424 (N_424,In_407,In_1947);
nor U425 (N_425,In_549,In_808);
xnor U426 (N_426,N_60,In_239);
nor U427 (N_427,In_421,In_1966);
nor U428 (N_428,In_252,In_1907);
nor U429 (N_429,In_504,In_110);
nor U430 (N_430,In_373,In_813);
nand U431 (N_431,In_467,N_104);
or U432 (N_432,In_1835,In_1663);
nor U433 (N_433,In_1006,In_840);
and U434 (N_434,In_1154,In_188);
nand U435 (N_435,In_679,In_1367);
nand U436 (N_436,In_838,In_1546);
xor U437 (N_437,N_228,N_93);
nand U438 (N_438,In_659,N_208);
nand U439 (N_439,In_1513,In_1545);
or U440 (N_440,In_887,In_293);
nor U441 (N_441,In_1490,In_1873);
and U442 (N_442,In_793,In_1712);
or U443 (N_443,In_1634,In_1615);
or U444 (N_444,In_231,In_61);
or U445 (N_445,In_1228,In_382);
xnor U446 (N_446,In_1334,In_999);
or U447 (N_447,N_240,In_1481);
nor U448 (N_448,In_861,In_9);
nand U449 (N_449,In_623,In_919);
xnor U450 (N_450,In_976,In_1900);
or U451 (N_451,In_1648,In_725);
or U452 (N_452,In_1558,In_323);
and U453 (N_453,In_1840,In_644);
or U454 (N_454,In_871,In_1919);
nor U455 (N_455,In_1695,In_1629);
or U456 (N_456,In_1161,In_1701);
xnor U457 (N_457,In_1702,In_780);
or U458 (N_458,In_1518,In_944);
and U459 (N_459,In_1387,In_1116);
and U460 (N_460,In_661,In_1461);
nand U461 (N_461,In_778,In_1139);
nand U462 (N_462,In_642,In_157);
or U463 (N_463,N_61,In_1349);
xor U464 (N_464,In_738,In_946);
xnor U465 (N_465,In_1250,In_121);
nor U466 (N_466,In_581,In_1525);
nor U467 (N_467,In_1110,In_1094);
and U468 (N_468,In_1740,In_671);
nand U469 (N_469,In_619,In_1539);
nand U470 (N_470,In_390,In_988);
xnor U471 (N_471,In_1953,N_70);
nor U472 (N_472,In_222,In_1486);
or U473 (N_473,In_1020,In_416);
nor U474 (N_474,In_132,N_46);
or U475 (N_475,N_16,In_1062);
nand U476 (N_476,In_924,In_558);
or U477 (N_477,In_917,In_223);
and U478 (N_478,In_1711,In_1636);
nor U479 (N_479,In_1080,In_934);
xor U480 (N_480,In_1130,In_1842);
xor U481 (N_481,In_1066,In_910);
xnor U482 (N_482,In_1304,In_792);
nor U483 (N_483,N_167,In_24);
and U484 (N_484,In_1603,In_1412);
nor U485 (N_485,In_594,In_754);
nand U486 (N_486,In_878,In_1200);
or U487 (N_487,In_1575,In_1851);
nand U488 (N_488,In_1433,In_711);
nand U489 (N_489,In_173,N_187);
or U490 (N_490,In_1656,In_1124);
and U491 (N_491,In_128,In_1837);
and U492 (N_492,In_52,N_34);
xor U493 (N_493,In_131,In_687);
nand U494 (N_494,In_1088,N_234);
xnor U495 (N_495,In_1114,N_4);
nand U496 (N_496,In_1641,In_1645);
or U497 (N_497,In_516,In_542);
xnor U498 (N_498,In_1270,N_247);
xnor U499 (N_499,In_290,In_1286);
nand U500 (N_500,N_382,In_1413);
nor U501 (N_501,In_1398,In_715);
or U502 (N_502,In_404,N_265);
nor U503 (N_503,N_164,In_392);
nand U504 (N_504,In_260,In_700);
and U505 (N_505,In_271,N_188);
and U506 (N_506,In_141,In_1800);
nand U507 (N_507,In_1675,In_359);
or U508 (N_508,In_1896,In_113);
nand U509 (N_509,In_812,N_403);
nand U510 (N_510,In_954,In_1862);
nor U511 (N_511,N_308,In_1408);
nor U512 (N_512,In_97,N_168);
and U513 (N_513,In_1626,In_669);
nand U514 (N_514,In_702,In_464);
nand U515 (N_515,In_585,N_459);
and U516 (N_516,In_1520,In_1921);
nor U517 (N_517,In_92,In_698);
and U518 (N_518,In_1158,In_26);
xor U519 (N_519,N_324,In_1760);
nor U520 (N_520,In_951,In_1003);
or U521 (N_521,N_358,In_1330);
nor U522 (N_522,In_859,In_1274);
nand U523 (N_523,N_493,In_1429);
and U524 (N_524,In_1240,In_460);
nand U525 (N_525,In_50,In_1540);
nand U526 (N_526,In_1179,In_849);
or U527 (N_527,In_534,In_158);
or U528 (N_528,N_5,In_723);
nor U529 (N_529,In_1134,In_1446);
nand U530 (N_530,In_142,N_157);
or U531 (N_531,In_1385,In_1729);
and U532 (N_532,In_432,In_1723);
nand U533 (N_533,In_1986,N_350);
or U534 (N_534,In_1499,In_347);
xnor U535 (N_535,N_290,In_322);
nand U536 (N_536,In_345,In_1204);
nand U537 (N_537,In_453,In_1314);
and U538 (N_538,In_85,In_1278);
nor U539 (N_539,In_566,In_617);
nand U540 (N_540,In_1578,N_450);
nor U541 (N_541,N_178,N_10);
or U542 (N_542,In_1619,In_185);
xnor U543 (N_543,In_1795,N_483);
nor U544 (N_544,In_1580,N_449);
and U545 (N_545,In_1120,In_413);
nand U546 (N_546,In_1115,In_602);
nand U547 (N_547,In_1255,N_475);
or U548 (N_548,In_900,N_22);
nor U549 (N_549,N_231,N_269);
nand U550 (N_550,In_681,In_583);
and U551 (N_551,In_853,In_98);
xnor U552 (N_552,In_1028,In_1039);
and U553 (N_553,In_1483,In_1950);
and U554 (N_554,N_64,N_415);
or U555 (N_555,In_1550,In_1893);
or U556 (N_556,In_637,N_179);
xnor U557 (N_557,N_68,In_381);
nand U558 (N_558,N_333,N_166);
or U559 (N_559,N_86,In_66);
xnor U560 (N_560,In_977,In_1098);
xor U561 (N_561,N_82,In_242);
nor U562 (N_562,In_306,In_805);
nor U563 (N_563,N_210,N_201);
xnor U564 (N_564,In_1000,In_902);
nor U565 (N_565,N_444,In_1544);
or U566 (N_566,In_492,In_1138);
nor U567 (N_567,In_1021,In_1448);
and U568 (N_568,In_618,In_36);
or U569 (N_569,In_1389,In_1283);
and U570 (N_570,N_116,In_393);
or U571 (N_571,In_1455,In_757);
or U572 (N_572,In_430,In_846);
and U573 (N_573,N_347,N_259);
nand U574 (N_574,N_91,In_1980);
nand U575 (N_575,In_135,In_112);
and U576 (N_576,N_476,N_396);
or U577 (N_577,In_1353,In_54);
and U578 (N_578,In_1761,In_1346);
nor U579 (N_579,In_245,In_578);
nor U580 (N_580,In_1177,In_65);
nor U581 (N_581,In_1562,In_803);
or U582 (N_582,N_470,N_202);
nand U583 (N_583,N_296,In_525);
nand U584 (N_584,In_983,In_1199);
and U585 (N_585,In_1850,In_1180);
nand U586 (N_586,N_405,In_1608);
nor U587 (N_587,N_62,In_456);
nor U588 (N_588,N_233,N_42);
xor U589 (N_589,In_628,N_311);
nand U590 (N_590,In_1844,In_1843);
nand U591 (N_591,N_217,In_343);
or U592 (N_592,In_599,In_682);
xnor U593 (N_593,In_1789,In_1253);
nor U594 (N_594,N_235,In_1982);
and U595 (N_595,N_408,In_1624);
nor U596 (N_596,In_1260,In_1261);
or U597 (N_597,N_56,In_555);
nand U598 (N_598,In_1808,In_514);
and U599 (N_599,N_477,In_1236);
and U600 (N_600,In_199,In_1254);
or U601 (N_601,In_817,N_184);
and U602 (N_602,In_1193,In_1825);
or U603 (N_603,In_44,In_1480);
nor U604 (N_604,In_529,In_443);
nor U605 (N_605,In_1688,In_1047);
nor U606 (N_606,N_487,In_1060);
and U607 (N_607,N_94,In_183);
nor U608 (N_608,N_386,N_9);
and U609 (N_609,In_1915,In_1495);
nand U610 (N_610,In_1537,In_799);
and U611 (N_611,In_469,In_1277);
and U612 (N_612,N_239,In_863);
nor U613 (N_613,In_281,In_720);
or U614 (N_614,N_343,In_107);
nand U615 (N_615,In_1307,N_272);
or U616 (N_616,N_289,In_1225);
xor U617 (N_617,N_260,In_1058);
xnor U618 (N_618,In_854,In_269);
xor U619 (N_619,In_502,N_83);
nand U620 (N_620,In_507,In_1421);
or U621 (N_621,In_1958,In_1342);
nor U622 (N_622,N_425,In_759);
and U623 (N_623,In_358,N_127);
or U624 (N_624,In_770,In_1597);
xor U625 (N_625,In_124,In_367);
or U626 (N_626,In_1091,In_560);
nand U627 (N_627,In_1992,In_1633);
and U628 (N_628,In_328,In_1109);
nand U629 (N_629,In_1497,In_1882);
xnor U630 (N_630,In_1033,In_755);
or U631 (N_631,In_771,In_1705);
or U632 (N_632,In_1736,In_1449);
nor U633 (N_633,In_1086,In_1752);
nand U634 (N_634,In_743,In_727);
and U635 (N_635,In_40,In_798);
or U636 (N_636,In_1467,N_119);
nand U637 (N_637,In_1163,In_99);
nand U638 (N_638,N_244,N_372);
nand U639 (N_639,In_11,In_731);
or U640 (N_640,N_463,In_350);
nor U641 (N_641,In_374,In_397);
or U642 (N_642,N_410,In_1037);
nand U643 (N_643,In_1771,In_1642);
and U644 (N_644,In_1496,N_378);
nor U645 (N_645,In_1942,In_395);
nor U646 (N_646,N_251,In_307);
and U647 (N_647,In_1024,N_268);
nand U648 (N_648,In_1878,In_1854);
nor U649 (N_649,In_1674,In_1592);
or U650 (N_650,N_394,N_374);
nor U651 (N_651,In_1514,N_197);
nand U652 (N_652,In_1379,N_313);
nor U653 (N_653,In_1699,In_608);
xor U654 (N_654,In_833,In_1220);
or U655 (N_655,In_748,N_423);
and U656 (N_656,N_258,N_469);
nor U657 (N_657,In_1751,N_387);
xnor U658 (N_658,In_884,In_613);
nor U659 (N_659,In_1185,In_1196);
nand U660 (N_660,In_495,In_1263);
and U661 (N_661,N_142,N_190);
or U662 (N_662,N_432,In_1416);
xnor U663 (N_663,N_139,N_14);
xor U664 (N_664,In_1897,In_1534);
or U665 (N_665,In_1362,In_1184);
nor U666 (N_666,In_512,In_633);
and U667 (N_667,In_425,In_1311);
or U668 (N_668,In_1071,In_1287);
nor U669 (N_669,In_1998,N_312);
nor U670 (N_670,N_165,In_1371);
and U671 (N_671,In_787,In_317);
and U672 (N_672,N_490,In_1742);
nand U673 (N_673,N_327,N_440);
nor U674 (N_674,In_1981,In_797);
nand U675 (N_675,N_414,N_198);
nand U676 (N_676,In_150,N_401);
nand U677 (N_677,In_1933,In_1005);
and U678 (N_678,In_1194,N_306);
nor U679 (N_679,In_60,In_498);
nor U680 (N_680,N_428,In_1233);
and U681 (N_681,In_1605,N_192);
or U682 (N_682,In_1279,In_1063);
or U683 (N_683,N_456,In_796);
xnor U684 (N_684,In_96,In_1599);
and U685 (N_685,In_1572,N_32);
xnor U686 (N_686,In_255,In_1793);
nor U687 (N_687,In_1813,In_741);
xnor U688 (N_688,In_1502,In_1291);
and U689 (N_689,In_478,In_0);
nor U690 (N_690,N_320,In_903);
nor U691 (N_691,In_1172,N_294);
nand U692 (N_692,In_1725,N_57);
nand U693 (N_693,N_281,In_1122);
or U694 (N_694,In_639,N_220);
and U695 (N_695,In_1833,In_819);
nor U696 (N_696,N_137,In_1321);
and U697 (N_697,In_1155,In_557);
xnor U698 (N_698,N_309,In_1325);
and U699 (N_699,In_1390,In_942);
or U700 (N_700,In_1635,In_1911);
nor U701 (N_701,In_276,In_1775);
or U702 (N_702,N_158,In_1568);
and U703 (N_703,In_1902,In_76);
nor U704 (N_704,N_419,In_1627);
xnor U705 (N_705,In_1617,In_621);
xnor U706 (N_706,In_1391,In_732);
xor U707 (N_707,In_745,In_1017);
nand U708 (N_708,N_130,In_1750);
nor U709 (N_709,N_341,N_286);
nand U710 (N_710,N_325,N_176);
and U711 (N_711,In_1860,In_193);
nand U712 (N_712,In_1936,N_400);
xor U713 (N_713,In_1926,In_1639);
nand U714 (N_714,In_1403,In_1121);
nor U715 (N_715,N_123,In_1393);
xnor U716 (N_716,N_431,In_1560);
nand U717 (N_717,In_102,In_749);
nand U718 (N_718,N_445,N_181);
nand U719 (N_719,In_1151,N_399);
xnor U720 (N_720,N_85,In_88);
xnor U721 (N_721,In_1689,N_15);
or U722 (N_722,In_402,In_1587);
or U723 (N_723,In_692,In_1823);
xor U724 (N_724,In_1223,In_1886);
nor U725 (N_725,In_956,N_488);
nand U726 (N_726,N_2,N_131);
nor U727 (N_727,In_126,N_58);
nor U728 (N_728,In_45,In_1960);
and U729 (N_729,N_41,In_1386);
nand U730 (N_730,N_424,N_413);
and U731 (N_731,In_1691,N_340);
or U732 (N_732,N_393,N_395);
nor U733 (N_733,In_1485,In_1264);
or U734 (N_734,In_274,N_134);
or U735 (N_735,In_278,In_824);
xor U736 (N_736,N_375,In_1262);
xor U737 (N_737,N_214,In_163);
and U738 (N_738,In_1786,N_237);
nand U739 (N_739,In_352,N_391);
or U740 (N_740,N_216,In_1746);
nor U741 (N_741,In_481,In_215);
nand U742 (N_742,In_362,In_718);
or U743 (N_743,In_283,In_1451);
or U744 (N_744,N_40,N_99);
nand U745 (N_745,In_427,N_229);
nand U746 (N_746,In_1167,In_1830);
nor U747 (N_747,In_1189,N_293);
nand U748 (N_748,In_1822,In_1853);
and U749 (N_749,In_674,In_1026);
and U750 (N_750,N_111,In_167);
and U751 (N_751,In_3,In_1051);
or U752 (N_752,N_307,N_397);
nand U753 (N_753,In_686,In_1647);
nand U754 (N_754,In_1669,In_643);
or U755 (N_755,N_548,In_101);
xor U756 (N_756,In_765,In_1242);
or U757 (N_757,In_238,In_216);
nand U758 (N_758,N_697,In_227);
nor U759 (N_759,N_516,N_368);
or U760 (N_760,N_710,N_128);
and U761 (N_761,N_629,In_383);
nand U762 (N_762,N_108,N_145);
xnor U763 (N_763,In_1140,In_1614);
or U764 (N_764,In_1384,N_285);
or U765 (N_765,In_1400,In_1637);
nand U766 (N_766,N_737,In_1508);
or U767 (N_767,N_663,N_623);
and U768 (N_768,In_746,N_148);
nand U769 (N_769,N_411,In_1217);
xor U770 (N_770,N_577,In_1476);
and U771 (N_771,N_156,In_835);
or U772 (N_772,In_366,In_466);
nor U773 (N_773,In_251,N_452);
xnor U774 (N_774,In_1707,In_1970);
and U775 (N_775,In_1770,N_719);
and U776 (N_776,N_282,In_781);
nor U777 (N_777,N_566,N_506);
or U778 (N_778,N_172,N_250);
nand U779 (N_779,In_744,N_352);
or U780 (N_780,N_518,In_1905);
nor U781 (N_781,N_665,In_1317);
nor U782 (N_782,N_455,N_591);
nand U783 (N_783,N_367,N_261);
or U784 (N_784,In_1203,In_519);
and U785 (N_785,In_893,In_363);
nand U786 (N_786,N_462,In_789);
xnor U787 (N_787,In_1536,In_978);
and U788 (N_788,In_941,In_15);
nor U789 (N_789,In_1191,In_1653);
nor U790 (N_790,N_389,N_647);
and U791 (N_791,In_133,In_1779);
and U792 (N_792,In_1077,N_485);
nor U793 (N_793,In_1979,In_963);
nor U794 (N_794,In_506,N_252);
and U795 (N_795,N_586,In_1944);
or U796 (N_796,N_662,In_1512);
or U797 (N_797,N_426,In_839);
and U798 (N_798,In_760,In_784);
xor U799 (N_799,In_1178,N_738);
nand U800 (N_800,N_441,N_551);
xnor U801 (N_801,In_1934,N_301);
nand U802 (N_802,N_189,In_315);
and U803 (N_803,In_722,N_195);
xor U804 (N_804,In_645,N_667);
or U805 (N_805,In_993,N_427);
nor U806 (N_806,N_384,N_749);
and U807 (N_807,N_645,In_296);
nor U808 (N_808,In_440,N_669);
xor U809 (N_809,N_78,N_740);
nand U810 (N_810,N_741,In_192);
xor U811 (N_811,N_182,In_149);
and U812 (N_812,N_701,N_443);
nand U813 (N_813,N_515,N_734);
and U814 (N_814,N_576,In_1652);
and U815 (N_815,N_472,In_1355);
nand U816 (N_816,N_486,In_160);
nor U817 (N_817,N_105,In_869);
nor U818 (N_818,N_315,N_568);
nor U819 (N_819,In_339,In_740);
xnor U820 (N_820,In_1107,In_653);
or U821 (N_821,N_339,In_1987);
nand U822 (N_822,In_1929,N_545);
nand U823 (N_823,In_1256,In_63);
nor U824 (N_824,In_1890,In_1791);
xor U825 (N_825,N_430,N_53);
nand U826 (N_826,N_334,In_1350);
nand U827 (N_827,In_886,N_507);
and U828 (N_828,In_1238,N_464);
and U829 (N_829,In_543,N_409);
or U830 (N_830,In_186,N_595);
xor U831 (N_831,N_708,N_553);
nor U832 (N_832,In_42,In_564);
nor U833 (N_833,In_801,N_605);
nand U834 (N_834,N_658,N_674);
nor U835 (N_835,N_554,In_624);
nand U836 (N_836,N_511,In_1817);
xnor U837 (N_837,N_354,N_110);
nand U838 (N_838,In_1284,In_1646);
nor U839 (N_839,N_668,N_366);
nor U840 (N_840,N_361,In_1922);
and U841 (N_841,In_246,In_858);
xor U842 (N_842,In_1683,In_1869);
and U843 (N_843,N_528,N_448);
nor U844 (N_844,In_990,N_521);
xor U845 (N_845,In_1072,In_522);
and U846 (N_846,In_850,N_364);
xor U847 (N_847,N_11,In_32);
nand U848 (N_848,N_538,In_1186);
and U849 (N_849,In_156,N_688);
nor U850 (N_850,N_689,N_542);
or U851 (N_851,In_1954,N_263);
nor U852 (N_852,In_929,In_579);
nand U853 (N_853,In_100,In_1361);
nor U854 (N_854,N_549,In_299);
nand U855 (N_855,N_565,N_207);
nand U856 (N_856,N_481,N_254);
nor U857 (N_857,In_697,N_322);
xnor U858 (N_858,In_1820,In_477);
xnor U859 (N_859,N_614,N_656);
and U860 (N_860,N_300,In_933);
or U861 (N_861,N_421,In_1057);
nand U862 (N_862,In_316,In_1336);
xnor U863 (N_863,N_365,In_67);
nor U864 (N_864,In_1962,N_318);
nor U865 (N_865,N_541,In_1618);
and U866 (N_866,In_1376,N_468);
or U867 (N_867,In_6,In_237);
nor U868 (N_868,N_590,N_329);
nand U869 (N_869,N_607,In_1046);
and U870 (N_870,N_336,In_1564);
nor U871 (N_871,In_1323,In_1576);
nand U872 (N_872,In_847,N_597);
xor U873 (N_873,N_652,In_827);
nor U874 (N_874,N_660,In_1978);
nand U875 (N_875,N_439,In_610);
nand U876 (N_876,N_114,N_6);
and U877 (N_877,In_528,In_70);
nor U878 (N_878,In_284,In_1559);
nand U879 (N_879,N_433,N_735);
nor U880 (N_880,N_712,In_1394);
nand U881 (N_881,In_48,In_311);
and U882 (N_882,In_1357,In_1549);
nand U883 (N_883,In_1876,In_147);
xor U884 (N_884,In_257,N_302);
nor U885 (N_885,In_1043,N_371);
nand U886 (N_886,N_723,N_319);
nand U887 (N_887,In_208,In_728);
and U888 (N_888,N_489,In_979);
or U889 (N_889,N_146,In_1022);
or U890 (N_890,In_582,In_95);
and U891 (N_891,N_583,N_703);
nand U892 (N_892,In_818,In_1494);
nor U893 (N_893,In_1092,In_961);
and U894 (N_894,In_1344,N_696);
or U895 (N_895,In_354,In_1847);
or U896 (N_896,In_1654,N_479);
xnor U897 (N_897,N_303,In_957);
and U898 (N_898,N_77,In_1395);
xnor U899 (N_899,In_865,N_160);
and U900 (N_900,In_518,N_51);
and U901 (N_901,N_88,N_18);
xor U902 (N_902,N_348,N_180);
nor U903 (N_903,N_679,N_159);
xor U904 (N_904,N_402,N_609);
nand U905 (N_905,N_291,In_773);
nor U906 (N_906,In_1034,N_608);
or U907 (N_907,N_248,In_1013);
nand U908 (N_908,In_652,In_437);
or U909 (N_909,In_631,In_16);
nand U910 (N_910,N_580,N_471);
nand U911 (N_911,In_225,N_509);
nor U912 (N_912,N_598,In_548);
and U913 (N_913,N_681,In_1590);
or U914 (N_914,In_1583,N_641);
and U915 (N_915,N_638,In_247);
or U916 (N_916,In_406,In_1142);
xnor U917 (N_917,In_551,In_1248);
nand U918 (N_918,N_569,N_278);
xnor U919 (N_919,In_683,In_945);
or U920 (N_920,In_408,In_572);
nand U921 (N_921,In_1660,In_1009);
or U922 (N_922,N_513,N_527);
nor U923 (N_923,N_349,N_606);
nor U924 (N_924,N_241,In_677);
or U925 (N_925,N_550,N_547);
or U926 (N_926,N_512,In_1025);
xnor U927 (N_927,In_297,N_559);
nor U928 (N_928,N_226,In_442);
nor U929 (N_929,In_1644,In_1373);
nand U930 (N_930,N_398,In_1491);
and U931 (N_931,In_189,In_989);
xnor U932 (N_932,In_143,N_274);
or U933 (N_933,In_270,In_360);
nor U934 (N_934,In_431,In_1766);
nor U935 (N_935,N_574,In_1567);
nand U936 (N_936,In_1160,N_29);
xnor U937 (N_937,N_152,N_685);
nand U938 (N_938,In_180,N_380);
xor U939 (N_939,In_660,N_579);
nor U940 (N_940,N_407,N_709);
xor U941 (N_941,In_178,In_1529);
nand U942 (N_942,In_1569,N_496);
nor U943 (N_943,N_539,In_524);
xor U944 (N_944,In_1676,In_179);
xor U945 (N_945,In_636,In_1208);
and U946 (N_946,In_1127,In_713);
nand U947 (N_947,In_1232,In_197);
xor U948 (N_948,N_716,In_1577);
nand U949 (N_949,N_149,N_288);
nand U950 (N_950,In_556,N_262);
and U951 (N_951,In_1866,N_594);
nor U952 (N_952,In_823,N_219);
nor U953 (N_953,N_731,In_1351);
xor U954 (N_954,In_1511,In_1419);
or U955 (N_955,N_342,In_1439);
and U956 (N_956,N_236,N_555);
nand U957 (N_957,N_721,N_121);
nor U958 (N_958,N_746,In_261);
or U959 (N_959,In_319,N_39);
nor U960 (N_960,In_1664,In_1111);
and U961 (N_961,N_643,N_264);
and U962 (N_962,In_1482,In_91);
xor U963 (N_963,N_648,In_1589);
or U964 (N_964,In_445,In_814);
and U965 (N_965,In_318,N_363);
nor U966 (N_966,N_270,In_995);
or U967 (N_967,N_619,In_117);
nor U968 (N_968,N_584,In_938);
nor U969 (N_969,In_1405,In_1754);
nor U970 (N_970,N_321,In_712);
or U971 (N_971,N_540,N_622);
and U972 (N_972,In_905,In_1625);
xor U973 (N_973,In_1983,In_380);
nor U974 (N_974,In_1027,N_267);
and U975 (N_975,In_457,In_1205);
nor U976 (N_976,In_845,In_1698);
or U977 (N_977,In_1547,N_694);
nand U978 (N_978,N_326,In_509);
nand U979 (N_979,N_376,In_351);
nand U980 (N_980,N_714,In_546);
nor U981 (N_981,N_356,In_1756);
xor U982 (N_982,In_480,In_1195);
or U983 (N_983,N_642,N_143);
nor U984 (N_984,In_1894,In_1828);
nand U985 (N_985,N_640,In_1259);
and U986 (N_986,In_783,N_733);
nand U987 (N_987,In_779,N_562);
or U988 (N_988,In_1322,In_1516);
nor U989 (N_989,In_1410,In_462);
nor U990 (N_990,In_1460,N_573);
xnor U991 (N_991,In_1084,N_492);
and U992 (N_992,N_242,In_635);
or U993 (N_993,In_1662,In_1440);
nand U994 (N_994,In_673,In_1401);
nand U995 (N_995,N_429,N_390);
nand U996 (N_996,In_1019,N_501);
nand U997 (N_997,N_193,N_388);
nand U998 (N_998,N_561,In_1049);
or U999 (N_999,In_1685,In_1694);
and U1000 (N_1000,In_53,N_406);
xor U1001 (N_1001,In_1308,N_498);
xnor U1002 (N_1002,N_815,N_255);
xor U1003 (N_1003,In_868,In_1871);
nand U1004 (N_1004,In_1579,N_693);
xor U1005 (N_1005,N_497,N_212);
xnor U1006 (N_1006,In_1824,N_238);
or U1007 (N_1007,In_1845,N_466);
nand U1008 (N_1008,N_841,N_37);
xnor U1009 (N_1009,N_924,In_1212);
nor U1010 (N_1010,N_373,In_1404);
xor U1011 (N_1011,N_533,N_338);
or U1012 (N_1012,In_388,In_1464);
nand U1013 (N_1013,In_1312,N_759);
or U1014 (N_1014,N_718,N_564);
nor U1015 (N_1015,In_1309,N_921);
or U1016 (N_1016,N_690,N_926);
or U1017 (N_1017,N_951,N_81);
and U1018 (N_1018,N_90,N_557);
and U1019 (N_1019,In_1041,In_1655);
nor U1020 (N_1020,In_1426,In_376);
nand U1021 (N_1021,N_726,In_1737);
nand U1022 (N_1022,N_965,In_265);
and U1023 (N_1023,In_1968,In_151);
nor U1024 (N_1024,N_934,N_906);
nor U1025 (N_1025,N_460,N_908);
and U1026 (N_1026,N_880,In_1056);
nor U1027 (N_1027,In_1601,N_986);
or U1028 (N_1028,In_717,In_371);
and U1029 (N_1029,N_331,In_194);
nand U1030 (N_1030,N_33,N_946);
xor U1031 (N_1031,N_980,N_764);
or U1032 (N_1032,In_470,In_1984);
nor U1033 (N_1033,In_605,N_295);
or U1034 (N_1034,N_437,N_911);
or U1035 (N_1035,In_1348,N_310);
xor U1036 (N_1036,In_267,N_812);
nor U1037 (N_1037,In_80,N_773);
nor U1038 (N_1038,N_297,N_385);
or U1039 (N_1039,N_474,In_1839);
and U1040 (N_1040,N_953,In_570);
or U1041 (N_1041,In_334,In_739);
xor U1042 (N_1042,In_973,In_1916);
nand U1043 (N_1043,N_994,In_435);
nor U1044 (N_1044,In_866,N_66);
and U1045 (N_1045,N_932,N_757);
nor U1046 (N_1046,In_1852,N_919);
nand U1047 (N_1047,N_950,N_677);
and U1048 (N_1048,In_1762,N_852);
or U1049 (N_1049,In_1148,N_634);
nand U1050 (N_1050,N_107,N_659);
or U1051 (N_1051,N_915,N_977);
nor U1052 (N_1052,In_800,N_675);
nor U1053 (N_1053,N_191,In_804);
nor U1054 (N_1054,N_886,In_1649);
and U1055 (N_1055,N_628,In_1821);
xnor U1056 (N_1056,N_581,In_756);
nor U1057 (N_1057,In_310,In_1210);
xor U1058 (N_1058,In_1602,N_353);
nand U1059 (N_1059,In_1747,N_631);
xnor U1060 (N_1060,N_535,N_844);
nor U1061 (N_1061,In_175,In_8);
nor U1062 (N_1062,N_480,In_1696);
nor U1063 (N_1063,In_1146,In_622);
nor U1064 (N_1064,N_728,N_896);
nor U1065 (N_1065,N_357,In_1794);
xnor U1066 (N_1066,In_1543,N_670);
or U1067 (N_1067,In_998,N_879);
nor U1068 (N_1068,N_791,N_21);
nand U1069 (N_1069,N_337,In_1759);
and U1070 (N_1070,N_266,N_552);
nor U1071 (N_1071,N_345,In_1420);
nand U1072 (N_1072,In_950,N_273);
and U1073 (N_1073,N_196,N_362);
and U1074 (N_1074,In_505,In_1721);
nand U1075 (N_1075,N_621,In_355);
nor U1076 (N_1076,N_12,In_368);
nand U1077 (N_1077,In_520,In_19);
xor U1078 (N_1078,In_439,N_461);
xnor U1079 (N_1079,N_784,In_1016);
nor U1080 (N_1080,In_531,N_936);
or U1081 (N_1081,N_769,N_494);
nor U1082 (N_1082,N_698,In_896);
and U1083 (N_1083,In_719,In_417);
nand U1084 (N_1084,N_861,N_624);
nand U1085 (N_1085,In_1280,N_109);
nand U1086 (N_1086,N_627,In_329);
xnor U1087 (N_1087,N_536,In_1532);
nand U1088 (N_1088,N_314,In_1782);
xnor U1089 (N_1089,In_68,In_894);
xnor U1090 (N_1090,N_739,N_447);
nor U1091 (N_1091,In_553,N_611);
nand U1092 (N_1092,In_1079,N_360);
xnor U1093 (N_1093,N_992,In_895);
nand U1094 (N_1094,N_695,In_51);
or U1095 (N_1095,In_726,N_484);
and U1096 (N_1096,N_453,N_525);
nor U1097 (N_1097,In_688,N_866);
and U1098 (N_1098,In_1777,In_616);
and U1099 (N_1099,N_560,N_585);
nor U1100 (N_1100,N_885,N_955);
or U1101 (N_1101,N_772,N_730);
or U1102 (N_1102,N_556,N_650);
xor U1103 (N_1103,N_813,In_668);
nand U1104 (N_1104,In_1008,In_1434);
or U1105 (N_1105,N_438,In_1479);
nor U1106 (N_1106,In_1834,In_454);
xor U1107 (N_1107,N_958,In_916);
or U1108 (N_1108,N_910,In_1375);
nand U1109 (N_1109,N_949,In_1251);
xor U1110 (N_1110,N_478,N_969);
and U1111 (N_1111,N_204,N_304);
nand U1112 (N_1112,In_1249,In_335);
nor U1113 (N_1113,In_1218,In_217);
nor U1114 (N_1114,N_747,N_95);
nor U1115 (N_1115,N_783,N_931);
nand U1116 (N_1116,N_822,N_801);
xor U1117 (N_1117,N_3,In_1535);
nand U1118 (N_1118,N_587,N_558);
nand U1119 (N_1119,In_857,In_791);
and U1120 (N_1120,In_1899,In_353);
nand U1121 (N_1121,N_922,N_126);
nor U1122 (N_1122,N_524,N_761);
or U1123 (N_1123,In_1466,In_1012);
nor U1124 (N_1124,N_793,In_1418);
nor U1125 (N_1125,N_519,N_963);
xor U1126 (N_1126,N_970,In_1973);
and U1127 (N_1127,N_891,N_790);
or U1128 (N_1128,N_989,N_993);
nand U1129 (N_1129,N_636,N_346);
nand U1130 (N_1130,In_1538,N_850);
or U1131 (N_1131,In_475,N_763);
xor U1132 (N_1132,N_745,In_1370);
or U1133 (N_1133,N_625,N_704);
or U1134 (N_1134,N_952,In_1144);
xor U1135 (N_1135,In_834,In_632);
nor U1136 (N_1136,N_988,In_292);
nand U1137 (N_1137,In_418,In_1677);
nand U1138 (N_1138,N_224,In_1667);
and U1139 (N_1139,In_27,In_1517);
and U1140 (N_1140,In_1561,In_607);
nor U1141 (N_1141,N_707,N_416);
nand U1142 (N_1142,N_63,In_721);
nor U1143 (N_1143,N_916,N_305);
or U1144 (N_1144,N_699,In_785);
xor U1145 (N_1145,In_690,In_1230);
xor U1146 (N_1146,N_504,In_1666);
or U1147 (N_1147,In_980,In_830);
nand U1148 (N_1148,N_754,In_820);
xnor U1149 (N_1149,N_853,N_810);
or U1150 (N_1150,In_603,In_521);
xnor U1151 (N_1151,In_921,N_945);
nor U1152 (N_1152,In_997,In_786);
xor U1153 (N_1153,N_635,N_680);
and U1154 (N_1154,N_615,In_1861);
nand U1155 (N_1155,In_1671,N_942);
nor U1156 (N_1156,N_918,N_355);
nor U1157 (N_1157,N_998,N_775);
nand U1158 (N_1158,N_770,N_626);
nand U1159 (N_1159,N_616,N_482);
nand U1160 (N_1160,In_1818,N_678);
and U1161 (N_1161,In_321,In_1920);
nor U1162 (N_1162,N_691,N_292);
nand U1163 (N_1163,N_930,N_222);
xnor U1164 (N_1164,In_1773,N_661);
xor U1165 (N_1165,N_987,In_1957);
or U1166 (N_1166,N_211,In_1002);
and U1167 (N_1167,N_617,In_436);
nor U1168 (N_1168,N_644,In_1147);
nor U1169 (N_1169,In_880,In_1435);
and U1170 (N_1170,In_1787,N_232);
nand U1171 (N_1171,In_1145,N_655);
or U1172 (N_1172,N_370,In_912);
or U1173 (N_1173,In_611,In_1382);
or U1174 (N_1174,N_543,N_620);
or U1175 (N_1175,N_84,N_858);
nor U1176 (N_1176,In_72,In_883);
or U1177 (N_1177,In_627,In_1521);
nor U1178 (N_1178,In_1358,N_436);
or U1179 (N_1179,N_960,In_1102);
nand U1180 (N_1180,N_887,N_847);
and U1181 (N_1181,In_449,N_865);
or U1182 (N_1182,N_755,N_578);
xnor U1183 (N_1183,N_526,N_954);
or U1184 (N_1184,In_1472,N_743);
nor U1185 (N_1185,N_837,N_900);
nand U1186 (N_1186,In_736,N_742);
nor U1187 (N_1187,In_672,In_960);
nor U1188 (N_1188,In_882,N_898);
nand U1189 (N_1189,In_415,N_317);
or U1190 (N_1190,In_1059,N_848);
xnor U1191 (N_1191,In_693,In_162);
and U1192 (N_1192,In_1333,N_736);
nand U1193 (N_1193,In_1708,N_125);
nand U1194 (N_1194,N_630,N_768);
nand U1195 (N_1195,N_713,N_944);
and U1196 (N_1196,N_927,N_392);
nor U1197 (N_1197,In_1504,N_653);
or U1198 (N_1198,In_1730,N_711);
xnor U1199 (N_1199,In_170,In_1176);
and U1200 (N_1200,N_800,N_442);
nor U1201 (N_1201,N_839,N_725);
or U1202 (N_1202,In_1126,N_256);
xnor U1203 (N_1203,In_1875,N_13);
nand U1204 (N_1204,N_758,N_563);
and U1205 (N_1205,In_108,In_966);
nor U1206 (N_1206,In_401,In_1131);
nor U1207 (N_1207,N_103,N_873);
xnor U1208 (N_1208,N_588,N_717);
nor U1209 (N_1209,In_1700,N_687);
xnor U1210 (N_1210,N_277,N_818);
or U1211 (N_1211,N_646,In_1339);
or U1212 (N_1212,In_46,In_249);
xor U1213 (N_1213,N_840,N_855);
nor U1214 (N_1214,N_832,In_1169);
xor U1215 (N_1215,In_1734,N_975);
or U1216 (N_1216,N_604,N_572);
xor U1217 (N_1217,In_774,In_571);
nor U1218 (N_1218,N_825,N_824);
and U1219 (N_1219,In_333,In_1143);
xor U1220 (N_1220,N_682,In_152);
nor U1221 (N_1221,N_846,In_1293);
or U1222 (N_1222,N_787,In_1872);
nand U1223 (N_1223,N_457,N_499);
nand U1224 (N_1224,N_732,In_1112);
xor U1225 (N_1225,In_1310,In_258);
and U1226 (N_1226,In_191,N_888);
xnor U1227 (N_1227,In_962,N_55);
nor U1228 (N_1228,N_335,N_947);
nor U1229 (N_1229,In_138,N_849);
and U1230 (N_1230,N_882,In_485);
and U1231 (N_1231,In_13,In_134);
xor U1232 (N_1232,N_249,N_914);
and U1233 (N_1233,N_766,In_1257);
and U1234 (N_1234,N_20,N_218);
nor U1235 (N_1235,In_1266,In_172);
xor U1236 (N_1236,In_1135,In_1784);
nand U1237 (N_1237,In_772,N_316);
or U1238 (N_1238,In_913,In_1965);
and U1239 (N_1239,In_1991,N_213);
nand U1240 (N_1240,N_28,N_603);
xor U1241 (N_1241,In_974,In_256);
nand U1242 (N_1242,In_1735,N_895);
xor U1243 (N_1243,N_330,In_384);
or U1244 (N_1244,N_933,In_1552);
nand U1245 (N_1245,In_568,In_513);
nor U1246 (N_1246,N_514,In_1216);
or U1247 (N_1247,In_1332,N_829);
and U1248 (N_1248,N_870,N_48);
xnor U1249 (N_1249,In_324,In_1571);
xnor U1250 (N_1250,N_118,N_820);
and U1251 (N_1251,In_1769,N_1119);
xor U1252 (N_1252,N_1174,N_418);
or U1253 (N_1253,N_1006,N_253);
or U1254 (N_1254,N_279,In_344);
or U1255 (N_1255,In_148,N_651);
nand U1256 (N_1256,In_455,N_1110);
nor U1257 (N_1257,In_1790,N_1023);
and U1258 (N_1258,N_1146,N_981);
nand U1259 (N_1259,In_1620,N_781);
nand U1260 (N_1260,N_1053,N_1200);
and U1261 (N_1261,N_1032,N_923);
xnor U1262 (N_1262,In_1604,N_881);
or U1263 (N_1263,N_1173,N_828);
and U1264 (N_1264,N_1092,N_215);
or U1265 (N_1265,In_1503,N_715);
nand U1266 (N_1266,N_1060,N_779);
nand U1267 (N_1267,N_1050,N_141);
nand U1268 (N_1268,N_1212,In_1381);
xor U1269 (N_1269,N_65,In_1136);
xor U1270 (N_1270,In_1258,N_1164);
and U1271 (N_1271,In_716,N_1135);
nor U1272 (N_1272,N_1215,N_1096);
and U1273 (N_1273,N_673,In_1465);
and U1274 (N_1274,N_973,N_806);
or U1275 (N_1275,N_610,In_811);
nand U1276 (N_1276,N_1090,In_1352);
xor U1277 (N_1277,N_1176,In_78);
xor U1278 (N_1278,N_537,N_298);
or U1279 (N_1279,N_52,N_1087);
nand U1280 (N_1280,N_1150,In_1846);
and U1281 (N_1281,N_903,N_996);
or U1282 (N_1282,N_133,N_851);
xor U1283 (N_1283,N_1036,N_913);
nand U1284 (N_1284,N_1045,In_911);
and U1285 (N_1285,In_536,N_257);
or U1286 (N_1286,In_1055,N_1038);
xnor U1287 (N_1287,N_144,N_0);
nand U1288 (N_1288,N_974,N_1148);
xnor U1289 (N_1289,N_1161,N_1001);
or U1290 (N_1290,N_1192,N_1179);
xnor U1291 (N_1291,N_420,In_1657);
nor U1292 (N_1292,In_1298,N_1228);
nor U1293 (N_1293,N_534,N_948);
and U1294 (N_1294,In_1295,N_1039);
nor U1295 (N_1295,In_1173,N_1208);
xor U1296 (N_1296,N_1057,In_634);
or U1297 (N_1297,In_1874,N_756);
xor U1298 (N_1298,N_664,N_1095);
or U1299 (N_1299,N_1120,N_1028);
and U1300 (N_1300,N_454,N_1015);
nand U1301 (N_1301,In_1940,In_1488);
and U1302 (N_1302,In_1570,N_505);
and U1303 (N_1303,In_331,N_894);
and U1304 (N_1304,N_854,In_129);
nand U1305 (N_1305,N_1071,In_332);
nor U1306 (N_1306,N_786,In_1985);
xnor U1307 (N_1307,N_686,N_982);
nor U1308 (N_1308,N_883,In_1574);
xor U1309 (N_1309,N_544,N_961);
nor U1310 (N_1310,N_819,N_1027);
and U1311 (N_1311,N_1112,In_651);
nor U1312 (N_1312,N_929,N_283);
and U1313 (N_1313,N_612,N_856);
and U1314 (N_1314,N_132,N_589);
xnor U1315 (N_1315,In_836,In_909);
xor U1316 (N_1316,In_201,N_1155);
xor U1317 (N_1317,N_1218,In_764);
xor U1318 (N_1318,N_1242,N_809);
and U1319 (N_1319,N_972,N_1127);
and U1320 (N_1320,N_417,N_1160);
and U1321 (N_1321,N_750,In_1913);
nor U1322 (N_1322,N_794,N_1205);
xnor U1323 (N_1323,N_502,N_869);
and U1324 (N_1324,N_722,In_1366);
nor U1325 (N_1325,N_920,In_1378);
and U1326 (N_1326,N_1075,N_672);
and U1327 (N_1327,In_82,N_1131);
and U1328 (N_1328,N_1193,N_744);
or U1329 (N_1329,N_1213,N_939);
and U1330 (N_1330,N_1147,N_531);
nand U1331 (N_1331,N_1073,N_666);
nand U1332 (N_1332,N_503,N_1046);
and U1333 (N_1333,In_263,N_45);
nand U1334 (N_1334,N_683,In_1360);
nor U1335 (N_1335,In_200,N_1206);
xor U1336 (N_1336,In_1743,N_1126);
nor U1337 (N_1337,N_434,In_210);
nand U1338 (N_1338,N_1033,N_1217);
or U1339 (N_1339,In_268,In_790);
and U1340 (N_1340,In_438,In_1032);
nor U1341 (N_1341,In_510,N_1158);
nand U1342 (N_1342,In_707,N_1064);
nand U1343 (N_1343,N_802,N_1151);
nor U1344 (N_1344,N_765,N_1198);
and U1345 (N_1345,N_446,In_287);
or U1346 (N_1346,N_1072,N_1044);
nand U1347 (N_1347,N_602,In_1050);
nor U1348 (N_1348,N_1184,N_1247);
nor U1349 (N_1349,In_584,N_966);
xnor U1350 (N_1350,N_1076,N_500);
or U1351 (N_1351,N_1108,N_633);
xnor U1352 (N_1352,N_1171,N_777);
xnor U1353 (N_1353,N_999,In_544);
nand U1354 (N_1354,N_1098,N_874);
nor U1355 (N_1355,N_54,N_36);
or U1356 (N_1356,N_1139,N_412);
and U1357 (N_1357,N_163,N_860);
nand U1358 (N_1358,In_434,N_1144);
and U1359 (N_1359,N_859,N_1041);
nand U1360 (N_1360,N_1105,N_814);
nor U1361 (N_1361,N_1180,N_976);
nand U1362 (N_1362,In_86,In_1809);
nor U1363 (N_1363,N_1113,N_523);
nor U1364 (N_1364,N_1025,N_31);
or U1365 (N_1365,N_1012,N_1037);
nor U1366 (N_1366,N_968,N_795);
xor U1367 (N_1367,In_1554,In_761);
nor U1368 (N_1368,In_776,In_1767);
nor U1369 (N_1369,N_940,N_943);
nand U1370 (N_1370,N_1009,In_1758);
or U1371 (N_1371,N_323,In_165);
nand U1372 (N_1372,In_1101,In_1898);
xor U1373 (N_1373,In_405,N_979);
xor U1374 (N_1374,N_978,N_1034);
nand U1375 (N_1375,N_796,N_1074);
or U1376 (N_1376,In_1573,N_884);
nor U1377 (N_1377,N_767,In_57);
xor U1378 (N_1378,N_785,In_735);
or U1379 (N_1379,N_1070,N_1052);
nand U1380 (N_1380,N_845,In_766);
or U1381 (N_1381,In_1515,N_1142);
xnor U1382 (N_1382,In_1623,N_613);
xor U1383 (N_1383,N_632,N_657);
xor U1384 (N_1384,N_1104,N_1022);
or U1385 (N_1385,In_1097,N_1141);
nand U1386 (N_1386,In_198,N_676);
nand U1387 (N_1387,N_328,N_1083);
and U1388 (N_1388,N_1040,N_760);
and U1389 (N_1389,In_872,N_1062);
nand U1390 (N_1390,N_1220,N_1190);
or U1391 (N_1391,N_1224,N_592);
xnor U1392 (N_1392,N_995,In_1507);
xnor U1393 (N_1393,N_1223,N_1154);
xor U1394 (N_1394,In_153,N_491);
and U1395 (N_1395,N_174,In_1229);
and U1396 (N_1396,N_1202,N_816);
and U1397 (N_1397,N_835,N_706);
nand U1398 (N_1398,N_778,N_1196);
or U1399 (N_1399,N_151,N_1048);
and U1400 (N_1400,N_984,N_287);
nand U1401 (N_1401,N_276,N_705);
or U1402 (N_1402,In_1471,N_1140);
xor U1403 (N_1403,N_827,In_1686);
or U1404 (N_1404,N_788,N_1232);
nor U1405 (N_1405,N_567,In_648);
xnor U1406 (N_1406,N_1226,N_162);
xor U1407 (N_1407,In_1201,N_1065);
xor U1408 (N_1408,N_38,N_1067);
or U1409 (N_1409,In_1359,N_1085);
or U1410 (N_1410,N_1097,N_1047);
xnor U1411 (N_1411,N_1031,N_1238);
xnor U1412 (N_1412,N_1229,N_44);
or U1413 (N_1413,N_596,In_767);
and U1414 (N_1414,In_1870,N_1243);
nor U1415 (N_1415,N_1014,N_271);
and U1416 (N_1416,N_1086,In_489);
or U1417 (N_1417,N_857,In_451);
and U1418 (N_1418,N_774,N_956);
nor U1419 (N_1419,N_909,N_751);
nor U1420 (N_1420,N_1118,N_834);
nor U1421 (N_1421,N_575,N_782);
nand U1422 (N_1422,N_1203,N_1000);
xor U1423 (N_1423,N_1167,N_1016);
xnor U1424 (N_1424,N_522,N_1166);
or U1425 (N_1425,N_1055,N_1170);
nand U1426 (N_1426,In_496,N_299);
nand U1427 (N_1427,N_517,N_510);
xor U1428 (N_1428,In_1104,In_928);
xnor U1429 (N_1429,In_115,N_1068);
or U1430 (N_1430,N_1079,N_762);
or U1431 (N_1431,N_938,N_530);
or U1432 (N_1432,N_872,N_243);
or U1433 (N_1433,N_753,N_1143);
and U1434 (N_1434,N_1063,N_1207);
xnor U1435 (N_1435,N_1201,N_1177);
xor U1436 (N_1436,N_1010,N_1239);
xor U1437 (N_1437,N_889,N_1005);
xor U1438 (N_1438,N_8,N_864);
xor U1439 (N_1439,N_135,In_1836);
xnor U1440 (N_1440,In_1802,N_1102);
and U1441 (N_1441,N_1245,N_1175);
nand U1442 (N_1442,N_520,In_1030);
or U1443 (N_1443,N_1227,In_620);
nand U1444 (N_1444,N_1162,N_897);
xor U1445 (N_1445,In_174,N_805);
nor U1446 (N_1446,In_18,N_1029);
or U1447 (N_1447,In_59,N_1081);
nor U1448 (N_1448,N_877,N_797);
nor U1449 (N_1449,N_649,N_1156);
and U1450 (N_1450,In_1267,N_1136);
and U1451 (N_1451,N_1043,In_1343);
xnor U1452 (N_1452,N_997,N_69);
nand U1453 (N_1453,In_1374,N_907);
or U1454 (N_1454,N_727,In_73);
nor U1455 (N_1455,N_435,N_1165);
and U1456 (N_1456,N_369,N_826);
and U1457 (N_1457,N_1115,N_671);
nand U1458 (N_1458,N_1159,N_962);
nand U1459 (N_1459,N_1082,N_1019);
and U1460 (N_1460,N_383,In_1924);
and U1461 (N_1461,N_1011,N_1109);
nor U1462 (N_1462,N_359,In_250);
xnor U1463 (N_1463,N_1149,N_771);
nand U1464 (N_1464,In_490,In_286);
nand U1465 (N_1465,N_1172,N_1133);
xor U1466 (N_1466,N_1153,In_1213);
and U1467 (N_1467,In_918,N_1099);
and U1468 (N_1468,N_381,In_1168);
xnor U1469 (N_1469,N_1013,N_821);
and U1470 (N_1470,N_899,In_1045);
and U1471 (N_1471,In_802,N_1026);
nand U1472 (N_1472,N_153,N_684);
or U1473 (N_1473,In_1406,N_1186);
nor U1474 (N_1474,N_451,In_1972);
xor U1475 (N_1475,In_341,N_729);
and U1476 (N_1476,In_1939,N_1002);
and U1477 (N_1477,N_1122,In_870);
nand U1478 (N_1478,N_862,N_1194);
nor U1479 (N_1479,N_50,N_905);
xor U1480 (N_1480,N_878,N_351);
nand U1481 (N_1481,In_1584,In_1807);
nand U1482 (N_1482,N_971,N_1084);
and U1483 (N_1483,N_106,In_1294);
and U1484 (N_1484,N_206,In_1065);
xnor U1485 (N_1485,In_1431,In_340);
or U1486 (N_1486,In_1170,N_1248);
xnor U1487 (N_1487,N_508,N_990);
xor U1488 (N_1488,In_971,In_795);
xor U1489 (N_1489,N_532,N_1195);
nand U1490 (N_1490,N_1042,N_639);
or U1491 (N_1491,In_891,In_1906);
nand U1492 (N_1492,N_892,N_379);
nor U1493 (N_1493,N_1134,N_902);
nor U1494 (N_1494,N_571,In_1149);
nor U1495 (N_1495,In_1129,N_863);
or U1496 (N_1496,N_1061,In_947);
nor U1497 (N_1497,In_1423,In_691);
nor U1498 (N_1498,N_1216,In_856);
and U1499 (N_1499,In_867,N_808);
nand U1500 (N_1500,N_1130,N_1357);
nor U1501 (N_1501,N_1386,N_1335);
and U1502 (N_1502,N_1296,N_1415);
nand U1503 (N_1503,N_1305,In_662);
nor U1504 (N_1504,N_1401,N_1449);
nor U1505 (N_1505,N_1094,N_1469);
or U1506 (N_1506,N_600,In_348);
xor U1507 (N_1507,N_1459,N_1480);
or U1508 (N_1508,N_1297,N_1418);
nor U1509 (N_1509,N_1222,N_1413);
or U1510 (N_1510,In_1095,N_1365);
or U1511 (N_1511,N_1157,N_1484);
nand U1512 (N_1512,N_823,In_493);
nand U1513 (N_1513,N_1138,In_981);
or U1514 (N_1514,N_1286,N_912);
and U1515 (N_1515,N_1101,N_1030);
xor U1516 (N_1516,N_1258,N_1467);
and U1517 (N_1517,N_1390,N_1356);
and U1518 (N_1518,N_47,N_1313);
or U1519 (N_1519,N_1451,N_1283);
or U1520 (N_1520,N_1008,N_1107);
and U1521 (N_1521,N_1051,N_1462);
or U1522 (N_1522,N_1406,N_1351);
nand U1523 (N_1523,N_1211,N_1331);
nand U1524 (N_1524,N_1182,N_1358);
xnor U1525 (N_1525,N_1091,In_1392);
or U1526 (N_1526,N_1293,In_927);
or U1527 (N_1527,N_112,N_404);
xor U1528 (N_1528,N_1450,N_1474);
and U1529 (N_1529,N_1470,N_1330);
xnor U1530 (N_1530,N_1319,N_1244);
xnor U1531 (N_1531,In_155,In_1430);
or U1532 (N_1532,In_768,N_1191);
nand U1533 (N_1533,N_1400,N_1306);
nand U1534 (N_1534,N_1264,N_983);
and U1535 (N_1535,In_1004,N_1121);
and U1536 (N_1536,N_1421,N_838);
and U1537 (N_1537,N_1377,N_1361);
and U1538 (N_1538,In_273,In_202);
nor U1539 (N_1539,In_1282,N_1487);
nor U1540 (N_1540,N_1349,N_1431);
or U1541 (N_1541,N_1442,In_1682);
xnor U1542 (N_1542,N_875,In_1447);
xor U1543 (N_1543,N_582,N_1254);
or U1544 (N_1544,N_1233,N_1396);
or U1545 (N_1545,N_1333,N_1281);
nand U1546 (N_1546,N_1219,N_1236);
and U1547 (N_1547,N_599,N_692);
and U1548 (N_1548,N_74,In_1324);
xor U1549 (N_1549,N_473,N_1277);
or U1550 (N_1550,N_1394,N_1366);
and U1551 (N_1551,N_1007,N_1326);
xnor U1552 (N_1552,N_1298,N_1443);
xor U1553 (N_1553,N_1252,N_1417);
xnor U1554 (N_1554,In_232,In_1925);
xnor U1555 (N_1555,N_1494,N_1285);
or U1556 (N_1556,In_23,N_1250);
nand U1557 (N_1557,N_1425,N_1301);
nor U1558 (N_1558,In_901,N_868);
nor U1559 (N_1559,N_1441,N_1472);
nor U1560 (N_1560,N_1473,N_275);
xnor U1561 (N_1561,N_1246,N_1493);
nand U1562 (N_1562,N_1477,N_1332);
xnor U1563 (N_1563,N_1380,N_917);
xnor U1564 (N_1564,In_1364,N_1446);
xnor U1565 (N_1565,N_904,N_1476);
xnor U1566 (N_1566,N_1381,In_144);
and U1567 (N_1567,N_1453,In_538);
xor U1568 (N_1568,N_935,N_1255);
nor U1569 (N_1569,N_546,N_1342);
nand U1570 (N_1570,N_1428,In_1067);
and U1571 (N_1571,In_1596,In_904);
or U1572 (N_1572,N_1374,N_1435);
nand U1573 (N_1573,N_843,N_1452);
nand U1574 (N_1574,N_1163,N_1169);
and U1575 (N_1575,In_708,N_1266);
and U1576 (N_1576,N_1486,N_1178);
or U1577 (N_1577,N_959,N_1398);
and U1578 (N_1578,N_1290,N_1391);
xnor U1579 (N_1579,N_836,In_837);
xor U1580 (N_1580,N_1265,N_1465);
and U1581 (N_1581,N_1320,N_1346);
or U1582 (N_1582,N_1350,N_1273);
and U1583 (N_1583,N_601,N_1270);
nand U1584 (N_1584,In_1527,In_1990);
nor U1585 (N_1585,In_1956,N_957);
and U1586 (N_1586,N_1234,N_1237);
xnor U1587 (N_1587,N_1369,N_1137);
or U1588 (N_1588,N_1230,In_593);
nor U1589 (N_1589,N_748,In_385);
and U1590 (N_1590,N_1455,N_1318);
or U1591 (N_1591,N_1309,N_1389);
or U1592 (N_1592,N_804,N_1321);
and U1593 (N_1593,N_1199,N_225);
nand U1594 (N_1594,N_1399,N_871);
nor U1595 (N_1595,N_1235,N_1385);
or U1596 (N_1596,N_1307,N_1325);
xor U1597 (N_1597,N_467,In_1215);
nor U1598 (N_1598,N_1371,N_1491);
or U1599 (N_1599,N_776,N_1189);
and U1600 (N_1600,N_155,N_1372);
xor U1601 (N_1601,N_1495,N_1225);
xor U1602 (N_1602,In_338,In_1621);
nor U1603 (N_1603,N_1249,In_1296);
or U1604 (N_1604,N_1353,N_1498);
nand U1605 (N_1605,N_1403,N_1379);
and U1606 (N_1606,In_1320,N_1308);
xor U1607 (N_1607,N_1024,In_1276);
or U1608 (N_1608,N_1383,In_203);
xnor U1609 (N_1609,N_570,N_1479);
or U1610 (N_1610,N_1355,N_1089);
or U1611 (N_1611,N_1183,N_1289);
xnor U1612 (N_1612,N_1221,N_1341);
or U1613 (N_1613,N_1058,N_1338);
nand U1614 (N_1614,N_1059,N_1395);
xnor U1615 (N_1615,N_1466,N_1460);
nand U1616 (N_1616,N_1420,N_280);
nor U1617 (N_1617,N_1316,N_1483);
and U1618 (N_1618,N_1416,N_1481);
or U1619 (N_1619,N_789,N_1328);
and U1620 (N_1620,N_422,N_529);
xnor U1621 (N_1621,In_474,N_811);
nor U1622 (N_1622,N_1433,N_1388);
nor U1623 (N_1623,In_704,N_1314);
nor U1624 (N_1624,N_1344,N_1303);
xnor U1625 (N_1625,N_1125,N_1497);
nor U1626 (N_1626,N_284,N_1124);
nand U1627 (N_1627,N_1021,N_1257);
or U1628 (N_1628,N_1387,N_1304);
nor U1629 (N_1629,N_967,N_1375);
and U1630 (N_1630,N_80,N_1410);
nand U1631 (N_1631,N_129,N_1269);
or U1632 (N_1632,N_377,N_1384);
or U1633 (N_1633,N_1251,In_94);
and U1634 (N_1634,N_1204,N_344);
nor U1635 (N_1635,N_35,N_1444);
xor U1636 (N_1636,N_1376,N_1188);
and U1637 (N_1637,N_1327,In_1206);
and U1638 (N_1638,In_885,N_1368);
and U1639 (N_1639,N_1294,N_1187);
nor U1640 (N_1640,In_21,N_1426);
nand U1641 (N_1641,N_1276,N_702);
and U1642 (N_1642,N_1348,N_1323);
nor U1643 (N_1643,In_1014,N_792);
or U1644 (N_1644,In_1877,In_1952);
xnor U1645 (N_1645,N_1334,N_1448);
xor U1646 (N_1646,N_893,N_1440);
or U1647 (N_1647,N_1069,N_1492);
nand U1648 (N_1648,N_901,In_209);
xor U1649 (N_1649,N_1049,N_1412);
or U1650 (N_1650,N_1363,N_1329);
xor U1651 (N_1651,N_618,N_1409);
nand U1652 (N_1652,In_56,N_752);
xor U1653 (N_1653,In_81,N_1185);
or U1654 (N_1654,N_1132,In_1651);
nand U1655 (N_1655,N_458,N_925);
and U1656 (N_1656,N_1439,N_1461);
or U1657 (N_1657,N_1100,In_532);
xor U1658 (N_1658,N_1103,N_831);
and U1659 (N_1659,N_1370,N_1468);
nor U1660 (N_1660,N_1272,N_1017);
nor U1661 (N_1661,N_1367,N_1434);
and U1662 (N_1662,N_833,N_1231);
and U1663 (N_1663,N_1437,N_1463);
xnor U1664 (N_1664,N_1430,N_817);
and U1665 (N_1665,N_1111,N_1364);
nand U1666 (N_1666,N_1457,N_1106);
and U1667 (N_1667,N_1490,N_1145);
and U1668 (N_1668,N_1478,In_1007);
nand U1669 (N_1669,N_1129,N_807);
or U1670 (N_1670,N_985,N_1279);
or U1671 (N_1671,N_1422,N_1056);
nor U1672 (N_1672,N_1339,N_1456);
nor U1673 (N_1673,N_1458,In_742);
xor U1674 (N_1674,N_1317,N_1436);
or U1675 (N_1675,N_1287,N_1210);
xnor U1676 (N_1676,N_1343,N_780);
nor U1677 (N_1677,In_1313,N_1496);
and U1678 (N_1678,N_1354,In_1757);
or U1679 (N_1679,N_876,N_941);
nor U1680 (N_1680,N_1078,N_43);
or U1681 (N_1681,N_1392,N_1360);
nand U1682 (N_1682,N_654,N_1340);
nand U1683 (N_1683,N_1080,N_1280);
and U1684 (N_1684,N_1429,In_1327);
nand U1685 (N_1685,In_5,N_1241);
nor U1686 (N_1686,N_1324,N_1197);
and U1687 (N_1687,N_1352,N_1402);
or U1688 (N_1688,N_1291,N_1093);
nand U1689 (N_1689,N_1117,N_1152);
nor U1690 (N_1690,N_1482,N_1004);
nor U1691 (N_1691,In_75,In_465);
xnor U1692 (N_1692,N_1256,N_1438);
nor U1693 (N_1693,N_1312,N_1077);
or U1694 (N_1694,In_762,N_1310);
and U1695 (N_1695,N_1263,N_332);
or U1696 (N_1696,N_1336,N_1123);
xor U1697 (N_1697,N_1378,N_867);
nand U1698 (N_1698,N_1489,N_1274);
and U1699 (N_1699,N_495,N_593);
nor U1700 (N_1700,N_1214,N_928);
nand U1701 (N_1701,N_1299,N_1018);
or U1702 (N_1702,In_64,N_1407);
xor U1703 (N_1703,In_1165,In_1785);
nand U1704 (N_1704,N_798,In_1884);
and U1705 (N_1705,N_842,N_1054);
xor U1706 (N_1706,N_1088,N_890);
nand U1707 (N_1707,N_1240,N_1271);
and U1708 (N_1708,N_1315,N_1302);
or U1709 (N_1709,N_1288,N_1275);
nor U1710 (N_1710,In_1542,N_1427);
xor U1711 (N_1711,N_124,N_964);
and U1712 (N_1712,N_1003,N_227);
and U1713 (N_1713,In_471,N_1419);
nor U1714 (N_1714,N_1414,N_1404);
xnor U1715 (N_1715,N_1300,In_378);
xor U1716 (N_1716,N_937,N_1337);
or U1717 (N_1717,N_1181,N_1411);
xnor U1718 (N_1718,N_1382,N_1373);
nor U1719 (N_1719,In_1452,N_1405);
nand U1720 (N_1720,N_1278,N_1020);
nor U1721 (N_1721,In_1300,N_1423);
nand U1722 (N_1722,In_873,N_1209);
and U1723 (N_1723,N_1282,N_1397);
xnor U1724 (N_1724,N_1432,N_1066);
xor U1725 (N_1725,N_1447,N_1445);
or U1726 (N_1726,N_1362,N_1408);
or U1727 (N_1727,N_637,In_1118);
xor U1728 (N_1728,N_1262,N_1347);
nand U1729 (N_1729,N_1035,N_1475);
nor U1730 (N_1730,N_1114,N_138);
nand U1731 (N_1731,N_1311,N_465);
nor U1732 (N_1732,In_254,N_991);
and U1733 (N_1733,N_720,N_1499);
nand U1734 (N_1734,N_803,N_1345);
and U1735 (N_1735,N_1359,N_1464);
or U1736 (N_1736,N_1295,In_1679);
or U1737 (N_1737,N_1454,N_1267);
nand U1738 (N_1738,N_1128,N_1168);
xnor U1739 (N_1739,N_1393,N_724);
xor U1740 (N_1740,N_700,N_1424);
and U1741 (N_1741,N_1488,In_1553);
xor U1742 (N_1742,N_1116,N_1253);
nand U1743 (N_1743,N_1259,N_1292);
and U1744 (N_1744,In_914,N_1322);
and U1745 (N_1745,In_710,N_1268);
xnor U1746 (N_1746,N_1471,N_1261);
nand U1747 (N_1747,N_799,N_830);
nor U1748 (N_1748,N_1260,N_1284);
or U1749 (N_1749,N_1485,N_102);
nor U1750 (N_1750,N_1558,N_1610);
nand U1751 (N_1751,N_1561,N_1594);
or U1752 (N_1752,N_1501,N_1741);
or U1753 (N_1753,N_1623,N_1596);
or U1754 (N_1754,N_1681,N_1582);
and U1755 (N_1755,N_1658,N_1527);
and U1756 (N_1756,N_1644,N_1615);
nor U1757 (N_1757,N_1735,N_1722);
and U1758 (N_1758,N_1673,N_1567);
or U1759 (N_1759,N_1647,N_1670);
xor U1760 (N_1760,N_1534,N_1740);
or U1761 (N_1761,N_1518,N_1713);
and U1762 (N_1762,N_1694,N_1607);
and U1763 (N_1763,N_1731,N_1618);
nand U1764 (N_1764,N_1676,N_1506);
nor U1765 (N_1765,N_1540,N_1746);
nor U1766 (N_1766,N_1630,N_1634);
xnor U1767 (N_1767,N_1662,N_1749);
nor U1768 (N_1768,N_1563,N_1507);
nand U1769 (N_1769,N_1698,N_1545);
and U1770 (N_1770,N_1584,N_1649);
and U1771 (N_1771,N_1668,N_1743);
nand U1772 (N_1772,N_1717,N_1583);
nor U1773 (N_1773,N_1553,N_1627);
nor U1774 (N_1774,N_1748,N_1712);
nand U1775 (N_1775,N_1577,N_1564);
nand U1776 (N_1776,N_1631,N_1654);
or U1777 (N_1777,N_1544,N_1529);
or U1778 (N_1778,N_1535,N_1747);
xnor U1779 (N_1779,N_1517,N_1559);
xnor U1780 (N_1780,N_1657,N_1692);
or U1781 (N_1781,N_1624,N_1711);
or U1782 (N_1782,N_1547,N_1639);
xor U1783 (N_1783,N_1680,N_1683);
and U1784 (N_1784,N_1736,N_1508);
nor U1785 (N_1785,N_1656,N_1520);
nor U1786 (N_1786,N_1591,N_1589);
and U1787 (N_1787,N_1605,N_1643);
nor U1788 (N_1788,N_1664,N_1744);
or U1789 (N_1789,N_1542,N_1661);
or U1790 (N_1790,N_1732,N_1652);
or U1791 (N_1791,N_1593,N_1574);
nor U1792 (N_1792,N_1504,N_1704);
and U1793 (N_1793,N_1580,N_1587);
and U1794 (N_1794,N_1539,N_1515);
and U1795 (N_1795,N_1679,N_1620);
or U1796 (N_1796,N_1629,N_1588);
nor U1797 (N_1797,N_1628,N_1665);
and U1798 (N_1798,N_1667,N_1617);
and U1799 (N_1799,N_1669,N_1636);
nor U1800 (N_1800,N_1666,N_1640);
or U1801 (N_1801,N_1682,N_1733);
and U1802 (N_1802,N_1590,N_1715);
or U1803 (N_1803,N_1659,N_1604);
nor U1804 (N_1804,N_1695,N_1536);
and U1805 (N_1805,N_1725,N_1608);
nor U1806 (N_1806,N_1560,N_1551);
xnor U1807 (N_1807,N_1609,N_1660);
and U1808 (N_1808,N_1510,N_1606);
and U1809 (N_1809,N_1718,N_1601);
or U1810 (N_1810,N_1557,N_1663);
nand U1811 (N_1811,N_1635,N_1730);
xor U1812 (N_1812,N_1648,N_1696);
nand U1813 (N_1813,N_1651,N_1500);
nor U1814 (N_1814,N_1552,N_1709);
nor U1815 (N_1815,N_1650,N_1576);
xor U1816 (N_1816,N_1546,N_1548);
nand U1817 (N_1817,N_1614,N_1622);
nand U1818 (N_1818,N_1688,N_1710);
nor U1819 (N_1819,N_1701,N_1505);
nor U1820 (N_1820,N_1519,N_1729);
or U1821 (N_1821,N_1565,N_1572);
nand U1822 (N_1822,N_1503,N_1646);
xor U1823 (N_1823,N_1602,N_1697);
nor U1824 (N_1824,N_1687,N_1599);
xor U1825 (N_1825,N_1714,N_1562);
nor U1826 (N_1826,N_1685,N_1674);
xnor U1827 (N_1827,N_1734,N_1638);
nand U1828 (N_1828,N_1525,N_1677);
xnor U1829 (N_1829,N_1700,N_1523);
nor U1830 (N_1830,N_1675,N_1611);
and U1831 (N_1831,N_1702,N_1616);
nand U1832 (N_1832,N_1653,N_1541);
xor U1833 (N_1833,N_1579,N_1726);
nor U1834 (N_1834,N_1693,N_1569);
xor U1835 (N_1835,N_1516,N_1691);
and U1836 (N_1836,N_1621,N_1571);
or U1837 (N_1837,N_1633,N_1502);
xor U1838 (N_1838,N_1678,N_1641);
and U1839 (N_1839,N_1556,N_1742);
xnor U1840 (N_1840,N_1655,N_1514);
nand U1841 (N_1841,N_1530,N_1671);
or U1842 (N_1842,N_1524,N_1739);
and U1843 (N_1843,N_1619,N_1521);
xor U1844 (N_1844,N_1566,N_1690);
nor U1845 (N_1845,N_1531,N_1684);
xnor U1846 (N_1846,N_1728,N_1745);
or U1847 (N_1847,N_1570,N_1511);
nor U1848 (N_1848,N_1554,N_1632);
nor U1849 (N_1849,N_1522,N_1600);
and U1850 (N_1850,N_1737,N_1586);
and U1851 (N_1851,N_1672,N_1707);
xnor U1852 (N_1852,N_1513,N_1724);
nand U1853 (N_1853,N_1719,N_1689);
and U1854 (N_1854,N_1720,N_1549);
xnor U1855 (N_1855,N_1568,N_1537);
nor U1856 (N_1856,N_1538,N_1526);
nor U1857 (N_1857,N_1625,N_1727);
and U1858 (N_1858,N_1716,N_1528);
nor U1859 (N_1859,N_1509,N_1626);
and U1860 (N_1860,N_1585,N_1578);
and U1861 (N_1861,N_1512,N_1533);
or U1862 (N_1862,N_1612,N_1723);
and U1863 (N_1863,N_1532,N_1721);
nand U1864 (N_1864,N_1597,N_1699);
nand U1865 (N_1865,N_1595,N_1598);
nor U1866 (N_1866,N_1603,N_1555);
xnor U1867 (N_1867,N_1738,N_1543);
nor U1868 (N_1868,N_1550,N_1705);
and U1869 (N_1869,N_1613,N_1686);
and U1870 (N_1870,N_1573,N_1708);
xnor U1871 (N_1871,N_1642,N_1645);
nand U1872 (N_1872,N_1575,N_1706);
xor U1873 (N_1873,N_1637,N_1592);
nor U1874 (N_1874,N_1703,N_1581);
and U1875 (N_1875,N_1642,N_1550);
nor U1876 (N_1876,N_1577,N_1631);
and U1877 (N_1877,N_1676,N_1568);
nor U1878 (N_1878,N_1643,N_1697);
or U1879 (N_1879,N_1608,N_1580);
or U1880 (N_1880,N_1601,N_1697);
nand U1881 (N_1881,N_1553,N_1633);
xor U1882 (N_1882,N_1707,N_1622);
nand U1883 (N_1883,N_1519,N_1739);
and U1884 (N_1884,N_1634,N_1595);
nand U1885 (N_1885,N_1660,N_1518);
nor U1886 (N_1886,N_1509,N_1698);
and U1887 (N_1887,N_1707,N_1521);
and U1888 (N_1888,N_1551,N_1600);
xnor U1889 (N_1889,N_1720,N_1583);
or U1890 (N_1890,N_1607,N_1535);
nor U1891 (N_1891,N_1669,N_1548);
and U1892 (N_1892,N_1558,N_1709);
or U1893 (N_1893,N_1577,N_1590);
xor U1894 (N_1894,N_1670,N_1642);
xor U1895 (N_1895,N_1520,N_1544);
xor U1896 (N_1896,N_1573,N_1591);
and U1897 (N_1897,N_1560,N_1737);
and U1898 (N_1898,N_1703,N_1732);
xnor U1899 (N_1899,N_1706,N_1514);
and U1900 (N_1900,N_1647,N_1611);
or U1901 (N_1901,N_1605,N_1676);
nand U1902 (N_1902,N_1719,N_1625);
and U1903 (N_1903,N_1553,N_1649);
or U1904 (N_1904,N_1644,N_1610);
nand U1905 (N_1905,N_1738,N_1606);
xor U1906 (N_1906,N_1718,N_1603);
and U1907 (N_1907,N_1509,N_1708);
nor U1908 (N_1908,N_1605,N_1721);
and U1909 (N_1909,N_1604,N_1571);
xor U1910 (N_1910,N_1726,N_1633);
and U1911 (N_1911,N_1727,N_1571);
or U1912 (N_1912,N_1731,N_1544);
xor U1913 (N_1913,N_1603,N_1613);
or U1914 (N_1914,N_1587,N_1619);
nor U1915 (N_1915,N_1749,N_1591);
xor U1916 (N_1916,N_1661,N_1639);
nor U1917 (N_1917,N_1546,N_1611);
nor U1918 (N_1918,N_1631,N_1549);
or U1919 (N_1919,N_1520,N_1566);
nor U1920 (N_1920,N_1541,N_1638);
xnor U1921 (N_1921,N_1643,N_1662);
nand U1922 (N_1922,N_1706,N_1687);
or U1923 (N_1923,N_1605,N_1730);
nand U1924 (N_1924,N_1671,N_1637);
nor U1925 (N_1925,N_1661,N_1561);
and U1926 (N_1926,N_1731,N_1589);
and U1927 (N_1927,N_1504,N_1502);
xor U1928 (N_1928,N_1581,N_1544);
nor U1929 (N_1929,N_1570,N_1683);
nor U1930 (N_1930,N_1579,N_1692);
and U1931 (N_1931,N_1635,N_1525);
and U1932 (N_1932,N_1730,N_1676);
and U1933 (N_1933,N_1613,N_1539);
nand U1934 (N_1934,N_1561,N_1625);
and U1935 (N_1935,N_1685,N_1696);
and U1936 (N_1936,N_1716,N_1728);
nor U1937 (N_1937,N_1665,N_1601);
nor U1938 (N_1938,N_1719,N_1653);
or U1939 (N_1939,N_1531,N_1686);
or U1940 (N_1940,N_1700,N_1702);
xor U1941 (N_1941,N_1700,N_1703);
nand U1942 (N_1942,N_1611,N_1707);
nand U1943 (N_1943,N_1626,N_1584);
nand U1944 (N_1944,N_1521,N_1633);
and U1945 (N_1945,N_1560,N_1572);
nor U1946 (N_1946,N_1673,N_1560);
nand U1947 (N_1947,N_1747,N_1513);
and U1948 (N_1948,N_1713,N_1549);
and U1949 (N_1949,N_1538,N_1632);
nand U1950 (N_1950,N_1650,N_1504);
nor U1951 (N_1951,N_1632,N_1667);
nand U1952 (N_1952,N_1682,N_1557);
and U1953 (N_1953,N_1736,N_1632);
or U1954 (N_1954,N_1562,N_1729);
xnor U1955 (N_1955,N_1512,N_1538);
xnor U1956 (N_1956,N_1692,N_1739);
or U1957 (N_1957,N_1652,N_1687);
nor U1958 (N_1958,N_1527,N_1587);
and U1959 (N_1959,N_1608,N_1507);
xor U1960 (N_1960,N_1696,N_1579);
and U1961 (N_1961,N_1700,N_1543);
nor U1962 (N_1962,N_1558,N_1604);
or U1963 (N_1963,N_1552,N_1690);
nand U1964 (N_1964,N_1577,N_1687);
nand U1965 (N_1965,N_1746,N_1533);
and U1966 (N_1966,N_1536,N_1660);
nand U1967 (N_1967,N_1730,N_1678);
nand U1968 (N_1968,N_1549,N_1712);
nand U1969 (N_1969,N_1522,N_1603);
and U1970 (N_1970,N_1737,N_1716);
and U1971 (N_1971,N_1647,N_1570);
nand U1972 (N_1972,N_1544,N_1727);
xnor U1973 (N_1973,N_1688,N_1697);
nor U1974 (N_1974,N_1542,N_1626);
nor U1975 (N_1975,N_1747,N_1684);
and U1976 (N_1976,N_1748,N_1641);
xor U1977 (N_1977,N_1700,N_1729);
and U1978 (N_1978,N_1740,N_1620);
xnor U1979 (N_1979,N_1536,N_1598);
and U1980 (N_1980,N_1618,N_1544);
xnor U1981 (N_1981,N_1636,N_1537);
nor U1982 (N_1982,N_1713,N_1659);
and U1983 (N_1983,N_1612,N_1579);
xnor U1984 (N_1984,N_1662,N_1670);
and U1985 (N_1985,N_1586,N_1595);
nor U1986 (N_1986,N_1524,N_1720);
or U1987 (N_1987,N_1716,N_1672);
and U1988 (N_1988,N_1583,N_1552);
or U1989 (N_1989,N_1723,N_1620);
and U1990 (N_1990,N_1674,N_1645);
xor U1991 (N_1991,N_1605,N_1616);
xnor U1992 (N_1992,N_1547,N_1597);
nor U1993 (N_1993,N_1575,N_1677);
or U1994 (N_1994,N_1548,N_1509);
and U1995 (N_1995,N_1506,N_1537);
and U1996 (N_1996,N_1645,N_1708);
nor U1997 (N_1997,N_1538,N_1569);
xor U1998 (N_1998,N_1523,N_1564);
xnor U1999 (N_1999,N_1547,N_1576);
and U2000 (N_2000,N_1992,N_1932);
xor U2001 (N_2001,N_1885,N_1809);
nor U2002 (N_2002,N_1990,N_1834);
nor U2003 (N_2003,N_1830,N_1897);
and U2004 (N_2004,N_1956,N_1882);
or U2005 (N_2005,N_1775,N_1979);
nand U2006 (N_2006,N_1850,N_1890);
nor U2007 (N_2007,N_1963,N_1957);
and U2008 (N_2008,N_1887,N_1792);
nand U2009 (N_2009,N_1759,N_1876);
nand U2010 (N_2010,N_1863,N_1845);
or U2011 (N_2011,N_1753,N_1823);
nand U2012 (N_2012,N_1942,N_1819);
nor U2013 (N_2013,N_1812,N_1991);
nand U2014 (N_2014,N_1790,N_1921);
xor U2015 (N_2015,N_1805,N_1813);
and U2016 (N_2016,N_1842,N_1922);
nand U2017 (N_2017,N_1877,N_1855);
nor U2018 (N_2018,N_1778,N_1904);
nand U2019 (N_2019,N_1983,N_1886);
nor U2020 (N_2020,N_1901,N_1782);
nor U2021 (N_2021,N_1961,N_1797);
or U2022 (N_2022,N_1950,N_1953);
nand U2023 (N_2023,N_1948,N_1865);
nor U2024 (N_2024,N_1879,N_1803);
or U2025 (N_2025,N_1935,N_1905);
and U2026 (N_2026,N_1980,N_1984);
nor U2027 (N_2027,N_1985,N_1978);
nor U2028 (N_2028,N_1930,N_1927);
nand U2029 (N_2029,N_1958,N_1915);
and U2030 (N_2030,N_1971,N_1808);
or U2031 (N_2031,N_1954,N_1784);
nor U2032 (N_2032,N_1928,N_1820);
or U2033 (N_2033,N_1866,N_1936);
nand U2034 (N_2034,N_1997,N_1777);
or U2035 (N_2035,N_1994,N_1947);
nor U2036 (N_2036,N_1924,N_1872);
and U2037 (N_2037,N_1796,N_1814);
nor U2038 (N_2038,N_1986,N_1829);
nor U2039 (N_2039,N_1795,N_1860);
and U2040 (N_2040,N_1919,N_1889);
nor U2041 (N_2041,N_1831,N_1825);
xor U2042 (N_2042,N_1940,N_1938);
nand U2043 (N_2043,N_1851,N_1896);
nor U2044 (N_2044,N_1780,N_1955);
nand U2045 (N_2045,N_1873,N_1756);
nor U2046 (N_2046,N_1828,N_1970);
nor U2047 (N_2047,N_1835,N_1871);
nand U2048 (N_2048,N_1769,N_1982);
or U2049 (N_2049,N_1976,N_1960);
and U2050 (N_2050,N_1996,N_1761);
xor U2051 (N_2051,N_1964,N_1969);
and U2052 (N_2052,N_1802,N_1859);
and U2053 (N_2053,N_1815,N_1962);
xor U2054 (N_2054,N_1826,N_1849);
nor U2055 (N_2055,N_1766,N_1917);
nand U2056 (N_2056,N_1848,N_1788);
nor U2057 (N_2057,N_1952,N_1906);
and U2058 (N_2058,N_1895,N_1837);
and U2059 (N_2059,N_1911,N_1843);
xnor U2060 (N_2060,N_1937,N_1852);
and U2061 (N_2061,N_1858,N_1838);
or U2062 (N_2062,N_1977,N_1884);
xnor U2063 (N_2063,N_1900,N_1910);
xnor U2064 (N_2064,N_1894,N_1998);
xor U2065 (N_2065,N_1781,N_1791);
xor U2066 (N_2066,N_1951,N_1916);
nand U2067 (N_2067,N_1836,N_1869);
nand U2068 (N_2068,N_1801,N_1888);
xnor U2069 (N_2069,N_1763,N_1966);
and U2070 (N_2070,N_1817,N_1883);
xor U2071 (N_2071,N_1908,N_1870);
nor U2072 (N_2072,N_1841,N_1768);
xnor U2073 (N_2073,N_1891,N_1989);
or U2074 (N_2074,N_1839,N_1974);
xor U2075 (N_2075,N_1776,N_1893);
nor U2076 (N_2076,N_1912,N_1907);
nor U2077 (N_2077,N_1750,N_1767);
and U2078 (N_2078,N_1965,N_1903);
or U2079 (N_2079,N_1810,N_1993);
and U2080 (N_2080,N_1968,N_1799);
nand U2081 (N_2081,N_1793,N_1755);
nand U2082 (N_2082,N_1967,N_1939);
nor U2083 (N_2083,N_1785,N_1923);
xnor U2084 (N_2084,N_1816,N_1945);
nand U2085 (N_2085,N_1874,N_1760);
and U2086 (N_2086,N_1875,N_1868);
or U2087 (N_2087,N_1827,N_1818);
and U2088 (N_2088,N_1757,N_1806);
or U2089 (N_2089,N_1765,N_1909);
or U2090 (N_2090,N_1867,N_1880);
nand U2091 (N_2091,N_1846,N_1856);
or U2092 (N_2092,N_1861,N_1931);
nor U2093 (N_2093,N_1847,N_1832);
or U2094 (N_2094,N_1786,N_1881);
and U2095 (N_2095,N_1764,N_1773);
nor U2096 (N_2096,N_1787,N_1771);
and U2097 (N_2097,N_1772,N_1944);
xor U2098 (N_2098,N_1914,N_1975);
nor U2099 (N_2099,N_1857,N_1934);
or U2100 (N_2100,N_1902,N_1822);
nor U2101 (N_2101,N_1821,N_1981);
or U2102 (N_2102,N_1920,N_1804);
or U2103 (N_2103,N_1941,N_1898);
xor U2104 (N_2104,N_1840,N_1824);
nor U2105 (N_2105,N_1758,N_1959);
and U2106 (N_2106,N_1913,N_1862);
and U2107 (N_2107,N_1752,N_1853);
or U2108 (N_2108,N_1751,N_1949);
nand U2109 (N_2109,N_1789,N_1754);
nand U2110 (N_2110,N_1943,N_1988);
or U2111 (N_2111,N_1929,N_1892);
and U2112 (N_2112,N_1933,N_1783);
xor U2113 (N_2113,N_1926,N_1854);
and U2114 (N_2114,N_1999,N_1762);
nand U2115 (N_2115,N_1798,N_1774);
or U2116 (N_2116,N_1779,N_1878);
nand U2117 (N_2117,N_1925,N_1794);
nand U2118 (N_2118,N_1807,N_1844);
nand U2119 (N_2119,N_1918,N_1800);
nand U2120 (N_2120,N_1899,N_1946);
nor U2121 (N_2121,N_1995,N_1972);
and U2122 (N_2122,N_1987,N_1864);
xor U2123 (N_2123,N_1770,N_1973);
or U2124 (N_2124,N_1833,N_1811);
or U2125 (N_2125,N_1809,N_1891);
xor U2126 (N_2126,N_1956,N_1793);
nand U2127 (N_2127,N_1862,N_1826);
xnor U2128 (N_2128,N_1823,N_1954);
or U2129 (N_2129,N_1819,N_1825);
xnor U2130 (N_2130,N_1838,N_1965);
xnor U2131 (N_2131,N_1818,N_1911);
nor U2132 (N_2132,N_1757,N_1949);
nand U2133 (N_2133,N_1768,N_1814);
and U2134 (N_2134,N_1800,N_1911);
xor U2135 (N_2135,N_1985,N_1824);
nand U2136 (N_2136,N_1939,N_1923);
xnor U2137 (N_2137,N_1940,N_1946);
nand U2138 (N_2138,N_1863,N_1972);
or U2139 (N_2139,N_1948,N_1946);
nand U2140 (N_2140,N_1796,N_1863);
or U2141 (N_2141,N_1915,N_1776);
xnor U2142 (N_2142,N_1861,N_1803);
and U2143 (N_2143,N_1991,N_1853);
nor U2144 (N_2144,N_1992,N_1931);
xor U2145 (N_2145,N_1999,N_1771);
and U2146 (N_2146,N_1911,N_1952);
or U2147 (N_2147,N_1877,N_1964);
and U2148 (N_2148,N_1765,N_1826);
and U2149 (N_2149,N_1978,N_1750);
nor U2150 (N_2150,N_1979,N_1773);
or U2151 (N_2151,N_1827,N_1931);
or U2152 (N_2152,N_1836,N_1993);
xnor U2153 (N_2153,N_1877,N_1828);
or U2154 (N_2154,N_1796,N_1949);
xor U2155 (N_2155,N_1958,N_1845);
xnor U2156 (N_2156,N_1845,N_1828);
xor U2157 (N_2157,N_1944,N_1888);
xor U2158 (N_2158,N_1774,N_1814);
and U2159 (N_2159,N_1978,N_1791);
or U2160 (N_2160,N_1838,N_1974);
and U2161 (N_2161,N_1985,N_1962);
nor U2162 (N_2162,N_1948,N_1835);
xor U2163 (N_2163,N_1921,N_1791);
or U2164 (N_2164,N_1967,N_1863);
or U2165 (N_2165,N_1950,N_1927);
nand U2166 (N_2166,N_1789,N_1951);
xor U2167 (N_2167,N_1835,N_1834);
and U2168 (N_2168,N_1769,N_1974);
xor U2169 (N_2169,N_1922,N_1815);
nor U2170 (N_2170,N_1881,N_1890);
xnor U2171 (N_2171,N_1833,N_1858);
xor U2172 (N_2172,N_1955,N_1858);
nor U2173 (N_2173,N_1831,N_1910);
nor U2174 (N_2174,N_1930,N_1791);
nand U2175 (N_2175,N_1771,N_1951);
or U2176 (N_2176,N_1816,N_1836);
nor U2177 (N_2177,N_1766,N_1930);
nor U2178 (N_2178,N_1807,N_1999);
nor U2179 (N_2179,N_1756,N_1892);
and U2180 (N_2180,N_1969,N_1925);
nand U2181 (N_2181,N_1862,N_1846);
nor U2182 (N_2182,N_1809,N_1930);
nor U2183 (N_2183,N_1809,N_1965);
nand U2184 (N_2184,N_1934,N_1825);
nand U2185 (N_2185,N_1876,N_1772);
or U2186 (N_2186,N_1756,N_1932);
nor U2187 (N_2187,N_1889,N_1806);
or U2188 (N_2188,N_1907,N_1915);
nand U2189 (N_2189,N_1958,N_1781);
nand U2190 (N_2190,N_1946,N_1999);
and U2191 (N_2191,N_1788,N_1839);
nand U2192 (N_2192,N_1846,N_1854);
and U2193 (N_2193,N_1952,N_1842);
and U2194 (N_2194,N_1873,N_1961);
nand U2195 (N_2195,N_1936,N_1853);
nor U2196 (N_2196,N_1778,N_1761);
or U2197 (N_2197,N_1987,N_1853);
or U2198 (N_2198,N_1908,N_1760);
nand U2199 (N_2199,N_1943,N_1761);
nor U2200 (N_2200,N_1855,N_1852);
nand U2201 (N_2201,N_1867,N_1937);
xor U2202 (N_2202,N_1865,N_1961);
nor U2203 (N_2203,N_1891,N_1826);
and U2204 (N_2204,N_1950,N_1986);
or U2205 (N_2205,N_1924,N_1906);
and U2206 (N_2206,N_1887,N_1991);
xor U2207 (N_2207,N_1906,N_1855);
and U2208 (N_2208,N_1750,N_1753);
or U2209 (N_2209,N_1987,N_1984);
or U2210 (N_2210,N_1879,N_1835);
or U2211 (N_2211,N_1899,N_1952);
and U2212 (N_2212,N_1889,N_1793);
xnor U2213 (N_2213,N_1757,N_1785);
nor U2214 (N_2214,N_1851,N_1766);
nor U2215 (N_2215,N_1986,N_1967);
nor U2216 (N_2216,N_1875,N_1807);
xor U2217 (N_2217,N_1822,N_1922);
or U2218 (N_2218,N_1758,N_1989);
xor U2219 (N_2219,N_1961,N_1819);
or U2220 (N_2220,N_1777,N_1912);
and U2221 (N_2221,N_1961,N_1945);
or U2222 (N_2222,N_1953,N_1834);
or U2223 (N_2223,N_1961,N_1866);
and U2224 (N_2224,N_1959,N_1810);
or U2225 (N_2225,N_1986,N_1956);
nand U2226 (N_2226,N_1967,N_1990);
and U2227 (N_2227,N_1818,N_1782);
nor U2228 (N_2228,N_1792,N_1981);
xor U2229 (N_2229,N_1982,N_1974);
xor U2230 (N_2230,N_1834,N_1840);
nand U2231 (N_2231,N_1877,N_1994);
and U2232 (N_2232,N_1806,N_1768);
xor U2233 (N_2233,N_1944,N_1959);
nand U2234 (N_2234,N_1846,N_1849);
and U2235 (N_2235,N_1865,N_1887);
xor U2236 (N_2236,N_1892,N_1973);
nand U2237 (N_2237,N_1936,N_1833);
or U2238 (N_2238,N_1971,N_1786);
and U2239 (N_2239,N_1855,N_1965);
and U2240 (N_2240,N_1894,N_1890);
nor U2241 (N_2241,N_1788,N_1889);
xor U2242 (N_2242,N_1948,N_1944);
nor U2243 (N_2243,N_1969,N_1915);
and U2244 (N_2244,N_1817,N_1752);
nor U2245 (N_2245,N_1905,N_1911);
or U2246 (N_2246,N_1911,N_1826);
nor U2247 (N_2247,N_1854,N_1921);
and U2248 (N_2248,N_1775,N_1893);
and U2249 (N_2249,N_1957,N_1994);
nor U2250 (N_2250,N_2152,N_2098);
xor U2251 (N_2251,N_2001,N_2208);
nor U2252 (N_2252,N_2084,N_2223);
nor U2253 (N_2253,N_2027,N_2034);
or U2254 (N_2254,N_2144,N_2184);
or U2255 (N_2255,N_2062,N_2042);
nand U2256 (N_2256,N_2224,N_2159);
xor U2257 (N_2257,N_2226,N_2036);
xnor U2258 (N_2258,N_2164,N_2232);
nand U2259 (N_2259,N_2217,N_2123);
nand U2260 (N_2260,N_2017,N_2068);
and U2261 (N_2261,N_2190,N_2227);
xor U2262 (N_2262,N_2135,N_2048);
nor U2263 (N_2263,N_2120,N_2161);
nand U2264 (N_2264,N_2012,N_2213);
or U2265 (N_2265,N_2193,N_2032);
nand U2266 (N_2266,N_2040,N_2009);
xnor U2267 (N_2267,N_2006,N_2245);
xor U2268 (N_2268,N_2127,N_2172);
xor U2269 (N_2269,N_2030,N_2011);
nand U2270 (N_2270,N_2079,N_2129);
and U2271 (N_2271,N_2216,N_2151);
nand U2272 (N_2272,N_2138,N_2233);
nor U2273 (N_2273,N_2142,N_2115);
nand U2274 (N_2274,N_2178,N_2220);
and U2275 (N_2275,N_2039,N_2185);
xnor U2276 (N_2276,N_2015,N_2195);
nand U2277 (N_2277,N_2225,N_2108);
or U2278 (N_2278,N_2126,N_2075);
nand U2279 (N_2279,N_2202,N_2081);
xor U2280 (N_2280,N_2106,N_2206);
or U2281 (N_2281,N_2072,N_2066);
and U2282 (N_2282,N_2189,N_2182);
or U2283 (N_2283,N_2124,N_2136);
or U2284 (N_2284,N_2071,N_2181);
xnor U2285 (N_2285,N_2060,N_2035);
xnor U2286 (N_2286,N_2024,N_2014);
nor U2287 (N_2287,N_2078,N_2050);
and U2288 (N_2288,N_2004,N_2209);
and U2289 (N_2289,N_2241,N_2218);
xor U2290 (N_2290,N_2038,N_2114);
and U2291 (N_2291,N_2155,N_2061);
nor U2292 (N_2292,N_2237,N_2097);
and U2293 (N_2293,N_2148,N_2064);
nor U2294 (N_2294,N_2083,N_2179);
nor U2295 (N_2295,N_2057,N_2021);
xor U2296 (N_2296,N_2246,N_2247);
nor U2297 (N_2297,N_2105,N_2243);
or U2298 (N_2298,N_2101,N_2240);
nor U2299 (N_2299,N_2049,N_2067);
xor U2300 (N_2300,N_2054,N_2056);
xor U2301 (N_2301,N_2249,N_2139);
nor U2302 (N_2302,N_2150,N_2191);
nand U2303 (N_2303,N_2082,N_2230);
or U2304 (N_2304,N_2134,N_2010);
and U2305 (N_2305,N_2215,N_2053);
nor U2306 (N_2306,N_2204,N_2087);
xnor U2307 (N_2307,N_2186,N_2093);
xor U2308 (N_2308,N_2007,N_2154);
xnor U2309 (N_2309,N_2005,N_2211);
xor U2310 (N_2310,N_2052,N_2096);
nand U2311 (N_2311,N_2132,N_2166);
and U2312 (N_2312,N_2045,N_2163);
and U2313 (N_2313,N_2137,N_2095);
nand U2314 (N_2314,N_2175,N_2133);
or U2315 (N_2315,N_2194,N_2157);
nor U2316 (N_2316,N_2167,N_2031);
nor U2317 (N_2317,N_2125,N_2076);
nand U2318 (N_2318,N_2090,N_2002);
nor U2319 (N_2319,N_2140,N_2029);
and U2320 (N_2320,N_2171,N_2234);
nor U2321 (N_2321,N_2146,N_2188);
nor U2322 (N_2322,N_2055,N_2174);
nand U2323 (N_2323,N_2153,N_2228);
xor U2324 (N_2324,N_2173,N_2122);
nand U2325 (N_2325,N_2210,N_2168);
nor U2326 (N_2326,N_2200,N_2117);
and U2327 (N_2327,N_2089,N_2019);
nor U2328 (N_2328,N_2201,N_2110);
nor U2329 (N_2329,N_2116,N_2205);
and U2330 (N_2330,N_2121,N_2149);
xnor U2331 (N_2331,N_2197,N_2069);
xnor U2332 (N_2332,N_2219,N_2239);
nand U2333 (N_2333,N_2088,N_2203);
and U2334 (N_2334,N_2091,N_2085);
xor U2335 (N_2335,N_2199,N_2016);
xnor U2336 (N_2336,N_2063,N_2196);
xor U2337 (N_2337,N_2099,N_2086);
xnor U2338 (N_2338,N_2242,N_2180);
nand U2339 (N_2339,N_2109,N_2162);
nand U2340 (N_2340,N_2131,N_2103);
and U2341 (N_2341,N_2118,N_2013);
nor U2342 (N_2342,N_2028,N_2187);
xor U2343 (N_2343,N_2207,N_2047);
nor U2344 (N_2344,N_2065,N_2119);
or U2345 (N_2345,N_2183,N_2192);
xor U2346 (N_2346,N_2222,N_2018);
or U2347 (N_2347,N_2165,N_2022);
and U2348 (N_2348,N_2170,N_2158);
nand U2349 (N_2349,N_2111,N_2059);
or U2350 (N_2350,N_2198,N_2169);
nor U2351 (N_2351,N_2244,N_2145);
nand U2352 (N_2352,N_2104,N_2043);
nand U2353 (N_2353,N_2044,N_2026);
xnor U2354 (N_2354,N_2023,N_2008);
or U2355 (N_2355,N_2229,N_2177);
or U2356 (N_2356,N_2214,N_2147);
or U2357 (N_2357,N_2046,N_2130);
nor U2358 (N_2358,N_2235,N_2160);
or U2359 (N_2359,N_2020,N_2212);
and U2360 (N_2360,N_2074,N_2037);
nand U2361 (N_2361,N_2100,N_2238);
nor U2362 (N_2362,N_2176,N_2221);
nand U2363 (N_2363,N_2128,N_2112);
and U2364 (N_2364,N_2102,N_2156);
or U2365 (N_2365,N_2033,N_2070);
xor U2366 (N_2366,N_2236,N_2113);
and U2367 (N_2367,N_2003,N_2041);
nor U2368 (N_2368,N_2025,N_2077);
xnor U2369 (N_2369,N_2141,N_2092);
nand U2370 (N_2370,N_2073,N_2051);
nor U2371 (N_2371,N_2080,N_2000);
nand U2372 (N_2372,N_2248,N_2143);
xnor U2373 (N_2373,N_2107,N_2058);
xnor U2374 (N_2374,N_2231,N_2094);
and U2375 (N_2375,N_2201,N_2140);
nor U2376 (N_2376,N_2117,N_2246);
nor U2377 (N_2377,N_2102,N_2138);
and U2378 (N_2378,N_2239,N_2102);
nor U2379 (N_2379,N_2090,N_2235);
xor U2380 (N_2380,N_2221,N_2070);
or U2381 (N_2381,N_2126,N_2180);
nand U2382 (N_2382,N_2053,N_2192);
or U2383 (N_2383,N_2094,N_2051);
and U2384 (N_2384,N_2039,N_2013);
nor U2385 (N_2385,N_2247,N_2131);
nor U2386 (N_2386,N_2182,N_2229);
nand U2387 (N_2387,N_2100,N_2137);
nor U2388 (N_2388,N_2117,N_2176);
nand U2389 (N_2389,N_2117,N_2039);
or U2390 (N_2390,N_2155,N_2015);
and U2391 (N_2391,N_2125,N_2095);
nand U2392 (N_2392,N_2005,N_2012);
or U2393 (N_2393,N_2186,N_2234);
nor U2394 (N_2394,N_2242,N_2165);
or U2395 (N_2395,N_2147,N_2240);
nand U2396 (N_2396,N_2164,N_2182);
and U2397 (N_2397,N_2069,N_2083);
xnor U2398 (N_2398,N_2027,N_2061);
and U2399 (N_2399,N_2009,N_2041);
xnor U2400 (N_2400,N_2113,N_2215);
xor U2401 (N_2401,N_2244,N_2200);
xor U2402 (N_2402,N_2135,N_2014);
xor U2403 (N_2403,N_2242,N_2059);
nand U2404 (N_2404,N_2176,N_2046);
nand U2405 (N_2405,N_2065,N_2243);
nand U2406 (N_2406,N_2074,N_2026);
and U2407 (N_2407,N_2125,N_2109);
and U2408 (N_2408,N_2155,N_2125);
nand U2409 (N_2409,N_2000,N_2247);
nand U2410 (N_2410,N_2233,N_2089);
nand U2411 (N_2411,N_2024,N_2243);
and U2412 (N_2412,N_2046,N_2105);
and U2413 (N_2413,N_2223,N_2234);
nand U2414 (N_2414,N_2143,N_2064);
and U2415 (N_2415,N_2224,N_2115);
and U2416 (N_2416,N_2206,N_2246);
xor U2417 (N_2417,N_2027,N_2224);
and U2418 (N_2418,N_2161,N_2249);
nand U2419 (N_2419,N_2137,N_2115);
xnor U2420 (N_2420,N_2051,N_2151);
nor U2421 (N_2421,N_2185,N_2108);
nor U2422 (N_2422,N_2037,N_2161);
nor U2423 (N_2423,N_2130,N_2105);
nor U2424 (N_2424,N_2078,N_2219);
and U2425 (N_2425,N_2231,N_2247);
nand U2426 (N_2426,N_2150,N_2017);
and U2427 (N_2427,N_2178,N_2118);
nand U2428 (N_2428,N_2007,N_2012);
or U2429 (N_2429,N_2055,N_2073);
and U2430 (N_2430,N_2183,N_2165);
nor U2431 (N_2431,N_2032,N_2072);
nor U2432 (N_2432,N_2002,N_2000);
or U2433 (N_2433,N_2035,N_2007);
nor U2434 (N_2434,N_2169,N_2099);
or U2435 (N_2435,N_2024,N_2210);
nor U2436 (N_2436,N_2129,N_2203);
xor U2437 (N_2437,N_2211,N_2191);
nor U2438 (N_2438,N_2234,N_2196);
xnor U2439 (N_2439,N_2238,N_2140);
nor U2440 (N_2440,N_2100,N_2244);
xor U2441 (N_2441,N_2077,N_2011);
xor U2442 (N_2442,N_2016,N_2197);
nor U2443 (N_2443,N_2028,N_2057);
nor U2444 (N_2444,N_2121,N_2226);
nor U2445 (N_2445,N_2134,N_2067);
nor U2446 (N_2446,N_2043,N_2188);
nand U2447 (N_2447,N_2199,N_2185);
and U2448 (N_2448,N_2144,N_2085);
xor U2449 (N_2449,N_2185,N_2043);
xor U2450 (N_2450,N_2058,N_2040);
nand U2451 (N_2451,N_2149,N_2019);
nand U2452 (N_2452,N_2079,N_2112);
and U2453 (N_2453,N_2184,N_2004);
and U2454 (N_2454,N_2073,N_2019);
nand U2455 (N_2455,N_2139,N_2154);
nand U2456 (N_2456,N_2048,N_2010);
and U2457 (N_2457,N_2216,N_2157);
or U2458 (N_2458,N_2025,N_2000);
and U2459 (N_2459,N_2039,N_2103);
xor U2460 (N_2460,N_2002,N_2143);
nand U2461 (N_2461,N_2158,N_2013);
and U2462 (N_2462,N_2195,N_2173);
nor U2463 (N_2463,N_2197,N_2012);
or U2464 (N_2464,N_2031,N_2091);
or U2465 (N_2465,N_2069,N_2092);
or U2466 (N_2466,N_2141,N_2135);
or U2467 (N_2467,N_2016,N_2027);
nor U2468 (N_2468,N_2037,N_2140);
nor U2469 (N_2469,N_2071,N_2167);
and U2470 (N_2470,N_2144,N_2149);
nand U2471 (N_2471,N_2045,N_2006);
and U2472 (N_2472,N_2197,N_2169);
and U2473 (N_2473,N_2197,N_2129);
or U2474 (N_2474,N_2058,N_2217);
or U2475 (N_2475,N_2073,N_2211);
nor U2476 (N_2476,N_2047,N_2059);
nand U2477 (N_2477,N_2052,N_2042);
nand U2478 (N_2478,N_2047,N_2100);
nor U2479 (N_2479,N_2122,N_2240);
xor U2480 (N_2480,N_2221,N_2095);
nor U2481 (N_2481,N_2077,N_2159);
nand U2482 (N_2482,N_2037,N_2201);
nor U2483 (N_2483,N_2183,N_2071);
nor U2484 (N_2484,N_2058,N_2056);
nor U2485 (N_2485,N_2045,N_2064);
or U2486 (N_2486,N_2056,N_2247);
and U2487 (N_2487,N_2202,N_2042);
nand U2488 (N_2488,N_2136,N_2180);
xor U2489 (N_2489,N_2168,N_2113);
xor U2490 (N_2490,N_2069,N_2143);
nor U2491 (N_2491,N_2004,N_2096);
nand U2492 (N_2492,N_2152,N_2126);
xor U2493 (N_2493,N_2012,N_2225);
or U2494 (N_2494,N_2117,N_2173);
nand U2495 (N_2495,N_2068,N_2191);
xor U2496 (N_2496,N_2186,N_2068);
and U2497 (N_2497,N_2159,N_2217);
nand U2498 (N_2498,N_2208,N_2227);
or U2499 (N_2499,N_2156,N_2197);
or U2500 (N_2500,N_2421,N_2300);
xnor U2501 (N_2501,N_2262,N_2457);
and U2502 (N_2502,N_2385,N_2437);
nor U2503 (N_2503,N_2287,N_2475);
xnor U2504 (N_2504,N_2261,N_2402);
and U2505 (N_2505,N_2382,N_2363);
nor U2506 (N_2506,N_2389,N_2391);
nor U2507 (N_2507,N_2376,N_2408);
or U2508 (N_2508,N_2289,N_2304);
xnor U2509 (N_2509,N_2463,N_2340);
and U2510 (N_2510,N_2331,N_2336);
and U2511 (N_2511,N_2252,N_2413);
or U2512 (N_2512,N_2430,N_2405);
nand U2513 (N_2513,N_2418,N_2316);
or U2514 (N_2514,N_2293,N_2444);
xnor U2515 (N_2515,N_2335,N_2360);
xnor U2516 (N_2516,N_2428,N_2443);
xnor U2517 (N_2517,N_2283,N_2373);
and U2518 (N_2518,N_2411,N_2407);
nor U2519 (N_2519,N_2260,N_2442);
or U2520 (N_2520,N_2352,N_2476);
or U2521 (N_2521,N_2267,N_2447);
nand U2522 (N_2522,N_2270,N_2333);
nand U2523 (N_2523,N_2455,N_2327);
nor U2524 (N_2524,N_2341,N_2461);
and U2525 (N_2525,N_2364,N_2257);
or U2526 (N_2526,N_2375,N_2349);
or U2527 (N_2527,N_2435,N_2434);
nor U2528 (N_2528,N_2305,N_2296);
and U2529 (N_2529,N_2273,N_2308);
nand U2530 (N_2530,N_2483,N_2351);
or U2531 (N_2531,N_2330,N_2344);
nand U2532 (N_2532,N_2431,N_2275);
xor U2533 (N_2533,N_2496,N_2282);
or U2534 (N_2534,N_2271,N_2387);
and U2535 (N_2535,N_2479,N_2350);
nand U2536 (N_2536,N_2306,N_2436);
nand U2537 (N_2537,N_2315,N_2301);
and U2538 (N_2538,N_2494,N_2460);
xor U2539 (N_2539,N_2386,N_2313);
and U2540 (N_2540,N_2467,N_2397);
nand U2541 (N_2541,N_2338,N_2464);
or U2542 (N_2542,N_2481,N_2498);
and U2543 (N_2543,N_2365,N_2297);
and U2544 (N_2544,N_2474,N_2319);
or U2545 (N_2545,N_2497,N_2491);
or U2546 (N_2546,N_2379,N_2450);
or U2547 (N_2547,N_2312,N_2309);
and U2548 (N_2548,N_2265,N_2291);
nor U2549 (N_2549,N_2290,N_2406);
and U2550 (N_2550,N_2310,N_2369);
and U2551 (N_2551,N_2318,N_2342);
nor U2552 (N_2552,N_2356,N_2445);
nor U2553 (N_2553,N_2307,N_2250);
or U2554 (N_2554,N_2264,N_2394);
or U2555 (N_2555,N_2285,N_2414);
nand U2556 (N_2556,N_2492,N_2393);
nor U2557 (N_2557,N_2490,N_2347);
and U2558 (N_2558,N_2371,N_2272);
or U2559 (N_2559,N_2343,N_2355);
nand U2560 (N_2560,N_2328,N_2326);
nor U2561 (N_2561,N_2357,N_2302);
nor U2562 (N_2562,N_2398,N_2468);
xnor U2563 (N_2563,N_2322,N_2495);
xor U2564 (N_2564,N_2303,N_2256);
and U2565 (N_2565,N_2324,N_2419);
and U2566 (N_2566,N_2339,N_2493);
or U2567 (N_2567,N_2484,N_2459);
nand U2568 (N_2568,N_2451,N_2359);
and U2569 (N_2569,N_2294,N_2456);
xnor U2570 (N_2570,N_2337,N_2288);
and U2571 (N_2571,N_2281,N_2254);
nand U2572 (N_2572,N_2346,N_2486);
and U2573 (N_2573,N_2284,N_2478);
nand U2574 (N_2574,N_2329,N_2390);
or U2575 (N_2575,N_2269,N_2427);
xor U2576 (N_2576,N_2489,N_2470);
nor U2577 (N_2577,N_2263,N_2392);
or U2578 (N_2578,N_2404,N_2417);
or U2579 (N_2579,N_2440,N_2278);
xor U2580 (N_2580,N_2454,N_2266);
nor U2581 (N_2581,N_2368,N_2251);
or U2582 (N_2582,N_2433,N_2345);
nor U2583 (N_2583,N_2401,N_2311);
and U2584 (N_2584,N_2465,N_2426);
and U2585 (N_2585,N_2448,N_2416);
xor U2586 (N_2586,N_2292,N_2258);
or U2587 (N_2587,N_2314,N_2362);
or U2588 (N_2588,N_2370,N_2466);
and U2589 (N_2589,N_2323,N_2432);
and U2590 (N_2590,N_2499,N_2449);
xor U2591 (N_2591,N_2480,N_2268);
and U2592 (N_2592,N_2395,N_2353);
nand U2593 (N_2593,N_2399,N_2274);
and U2594 (N_2594,N_2400,N_2423);
and U2595 (N_2595,N_2299,N_2381);
nor U2596 (N_2596,N_2280,N_2334);
xor U2597 (N_2597,N_2403,N_2380);
nand U2598 (N_2598,N_2425,N_2453);
and U2599 (N_2599,N_2488,N_2422);
xor U2600 (N_2600,N_2320,N_2361);
and U2601 (N_2601,N_2358,N_2366);
nor U2602 (N_2602,N_2259,N_2429);
nand U2603 (N_2603,N_2458,N_2438);
nor U2604 (N_2604,N_2462,N_2482);
or U2605 (N_2605,N_2253,N_2348);
and U2606 (N_2606,N_2279,N_2412);
or U2607 (N_2607,N_2396,N_2298);
nor U2608 (N_2608,N_2255,N_2477);
or U2609 (N_2609,N_2410,N_2469);
nor U2610 (N_2610,N_2471,N_2487);
nand U2611 (N_2611,N_2485,N_2276);
nor U2612 (N_2612,N_2317,N_2295);
nor U2613 (N_2613,N_2374,N_2415);
nor U2614 (N_2614,N_2388,N_2409);
nand U2615 (N_2615,N_2277,N_2325);
nand U2616 (N_2616,N_2424,N_2473);
nor U2617 (N_2617,N_2332,N_2321);
nand U2618 (N_2618,N_2377,N_2446);
nor U2619 (N_2619,N_2354,N_2384);
xor U2620 (N_2620,N_2452,N_2441);
nor U2621 (N_2621,N_2420,N_2372);
nor U2622 (N_2622,N_2378,N_2367);
nor U2623 (N_2623,N_2286,N_2472);
xnor U2624 (N_2624,N_2439,N_2383);
nand U2625 (N_2625,N_2424,N_2353);
nand U2626 (N_2626,N_2416,N_2397);
or U2627 (N_2627,N_2262,N_2411);
xor U2628 (N_2628,N_2252,N_2457);
xnor U2629 (N_2629,N_2422,N_2438);
and U2630 (N_2630,N_2422,N_2270);
xor U2631 (N_2631,N_2470,N_2490);
or U2632 (N_2632,N_2362,N_2379);
xnor U2633 (N_2633,N_2484,N_2279);
and U2634 (N_2634,N_2370,N_2440);
xor U2635 (N_2635,N_2499,N_2481);
or U2636 (N_2636,N_2356,N_2276);
nand U2637 (N_2637,N_2381,N_2366);
nor U2638 (N_2638,N_2446,N_2423);
nand U2639 (N_2639,N_2403,N_2348);
nor U2640 (N_2640,N_2269,N_2314);
xnor U2641 (N_2641,N_2277,N_2414);
xnor U2642 (N_2642,N_2295,N_2479);
xnor U2643 (N_2643,N_2337,N_2369);
nand U2644 (N_2644,N_2355,N_2379);
and U2645 (N_2645,N_2354,N_2396);
and U2646 (N_2646,N_2408,N_2323);
nor U2647 (N_2647,N_2396,N_2364);
or U2648 (N_2648,N_2462,N_2281);
or U2649 (N_2649,N_2355,N_2255);
or U2650 (N_2650,N_2450,N_2472);
and U2651 (N_2651,N_2396,N_2474);
nor U2652 (N_2652,N_2299,N_2441);
nor U2653 (N_2653,N_2420,N_2278);
nand U2654 (N_2654,N_2291,N_2306);
xnor U2655 (N_2655,N_2336,N_2357);
or U2656 (N_2656,N_2418,N_2288);
or U2657 (N_2657,N_2380,N_2357);
nand U2658 (N_2658,N_2369,N_2309);
xor U2659 (N_2659,N_2268,N_2328);
nand U2660 (N_2660,N_2341,N_2406);
and U2661 (N_2661,N_2283,N_2450);
nand U2662 (N_2662,N_2476,N_2270);
or U2663 (N_2663,N_2366,N_2280);
xor U2664 (N_2664,N_2443,N_2466);
xnor U2665 (N_2665,N_2305,N_2261);
and U2666 (N_2666,N_2336,N_2473);
or U2667 (N_2667,N_2458,N_2481);
nand U2668 (N_2668,N_2267,N_2496);
and U2669 (N_2669,N_2264,N_2377);
and U2670 (N_2670,N_2398,N_2481);
xnor U2671 (N_2671,N_2271,N_2395);
nand U2672 (N_2672,N_2455,N_2343);
xnor U2673 (N_2673,N_2414,N_2439);
and U2674 (N_2674,N_2294,N_2305);
or U2675 (N_2675,N_2422,N_2449);
and U2676 (N_2676,N_2413,N_2474);
or U2677 (N_2677,N_2328,N_2320);
xnor U2678 (N_2678,N_2385,N_2393);
xnor U2679 (N_2679,N_2284,N_2394);
and U2680 (N_2680,N_2396,N_2336);
or U2681 (N_2681,N_2479,N_2374);
or U2682 (N_2682,N_2485,N_2402);
nand U2683 (N_2683,N_2427,N_2461);
or U2684 (N_2684,N_2313,N_2250);
nand U2685 (N_2685,N_2417,N_2483);
and U2686 (N_2686,N_2381,N_2405);
xnor U2687 (N_2687,N_2441,N_2454);
or U2688 (N_2688,N_2436,N_2325);
or U2689 (N_2689,N_2396,N_2401);
or U2690 (N_2690,N_2467,N_2281);
and U2691 (N_2691,N_2251,N_2385);
or U2692 (N_2692,N_2431,N_2408);
nand U2693 (N_2693,N_2262,N_2281);
nor U2694 (N_2694,N_2356,N_2254);
nand U2695 (N_2695,N_2408,N_2421);
or U2696 (N_2696,N_2294,N_2381);
and U2697 (N_2697,N_2361,N_2371);
xnor U2698 (N_2698,N_2290,N_2468);
nor U2699 (N_2699,N_2362,N_2357);
nand U2700 (N_2700,N_2409,N_2436);
nand U2701 (N_2701,N_2261,N_2374);
or U2702 (N_2702,N_2447,N_2493);
or U2703 (N_2703,N_2276,N_2320);
xor U2704 (N_2704,N_2335,N_2268);
xnor U2705 (N_2705,N_2358,N_2313);
and U2706 (N_2706,N_2469,N_2400);
and U2707 (N_2707,N_2464,N_2493);
xnor U2708 (N_2708,N_2283,N_2410);
nor U2709 (N_2709,N_2317,N_2412);
nand U2710 (N_2710,N_2493,N_2351);
xor U2711 (N_2711,N_2353,N_2382);
and U2712 (N_2712,N_2426,N_2357);
nand U2713 (N_2713,N_2433,N_2395);
nor U2714 (N_2714,N_2423,N_2310);
and U2715 (N_2715,N_2456,N_2437);
nand U2716 (N_2716,N_2275,N_2419);
nor U2717 (N_2717,N_2290,N_2278);
xor U2718 (N_2718,N_2339,N_2439);
xor U2719 (N_2719,N_2451,N_2477);
and U2720 (N_2720,N_2427,N_2446);
nor U2721 (N_2721,N_2346,N_2272);
and U2722 (N_2722,N_2272,N_2468);
and U2723 (N_2723,N_2348,N_2462);
or U2724 (N_2724,N_2421,N_2382);
nor U2725 (N_2725,N_2350,N_2358);
xnor U2726 (N_2726,N_2272,N_2268);
xnor U2727 (N_2727,N_2466,N_2299);
nand U2728 (N_2728,N_2382,N_2444);
and U2729 (N_2729,N_2424,N_2289);
nor U2730 (N_2730,N_2490,N_2328);
or U2731 (N_2731,N_2422,N_2337);
nor U2732 (N_2732,N_2372,N_2307);
and U2733 (N_2733,N_2414,N_2454);
nor U2734 (N_2734,N_2440,N_2455);
xor U2735 (N_2735,N_2330,N_2292);
or U2736 (N_2736,N_2316,N_2411);
nor U2737 (N_2737,N_2389,N_2385);
and U2738 (N_2738,N_2413,N_2346);
and U2739 (N_2739,N_2419,N_2293);
and U2740 (N_2740,N_2421,N_2480);
or U2741 (N_2741,N_2380,N_2279);
nand U2742 (N_2742,N_2261,N_2264);
or U2743 (N_2743,N_2302,N_2434);
nor U2744 (N_2744,N_2283,N_2306);
nor U2745 (N_2745,N_2490,N_2437);
and U2746 (N_2746,N_2264,N_2294);
nor U2747 (N_2747,N_2416,N_2486);
xnor U2748 (N_2748,N_2464,N_2360);
or U2749 (N_2749,N_2254,N_2463);
and U2750 (N_2750,N_2711,N_2723);
nand U2751 (N_2751,N_2570,N_2636);
nor U2752 (N_2752,N_2568,N_2676);
or U2753 (N_2753,N_2655,N_2733);
nor U2754 (N_2754,N_2542,N_2567);
nor U2755 (N_2755,N_2700,N_2574);
or U2756 (N_2756,N_2521,N_2526);
or U2757 (N_2757,N_2531,N_2598);
nor U2758 (N_2758,N_2675,N_2706);
nor U2759 (N_2759,N_2619,N_2522);
and U2760 (N_2760,N_2569,N_2688);
or U2761 (N_2761,N_2566,N_2629);
and U2762 (N_2762,N_2677,N_2687);
xor U2763 (N_2763,N_2633,N_2565);
nand U2764 (N_2764,N_2593,N_2620);
nand U2765 (N_2765,N_2614,N_2735);
and U2766 (N_2766,N_2651,N_2606);
nor U2767 (N_2767,N_2518,N_2690);
or U2768 (N_2768,N_2670,N_2539);
or U2769 (N_2769,N_2552,N_2635);
nor U2770 (N_2770,N_2543,N_2685);
nand U2771 (N_2771,N_2587,N_2578);
and U2772 (N_2772,N_2680,N_2624);
or U2773 (N_2773,N_2725,N_2746);
and U2774 (N_2774,N_2645,N_2715);
nand U2775 (N_2775,N_2638,N_2729);
xnor U2776 (N_2776,N_2724,N_2601);
and U2777 (N_2777,N_2741,N_2692);
and U2778 (N_2778,N_2513,N_2653);
nor U2779 (N_2779,N_2661,N_2643);
or U2780 (N_2780,N_2644,N_2699);
and U2781 (N_2781,N_2622,N_2730);
and U2782 (N_2782,N_2697,N_2748);
and U2783 (N_2783,N_2667,N_2659);
nor U2784 (N_2784,N_2732,N_2671);
or U2785 (N_2785,N_2535,N_2580);
xor U2786 (N_2786,N_2538,N_2616);
and U2787 (N_2787,N_2689,N_2737);
and U2788 (N_2788,N_2739,N_2610);
xor U2789 (N_2789,N_2602,N_2517);
xnor U2790 (N_2790,N_2743,N_2533);
xor U2791 (N_2791,N_2684,N_2586);
or U2792 (N_2792,N_2530,N_2681);
and U2793 (N_2793,N_2537,N_2704);
nand U2794 (N_2794,N_2731,N_2658);
nor U2795 (N_2795,N_2703,N_2506);
or U2796 (N_2796,N_2716,N_2525);
or U2797 (N_2797,N_2632,N_2502);
xor U2798 (N_2798,N_2654,N_2665);
or U2799 (N_2799,N_2612,N_2548);
or U2800 (N_2800,N_2503,N_2701);
and U2801 (N_2801,N_2603,N_2590);
nor U2802 (N_2802,N_2696,N_2510);
nor U2803 (N_2803,N_2617,N_2718);
or U2804 (N_2804,N_2634,N_2507);
nor U2805 (N_2805,N_2694,N_2550);
and U2806 (N_2806,N_2597,N_2747);
xnor U2807 (N_2807,N_2693,N_2556);
xnor U2808 (N_2808,N_2663,N_2583);
xor U2809 (N_2809,N_2664,N_2674);
xnor U2810 (N_2810,N_2501,N_2734);
or U2811 (N_2811,N_2563,N_2541);
nand U2812 (N_2812,N_2599,N_2744);
xnor U2813 (N_2813,N_2631,N_2719);
xor U2814 (N_2814,N_2536,N_2666);
nor U2815 (N_2815,N_2547,N_2554);
xor U2816 (N_2816,N_2560,N_2577);
xnor U2817 (N_2817,N_2551,N_2717);
nor U2818 (N_2818,N_2649,N_2740);
or U2819 (N_2819,N_2630,N_2613);
and U2820 (N_2820,N_2527,N_2709);
xnor U2821 (N_2821,N_2600,N_2596);
xnor U2822 (N_2822,N_2673,N_2691);
and U2823 (N_2823,N_2575,N_2608);
or U2824 (N_2824,N_2648,N_2558);
nor U2825 (N_2825,N_2529,N_2652);
or U2826 (N_2826,N_2628,N_2572);
xor U2827 (N_2827,N_2686,N_2656);
nand U2828 (N_2828,N_2545,N_2534);
xor U2829 (N_2829,N_2520,N_2720);
nor U2830 (N_2830,N_2657,N_2627);
xor U2831 (N_2831,N_2509,N_2504);
and U2832 (N_2832,N_2579,N_2607);
xnor U2833 (N_2833,N_2708,N_2705);
nand U2834 (N_2834,N_2557,N_2738);
nor U2835 (N_2835,N_2515,N_2588);
xor U2836 (N_2836,N_2742,N_2721);
or U2837 (N_2837,N_2508,N_2516);
or U2838 (N_2838,N_2562,N_2555);
and U2839 (N_2839,N_2609,N_2668);
xnor U2840 (N_2840,N_2710,N_2546);
or U2841 (N_2841,N_2559,N_2500);
xor U2842 (N_2842,N_2745,N_2637);
nand U2843 (N_2843,N_2561,N_2736);
or U2844 (N_2844,N_2726,N_2611);
xnor U2845 (N_2845,N_2591,N_2695);
nor U2846 (N_2846,N_2514,N_2511);
and U2847 (N_2847,N_2576,N_2679);
or U2848 (N_2848,N_2528,N_2519);
xnor U2849 (N_2849,N_2714,N_2589);
xnor U2850 (N_2850,N_2582,N_2683);
or U2851 (N_2851,N_2553,N_2728);
nand U2852 (N_2852,N_2604,N_2650);
or U2853 (N_2853,N_2571,N_2641);
xor U2854 (N_2854,N_2669,N_2640);
nand U2855 (N_2855,N_2615,N_2698);
or U2856 (N_2856,N_2581,N_2505);
or U2857 (N_2857,N_2512,N_2660);
nor U2858 (N_2858,N_2749,N_2639);
and U2859 (N_2859,N_2592,N_2625);
or U2860 (N_2860,N_2712,N_2702);
and U2861 (N_2861,N_2707,N_2524);
nand U2862 (N_2862,N_2626,N_2618);
and U2863 (N_2863,N_2584,N_2564);
nor U2864 (N_2864,N_2722,N_2544);
or U2865 (N_2865,N_2540,N_2621);
nor U2866 (N_2866,N_2523,N_2585);
xnor U2867 (N_2867,N_2642,N_2623);
nand U2868 (N_2868,N_2727,N_2672);
nor U2869 (N_2869,N_2682,N_2713);
and U2870 (N_2870,N_2678,N_2573);
nor U2871 (N_2871,N_2549,N_2532);
nor U2872 (N_2872,N_2662,N_2647);
and U2873 (N_2873,N_2594,N_2605);
xor U2874 (N_2874,N_2646,N_2595);
xor U2875 (N_2875,N_2649,N_2639);
nand U2876 (N_2876,N_2586,N_2507);
and U2877 (N_2877,N_2705,N_2704);
xor U2878 (N_2878,N_2615,N_2687);
and U2879 (N_2879,N_2651,N_2556);
nand U2880 (N_2880,N_2659,N_2587);
nor U2881 (N_2881,N_2660,N_2676);
nor U2882 (N_2882,N_2730,N_2740);
and U2883 (N_2883,N_2525,N_2552);
nand U2884 (N_2884,N_2672,N_2631);
or U2885 (N_2885,N_2592,N_2648);
and U2886 (N_2886,N_2719,N_2706);
or U2887 (N_2887,N_2682,N_2603);
and U2888 (N_2888,N_2611,N_2604);
nand U2889 (N_2889,N_2727,N_2545);
nor U2890 (N_2890,N_2740,N_2684);
or U2891 (N_2891,N_2563,N_2678);
nor U2892 (N_2892,N_2517,N_2728);
and U2893 (N_2893,N_2533,N_2669);
nor U2894 (N_2894,N_2745,N_2513);
and U2895 (N_2895,N_2646,N_2697);
nor U2896 (N_2896,N_2671,N_2657);
and U2897 (N_2897,N_2720,N_2673);
xnor U2898 (N_2898,N_2639,N_2512);
nand U2899 (N_2899,N_2665,N_2747);
and U2900 (N_2900,N_2656,N_2689);
xor U2901 (N_2901,N_2672,N_2635);
nor U2902 (N_2902,N_2571,N_2651);
nor U2903 (N_2903,N_2710,N_2686);
nor U2904 (N_2904,N_2721,N_2549);
xnor U2905 (N_2905,N_2522,N_2539);
and U2906 (N_2906,N_2683,N_2668);
xnor U2907 (N_2907,N_2607,N_2569);
nand U2908 (N_2908,N_2543,N_2613);
and U2909 (N_2909,N_2705,N_2592);
nand U2910 (N_2910,N_2594,N_2642);
nor U2911 (N_2911,N_2730,N_2538);
nand U2912 (N_2912,N_2552,N_2638);
xor U2913 (N_2913,N_2650,N_2584);
or U2914 (N_2914,N_2734,N_2537);
nor U2915 (N_2915,N_2678,N_2700);
or U2916 (N_2916,N_2630,N_2692);
nor U2917 (N_2917,N_2656,N_2619);
and U2918 (N_2918,N_2640,N_2720);
or U2919 (N_2919,N_2731,N_2737);
nand U2920 (N_2920,N_2666,N_2604);
and U2921 (N_2921,N_2598,N_2518);
xnor U2922 (N_2922,N_2500,N_2625);
xnor U2923 (N_2923,N_2530,N_2551);
and U2924 (N_2924,N_2522,N_2609);
or U2925 (N_2925,N_2594,N_2659);
xor U2926 (N_2926,N_2732,N_2683);
nand U2927 (N_2927,N_2547,N_2711);
or U2928 (N_2928,N_2547,N_2697);
and U2929 (N_2929,N_2744,N_2603);
xor U2930 (N_2930,N_2521,N_2706);
xnor U2931 (N_2931,N_2608,N_2559);
nor U2932 (N_2932,N_2584,N_2745);
nand U2933 (N_2933,N_2621,N_2742);
or U2934 (N_2934,N_2629,N_2582);
or U2935 (N_2935,N_2744,N_2601);
nand U2936 (N_2936,N_2506,N_2705);
or U2937 (N_2937,N_2717,N_2559);
xnor U2938 (N_2938,N_2632,N_2692);
or U2939 (N_2939,N_2515,N_2643);
xor U2940 (N_2940,N_2570,N_2707);
or U2941 (N_2941,N_2567,N_2596);
or U2942 (N_2942,N_2590,N_2699);
nor U2943 (N_2943,N_2559,N_2558);
nand U2944 (N_2944,N_2701,N_2633);
nor U2945 (N_2945,N_2645,N_2548);
xor U2946 (N_2946,N_2581,N_2702);
nand U2947 (N_2947,N_2513,N_2544);
or U2948 (N_2948,N_2578,N_2525);
and U2949 (N_2949,N_2704,N_2531);
and U2950 (N_2950,N_2590,N_2672);
nand U2951 (N_2951,N_2593,N_2507);
nand U2952 (N_2952,N_2612,N_2558);
xor U2953 (N_2953,N_2539,N_2638);
or U2954 (N_2954,N_2740,N_2569);
xnor U2955 (N_2955,N_2655,N_2517);
nand U2956 (N_2956,N_2618,N_2592);
or U2957 (N_2957,N_2562,N_2638);
nor U2958 (N_2958,N_2732,N_2700);
nor U2959 (N_2959,N_2628,N_2504);
xor U2960 (N_2960,N_2677,N_2592);
nand U2961 (N_2961,N_2731,N_2571);
nor U2962 (N_2962,N_2739,N_2578);
nand U2963 (N_2963,N_2602,N_2589);
and U2964 (N_2964,N_2603,N_2584);
or U2965 (N_2965,N_2640,N_2631);
nand U2966 (N_2966,N_2738,N_2570);
nand U2967 (N_2967,N_2716,N_2591);
xnor U2968 (N_2968,N_2635,N_2603);
nand U2969 (N_2969,N_2521,N_2577);
or U2970 (N_2970,N_2748,N_2514);
nand U2971 (N_2971,N_2571,N_2676);
nand U2972 (N_2972,N_2547,N_2572);
and U2973 (N_2973,N_2660,N_2692);
nor U2974 (N_2974,N_2545,N_2657);
nor U2975 (N_2975,N_2661,N_2655);
nand U2976 (N_2976,N_2533,N_2694);
nand U2977 (N_2977,N_2674,N_2510);
and U2978 (N_2978,N_2567,N_2686);
xnor U2979 (N_2979,N_2573,N_2660);
and U2980 (N_2980,N_2629,N_2553);
xnor U2981 (N_2981,N_2523,N_2553);
or U2982 (N_2982,N_2621,N_2572);
or U2983 (N_2983,N_2570,N_2516);
and U2984 (N_2984,N_2660,N_2576);
nand U2985 (N_2985,N_2609,N_2538);
or U2986 (N_2986,N_2721,N_2613);
and U2987 (N_2987,N_2605,N_2740);
nand U2988 (N_2988,N_2543,N_2515);
or U2989 (N_2989,N_2557,N_2631);
nor U2990 (N_2990,N_2598,N_2672);
nand U2991 (N_2991,N_2708,N_2619);
nor U2992 (N_2992,N_2573,N_2700);
and U2993 (N_2993,N_2550,N_2647);
or U2994 (N_2994,N_2596,N_2717);
nor U2995 (N_2995,N_2692,N_2739);
or U2996 (N_2996,N_2676,N_2507);
nor U2997 (N_2997,N_2661,N_2674);
and U2998 (N_2998,N_2573,N_2501);
nor U2999 (N_2999,N_2548,N_2573);
and U3000 (N_3000,N_2762,N_2976);
xor U3001 (N_3001,N_2754,N_2949);
and U3002 (N_3002,N_2755,N_2975);
and U3003 (N_3003,N_2787,N_2788);
nor U3004 (N_3004,N_2981,N_2957);
or U3005 (N_3005,N_2992,N_2919);
nand U3006 (N_3006,N_2966,N_2878);
and U3007 (N_3007,N_2900,N_2931);
or U3008 (N_3008,N_2830,N_2780);
xor U3009 (N_3009,N_2790,N_2761);
nand U3010 (N_3010,N_2808,N_2978);
or U3011 (N_3011,N_2873,N_2820);
nor U3012 (N_3012,N_2853,N_2983);
or U3013 (N_3013,N_2980,N_2944);
nor U3014 (N_3014,N_2963,N_2926);
and U3015 (N_3015,N_2922,N_2940);
nor U3016 (N_3016,N_2929,N_2846);
nor U3017 (N_3017,N_2807,N_2860);
xor U3018 (N_3018,N_2866,N_2991);
nand U3019 (N_3019,N_2801,N_2799);
nor U3020 (N_3020,N_2819,N_2773);
xnor U3021 (N_3021,N_2893,N_2890);
or U3022 (N_3022,N_2947,N_2886);
or U3023 (N_3023,N_2998,N_2862);
nor U3024 (N_3024,N_2906,N_2815);
xnor U3025 (N_3025,N_2812,N_2937);
nor U3026 (N_3026,N_2833,N_2989);
nor U3027 (N_3027,N_2885,N_2876);
or U3028 (N_3028,N_2924,N_2954);
nand U3029 (N_3029,N_2797,N_2881);
and U3030 (N_3030,N_2987,N_2865);
nor U3031 (N_3031,N_2794,N_2945);
xnor U3032 (N_3032,N_2850,N_2891);
nor U3033 (N_3033,N_2879,N_2767);
or U3034 (N_3034,N_2803,N_2813);
or U3035 (N_3035,N_2889,N_2760);
xnor U3036 (N_3036,N_2848,N_2766);
xnor U3037 (N_3037,N_2858,N_2824);
nand U3038 (N_3038,N_2840,N_2851);
or U3039 (N_3039,N_2832,N_2888);
and U3040 (N_3040,N_2943,N_2805);
or U3041 (N_3041,N_2814,N_2923);
nor U3042 (N_3042,N_2796,N_2758);
nand U3043 (N_3043,N_2964,N_2776);
or U3044 (N_3044,N_2962,N_2938);
or U3045 (N_3045,N_2870,N_2806);
nand U3046 (N_3046,N_2939,N_2765);
or U3047 (N_3047,N_2951,N_2977);
nand U3048 (N_3048,N_2775,N_2751);
nor U3049 (N_3049,N_2872,N_2867);
nand U3050 (N_3050,N_2882,N_2871);
xor U3051 (N_3051,N_2838,N_2917);
nand U3052 (N_3052,N_2956,N_2918);
xnor U3053 (N_3053,N_2823,N_2800);
and U3054 (N_3054,N_2909,N_2817);
xor U3055 (N_3055,N_2974,N_2841);
or U3056 (N_3056,N_2948,N_2935);
nand U3057 (N_3057,N_2955,N_2880);
and U3058 (N_3058,N_2884,N_2971);
xor U3059 (N_3059,N_2856,N_2855);
and U3060 (N_3060,N_2868,N_2854);
nand U3061 (N_3061,N_2986,N_2941);
and U3062 (N_3062,N_2916,N_2783);
and U3063 (N_3063,N_2928,N_2839);
xor U3064 (N_3064,N_2912,N_2932);
nand U3065 (N_3065,N_2990,N_2844);
nand U3066 (N_3066,N_2960,N_2915);
or U3067 (N_3067,N_2750,N_2999);
nand U3068 (N_3068,N_2911,N_2898);
nand U3069 (N_3069,N_2894,N_2753);
xnor U3070 (N_3070,N_2786,N_2863);
nand U3071 (N_3071,N_2843,N_2784);
xor U3072 (N_3072,N_2864,N_2979);
xnor U3073 (N_3073,N_2959,N_2822);
nand U3074 (N_3074,N_2904,N_2973);
xnor U3075 (N_3075,N_2920,N_2849);
or U3076 (N_3076,N_2965,N_2804);
nor U3077 (N_3077,N_2791,N_2847);
nand U3078 (N_3078,N_2899,N_2925);
and U3079 (N_3079,N_2771,N_2969);
or U3080 (N_3080,N_2927,N_2835);
nor U3081 (N_3081,N_2967,N_2934);
xor U3082 (N_3082,N_2988,N_2792);
nor U3083 (N_3083,N_2892,N_2897);
or U3084 (N_3084,N_2908,N_2985);
nor U3085 (N_3085,N_2764,N_2914);
nand U3086 (N_3086,N_2811,N_2769);
and U3087 (N_3087,N_2845,N_2997);
nand U3088 (N_3088,N_2795,N_2829);
and U3089 (N_3089,N_2993,N_2996);
nand U3090 (N_3090,N_2756,N_2887);
or U3091 (N_3091,N_2902,N_2968);
nand U3092 (N_3092,N_2861,N_2802);
nand U3093 (N_3093,N_2982,N_2809);
xnor U3094 (N_3094,N_2852,N_2768);
or U3095 (N_3095,N_2793,N_2877);
nor U3096 (N_3096,N_2875,N_2905);
nor U3097 (N_3097,N_2936,N_2910);
xor U3098 (N_3098,N_2930,N_2946);
xnor U3099 (N_3099,N_2836,N_2810);
and U3100 (N_3100,N_2757,N_2831);
nand U3101 (N_3101,N_2907,N_2895);
or U3102 (N_3102,N_2933,N_2995);
and U3103 (N_3103,N_2842,N_2821);
nor U3104 (N_3104,N_2772,N_2785);
nor U3105 (N_3105,N_2874,N_2816);
xnor U3106 (N_3106,N_2798,N_2970);
nand U3107 (N_3107,N_2953,N_2921);
nand U3108 (N_3108,N_2781,N_2826);
nor U3109 (N_3109,N_2958,N_2972);
or U3110 (N_3110,N_2789,N_2778);
and U3111 (N_3111,N_2782,N_2883);
or U3112 (N_3112,N_2950,N_2825);
nor U3113 (N_3113,N_2837,N_2984);
nor U3114 (N_3114,N_2869,N_2759);
and U3115 (N_3115,N_2901,N_2774);
nor U3116 (N_3116,N_2834,N_2827);
nand U3117 (N_3117,N_2828,N_2942);
nor U3118 (N_3118,N_2994,N_2961);
nor U3119 (N_3119,N_2859,N_2770);
or U3120 (N_3120,N_2752,N_2903);
or U3121 (N_3121,N_2896,N_2857);
nand U3122 (N_3122,N_2779,N_2913);
xnor U3123 (N_3123,N_2818,N_2952);
or U3124 (N_3124,N_2763,N_2777);
nand U3125 (N_3125,N_2778,N_2844);
nor U3126 (N_3126,N_2787,N_2963);
nor U3127 (N_3127,N_2784,N_2825);
nand U3128 (N_3128,N_2997,N_2827);
nor U3129 (N_3129,N_2928,N_2793);
nor U3130 (N_3130,N_2983,N_2793);
or U3131 (N_3131,N_2981,N_2868);
and U3132 (N_3132,N_2764,N_2971);
and U3133 (N_3133,N_2762,N_2963);
or U3134 (N_3134,N_2918,N_2882);
and U3135 (N_3135,N_2886,N_2975);
nand U3136 (N_3136,N_2764,N_2796);
nand U3137 (N_3137,N_2755,N_2764);
and U3138 (N_3138,N_2805,N_2844);
xor U3139 (N_3139,N_2837,N_2920);
xnor U3140 (N_3140,N_2793,N_2781);
nand U3141 (N_3141,N_2811,N_2968);
or U3142 (N_3142,N_2787,N_2831);
nor U3143 (N_3143,N_2887,N_2852);
nor U3144 (N_3144,N_2951,N_2875);
and U3145 (N_3145,N_2825,N_2982);
nand U3146 (N_3146,N_2846,N_2781);
nor U3147 (N_3147,N_2839,N_2976);
nand U3148 (N_3148,N_2792,N_2844);
and U3149 (N_3149,N_2896,N_2948);
xnor U3150 (N_3150,N_2883,N_2894);
xor U3151 (N_3151,N_2770,N_2964);
nand U3152 (N_3152,N_2929,N_2836);
nor U3153 (N_3153,N_2855,N_2895);
nand U3154 (N_3154,N_2751,N_2936);
and U3155 (N_3155,N_2863,N_2795);
nand U3156 (N_3156,N_2919,N_2771);
and U3157 (N_3157,N_2921,N_2840);
or U3158 (N_3158,N_2954,N_2905);
xnor U3159 (N_3159,N_2955,N_2972);
nor U3160 (N_3160,N_2774,N_2921);
and U3161 (N_3161,N_2808,N_2995);
and U3162 (N_3162,N_2810,N_2871);
or U3163 (N_3163,N_2794,N_2780);
or U3164 (N_3164,N_2873,N_2921);
xnor U3165 (N_3165,N_2796,N_2861);
nor U3166 (N_3166,N_2815,N_2826);
nor U3167 (N_3167,N_2754,N_2990);
xnor U3168 (N_3168,N_2888,N_2981);
nand U3169 (N_3169,N_2829,N_2751);
nand U3170 (N_3170,N_2879,N_2760);
nor U3171 (N_3171,N_2813,N_2849);
and U3172 (N_3172,N_2875,N_2808);
and U3173 (N_3173,N_2800,N_2899);
xor U3174 (N_3174,N_2899,N_2923);
or U3175 (N_3175,N_2995,N_2866);
and U3176 (N_3176,N_2784,N_2794);
nand U3177 (N_3177,N_2804,N_2808);
nor U3178 (N_3178,N_2933,N_2973);
nand U3179 (N_3179,N_2981,N_2816);
nor U3180 (N_3180,N_2868,N_2882);
xor U3181 (N_3181,N_2823,N_2976);
or U3182 (N_3182,N_2816,N_2771);
or U3183 (N_3183,N_2785,N_2931);
nor U3184 (N_3184,N_2936,N_2758);
nor U3185 (N_3185,N_2840,N_2927);
or U3186 (N_3186,N_2777,N_2946);
xor U3187 (N_3187,N_2826,N_2752);
nand U3188 (N_3188,N_2986,N_2782);
or U3189 (N_3189,N_2976,N_2898);
xnor U3190 (N_3190,N_2967,N_2830);
nor U3191 (N_3191,N_2839,N_2915);
nor U3192 (N_3192,N_2912,N_2877);
or U3193 (N_3193,N_2946,N_2936);
nand U3194 (N_3194,N_2907,N_2764);
nor U3195 (N_3195,N_2798,N_2768);
and U3196 (N_3196,N_2981,N_2849);
nor U3197 (N_3197,N_2817,N_2947);
xnor U3198 (N_3198,N_2766,N_2949);
xor U3199 (N_3199,N_2952,N_2816);
nand U3200 (N_3200,N_2923,N_2765);
nand U3201 (N_3201,N_2759,N_2925);
or U3202 (N_3202,N_2802,N_2797);
xor U3203 (N_3203,N_2857,N_2865);
or U3204 (N_3204,N_2990,N_2882);
or U3205 (N_3205,N_2883,N_2769);
or U3206 (N_3206,N_2962,N_2921);
nor U3207 (N_3207,N_2827,N_2885);
or U3208 (N_3208,N_2966,N_2881);
nor U3209 (N_3209,N_2846,N_2770);
or U3210 (N_3210,N_2860,N_2796);
nor U3211 (N_3211,N_2765,N_2769);
nor U3212 (N_3212,N_2836,N_2968);
nand U3213 (N_3213,N_2815,N_2836);
nor U3214 (N_3214,N_2966,N_2853);
nor U3215 (N_3215,N_2942,N_2813);
nand U3216 (N_3216,N_2867,N_2752);
or U3217 (N_3217,N_2960,N_2909);
xor U3218 (N_3218,N_2836,N_2764);
nor U3219 (N_3219,N_2766,N_2925);
and U3220 (N_3220,N_2917,N_2895);
or U3221 (N_3221,N_2901,N_2883);
and U3222 (N_3222,N_2783,N_2895);
nand U3223 (N_3223,N_2886,N_2976);
xnor U3224 (N_3224,N_2941,N_2775);
nor U3225 (N_3225,N_2785,N_2894);
or U3226 (N_3226,N_2992,N_2838);
nand U3227 (N_3227,N_2940,N_2941);
and U3228 (N_3228,N_2927,N_2842);
nand U3229 (N_3229,N_2820,N_2789);
or U3230 (N_3230,N_2918,N_2840);
nand U3231 (N_3231,N_2847,N_2757);
or U3232 (N_3232,N_2887,N_2876);
xor U3233 (N_3233,N_2830,N_2851);
nor U3234 (N_3234,N_2883,N_2996);
and U3235 (N_3235,N_2994,N_2822);
nor U3236 (N_3236,N_2928,N_2865);
or U3237 (N_3237,N_2926,N_2882);
or U3238 (N_3238,N_2833,N_2775);
or U3239 (N_3239,N_2784,N_2981);
xor U3240 (N_3240,N_2796,N_2809);
xor U3241 (N_3241,N_2799,N_2977);
nand U3242 (N_3242,N_2792,N_2976);
xnor U3243 (N_3243,N_2831,N_2947);
nor U3244 (N_3244,N_2929,N_2950);
nand U3245 (N_3245,N_2883,N_2788);
or U3246 (N_3246,N_2928,N_2762);
nor U3247 (N_3247,N_2957,N_2759);
nand U3248 (N_3248,N_2934,N_2762);
and U3249 (N_3249,N_2992,N_2943);
nand U3250 (N_3250,N_3240,N_3222);
nor U3251 (N_3251,N_3174,N_3171);
xnor U3252 (N_3252,N_3117,N_3113);
nand U3253 (N_3253,N_3056,N_3239);
nand U3254 (N_3254,N_3213,N_3017);
and U3255 (N_3255,N_3127,N_3125);
xnor U3256 (N_3256,N_3051,N_3235);
and U3257 (N_3257,N_3063,N_3236);
nor U3258 (N_3258,N_3142,N_3131);
xnor U3259 (N_3259,N_3134,N_3150);
xor U3260 (N_3260,N_3027,N_3154);
xor U3261 (N_3261,N_3192,N_3061);
or U3262 (N_3262,N_3159,N_3243);
or U3263 (N_3263,N_3225,N_3191);
and U3264 (N_3264,N_3234,N_3039);
or U3265 (N_3265,N_3210,N_3166);
xnor U3266 (N_3266,N_3123,N_3152);
nand U3267 (N_3267,N_3185,N_3137);
or U3268 (N_3268,N_3148,N_3032);
and U3269 (N_3269,N_3090,N_3048);
nand U3270 (N_3270,N_3057,N_3022);
xnor U3271 (N_3271,N_3217,N_3066);
or U3272 (N_3272,N_3093,N_3129);
nand U3273 (N_3273,N_3247,N_3206);
nand U3274 (N_3274,N_3141,N_3097);
and U3275 (N_3275,N_3145,N_3031);
and U3276 (N_3276,N_3077,N_3212);
nor U3277 (N_3277,N_3238,N_3168);
or U3278 (N_3278,N_3107,N_3079);
nand U3279 (N_3279,N_3038,N_3172);
xor U3280 (N_3280,N_3081,N_3099);
nand U3281 (N_3281,N_3101,N_3111);
xnor U3282 (N_3282,N_3053,N_3052);
nor U3283 (N_3283,N_3139,N_3012);
nand U3284 (N_3284,N_3041,N_3106);
and U3285 (N_3285,N_3028,N_3004);
xor U3286 (N_3286,N_3203,N_3018);
xnor U3287 (N_3287,N_3067,N_3064);
nor U3288 (N_3288,N_3085,N_3121);
or U3289 (N_3289,N_3233,N_3034);
xnor U3290 (N_3290,N_3180,N_3151);
or U3291 (N_3291,N_3195,N_3211);
and U3292 (N_3292,N_3074,N_3030);
nand U3293 (N_3293,N_3071,N_3136);
or U3294 (N_3294,N_3229,N_3226);
and U3295 (N_3295,N_3223,N_3157);
nor U3296 (N_3296,N_3199,N_3033);
xnor U3297 (N_3297,N_3242,N_3014);
nor U3298 (N_3298,N_3219,N_3116);
or U3299 (N_3299,N_3096,N_3007);
nand U3300 (N_3300,N_3047,N_3241);
and U3301 (N_3301,N_3050,N_3156);
nand U3302 (N_3302,N_3016,N_3059);
and U3303 (N_3303,N_3095,N_3089);
xnor U3304 (N_3304,N_3084,N_3146);
xnor U3305 (N_3305,N_3110,N_3153);
nand U3306 (N_3306,N_3193,N_3232);
xor U3307 (N_3307,N_3224,N_3037);
nand U3308 (N_3308,N_3013,N_3214);
xnor U3309 (N_3309,N_3122,N_3133);
and U3310 (N_3310,N_3023,N_3132);
nand U3311 (N_3311,N_3135,N_3036);
or U3312 (N_3312,N_3245,N_3204);
nand U3313 (N_3313,N_3227,N_3005);
and U3314 (N_3314,N_3175,N_3181);
nor U3315 (N_3315,N_3000,N_3147);
nand U3316 (N_3316,N_3114,N_3006);
or U3317 (N_3317,N_3044,N_3080);
or U3318 (N_3318,N_3078,N_3216);
and U3319 (N_3319,N_3112,N_3182);
nor U3320 (N_3320,N_3073,N_3248);
nor U3321 (N_3321,N_3008,N_3009);
nor U3322 (N_3322,N_3015,N_3177);
nand U3323 (N_3323,N_3091,N_3170);
xnor U3324 (N_3324,N_3184,N_3124);
nand U3325 (N_3325,N_3188,N_3045);
nor U3326 (N_3326,N_3200,N_3201);
nand U3327 (N_3327,N_3161,N_3138);
xnor U3328 (N_3328,N_3118,N_3207);
and U3329 (N_3329,N_3237,N_3179);
nand U3330 (N_3330,N_3231,N_3075);
nor U3331 (N_3331,N_3120,N_3163);
or U3332 (N_3332,N_3205,N_3183);
and U3333 (N_3333,N_3202,N_3144);
nand U3334 (N_3334,N_3046,N_3094);
nand U3335 (N_3335,N_3158,N_3162);
nand U3336 (N_3336,N_3070,N_3187);
nand U3337 (N_3337,N_3169,N_3190);
and U3338 (N_3338,N_3165,N_3221);
nor U3339 (N_3339,N_3230,N_3176);
or U3340 (N_3340,N_3209,N_3126);
nand U3341 (N_3341,N_3003,N_3186);
or U3342 (N_3342,N_3244,N_3143);
and U3343 (N_3343,N_3105,N_3011);
and U3344 (N_3344,N_3098,N_3020);
and U3345 (N_3345,N_3149,N_3021);
xor U3346 (N_3346,N_3082,N_3065);
nand U3347 (N_3347,N_3076,N_3068);
and U3348 (N_3348,N_3246,N_3215);
and U3349 (N_3349,N_3087,N_3019);
and U3350 (N_3350,N_3198,N_3173);
and U3351 (N_3351,N_3196,N_3102);
or U3352 (N_3352,N_3088,N_3100);
and U3353 (N_3353,N_3026,N_3218);
xnor U3354 (N_3354,N_3055,N_3130);
nand U3355 (N_3355,N_3197,N_3086);
or U3356 (N_3356,N_3001,N_3042);
nor U3357 (N_3357,N_3160,N_3072);
nor U3358 (N_3358,N_3119,N_3167);
xnor U3359 (N_3359,N_3083,N_3208);
and U3360 (N_3360,N_3043,N_3220);
nor U3361 (N_3361,N_3108,N_3062);
or U3362 (N_3362,N_3035,N_3060);
or U3363 (N_3363,N_3054,N_3049);
nand U3364 (N_3364,N_3103,N_3002);
nor U3365 (N_3365,N_3040,N_3109);
xor U3366 (N_3366,N_3128,N_3164);
and U3367 (N_3367,N_3069,N_3249);
nand U3368 (N_3368,N_3104,N_3155);
nand U3369 (N_3369,N_3024,N_3025);
xnor U3370 (N_3370,N_3189,N_3029);
nor U3371 (N_3371,N_3092,N_3010);
xor U3372 (N_3372,N_3228,N_3115);
and U3373 (N_3373,N_3140,N_3178);
and U3374 (N_3374,N_3058,N_3194);
nor U3375 (N_3375,N_3101,N_3032);
nand U3376 (N_3376,N_3025,N_3004);
nor U3377 (N_3377,N_3101,N_3106);
nand U3378 (N_3378,N_3164,N_3046);
nand U3379 (N_3379,N_3150,N_3235);
xor U3380 (N_3380,N_3159,N_3057);
nor U3381 (N_3381,N_3095,N_3010);
and U3382 (N_3382,N_3198,N_3189);
nor U3383 (N_3383,N_3220,N_3040);
nor U3384 (N_3384,N_3114,N_3039);
nand U3385 (N_3385,N_3130,N_3237);
xnor U3386 (N_3386,N_3018,N_3073);
nand U3387 (N_3387,N_3162,N_3010);
nor U3388 (N_3388,N_3201,N_3107);
or U3389 (N_3389,N_3105,N_3113);
and U3390 (N_3390,N_3249,N_3004);
nand U3391 (N_3391,N_3233,N_3141);
nor U3392 (N_3392,N_3084,N_3090);
or U3393 (N_3393,N_3115,N_3022);
nor U3394 (N_3394,N_3136,N_3099);
or U3395 (N_3395,N_3058,N_3064);
xor U3396 (N_3396,N_3171,N_3154);
and U3397 (N_3397,N_3008,N_3113);
and U3398 (N_3398,N_3160,N_3194);
nor U3399 (N_3399,N_3021,N_3037);
and U3400 (N_3400,N_3082,N_3185);
xor U3401 (N_3401,N_3225,N_3003);
nand U3402 (N_3402,N_3089,N_3098);
nand U3403 (N_3403,N_3115,N_3085);
and U3404 (N_3404,N_3241,N_3025);
or U3405 (N_3405,N_3140,N_3212);
or U3406 (N_3406,N_3196,N_3206);
xor U3407 (N_3407,N_3232,N_3247);
nor U3408 (N_3408,N_3205,N_3193);
or U3409 (N_3409,N_3158,N_3226);
nand U3410 (N_3410,N_3136,N_3075);
or U3411 (N_3411,N_3149,N_3074);
xnor U3412 (N_3412,N_3168,N_3169);
xnor U3413 (N_3413,N_3136,N_3061);
and U3414 (N_3414,N_3059,N_3081);
nor U3415 (N_3415,N_3175,N_3053);
xnor U3416 (N_3416,N_3115,N_3153);
nand U3417 (N_3417,N_3170,N_3061);
nor U3418 (N_3418,N_3025,N_3062);
nand U3419 (N_3419,N_3050,N_3186);
and U3420 (N_3420,N_3050,N_3142);
nor U3421 (N_3421,N_3192,N_3052);
xnor U3422 (N_3422,N_3200,N_3222);
and U3423 (N_3423,N_3241,N_3140);
and U3424 (N_3424,N_3091,N_3088);
nor U3425 (N_3425,N_3246,N_3057);
xnor U3426 (N_3426,N_3193,N_3012);
xnor U3427 (N_3427,N_3241,N_3204);
or U3428 (N_3428,N_3196,N_3226);
nand U3429 (N_3429,N_3190,N_3051);
and U3430 (N_3430,N_3028,N_3071);
nand U3431 (N_3431,N_3106,N_3024);
and U3432 (N_3432,N_3169,N_3173);
and U3433 (N_3433,N_3179,N_3083);
xor U3434 (N_3434,N_3213,N_3175);
nand U3435 (N_3435,N_3111,N_3108);
or U3436 (N_3436,N_3051,N_3215);
nand U3437 (N_3437,N_3201,N_3090);
and U3438 (N_3438,N_3101,N_3023);
nor U3439 (N_3439,N_3045,N_3185);
nand U3440 (N_3440,N_3227,N_3154);
or U3441 (N_3441,N_3055,N_3080);
or U3442 (N_3442,N_3042,N_3002);
and U3443 (N_3443,N_3061,N_3233);
or U3444 (N_3444,N_3223,N_3052);
xor U3445 (N_3445,N_3083,N_3213);
nand U3446 (N_3446,N_3161,N_3177);
and U3447 (N_3447,N_3186,N_3032);
xor U3448 (N_3448,N_3039,N_3073);
nand U3449 (N_3449,N_3155,N_3044);
xnor U3450 (N_3450,N_3134,N_3118);
nand U3451 (N_3451,N_3139,N_3138);
and U3452 (N_3452,N_3049,N_3075);
or U3453 (N_3453,N_3121,N_3086);
xnor U3454 (N_3454,N_3171,N_3100);
xor U3455 (N_3455,N_3069,N_3024);
nand U3456 (N_3456,N_3235,N_3086);
xnor U3457 (N_3457,N_3130,N_3185);
or U3458 (N_3458,N_3046,N_3071);
and U3459 (N_3459,N_3060,N_3236);
nor U3460 (N_3460,N_3016,N_3170);
and U3461 (N_3461,N_3177,N_3009);
nand U3462 (N_3462,N_3134,N_3126);
xor U3463 (N_3463,N_3223,N_3152);
nand U3464 (N_3464,N_3139,N_3123);
nand U3465 (N_3465,N_3180,N_3056);
nand U3466 (N_3466,N_3069,N_3098);
nand U3467 (N_3467,N_3226,N_3165);
and U3468 (N_3468,N_3246,N_3169);
or U3469 (N_3469,N_3053,N_3126);
or U3470 (N_3470,N_3020,N_3053);
xnor U3471 (N_3471,N_3211,N_3102);
or U3472 (N_3472,N_3199,N_3076);
xnor U3473 (N_3473,N_3022,N_3234);
nor U3474 (N_3474,N_3014,N_3228);
xor U3475 (N_3475,N_3130,N_3061);
nor U3476 (N_3476,N_3152,N_3159);
xor U3477 (N_3477,N_3131,N_3198);
xor U3478 (N_3478,N_3140,N_3071);
nor U3479 (N_3479,N_3015,N_3128);
nand U3480 (N_3480,N_3249,N_3059);
xnor U3481 (N_3481,N_3019,N_3193);
nor U3482 (N_3482,N_3239,N_3046);
nor U3483 (N_3483,N_3248,N_3095);
or U3484 (N_3484,N_3105,N_3059);
and U3485 (N_3485,N_3135,N_3011);
nor U3486 (N_3486,N_3037,N_3222);
xnor U3487 (N_3487,N_3129,N_3140);
nor U3488 (N_3488,N_3135,N_3107);
nor U3489 (N_3489,N_3222,N_3220);
nor U3490 (N_3490,N_3176,N_3165);
xor U3491 (N_3491,N_3049,N_3175);
nor U3492 (N_3492,N_3104,N_3044);
nand U3493 (N_3493,N_3126,N_3047);
xor U3494 (N_3494,N_3149,N_3102);
nor U3495 (N_3495,N_3046,N_3178);
and U3496 (N_3496,N_3014,N_3176);
xor U3497 (N_3497,N_3133,N_3126);
nand U3498 (N_3498,N_3035,N_3104);
and U3499 (N_3499,N_3040,N_3151);
xnor U3500 (N_3500,N_3342,N_3343);
xor U3501 (N_3501,N_3439,N_3384);
nand U3502 (N_3502,N_3442,N_3468);
nand U3503 (N_3503,N_3268,N_3317);
nor U3504 (N_3504,N_3345,N_3291);
and U3505 (N_3505,N_3318,N_3492);
nor U3506 (N_3506,N_3484,N_3408);
or U3507 (N_3507,N_3255,N_3454);
nand U3508 (N_3508,N_3420,N_3382);
or U3509 (N_3509,N_3341,N_3371);
nand U3510 (N_3510,N_3458,N_3433);
nand U3511 (N_3511,N_3426,N_3482);
or U3512 (N_3512,N_3322,N_3287);
and U3513 (N_3513,N_3479,N_3305);
xnor U3514 (N_3514,N_3309,N_3480);
nor U3515 (N_3515,N_3306,N_3279);
xnor U3516 (N_3516,N_3339,N_3412);
and U3517 (N_3517,N_3447,N_3378);
nor U3518 (N_3518,N_3374,N_3280);
nand U3519 (N_3519,N_3373,N_3301);
and U3520 (N_3520,N_3358,N_3366);
and U3521 (N_3521,N_3406,N_3489);
and U3522 (N_3522,N_3470,N_3375);
and U3523 (N_3523,N_3323,N_3302);
nor U3524 (N_3524,N_3485,N_3278);
nor U3525 (N_3525,N_3330,N_3367);
nor U3526 (N_3526,N_3423,N_3282);
xnor U3527 (N_3527,N_3385,N_3297);
and U3528 (N_3528,N_3274,N_3400);
nand U3529 (N_3529,N_3300,N_3498);
and U3530 (N_3530,N_3275,N_3263);
xor U3531 (N_3531,N_3258,N_3487);
nor U3532 (N_3532,N_3418,N_3348);
nor U3533 (N_3533,N_3281,N_3472);
and U3534 (N_3534,N_3466,N_3364);
xnor U3535 (N_3535,N_3356,N_3350);
xor U3536 (N_3536,N_3340,N_3303);
and U3537 (N_3537,N_3443,N_3370);
nor U3538 (N_3538,N_3486,N_3295);
or U3539 (N_3539,N_3383,N_3365);
nor U3540 (N_3540,N_3376,N_3308);
xnor U3541 (N_3541,N_3277,N_3267);
nand U3542 (N_3542,N_3438,N_3452);
and U3543 (N_3543,N_3349,N_3427);
nand U3544 (N_3544,N_3333,N_3455);
xnor U3545 (N_3545,N_3296,N_3284);
and U3546 (N_3546,N_3397,N_3490);
nand U3547 (N_3547,N_3362,N_3461);
and U3548 (N_3548,N_3276,N_3391);
and U3549 (N_3549,N_3425,N_3372);
or U3550 (N_3550,N_3437,N_3424);
nor U3551 (N_3551,N_3444,N_3446);
xnor U3552 (N_3552,N_3451,N_3257);
or U3553 (N_3553,N_3253,N_3394);
nand U3554 (N_3554,N_3273,N_3360);
nor U3555 (N_3555,N_3346,N_3448);
xor U3556 (N_3556,N_3459,N_3396);
xnor U3557 (N_3557,N_3256,N_3377);
xor U3558 (N_3558,N_3398,N_3422);
xnor U3559 (N_3559,N_3289,N_3411);
and U3560 (N_3560,N_3414,N_3270);
nor U3561 (N_3561,N_3285,N_3368);
nand U3562 (N_3562,N_3387,N_3460);
xor U3563 (N_3563,N_3336,N_3315);
and U3564 (N_3564,N_3338,N_3288);
nor U3565 (N_3565,N_3347,N_3344);
xor U3566 (N_3566,N_3319,N_3290);
and U3567 (N_3567,N_3413,N_3463);
and U3568 (N_3568,N_3250,N_3493);
or U3569 (N_3569,N_3326,N_3299);
xor U3570 (N_3570,N_3471,N_3393);
nor U3571 (N_3571,N_3252,N_3328);
and U3572 (N_3572,N_3475,N_3473);
nor U3573 (N_3573,N_3332,N_3395);
xor U3574 (N_3574,N_3316,N_3410);
xnor U3575 (N_3575,N_3497,N_3430);
and U3576 (N_3576,N_3416,N_3386);
nor U3577 (N_3577,N_3320,N_3251);
nand U3578 (N_3578,N_3264,N_3298);
or U3579 (N_3579,N_3381,N_3432);
nand U3580 (N_3580,N_3325,N_3494);
nor U3581 (N_3581,N_3478,N_3469);
xor U3582 (N_3582,N_3462,N_3421);
and U3583 (N_3583,N_3260,N_3457);
nor U3584 (N_3584,N_3335,N_3312);
xor U3585 (N_3585,N_3351,N_3453);
xnor U3586 (N_3586,N_3304,N_3441);
and U3587 (N_3587,N_3481,N_3265);
and U3588 (N_3588,N_3449,N_3474);
and U3589 (N_3589,N_3311,N_3405);
nand U3590 (N_3590,N_3283,N_3352);
nor U3591 (N_3591,N_3269,N_3399);
and U3592 (N_3592,N_3337,N_3262);
and U3593 (N_3593,N_3465,N_3379);
xor U3594 (N_3594,N_3272,N_3417);
or U3595 (N_3595,N_3401,N_3450);
nand U3596 (N_3596,N_3499,N_3271);
or U3597 (N_3597,N_3361,N_3409);
nand U3598 (N_3598,N_3436,N_3402);
nor U3599 (N_3599,N_3419,N_3254);
or U3600 (N_3600,N_3327,N_3331);
nand U3601 (N_3601,N_3390,N_3324);
or U3602 (N_3602,N_3431,N_3434);
or U3603 (N_3603,N_3321,N_3429);
nand U3604 (N_3604,N_3313,N_3380);
and U3605 (N_3605,N_3369,N_3363);
or U3606 (N_3606,N_3496,N_3261);
and U3607 (N_3607,N_3467,N_3314);
and U3608 (N_3608,N_3334,N_3357);
nand U3609 (N_3609,N_3464,N_3294);
nor U3610 (N_3610,N_3286,N_3404);
nand U3611 (N_3611,N_3415,N_3477);
xnor U3612 (N_3612,N_3407,N_3456);
nand U3613 (N_3613,N_3392,N_3359);
xor U3614 (N_3614,N_3491,N_3388);
nand U3615 (N_3615,N_3355,N_3495);
nand U3616 (N_3616,N_3488,N_3428);
and U3617 (N_3617,N_3476,N_3354);
or U3618 (N_3618,N_3389,N_3403);
and U3619 (N_3619,N_3435,N_3445);
nand U3620 (N_3620,N_3292,N_3329);
xnor U3621 (N_3621,N_3440,N_3483);
xor U3622 (N_3622,N_3310,N_3307);
and U3623 (N_3623,N_3293,N_3353);
or U3624 (N_3624,N_3259,N_3266);
and U3625 (N_3625,N_3349,N_3364);
or U3626 (N_3626,N_3308,N_3411);
or U3627 (N_3627,N_3425,N_3411);
and U3628 (N_3628,N_3368,N_3317);
xor U3629 (N_3629,N_3359,N_3415);
nand U3630 (N_3630,N_3375,N_3448);
nand U3631 (N_3631,N_3320,N_3348);
nand U3632 (N_3632,N_3345,N_3311);
or U3633 (N_3633,N_3323,N_3384);
nand U3634 (N_3634,N_3347,N_3309);
or U3635 (N_3635,N_3378,N_3309);
xor U3636 (N_3636,N_3365,N_3486);
and U3637 (N_3637,N_3308,N_3468);
nor U3638 (N_3638,N_3397,N_3341);
nor U3639 (N_3639,N_3268,N_3374);
or U3640 (N_3640,N_3472,N_3454);
nor U3641 (N_3641,N_3366,N_3411);
or U3642 (N_3642,N_3355,N_3316);
nor U3643 (N_3643,N_3421,N_3276);
xor U3644 (N_3644,N_3404,N_3333);
nand U3645 (N_3645,N_3494,N_3265);
nor U3646 (N_3646,N_3267,N_3410);
xnor U3647 (N_3647,N_3444,N_3344);
or U3648 (N_3648,N_3403,N_3329);
xnor U3649 (N_3649,N_3454,N_3315);
nor U3650 (N_3650,N_3382,N_3257);
or U3651 (N_3651,N_3271,N_3461);
xor U3652 (N_3652,N_3252,N_3319);
xnor U3653 (N_3653,N_3450,N_3256);
xor U3654 (N_3654,N_3393,N_3281);
nor U3655 (N_3655,N_3446,N_3327);
or U3656 (N_3656,N_3256,N_3314);
and U3657 (N_3657,N_3498,N_3484);
or U3658 (N_3658,N_3350,N_3339);
xor U3659 (N_3659,N_3251,N_3334);
and U3660 (N_3660,N_3275,N_3396);
nand U3661 (N_3661,N_3271,N_3494);
or U3662 (N_3662,N_3357,N_3265);
nand U3663 (N_3663,N_3358,N_3354);
xor U3664 (N_3664,N_3498,N_3441);
and U3665 (N_3665,N_3399,N_3268);
nor U3666 (N_3666,N_3359,N_3357);
or U3667 (N_3667,N_3328,N_3497);
or U3668 (N_3668,N_3267,N_3330);
or U3669 (N_3669,N_3463,N_3383);
xor U3670 (N_3670,N_3344,N_3263);
or U3671 (N_3671,N_3485,N_3265);
and U3672 (N_3672,N_3278,N_3258);
and U3673 (N_3673,N_3261,N_3319);
or U3674 (N_3674,N_3462,N_3471);
nand U3675 (N_3675,N_3401,N_3366);
and U3676 (N_3676,N_3296,N_3327);
and U3677 (N_3677,N_3471,N_3254);
and U3678 (N_3678,N_3276,N_3388);
and U3679 (N_3679,N_3463,N_3404);
nor U3680 (N_3680,N_3491,N_3302);
nand U3681 (N_3681,N_3457,N_3468);
nand U3682 (N_3682,N_3409,N_3472);
nand U3683 (N_3683,N_3351,N_3357);
nand U3684 (N_3684,N_3288,N_3344);
nor U3685 (N_3685,N_3404,N_3425);
and U3686 (N_3686,N_3293,N_3385);
and U3687 (N_3687,N_3441,N_3314);
xor U3688 (N_3688,N_3432,N_3301);
xnor U3689 (N_3689,N_3449,N_3441);
xnor U3690 (N_3690,N_3362,N_3354);
xor U3691 (N_3691,N_3406,N_3447);
nand U3692 (N_3692,N_3305,N_3301);
nand U3693 (N_3693,N_3258,N_3271);
xor U3694 (N_3694,N_3369,N_3443);
or U3695 (N_3695,N_3459,N_3399);
and U3696 (N_3696,N_3306,N_3413);
nor U3697 (N_3697,N_3482,N_3393);
xor U3698 (N_3698,N_3271,N_3451);
nand U3699 (N_3699,N_3481,N_3380);
or U3700 (N_3700,N_3444,N_3461);
xnor U3701 (N_3701,N_3422,N_3382);
or U3702 (N_3702,N_3446,N_3494);
nor U3703 (N_3703,N_3457,N_3325);
nor U3704 (N_3704,N_3257,N_3416);
nand U3705 (N_3705,N_3328,N_3403);
nand U3706 (N_3706,N_3495,N_3385);
nand U3707 (N_3707,N_3465,N_3287);
nand U3708 (N_3708,N_3397,N_3398);
nand U3709 (N_3709,N_3321,N_3293);
or U3710 (N_3710,N_3274,N_3354);
nor U3711 (N_3711,N_3398,N_3421);
nand U3712 (N_3712,N_3312,N_3404);
nand U3713 (N_3713,N_3446,N_3375);
nand U3714 (N_3714,N_3323,N_3401);
nor U3715 (N_3715,N_3250,N_3371);
xnor U3716 (N_3716,N_3276,N_3316);
nor U3717 (N_3717,N_3489,N_3323);
nand U3718 (N_3718,N_3302,N_3252);
nand U3719 (N_3719,N_3377,N_3458);
nand U3720 (N_3720,N_3443,N_3332);
nand U3721 (N_3721,N_3391,N_3268);
xnor U3722 (N_3722,N_3298,N_3252);
and U3723 (N_3723,N_3263,N_3476);
and U3724 (N_3724,N_3409,N_3473);
and U3725 (N_3725,N_3263,N_3323);
or U3726 (N_3726,N_3463,N_3380);
and U3727 (N_3727,N_3494,N_3492);
and U3728 (N_3728,N_3305,N_3467);
nor U3729 (N_3729,N_3480,N_3342);
and U3730 (N_3730,N_3328,N_3314);
nand U3731 (N_3731,N_3318,N_3490);
nand U3732 (N_3732,N_3466,N_3282);
and U3733 (N_3733,N_3441,N_3280);
and U3734 (N_3734,N_3423,N_3370);
and U3735 (N_3735,N_3371,N_3296);
or U3736 (N_3736,N_3335,N_3389);
xor U3737 (N_3737,N_3482,N_3272);
xnor U3738 (N_3738,N_3465,N_3404);
or U3739 (N_3739,N_3410,N_3279);
and U3740 (N_3740,N_3258,N_3422);
and U3741 (N_3741,N_3327,N_3274);
xnor U3742 (N_3742,N_3474,N_3274);
and U3743 (N_3743,N_3337,N_3490);
and U3744 (N_3744,N_3473,N_3302);
or U3745 (N_3745,N_3356,N_3441);
nand U3746 (N_3746,N_3488,N_3326);
nor U3747 (N_3747,N_3298,N_3466);
and U3748 (N_3748,N_3382,N_3425);
nand U3749 (N_3749,N_3348,N_3413);
and U3750 (N_3750,N_3519,N_3540);
or U3751 (N_3751,N_3686,N_3744);
nand U3752 (N_3752,N_3637,N_3517);
or U3753 (N_3753,N_3606,N_3716);
and U3754 (N_3754,N_3605,N_3592);
and U3755 (N_3755,N_3563,N_3653);
nand U3756 (N_3756,N_3589,N_3545);
nand U3757 (N_3757,N_3541,N_3630);
or U3758 (N_3758,N_3513,N_3565);
nand U3759 (N_3759,N_3511,N_3524);
and U3760 (N_3760,N_3733,N_3746);
nor U3761 (N_3761,N_3666,N_3556);
or U3762 (N_3762,N_3629,N_3646);
xor U3763 (N_3763,N_3594,N_3628);
and U3764 (N_3764,N_3564,N_3621);
nor U3765 (N_3765,N_3670,N_3701);
and U3766 (N_3766,N_3529,N_3662);
or U3767 (N_3767,N_3547,N_3546);
nor U3768 (N_3768,N_3729,N_3617);
or U3769 (N_3769,N_3510,N_3678);
nor U3770 (N_3770,N_3692,N_3591);
nor U3771 (N_3771,N_3571,N_3702);
or U3772 (N_3772,N_3580,N_3508);
or U3773 (N_3773,N_3554,N_3619);
and U3774 (N_3774,N_3694,N_3560);
or U3775 (N_3775,N_3635,N_3613);
and U3776 (N_3776,N_3588,N_3557);
nand U3777 (N_3777,N_3500,N_3640);
and U3778 (N_3778,N_3533,N_3674);
nand U3779 (N_3779,N_3639,N_3555);
and U3780 (N_3780,N_3722,N_3749);
xor U3781 (N_3781,N_3599,N_3717);
nor U3782 (N_3782,N_3544,N_3573);
nor U3783 (N_3783,N_3570,N_3514);
xor U3784 (N_3784,N_3721,N_3520);
and U3785 (N_3785,N_3699,N_3620);
nand U3786 (N_3786,N_3659,N_3743);
nand U3787 (N_3787,N_3608,N_3656);
nand U3788 (N_3788,N_3598,N_3723);
xor U3789 (N_3789,N_3603,N_3579);
nor U3790 (N_3790,N_3703,N_3668);
xnor U3791 (N_3791,N_3527,N_3568);
xor U3792 (N_3792,N_3607,N_3558);
or U3793 (N_3793,N_3731,N_3595);
or U3794 (N_3794,N_3574,N_3600);
nand U3795 (N_3795,N_3530,N_3676);
nor U3796 (N_3796,N_3633,N_3614);
or U3797 (N_3797,N_3632,N_3660);
or U3798 (N_3798,N_3679,N_3596);
and U3799 (N_3799,N_3661,N_3553);
xor U3800 (N_3800,N_3538,N_3691);
or U3801 (N_3801,N_3708,N_3652);
nand U3802 (N_3802,N_3685,N_3505);
or U3803 (N_3803,N_3569,N_3585);
nand U3804 (N_3804,N_3644,N_3502);
nand U3805 (N_3805,N_3503,N_3696);
nand U3806 (N_3806,N_3501,N_3531);
and U3807 (N_3807,N_3650,N_3738);
nor U3808 (N_3808,N_3586,N_3704);
nand U3809 (N_3809,N_3724,N_3618);
xnor U3810 (N_3810,N_3576,N_3597);
nand U3811 (N_3811,N_3682,N_3730);
and U3812 (N_3812,N_3638,N_3602);
and U3813 (N_3813,N_3705,N_3572);
nand U3814 (N_3814,N_3683,N_3714);
xnor U3815 (N_3815,N_3634,N_3673);
nand U3816 (N_3816,N_3623,N_3649);
or U3817 (N_3817,N_3518,N_3601);
nand U3818 (N_3818,N_3542,N_3551);
xor U3819 (N_3819,N_3507,N_3748);
nor U3820 (N_3820,N_3559,N_3710);
nor U3821 (N_3821,N_3698,N_3522);
xor U3822 (N_3822,N_3681,N_3713);
nor U3823 (N_3823,N_3526,N_3525);
and U3824 (N_3824,N_3735,N_3566);
nand U3825 (N_3825,N_3515,N_3669);
and U3826 (N_3826,N_3504,N_3709);
or U3827 (N_3827,N_3671,N_3578);
and U3828 (N_3828,N_3567,N_3593);
xnor U3829 (N_3829,N_3684,N_3658);
nor U3830 (N_3830,N_3624,N_3627);
and U3831 (N_3831,N_3667,N_3695);
and U3832 (N_3832,N_3745,N_3715);
and U3833 (N_3833,N_3711,N_3590);
nand U3834 (N_3834,N_3707,N_3610);
and U3835 (N_3835,N_3677,N_3626);
and U3836 (N_3836,N_3648,N_3725);
nand U3837 (N_3837,N_3697,N_3647);
xnor U3838 (N_3838,N_3616,N_3664);
xor U3839 (N_3839,N_3712,N_3612);
xnor U3840 (N_3840,N_3690,N_3536);
or U3841 (N_3841,N_3654,N_3611);
xor U3842 (N_3842,N_3506,N_3582);
and U3843 (N_3843,N_3562,N_3643);
and U3844 (N_3844,N_3625,N_3732);
nor U3845 (N_3845,N_3583,N_3651);
nor U3846 (N_3846,N_3577,N_3693);
nand U3847 (N_3847,N_3636,N_3747);
nand U3848 (N_3848,N_3641,N_3523);
and U3849 (N_3849,N_3740,N_3549);
nor U3850 (N_3850,N_3631,N_3561);
nand U3851 (N_3851,N_3689,N_3534);
nand U3852 (N_3852,N_3645,N_3655);
xor U3853 (N_3853,N_3736,N_3604);
nor U3854 (N_3854,N_3642,N_3584);
nand U3855 (N_3855,N_3609,N_3581);
and U3856 (N_3856,N_3739,N_3700);
and U3857 (N_3857,N_3718,N_3521);
xnor U3858 (N_3858,N_3675,N_3680);
xnor U3859 (N_3859,N_3734,N_3537);
nand U3860 (N_3860,N_3512,N_3535);
and U3861 (N_3861,N_3720,N_3737);
xor U3862 (N_3862,N_3532,N_3663);
nor U3863 (N_3863,N_3687,N_3543);
nor U3864 (N_3864,N_3539,N_3552);
nand U3865 (N_3865,N_3528,N_3509);
nand U3866 (N_3866,N_3719,N_3688);
xor U3867 (N_3867,N_3615,N_3665);
nand U3868 (N_3868,N_3657,N_3516);
or U3869 (N_3869,N_3742,N_3548);
and U3870 (N_3870,N_3672,N_3575);
nand U3871 (N_3871,N_3727,N_3550);
or U3872 (N_3872,N_3587,N_3706);
or U3873 (N_3873,N_3741,N_3726);
or U3874 (N_3874,N_3622,N_3728);
and U3875 (N_3875,N_3645,N_3708);
or U3876 (N_3876,N_3542,N_3666);
or U3877 (N_3877,N_3723,N_3707);
nand U3878 (N_3878,N_3598,N_3647);
or U3879 (N_3879,N_3724,N_3658);
xnor U3880 (N_3880,N_3711,N_3694);
and U3881 (N_3881,N_3661,N_3690);
nor U3882 (N_3882,N_3666,N_3505);
xor U3883 (N_3883,N_3714,N_3560);
xor U3884 (N_3884,N_3625,N_3734);
and U3885 (N_3885,N_3533,N_3578);
and U3886 (N_3886,N_3691,N_3656);
xnor U3887 (N_3887,N_3672,N_3522);
or U3888 (N_3888,N_3696,N_3740);
nor U3889 (N_3889,N_3581,N_3516);
or U3890 (N_3890,N_3640,N_3635);
and U3891 (N_3891,N_3748,N_3548);
or U3892 (N_3892,N_3709,N_3557);
nor U3893 (N_3893,N_3558,N_3502);
or U3894 (N_3894,N_3585,N_3700);
and U3895 (N_3895,N_3531,N_3525);
nor U3896 (N_3896,N_3635,N_3747);
xor U3897 (N_3897,N_3558,N_3654);
nand U3898 (N_3898,N_3695,N_3530);
or U3899 (N_3899,N_3699,N_3730);
xor U3900 (N_3900,N_3641,N_3688);
xnor U3901 (N_3901,N_3501,N_3652);
and U3902 (N_3902,N_3527,N_3549);
or U3903 (N_3903,N_3512,N_3704);
nor U3904 (N_3904,N_3744,N_3531);
nor U3905 (N_3905,N_3576,N_3637);
nor U3906 (N_3906,N_3669,N_3641);
nor U3907 (N_3907,N_3636,N_3526);
and U3908 (N_3908,N_3504,N_3732);
and U3909 (N_3909,N_3663,N_3740);
and U3910 (N_3910,N_3574,N_3627);
or U3911 (N_3911,N_3505,N_3724);
or U3912 (N_3912,N_3647,N_3511);
xnor U3913 (N_3913,N_3666,N_3528);
or U3914 (N_3914,N_3691,N_3509);
or U3915 (N_3915,N_3509,N_3689);
xnor U3916 (N_3916,N_3555,N_3553);
nor U3917 (N_3917,N_3557,N_3749);
and U3918 (N_3918,N_3612,N_3736);
or U3919 (N_3919,N_3598,N_3653);
or U3920 (N_3920,N_3655,N_3710);
xor U3921 (N_3921,N_3565,N_3508);
or U3922 (N_3922,N_3674,N_3675);
or U3923 (N_3923,N_3606,N_3597);
xnor U3924 (N_3924,N_3721,N_3691);
or U3925 (N_3925,N_3598,N_3543);
or U3926 (N_3926,N_3688,N_3590);
xnor U3927 (N_3927,N_3528,N_3746);
or U3928 (N_3928,N_3724,N_3712);
nor U3929 (N_3929,N_3681,N_3574);
and U3930 (N_3930,N_3619,N_3642);
or U3931 (N_3931,N_3638,N_3647);
nand U3932 (N_3932,N_3686,N_3688);
nand U3933 (N_3933,N_3672,N_3552);
or U3934 (N_3934,N_3630,N_3649);
or U3935 (N_3935,N_3701,N_3704);
nor U3936 (N_3936,N_3559,N_3557);
xnor U3937 (N_3937,N_3610,N_3552);
or U3938 (N_3938,N_3533,N_3550);
xor U3939 (N_3939,N_3631,N_3539);
nor U3940 (N_3940,N_3670,N_3548);
nor U3941 (N_3941,N_3684,N_3662);
or U3942 (N_3942,N_3684,N_3532);
nor U3943 (N_3943,N_3675,N_3684);
nor U3944 (N_3944,N_3548,N_3568);
and U3945 (N_3945,N_3654,N_3718);
and U3946 (N_3946,N_3545,N_3644);
and U3947 (N_3947,N_3694,N_3682);
or U3948 (N_3948,N_3615,N_3626);
or U3949 (N_3949,N_3661,N_3725);
and U3950 (N_3950,N_3538,N_3712);
xor U3951 (N_3951,N_3651,N_3740);
nand U3952 (N_3952,N_3712,N_3576);
or U3953 (N_3953,N_3706,N_3629);
xnor U3954 (N_3954,N_3641,N_3702);
and U3955 (N_3955,N_3668,N_3523);
or U3956 (N_3956,N_3685,N_3736);
nor U3957 (N_3957,N_3718,N_3734);
nand U3958 (N_3958,N_3627,N_3589);
or U3959 (N_3959,N_3744,N_3577);
and U3960 (N_3960,N_3721,N_3673);
or U3961 (N_3961,N_3693,N_3626);
and U3962 (N_3962,N_3601,N_3641);
nor U3963 (N_3963,N_3697,N_3538);
or U3964 (N_3964,N_3737,N_3593);
and U3965 (N_3965,N_3703,N_3564);
nand U3966 (N_3966,N_3629,N_3506);
nand U3967 (N_3967,N_3715,N_3726);
nor U3968 (N_3968,N_3711,N_3741);
nand U3969 (N_3969,N_3617,N_3745);
nand U3970 (N_3970,N_3714,N_3718);
nor U3971 (N_3971,N_3737,N_3677);
nor U3972 (N_3972,N_3632,N_3615);
and U3973 (N_3973,N_3663,N_3617);
or U3974 (N_3974,N_3741,N_3672);
xnor U3975 (N_3975,N_3710,N_3742);
nor U3976 (N_3976,N_3645,N_3682);
xor U3977 (N_3977,N_3708,N_3604);
nand U3978 (N_3978,N_3512,N_3671);
xor U3979 (N_3979,N_3733,N_3559);
nand U3980 (N_3980,N_3599,N_3709);
or U3981 (N_3981,N_3599,N_3582);
or U3982 (N_3982,N_3687,N_3532);
and U3983 (N_3983,N_3579,N_3556);
xnor U3984 (N_3984,N_3653,N_3656);
nand U3985 (N_3985,N_3739,N_3583);
or U3986 (N_3986,N_3700,N_3720);
and U3987 (N_3987,N_3693,N_3570);
and U3988 (N_3988,N_3501,N_3722);
nor U3989 (N_3989,N_3607,N_3550);
and U3990 (N_3990,N_3638,N_3511);
xor U3991 (N_3991,N_3741,N_3697);
xnor U3992 (N_3992,N_3628,N_3737);
or U3993 (N_3993,N_3687,N_3558);
nor U3994 (N_3994,N_3610,N_3680);
nor U3995 (N_3995,N_3736,N_3576);
xor U3996 (N_3996,N_3504,N_3575);
or U3997 (N_3997,N_3721,N_3517);
nor U3998 (N_3998,N_3727,N_3704);
nor U3999 (N_3999,N_3562,N_3523);
nor U4000 (N_4000,N_3997,N_3959);
nand U4001 (N_4001,N_3928,N_3946);
or U4002 (N_4002,N_3951,N_3896);
nor U4003 (N_4003,N_3802,N_3998);
or U4004 (N_4004,N_3907,N_3803);
xor U4005 (N_4005,N_3752,N_3850);
or U4006 (N_4006,N_3857,N_3984);
or U4007 (N_4007,N_3798,N_3860);
nand U4008 (N_4008,N_3847,N_3830);
or U4009 (N_4009,N_3804,N_3987);
xor U4010 (N_4010,N_3913,N_3911);
or U4011 (N_4011,N_3800,N_3983);
nor U4012 (N_4012,N_3968,N_3999);
nor U4013 (N_4013,N_3899,N_3880);
or U4014 (N_4014,N_3958,N_3975);
nor U4015 (N_4015,N_3866,N_3784);
nor U4016 (N_4016,N_3972,N_3827);
or U4017 (N_4017,N_3795,N_3807);
and U4018 (N_4018,N_3852,N_3960);
nor U4019 (N_4019,N_3937,N_3879);
xor U4020 (N_4020,N_3955,N_3853);
nand U4021 (N_4021,N_3816,N_3985);
or U4022 (N_4022,N_3772,N_3882);
and U4023 (N_4023,N_3868,N_3790);
or U4024 (N_4024,N_3856,N_3940);
nor U4025 (N_4025,N_3797,N_3819);
or U4026 (N_4026,N_3832,N_3978);
or U4027 (N_4027,N_3851,N_3858);
and U4028 (N_4028,N_3791,N_3967);
or U4029 (N_4029,N_3877,N_3986);
or U4030 (N_4030,N_3942,N_3924);
and U4031 (N_4031,N_3993,N_3874);
and U4032 (N_4032,N_3900,N_3750);
xor U4033 (N_4033,N_3815,N_3980);
nand U4034 (N_4034,N_3805,N_3822);
xor U4035 (N_4035,N_3915,N_3901);
nor U4036 (N_4036,N_3801,N_3898);
xnor U4037 (N_4037,N_3921,N_3758);
or U4038 (N_4038,N_3810,N_3962);
nor U4039 (N_4039,N_3887,N_3971);
and U4040 (N_4040,N_3761,N_3954);
xnor U4041 (N_4041,N_3825,N_3990);
and U4042 (N_4042,N_3957,N_3923);
or U4043 (N_4043,N_3792,N_3841);
and U4044 (N_4044,N_3884,N_3944);
xnor U4045 (N_4045,N_3994,N_3759);
xnor U4046 (N_4046,N_3861,N_3834);
xor U4047 (N_4047,N_3814,N_3891);
or U4048 (N_4048,N_3935,N_3931);
nor U4049 (N_4049,N_3903,N_3977);
or U4050 (N_4050,N_3775,N_3789);
nand U4051 (N_4051,N_3773,N_3920);
and U4052 (N_4052,N_3876,N_3873);
xnor U4053 (N_4053,N_3941,N_3893);
nand U4054 (N_4054,N_3979,N_3939);
nand U4055 (N_4055,N_3918,N_3849);
nand U4056 (N_4056,N_3767,N_3794);
xnor U4057 (N_4057,N_3904,N_3781);
and U4058 (N_4058,N_3966,N_3912);
nand U4059 (N_4059,N_3897,N_3870);
and U4060 (N_4060,N_3854,N_3836);
xnor U4061 (N_4061,N_3774,N_3890);
nand U4062 (N_4062,N_3906,N_3837);
or U4063 (N_4063,N_3845,N_3838);
xnor U4064 (N_4064,N_3964,N_3933);
nor U4065 (N_4065,N_3826,N_3864);
nor U4066 (N_4066,N_3925,N_3883);
or U4067 (N_4067,N_3885,N_3914);
and U4068 (N_4068,N_3757,N_3829);
or U4069 (N_4069,N_3872,N_3782);
and U4070 (N_4070,N_3763,N_3843);
nand U4071 (N_4071,N_3909,N_3776);
xnor U4072 (N_4072,N_3835,N_3756);
or U4073 (N_4073,N_3862,N_3976);
or U4074 (N_4074,N_3930,N_3934);
and U4075 (N_4075,N_3927,N_3974);
xor U4076 (N_4076,N_3840,N_3848);
nor U4077 (N_4077,N_3753,N_3808);
xor U4078 (N_4078,N_3821,N_3828);
xor U4079 (N_4079,N_3765,N_3770);
nand U4080 (N_4080,N_3865,N_3917);
or U4081 (N_4081,N_3796,N_3952);
nand U4082 (N_4082,N_3760,N_3833);
nand U4083 (N_4083,N_3751,N_3886);
xor U4084 (N_4084,N_3859,N_3844);
and U4085 (N_4085,N_3938,N_3842);
nor U4086 (N_4086,N_3813,N_3783);
or U4087 (N_4087,N_3996,N_3908);
nand U4088 (N_4088,N_3894,N_3786);
nor U4089 (N_4089,N_3910,N_3768);
nand U4090 (N_4090,N_3823,N_3764);
and U4091 (N_4091,N_3892,N_3875);
or U4092 (N_4092,N_3778,N_3995);
and U4093 (N_4093,N_3961,N_3855);
or U4094 (N_4094,N_3948,N_3777);
xnor U4095 (N_4095,N_3846,N_3956);
and U4096 (N_4096,N_3754,N_3793);
xnor U4097 (N_4097,N_3953,N_3945);
nand U4098 (N_4098,N_3839,N_3878);
and U4099 (N_4099,N_3963,N_3943);
nor U4100 (N_4100,N_3988,N_3869);
nand U4101 (N_4101,N_3762,N_3881);
and U4102 (N_4102,N_3970,N_3989);
nor U4103 (N_4103,N_3818,N_3831);
or U4104 (N_4104,N_3809,N_3863);
xor U4105 (N_4105,N_3982,N_3766);
xor U4106 (N_4106,N_3820,N_3824);
nor U4107 (N_4107,N_3926,N_3817);
nand U4108 (N_4108,N_3922,N_3888);
nor U4109 (N_4109,N_3992,N_3785);
nand U4110 (N_4110,N_3949,N_3780);
or U4111 (N_4111,N_3867,N_3779);
and U4112 (N_4112,N_3788,N_3965);
xor U4113 (N_4113,N_3787,N_3936);
nand U4114 (N_4114,N_3973,N_3981);
or U4115 (N_4115,N_3929,N_3889);
nor U4116 (N_4116,N_3806,N_3969);
nand U4117 (N_4117,N_3812,N_3947);
and U4118 (N_4118,N_3932,N_3991);
nand U4119 (N_4119,N_3950,N_3799);
nand U4120 (N_4120,N_3895,N_3916);
nor U4121 (N_4121,N_3905,N_3769);
and U4122 (N_4122,N_3871,N_3755);
or U4123 (N_4123,N_3771,N_3902);
nor U4124 (N_4124,N_3919,N_3811);
nor U4125 (N_4125,N_3947,N_3794);
and U4126 (N_4126,N_3962,N_3863);
xor U4127 (N_4127,N_3800,N_3948);
or U4128 (N_4128,N_3900,N_3936);
xor U4129 (N_4129,N_3860,N_3989);
nor U4130 (N_4130,N_3969,N_3973);
xor U4131 (N_4131,N_3810,N_3894);
or U4132 (N_4132,N_3856,N_3792);
and U4133 (N_4133,N_3935,N_3772);
nor U4134 (N_4134,N_3829,N_3898);
or U4135 (N_4135,N_3978,N_3769);
nand U4136 (N_4136,N_3864,N_3895);
or U4137 (N_4137,N_3770,N_3750);
xnor U4138 (N_4138,N_3845,N_3814);
nor U4139 (N_4139,N_3858,N_3939);
nor U4140 (N_4140,N_3875,N_3882);
or U4141 (N_4141,N_3788,N_3993);
xor U4142 (N_4142,N_3991,N_3850);
xor U4143 (N_4143,N_3799,N_3864);
nand U4144 (N_4144,N_3813,N_3969);
nand U4145 (N_4145,N_3786,N_3911);
nand U4146 (N_4146,N_3991,N_3916);
and U4147 (N_4147,N_3880,N_3763);
and U4148 (N_4148,N_3785,N_3919);
nand U4149 (N_4149,N_3754,N_3952);
and U4150 (N_4150,N_3819,N_3771);
and U4151 (N_4151,N_3867,N_3911);
nor U4152 (N_4152,N_3778,N_3794);
or U4153 (N_4153,N_3773,N_3983);
nand U4154 (N_4154,N_3990,N_3931);
and U4155 (N_4155,N_3949,N_3923);
nor U4156 (N_4156,N_3830,N_3894);
and U4157 (N_4157,N_3843,N_3801);
and U4158 (N_4158,N_3978,N_3850);
xnor U4159 (N_4159,N_3962,N_3905);
nand U4160 (N_4160,N_3990,N_3942);
xnor U4161 (N_4161,N_3889,N_3909);
and U4162 (N_4162,N_3991,N_3794);
xnor U4163 (N_4163,N_3997,N_3827);
and U4164 (N_4164,N_3803,N_3892);
nor U4165 (N_4165,N_3779,N_3998);
nor U4166 (N_4166,N_3783,N_3863);
or U4167 (N_4167,N_3947,N_3891);
or U4168 (N_4168,N_3873,N_3849);
or U4169 (N_4169,N_3995,N_3890);
xnor U4170 (N_4170,N_3956,N_3976);
nor U4171 (N_4171,N_3955,N_3949);
nor U4172 (N_4172,N_3940,N_3793);
xor U4173 (N_4173,N_3861,N_3967);
xnor U4174 (N_4174,N_3910,N_3893);
xnor U4175 (N_4175,N_3888,N_3821);
nor U4176 (N_4176,N_3786,N_3893);
nor U4177 (N_4177,N_3775,N_3877);
or U4178 (N_4178,N_3829,N_3882);
nor U4179 (N_4179,N_3949,N_3881);
nor U4180 (N_4180,N_3971,N_3799);
xnor U4181 (N_4181,N_3899,N_3828);
nor U4182 (N_4182,N_3859,N_3873);
xnor U4183 (N_4183,N_3840,N_3843);
nor U4184 (N_4184,N_3855,N_3859);
nand U4185 (N_4185,N_3899,N_3879);
nand U4186 (N_4186,N_3755,N_3992);
or U4187 (N_4187,N_3948,N_3968);
nor U4188 (N_4188,N_3882,N_3899);
nand U4189 (N_4189,N_3776,N_3940);
xor U4190 (N_4190,N_3857,N_3949);
and U4191 (N_4191,N_3825,N_3797);
nor U4192 (N_4192,N_3872,N_3959);
xor U4193 (N_4193,N_3911,N_3845);
or U4194 (N_4194,N_3809,N_3774);
nand U4195 (N_4195,N_3997,N_3918);
xnor U4196 (N_4196,N_3774,N_3833);
or U4197 (N_4197,N_3905,N_3776);
and U4198 (N_4198,N_3945,N_3968);
or U4199 (N_4199,N_3849,N_3927);
or U4200 (N_4200,N_3933,N_3762);
xor U4201 (N_4201,N_3777,N_3874);
or U4202 (N_4202,N_3811,N_3784);
xnor U4203 (N_4203,N_3826,N_3987);
nand U4204 (N_4204,N_3837,N_3847);
and U4205 (N_4205,N_3812,N_3962);
xnor U4206 (N_4206,N_3932,N_3946);
and U4207 (N_4207,N_3862,N_3790);
xnor U4208 (N_4208,N_3891,N_3872);
or U4209 (N_4209,N_3882,N_3815);
or U4210 (N_4210,N_3963,N_3844);
or U4211 (N_4211,N_3752,N_3920);
nand U4212 (N_4212,N_3869,N_3944);
xnor U4213 (N_4213,N_3897,N_3952);
nor U4214 (N_4214,N_3939,N_3818);
xnor U4215 (N_4215,N_3824,N_3861);
nand U4216 (N_4216,N_3798,N_3861);
and U4217 (N_4217,N_3991,N_3873);
nor U4218 (N_4218,N_3826,N_3838);
or U4219 (N_4219,N_3778,N_3872);
xor U4220 (N_4220,N_3851,N_3850);
nor U4221 (N_4221,N_3762,N_3922);
xor U4222 (N_4222,N_3968,N_3766);
nor U4223 (N_4223,N_3912,N_3889);
nand U4224 (N_4224,N_3777,N_3753);
nor U4225 (N_4225,N_3933,N_3751);
nand U4226 (N_4226,N_3821,N_3948);
nand U4227 (N_4227,N_3761,N_3943);
xnor U4228 (N_4228,N_3835,N_3861);
nor U4229 (N_4229,N_3924,N_3793);
nor U4230 (N_4230,N_3912,N_3901);
nand U4231 (N_4231,N_3844,N_3830);
xnor U4232 (N_4232,N_3956,N_3904);
or U4233 (N_4233,N_3892,N_3936);
and U4234 (N_4234,N_3829,N_3915);
or U4235 (N_4235,N_3935,N_3810);
or U4236 (N_4236,N_3944,N_3859);
nand U4237 (N_4237,N_3889,N_3844);
nor U4238 (N_4238,N_3866,N_3797);
xnor U4239 (N_4239,N_3770,N_3795);
nor U4240 (N_4240,N_3783,N_3908);
nand U4241 (N_4241,N_3791,N_3932);
xnor U4242 (N_4242,N_3797,N_3856);
nand U4243 (N_4243,N_3787,N_3980);
xor U4244 (N_4244,N_3978,N_3939);
and U4245 (N_4245,N_3784,N_3968);
nand U4246 (N_4246,N_3887,N_3883);
nand U4247 (N_4247,N_3852,N_3901);
nor U4248 (N_4248,N_3869,N_3926);
nand U4249 (N_4249,N_3967,N_3924);
xor U4250 (N_4250,N_4065,N_4133);
and U4251 (N_4251,N_4075,N_4022);
nand U4252 (N_4252,N_4063,N_4123);
and U4253 (N_4253,N_4197,N_4113);
xnor U4254 (N_4254,N_4137,N_4024);
and U4255 (N_4255,N_4033,N_4213);
nand U4256 (N_4256,N_4232,N_4187);
xnor U4257 (N_4257,N_4115,N_4010);
nor U4258 (N_4258,N_4122,N_4249);
xnor U4259 (N_4259,N_4156,N_4009);
nand U4260 (N_4260,N_4028,N_4098);
xor U4261 (N_4261,N_4214,N_4068);
nand U4262 (N_4262,N_4179,N_4185);
nand U4263 (N_4263,N_4078,N_4038);
xnor U4264 (N_4264,N_4086,N_4231);
or U4265 (N_4265,N_4008,N_4170);
and U4266 (N_4266,N_4007,N_4158);
xnor U4267 (N_4267,N_4169,N_4029);
or U4268 (N_4268,N_4106,N_4043);
nor U4269 (N_4269,N_4202,N_4215);
or U4270 (N_4270,N_4077,N_4200);
and U4271 (N_4271,N_4094,N_4136);
or U4272 (N_4272,N_4027,N_4092);
and U4273 (N_4273,N_4168,N_4052);
xnor U4274 (N_4274,N_4049,N_4247);
xnor U4275 (N_4275,N_4045,N_4109);
nand U4276 (N_4276,N_4039,N_4066);
and U4277 (N_4277,N_4223,N_4129);
or U4278 (N_4278,N_4153,N_4199);
nor U4279 (N_4279,N_4100,N_4054);
xor U4280 (N_4280,N_4062,N_4084);
xnor U4281 (N_4281,N_4093,N_4001);
nor U4282 (N_4282,N_4212,N_4099);
nor U4283 (N_4283,N_4015,N_4221);
nor U4284 (N_4284,N_4198,N_4102);
and U4285 (N_4285,N_4083,N_4161);
xor U4286 (N_4286,N_4004,N_4245);
nor U4287 (N_4287,N_4021,N_4151);
or U4288 (N_4288,N_4030,N_4186);
xnor U4289 (N_4289,N_4103,N_4229);
nor U4290 (N_4290,N_4206,N_4055);
nor U4291 (N_4291,N_4205,N_4108);
or U4292 (N_4292,N_4116,N_4165);
or U4293 (N_4293,N_4160,N_4163);
nand U4294 (N_4294,N_4020,N_4090);
nand U4295 (N_4295,N_4117,N_4145);
nand U4296 (N_4296,N_4208,N_4070);
nand U4297 (N_4297,N_4183,N_4047);
and U4298 (N_4298,N_4016,N_4104);
nand U4299 (N_4299,N_4235,N_4152);
or U4300 (N_4300,N_4142,N_4141);
xnor U4301 (N_4301,N_4224,N_4162);
or U4302 (N_4302,N_4079,N_4041);
or U4303 (N_4303,N_4080,N_4059);
xor U4304 (N_4304,N_4210,N_4037);
nor U4305 (N_4305,N_4204,N_4191);
nand U4306 (N_4306,N_4087,N_4225);
and U4307 (N_4307,N_4032,N_4174);
or U4308 (N_4308,N_4167,N_4000);
and U4309 (N_4309,N_4173,N_4110);
nor U4310 (N_4310,N_4230,N_4005);
or U4311 (N_4311,N_4073,N_4124);
nor U4312 (N_4312,N_4177,N_4067);
xor U4313 (N_4313,N_4201,N_4154);
or U4314 (N_4314,N_4132,N_4234);
nor U4315 (N_4315,N_4155,N_4175);
nor U4316 (N_4316,N_4040,N_4074);
and U4317 (N_4317,N_4188,N_4112);
or U4318 (N_4318,N_4081,N_4226);
nand U4319 (N_4319,N_4061,N_4166);
nand U4320 (N_4320,N_4120,N_4207);
and U4321 (N_4321,N_4196,N_4237);
nor U4322 (N_4322,N_4134,N_4118);
and U4323 (N_4323,N_4219,N_4222);
and U4324 (N_4324,N_4216,N_4144);
nor U4325 (N_4325,N_4189,N_4042);
nand U4326 (N_4326,N_4126,N_4046);
nand U4327 (N_4327,N_4119,N_4050);
xor U4328 (N_4328,N_4239,N_4044);
nand U4329 (N_4329,N_4060,N_4051);
or U4330 (N_4330,N_4082,N_4148);
nor U4331 (N_4331,N_4178,N_4088);
and U4332 (N_4332,N_4026,N_4019);
and U4333 (N_4333,N_4105,N_4233);
or U4334 (N_4334,N_4071,N_4125);
xnor U4335 (N_4335,N_4064,N_4171);
or U4336 (N_4336,N_4149,N_4036);
or U4337 (N_4337,N_4012,N_4180);
xor U4338 (N_4338,N_4246,N_4243);
and U4339 (N_4339,N_4031,N_4157);
xor U4340 (N_4340,N_4017,N_4211);
nor U4341 (N_4341,N_4018,N_4035);
nor U4342 (N_4342,N_4227,N_4218);
nand U4343 (N_4343,N_4182,N_4184);
and U4344 (N_4344,N_4193,N_4056);
xor U4345 (N_4345,N_4244,N_4135);
nand U4346 (N_4346,N_4013,N_4076);
nor U4347 (N_4347,N_4069,N_4128);
xor U4348 (N_4348,N_4101,N_4192);
and U4349 (N_4349,N_4023,N_4114);
xor U4350 (N_4350,N_4236,N_4002);
nand U4351 (N_4351,N_4238,N_4057);
and U4352 (N_4352,N_4209,N_4091);
xor U4353 (N_4353,N_4034,N_4127);
nand U4354 (N_4354,N_4089,N_4217);
and U4355 (N_4355,N_4195,N_4140);
xor U4356 (N_4356,N_4097,N_4048);
and U4357 (N_4357,N_4248,N_4181);
xnor U4358 (N_4358,N_4025,N_4203);
and U4359 (N_4359,N_4190,N_4150);
xor U4360 (N_4360,N_4096,N_4228);
nand U4361 (N_4361,N_4130,N_4014);
nor U4362 (N_4362,N_4085,N_4241);
nand U4363 (N_4363,N_4147,N_4107);
nand U4364 (N_4364,N_4164,N_4006);
or U4365 (N_4365,N_4194,N_4011);
nand U4366 (N_4366,N_4111,N_4138);
xnor U4367 (N_4367,N_4146,N_4159);
or U4368 (N_4368,N_4172,N_4220);
xor U4369 (N_4369,N_4058,N_4176);
nand U4370 (N_4370,N_4240,N_4121);
nor U4371 (N_4371,N_4072,N_4242);
and U4372 (N_4372,N_4143,N_4095);
xor U4373 (N_4373,N_4003,N_4053);
and U4374 (N_4374,N_4131,N_4139);
nor U4375 (N_4375,N_4017,N_4021);
nor U4376 (N_4376,N_4042,N_4109);
or U4377 (N_4377,N_4151,N_4205);
and U4378 (N_4378,N_4169,N_4067);
nor U4379 (N_4379,N_4041,N_4045);
nor U4380 (N_4380,N_4076,N_4056);
xor U4381 (N_4381,N_4191,N_4007);
nand U4382 (N_4382,N_4205,N_4206);
nand U4383 (N_4383,N_4026,N_4240);
and U4384 (N_4384,N_4043,N_4114);
or U4385 (N_4385,N_4141,N_4216);
xnor U4386 (N_4386,N_4150,N_4167);
nor U4387 (N_4387,N_4223,N_4236);
nand U4388 (N_4388,N_4012,N_4198);
xor U4389 (N_4389,N_4179,N_4096);
nand U4390 (N_4390,N_4121,N_4234);
and U4391 (N_4391,N_4187,N_4213);
nor U4392 (N_4392,N_4130,N_4142);
or U4393 (N_4393,N_4147,N_4171);
or U4394 (N_4394,N_4085,N_4144);
nand U4395 (N_4395,N_4075,N_4052);
nand U4396 (N_4396,N_4234,N_4129);
nand U4397 (N_4397,N_4028,N_4122);
and U4398 (N_4398,N_4055,N_4001);
or U4399 (N_4399,N_4093,N_4120);
nand U4400 (N_4400,N_4141,N_4203);
and U4401 (N_4401,N_4084,N_4091);
or U4402 (N_4402,N_4034,N_4198);
nand U4403 (N_4403,N_4008,N_4182);
and U4404 (N_4404,N_4094,N_4182);
and U4405 (N_4405,N_4216,N_4011);
and U4406 (N_4406,N_4155,N_4035);
or U4407 (N_4407,N_4145,N_4058);
xnor U4408 (N_4408,N_4063,N_4210);
xnor U4409 (N_4409,N_4048,N_4195);
nor U4410 (N_4410,N_4102,N_4158);
and U4411 (N_4411,N_4063,N_4083);
or U4412 (N_4412,N_4118,N_4055);
nor U4413 (N_4413,N_4234,N_4091);
and U4414 (N_4414,N_4094,N_4164);
xnor U4415 (N_4415,N_4015,N_4235);
nor U4416 (N_4416,N_4161,N_4160);
nor U4417 (N_4417,N_4079,N_4143);
and U4418 (N_4418,N_4045,N_4134);
nor U4419 (N_4419,N_4132,N_4005);
or U4420 (N_4420,N_4143,N_4085);
or U4421 (N_4421,N_4092,N_4043);
or U4422 (N_4422,N_4187,N_4170);
nand U4423 (N_4423,N_4064,N_4188);
xor U4424 (N_4424,N_4072,N_4039);
xor U4425 (N_4425,N_4134,N_4235);
nand U4426 (N_4426,N_4047,N_4155);
and U4427 (N_4427,N_4066,N_4055);
or U4428 (N_4428,N_4132,N_4225);
or U4429 (N_4429,N_4168,N_4220);
nor U4430 (N_4430,N_4087,N_4220);
and U4431 (N_4431,N_4168,N_4153);
and U4432 (N_4432,N_4020,N_4218);
xnor U4433 (N_4433,N_4076,N_4011);
nand U4434 (N_4434,N_4001,N_4002);
nand U4435 (N_4435,N_4084,N_4199);
or U4436 (N_4436,N_4214,N_4233);
nand U4437 (N_4437,N_4155,N_4150);
or U4438 (N_4438,N_4206,N_4190);
nand U4439 (N_4439,N_4038,N_4015);
nor U4440 (N_4440,N_4133,N_4103);
nor U4441 (N_4441,N_4134,N_4040);
xor U4442 (N_4442,N_4189,N_4237);
or U4443 (N_4443,N_4243,N_4003);
and U4444 (N_4444,N_4091,N_4129);
nand U4445 (N_4445,N_4175,N_4013);
nor U4446 (N_4446,N_4090,N_4200);
or U4447 (N_4447,N_4147,N_4034);
and U4448 (N_4448,N_4064,N_4108);
and U4449 (N_4449,N_4094,N_4194);
nor U4450 (N_4450,N_4098,N_4062);
xnor U4451 (N_4451,N_4028,N_4181);
xor U4452 (N_4452,N_4140,N_4154);
and U4453 (N_4453,N_4237,N_4229);
nor U4454 (N_4454,N_4016,N_4145);
nor U4455 (N_4455,N_4164,N_4029);
xnor U4456 (N_4456,N_4093,N_4097);
nand U4457 (N_4457,N_4072,N_4149);
xor U4458 (N_4458,N_4066,N_4131);
nor U4459 (N_4459,N_4148,N_4170);
and U4460 (N_4460,N_4052,N_4000);
nor U4461 (N_4461,N_4181,N_4161);
and U4462 (N_4462,N_4132,N_4242);
or U4463 (N_4463,N_4047,N_4163);
nor U4464 (N_4464,N_4227,N_4131);
or U4465 (N_4465,N_4053,N_4222);
xnor U4466 (N_4466,N_4244,N_4101);
nor U4467 (N_4467,N_4162,N_4068);
nor U4468 (N_4468,N_4050,N_4177);
xor U4469 (N_4469,N_4229,N_4174);
xnor U4470 (N_4470,N_4042,N_4184);
and U4471 (N_4471,N_4098,N_4017);
nand U4472 (N_4472,N_4159,N_4139);
nor U4473 (N_4473,N_4106,N_4065);
nand U4474 (N_4474,N_4199,N_4197);
nor U4475 (N_4475,N_4114,N_4214);
nor U4476 (N_4476,N_4106,N_4152);
nand U4477 (N_4477,N_4181,N_4243);
xor U4478 (N_4478,N_4232,N_4210);
nor U4479 (N_4479,N_4028,N_4172);
nand U4480 (N_4480,N_4036,N_4027);
nor U4481 (N_4481,N_4102,N_4173);
nor U4482 (N_4482,N_4060,N_4148);
and U4483 (N_4483,N_4164,N_4180);
xor U4484 (N_4484,N_4214,N_4029);
nand U4485 (N_4485,N_4139,N_4033);
nand U4486 (N_4486,N_4131,N_4191);
or U4487 (N_4487,N_4161,N_4184);
nor U4488 (N_4488,N_4145,N_4244);
nand U4489 (N_4489,N_4151,N_4123);
and U4490 (N_4490,N_4144,N_4108);
nor U4491 (N_4491,N_4141,N_4190);
xnor U4492 (N_4492,N_4216,N_4197);
nor U4493 (N_4493,N_4145,N_4028);
and U4494 (N_4494,N_4028,N_4042);
and U4495 (N_4495,N_4077,N_4083);
nor U4496 (N_4496,N_4124,N_4064);
xor U4497 (N_4497,N_4131,N_4244);
nor U4498 (N_4498,N_4120,N_4102);
nand U4499 (N_4499,N_4175,N_4248);
xor U4500 (N_4500,N_4482,N_4311);
and U4501 (N_4501,N_4451,N_4260);
nand U4502 (N_4502,N_4338,N_4373);
or U4503 (N_4503,N_4292,N_4360);
nor U4504 (N_4504,N_4405,N_4348);
nand U4505 (N_4505,N_4316,N_4267);
nand U4506 (N_4506,N_4328,N_4284);
nand U4507 (N_4507,N_4349,N_4372);
or U4508 (N_4508,N_4460,N_4361);
or U4509 (N_4509,N_4462,N_4371);
nor U4510 (N_4510,N_4445,N_4422);
nand U4511 (N_4511,N_4484,N_4258);
nand U4512 (N_4512,N_4305,N_4357);
nand U4513 (N_4513,N_4329,N_4404);
or U4514 (N_4514,N_4254,N_4483);
nor U4515 (N_4515,N_4307,N_4488);
xnor U4516 (N_4516,N_4467,N_4256);
xor U4517 (N_4517,N_4436,N_4417);
nand U4518 (N_4518,N_4286,N_4326);
nor U4519 (N_4519,N_4374,N_4293);
xor U4520 (N_4520,N_4476,N_4344);
nand U4521 (N_4521,N_4410,N_4345);
or U4522 (N_4522,N_4275,N_4428);
nand U4523 (N_4523,N_4498,N_4319);
and U4524 (N_4524,N_4459,N_4423);
nor U4525 (N_4525,N_4474,N_4489);
nand U4526 (N_4526,N_4418,N_4487);
nor U4527 (N_4527,N_4415,N_4313);
xnor U4528 (N_4528,N_4339,N_4294);
xor U4529 (N_4529,N_4325,N_4296);
nand U4530 (N_4530,N_4271,N_4407);
nand U4531 (N_4531,N_4340,N_4471);
nor U4532 (N_4532,N_4438,N_4359);
nand U4533 (N_4533,N_4479,N_4493);
or U4534 (N_4534,N_4457,N_4495);
and U4535 (N_4535,N_4285,N_4282);
nand U4536 (N_4536,N_4385,N_4367);
nand U4537 (N_4537,N_4399,N_4320);
and U4538 (N_4538,N_4424,N_4272);
or U4539 (N_4539,N_4448,N_4321);
and U4540 (N_4540,N_4295,N_4492);
xor U4541 (N_4541,N_4401,N_4446);
and U4542 (N_4542,N_4412,N_4378);
xnor U4543 (N_4543,N_4432,N_4334);
or U4544 (N_4544,N_4261,N_4465);
nor U4545 (N_4545,N_4379,N_4290);
and U4546 (N_4546,N_4420,N_4281);
nor U4547 (N_4547,N_4381,N_4337);
or U4548 (N_4548,N_4433,N_4478);
xor U4549 (N_4549,N_4464,N_4439);
or U4550 (N_4550,N_4306,N_4300);
xnor U4551 (N_4551,N_4310,N_4312);
nor U4552 (N_4552,N_4252,N_4463);
and U4553 (N_4553,N_4335,N_4315);
or U4554 (N_4554,N_4341,N_4461);
and U4555 (N_4555,N_4499,N_4481);
nor U4556 (N_4556,N_4416,N_4389);
nor U4557 (N_4557,N_4347,N_4466);
and U4558 (N_4558,N_4273,N_4301);
xor U4559 (N_4559,N_4473,N_4431);
xnor U4560 (N_4560,N_4332,N_4317);
nand U4561 (N_4561,N_4266,N_4425);
xnor U4562 (N_4562,N_4283,N_4268);
and U4563 (N_4563,N_4322,N_4350);
xor U4564 (N_4564,N_4270,N_4323);
nor U4565 (N_4565,N_4409,N_4362);
and U4566 (N_4566,N_4398,N_4278);
nor U4567 (N_4567,N_4336,N_4343);
nand U4568 (N_4568,N_4396,N_4355);
xor U4569 (N_4569,N_4490,N_4388);
nor U4570 (N_4570,N_4414,N_4299);
or U4571 (N_4571,N_4452,N_4380);
and U4572 (N_4572,N_4351,N_4429);
nand U4573 (N_4573,N_4434,N_4253);
xnor U4574 (N_4574,N_4472,N_4437);
or U4575 (N_4575,N_4314,N_4365);
xnor U4576 (N_4576,N_4382,N_4370);
or U4577 (N_4577,N_4443,N_4475);
and U4578 (N_4578,N_4368,N_4358);
nand U4579 (N_4579,N_4318,N_4411);
or U4580 (N_4580,N_4386,N_4259);
nor U4581 (N_4581,N_4387,N_4375);
and U4582 (N_4582,N_4384,N_4455);
or U4583 (N_4583,N_4469,N_4377);
xnor U4584 (N_4584,N_4397,N_4257);
nor U4585 (N_4585,N_4400,N_4291);
nand U4586 (N_4586,N_4426,N_4251);
nand U4587 (N_4587,N_4262,N_4255);
xor U4588 (N_4588,N_4480,N_4264);
or U4589 (N_4589,N_4496,N_4406);
xor U4590 (N_4590,N_4441,N_4279);
or U4591 (N_4591,N_4304,N_4468);
xor U4592 (N_4592,N_4477,N_4250);
xnor U4593 (N_4593,N_4390,N_4453);
nor U4594 (N_4594,N_4430,N_4308);
or U4595 (N_4595,N_4427,N_4444);
xor U4596 (N_4596,N_4302,N_4280);
and U4597 (N_4597,N_4376,N_4383);
xnor U4598 (N_4598,N_4485,N_4298);
or U4599 (N_4599,N_4470,N_4276);
or U4600 (N_4600,N_4408,N_4413);
and U4601 (N_4601,N_4277,N_4440);
and U4602 (N_4602,N_4352,N_4419);
nor U4603 (N_4603,N_4364,N_4297);
nor U4604 (N_4604,N_4342,N_4442);
or U4605 (N_4605,N_4309,N_4393);
xor U4606 (N_4606,N_4402,N_4288);
and U4607 (N_4607,N_4403,N_4353);
and U4608 (N_4608,N_4327,N_4274);
or U4609 (N_4609,N_4287,N_4486);
nand U4610 (N_4610,N_4369,N_4421);
and U4611 (N_4611,N_4324,N_4263);
nor U4612 (N_4612,N_4391,N_4435);
and U4613 (N_4613,N_4491,N_4331);
xor U4614 (N_4614,N_4449,N_4447);
and U4615 (N_4615,N_4333,N_4269);
nor U4616 (N_4616,N_4303,N_4366);
nor U4617 (N_4617,N_4497,N_4394);
and U4618 (N_4618,N_4494,N_4330);
and U4619 (N_4619,N_4346,N_4395);
xor U4620 (N_4620,N_4450,N_4356);
or U4621 (N_4621,N_4456,N_4265);
xnor U4622 (N_4622,N_4363,N_4354);
nand U4623 (N_4623,N_4458,N_4454);
xor U4624 (N_4624,N_4289,N_4392);
nand U4625 (N_4625,N_4414,N_4475);
xnor U4626 (N_4626,N_4386,N_4446);
and U4627 (N_4627,N_4368,N_4263);
xor U4628 (N_4628,N_4495,N_4358);
and U4629 (N_4629,N_4476,N_4352);
and U4630 (N_4630,N_4331,N_4478);
or U4631 (N_4631,N_4369,N_4351);
nand U4632 (N_4632,N_4395,N_4414);
nand U4633 (N_4633,N_4403,N_4380);
or U4634 (N_4634,N_4336,N_4411);
nor U4635 (N_4635,N_4465,N_4253);
or U4636 (N_4636,N_4362,N_4444);
and U4637 (N_4637,N_4435,N_4367);
or U4638 (N_4638,N_4372,N_4348);
or U4639 (N_4639,N_4379,N_4326);
and U4640 (N_4640,N_4452,N_4396);
xor U4641 (N_4641,N_4412,N_4263);
xor U4642 (N_4642,N_4372,N_4461);
or U4643 (N_4643,N_4275,N_4415);
nand U4644 (N_4644,N_4355,N_4412);
xor U4645 (N_4645,N_4277,N_4363);
xor U4646 (N_4646,N_4406,N_4349);
nor U4647 (N_4647,N_4384,N_4280);
or U4648 (N_4648,N_4270,N_4271);
nor U4649 (N_4649,N_4337,N_4312);
xnor U4650 (N_4650,N_4353,N_4420);
and U4651 (N_4651,N_4343,N_4310);
xor U4652 (N_4652,N_4371,N_4280);
nor U4653 (N_4653,N_4292,N_4490);
and U4654 (N_4654,N_4308,N_4490);
or U4655 (N_4655,N_4498,N_4317);
nor U4656 (N_4656,N_4394,N_4467);
or U4657 (N_4657,N_4250,N_4493);
xnor U4658 (N_4658,N_4352,N_4300);
xnor U4659 (N_4659,N_4382,N_4427);
nand U4660 (N_4660,N_4460,N_4459);
and U4661 (N_4661,N_4473,N_4254);
or U4662 (N_4662,N_4480,N_4451);
or U4663 (N_4663,N_4421,N_4278);
nor U4664 (N_4664,N_4349,N_4399);
nor U4665 (N_4665,N_4312,N_4413);
and U4666 (N_4666,N_4326,N_4396);
xnor U4667 (N_4667,N_4436,N_4353);
nand U4668 (N_4668,N_4363,N_4343);
or U4669 (N_4669,N_4452,N_4281);
or U4670 (N_4670,N_4418,N_4440);
nor U4671 (N_4671,N_4387,N_4418);
and U4672 (N_4672,N_4325,N_4254);
and U4673 (N_4673,N_4260,N_4397);
and U4674 (N_4674,N_4362,N_4342);
or U4675 (N_4675,N_4346,N_4382);
and U4676 (N_4676,N_4371,N_4392);
and U4677 (N_4677,N_4392,N_4399);
or U4678 (N_4678,N_4414,N_4419);
xnor U4679 (N_4679,N_4281,N_4448);
xor U4680 (N_4680,N_4425,N_4267);
or U4681 (N_4681,N_4455,N_4462);
nor U4682 (N_4682,N_4270,N_4263);
or U4683 (N_4683,N_4316,N_4436);
or U4684 (N_4684,N_4368,N_4408);
and U4685 (N_4685,N_4445,N_4305);
xnor U4686 (N_4686,N_4372,N_4354);
nand U4687 (N_4687,N_4494,N_4274);
and U4688 (N_4688,N_4301,N_4366);
xnor U4689 (N_4689,N_4425,N_4343);
or U4690 (N_4690,N_4422,N_4481);
nand U4691 (N_4691,N_4404,N_4298);
nor U4692 (N_4692,N_4483,N_4357);
or U4693 (N_4693,N_4419,N_4491);
nand U4694 (N_4694,N_4371,N_4428);
and U4695 (N_4695,N_4340,N_4339);
nor U4696 (N_4696,N_4271,N_4481);
xnor U4697 (N_4697,N_4335,N_4342);
or U4698 (N_4698,N_4347,N_4274);
xnor U4699 (N_4699,N_4306,N_4362);
nor U4700 (N_4700,N_4430,N_4429);
nand U4701 (N_4701,N_4295,N_4426);
or U4702 (N_4702,N_4292,N_4387);
nor U4703 (N_4703,N_4372,N_4306);
xor U4704 (N_4704,N_4481,N_4328);
xnor U4705 (N_4705,N_4498,N_4460);
and U4706 (N_4706,N_4438,N_4447);
xor U4707 (N_4707,N_4314,N_4400);
nand U4708 (N_4708,N_4395,N_4307);
and U4709 (N_4709,N_4418,N_4398);
and U4710 (N_4710,N_4392,N_4327);
nand U4711 (N_4711,N_4298,N_4365);
or U4712 (N_4712,N_4454,N_4376);
xnor U4713 (N_4713,N_4338,N_4366);
nor U4714 (N_4714,N_4295,N_4460);
or U4715 (N_4715,N_4425,N_4323);
or U4716 (N_4716,N_4258,N_4435);
or U4717 (N_4717,N_4411,N_4373);
xnor U4718 (N_4718,N_4323,N_4302);
nand U4719 (N_4719,N_4447,N_4371);
xor U4720 (N_4720,N_4398,N_4498);
xor U4721 (N_4721,N_4388,N_4323);
xnor U4722 (N_4722,N_4393,N_4476);
or U4723 (N_4723,N_4314,N_4288);
nand U4724 (N_4724,N_4442,N_4374);
xnor U4725 (N_4725,N_4364,N_4427);
or U4726 (N_4726,N_4449,N_4300);
and U4727 (N_4727,N_4332,N_4402);
xor U4728 (N_4728,N_4296,N_4361);
and U4729 (N_4729,N_4481,N_4287);
nand U4730 (N_4730,N_4481,N_4463);
nand U4731 (N_4731,N_4453,N_4430);
and U4732 (N_4732,N_4427,N_4366);
or U4733 (N_4733,N_4406,N_4495);
nor U4734 (N_4734,N_4468,N_4318);
nand U4735 (N_4735,N_4401,N_4254);
xor U4736 (N_4736,N_4380,N_4329);
and U4737 (N_4737,N_4344,N_4345);
nand U4738 (N_4738,N_4319,N_4418);
and U4739 (N_4739,N_4260,N_4464);
nand U4740 (N_4740,N_4418,N_4497);
nand U4741 (N_4741,N_4382,N_4405);
nor U4742 (N_4742,N_4333,N_4426);
nor U4743 (N_4743,N_4355,N_4381);
and U4744 (N_4744,N_4481,N_4424);
and U4745 (N_4745,N_4341,N_4369);
xor U4746 (N_4746,N_4268,N_4444);
or U4747 (N_4747,N_4496,N_4483);
xnor U4748 (N_4748,N_4387,N_4400);
nor U4749 (N_4749,N_4483,N_4477);
nor U4750 (N_4750,N_4557,N_4659);
and U4751 (N_4751,N_4649,N_4542);
xnor U4752 (N_4752,N_4566,N_4505);
nor U4753 (N_4753,N_4722,N_4726);
and U4754 (N_4754,N_4691,N_4708);
nor U4755 (N_4755,N_4547,N_4635);
xor U4756 (N_4756,N_4616,N_4551);
nor U4757 (N_4757,N_4657,N_4514);
xor U4758 (N_4758,N_4590,N_4730);
or U4759 (N_4759,N_4548,N_4723);
and U4760 (N_4760,N_4503,N_4540);
nor U4761 (N_4761,N_4625,N_4507);
nor U4762 (N_4762,N_4592,N_4633);
nand U4763 (N_4763,N_4574,N_4519);
or U4764 (N_4764,N_4604,N_4553);
nand U4765 (N_4765,N_4710,N_4586);
xor U4766 (N_4766,N_4632,N_4599);
or U4767 (N_4767,N_4588,N_4546);
nand U4768 (N_4768,N_4563,N_4677);
xnor U4769 (N_4769,N_4602,N_4748);
nand U4770 (N_4770,N_4567,N_4569);
nand U4771 (N_4771,N_4544,N_4713);
xor U4772 (N_4772,N_4656,N_4734);
nand U4773 (N_4773,N_4741,N_4539);
and U4774 (N_4774,N_4683,N_4728);
nand U4775 (N_4775,N_4512,N_4623);
and U4776 (N_4776,N_4528,N_4582);
or U4777 (N_4777,N_4555,N_4585);
nor U4778 (N_4778,N_4606,N_4716);
or U4779 (N_4779,N_4596,N_4502);
nand U4780 (N_4780,N_4605,N_4591);
and U4781 (N_4781,N_4711,N_4721);
or U4782 (N_4782,N_4676,N_4534);
xor U4783 (N_4783,N_4682,N_4658);
nor U4784 (N_4784,N_4646,N_4614);
xnor U4785 (N_4785,N_4529,N_4535);
nor U4786 (N_4786,N_4638,N_4583);
nand U4787 (N_4787,N_4695,N_4712);
or U4788 (N_4788,N_4675,N_4501);
or U4789 (N_4789,N_4550,N_4667);
xnor U4790 (N_4790,N_4742,N_4527);
xor U4791 (N_4791,N_4690,N_4597);
nor U4792 (N_4792,N_4747,N_4580);
xnor U4793 (N_4793,N_4593,N_4576);
or U4794 (N_4794,N_4707,N_4500);
nor U4795 (N_4795,N_4559,N_4587);
nand U4796 (N_4796,N_4626,N_4715);
nand U4797 (N_4797,N_4573,N_4686);
nand U4798 (N_4798,N_4729,N_4717);
nor U4799 (N_4799,N_4663,N_4692);
and U4800 (N_4800,N_4647,N_4669);
and U4801 (N_4801,N_4664,N_4584);
or U4802 (N_4802,N_4509,N_4738);
or U4803 (N_4803,N_4629,N_4680);
xnor U4804 (N_4804,N_4524,N_4517);
nand U4805 (N_4805,N_4615,N_4714);
and U4806 (N_4806,N_4654,N_4678);
nor U4807 (N_4807,N_4627,N_4624);
and U4808 (N_4808,N_4688,N_4732);
xor U4809 (N_4809,N_4526,N_4724);
and U4810 (N_4810,N_4725,N_4549);
nand U4811 (N_4811,N_4631,N_4653);
and U4812 (N_4812,N_4572,N_4685);
and U4813 (N_4813,N_4617,N_4666);
or U4814 (N_4814,N_4554,N_4508);
or U4815 (N_4815,N_4613,N_4515);
and U4816 (N_4816,N_4736,N_4518);
or U4817 (N_4817,N_4565,N_4536);
nand U4818 (N_4818,N_4608,N_4661);
nand U4819 (N_4819,N_4579,N_4578);
and U4820 (N_4820,N_4531,N_4668);
nand U4821 (N_4821,N_4611,N_4533);
nand U4822 (N_4822,N_4727,N_4739);
xor U4823 (N_4823,N_4621,N_4731);
xnor U4824 (N_4824,N_4581,N_4504);
xor U4825 (N_4825,N_4744,N_4709);
nand U4826 (N_4826,N_4648,N_4575);
nand U4827 (N_4827,N_4571,N_4705);
xor U4828 (N_4828,N_4543,N_4702);
nor U4829 (N_4829,N_4673,N_4640);
or U4830 (N_4830,N_4641,N_4639);
xor U4831 (N_4831,N_4525,N_4636);
and U4832 (N_4832,N_4718,N_4607);
nand U4833 (N_4833,N_4637,N_4630);
or U4834 (N_4834,N_4645,N_4589);
nor U4835 (N_4835,N_4516,N_4577);
xor U4836 (N_4836,N_4521,N_4552);
nand U4837 (N_4837,N_4693,N_4743);
xnor U4838 (N_4838,N_4749,N_4694);
or U4839 (N_4839,N_4520,N_4660);
or U4840 (N_4840,N_4541,N_4644);
xnor U4841 (N_4841,N_4684,N_4603);
or U4842 (N_4842,N_4701,N_4689);
nand U4843 (N_4843,N_4652,N_4687);
nand U4844 (N_4844,N_4532,N_4522);
or U4845 (N_4845,N_4619,N_4655);
or U4846 (N_4846,N_4530,N_4634);
nor U4847 (N_4847,N_4618,N_4538);
or U4848 (N_4848,N_4643,N_4506);
nor U4849 (N_4849,N_4601,N_4719);
nand U4850 (N_4850,N_4568,N_4700);
xnor U4851 (N_4851,N_4733,N_4513);
and U4852 (N_4852,N_4560,N_4697);
xor U4853 (N_4853,N_4679,N_4745);
and U4854 (N_4854,N_4703,N_4598);
nand U4855 (N_4855,N_4651,N_4564);
nor U4856 (N_4856,N_4510,N_4720);
nand U4857 (N_4857,N_4558,N_4698);
nor U4858 (N_4858,N_4523,N_4545);
nand U4859 (N_4859,N_4600,N_4746);
nor U4860 (N_4860,N_4612,N_4674);
and U4861 (N_4861,N_4672,N_4556);
xor U4862 (N_4862,N_4735,N_4595);
or U4863 (N_4863,N_4622,N_4699);
xnor U4864 (N_4864,N_4665,N_4704);
and U4865 (N_4865,N_4662,N_4610);
or U4866 (N_4866,N_4628,N_4681);
xor U4867 (N_4867,N_4609,N_4642);
nand U4868 (N_4868,N_4537,N_4670);
xor U4869 (N_4869,N_4671,N_4706);
and U4870 (N_4870,N_4737,N_4561);
xor U4871 (N_4871,N_4594,N_4650);
nand U4872 (N_4872,N_4562,N_4696);
and U4873 (N_4873,N_4511,N_4620);
and U4874 (N_4874,N_4570,N_4740);
nor U4875 (N_4875,N_4578,N_4656);
nor U4876 (N_4876,N_4556,N_4559);
or U4877 (N_4877,N_4589,N_4525);
xor U4878 (N_4878,N_4549,N_4705);
and U4879 (N_4879,N_4512,N_4515);
or U4880 (N_4880,N_4630,N_4599);
and U4881 (N_4881,N_4684,N_4580);
nand U4882 (N_4882,N_4566,N_4601);
nand U4883 (N_4883,N_4560,N_4527);
nor U4884 (N_4884,N_4595,N_4525);
nor U4885 (N_4885,N_4625,N_4577);
or U4886 (N_4886,N_4662,N_4507);
and U4887 (N_4887,N_4651,N_4590);
or U4888 (N_4888,N_4558,N_4655);
nand U4889 (N_4889,N_4734,N_4538);
xnor U4890 (N_4890,N_4516,N_4536);
or U4891 (N_4891,N_4555,N_4669);
nor U4892 (N_4892,N_4724,N_4506);
and U4893 (N_4893,N_4554,N_4603);
nor U4894 (N_4894,N_4676,N_4621);
and U4895 (N_4895,N_4676,N_4577);
nor U4896 (N_4896,N_4584,N_4558);
nor U4897 (N_4897,N_4705,N_4704);
nor U4898 (N_4898,N_4563,N_4601);
nor U4899 (N_4899,N_4720,N_4544);
and U4900 (N_4900,N_4714,N_4528);
xnor U4901 (N_4901,N_4562,N_4666);
nand U4902 (N_4902,N_4508,N_4704);
or U4903 (N_4903,N_4528,N_4583);
nand U4904 (N_4904,N_4520,N_4704);
nand U4905 (N_4905,N_4535,N_4583);
nor U4906 (N_4906,N_4527,N_4642);
or U4907 (N_4907,N_4719,N_4604);
or U4908 (N_4908,N_4666,N_4636);
nor U4909 (N_4909,N_4586,N_4564);
and U4910 (N_4910,N_4651,N_4610);
nand U4911 (N_4911,N_4542,N_4625);
xor U4912 (N_4912,N_4653,N_4502);
nand U4913 (N_4913,N_4648,N_4727);
nand U4914 (N_4914,N_4699,N_4687);
xnor U4915 (N_4915,N_4743,N_4641);
nand U4916 (N_4916,N_4634,N_4511);
xnor U4917 (N_4917,N_4523,N_4524);
xnor U4918 (N_4918,N_4688,N_4599);
nor U4919 (N_4919,N_4581,N_4602);
nand U4920 (N_4920,N_4632,N_4539);
or U4921 (N_4921,N_4584,N_4570);
nor U4922 (N_4922,N_4696,N_4549);
nor U4923 (N_4923,N_4556,N_4575);
xor U4924 (N_4924,N_4617,N_4714);
nand U4925 (N_4925,N_4656,N_4511);
nor U4926 (N_4926,N_4528,N_4696);
xnor U4927 (N_4927,N_4668,N_4698);
nor U4928 (N_4928,N_4716,N_4607);
nor U4929 (N_4929,N_4512,N_4704);
nand U4930 (N_4930,N_4620,N_4530);
nand U4931 (N_4931,N_4743,N_4529);
nand U4932 (N_4932,N_4652,N_4546);
nor U4933 (N_4933,N_4523,N_4697);
nand U4934 (N_4934,N_4731,N_4695);
and U4935 (N_4935,N_4512,N_4723);
xor U4936 (N_4936,N_4546,N_4523);
nand U4937 (N_4937,N_4650,N_4510);
and U4938 (N_4938,N_4727,N_4538);
and U4939 (N_4939,N_4627,N_4554);
nor U4940 (N_4940,N_4696,N_4500);
and U4941 (N_4941,N_4511,N_4584);
nand U4942 (N_4942,N_4520,N_4506);
nor U4943 (N_4943,N_4724,N_4720);
or U4944 (N_4944,N_4746,N_4565);
xor U4945 (N_4945,N_4518,N_4690);
nand U4946 (N_4946,N_4671,N_4719);
nand U4947 (N_4947,N_4583,N_4683);
xnor U4948 (N_4948,N_4535,N_4520);
and U4949 (N_4949,N_4526,N_4513);
nor U4950 (N_4950,N_4518,N_4705);
nand U4951 (N_4951,N_4511,N_4689);
and U4952 (N_4952,N_4734,N_4553);
or U4953 (N_4953,N_4542,N_4537);
and U4954 (N_4954,N_4636,N_4555);
nand U4955 (N_4955,N_4520,N_4563);
xor U4956 (N_4956,N_4711,N_4618);
nand U4957 (N_4957,N_4597,N_4626);
and U4958 (N_4958,N_4551,N_4722);
nor U4959 (N_4959,N_4657,N_4603);
xor U4960 (N_4960,N_4686,N_4636);
nand U4961 (N_4961,N_4522,N_4511);
nand U4962 (N_4962,N_4696,N_4659);
or U4963 (N_4963,N_4531,N_4630);
nand U4964 (N_4964,N_4685,N_4550);
nand U4965 (N_4965,N_4507,N_4747);
or U4966 (N_4966,N_4735,N_4671);
and U4967 (N_4967,N_4543,N_4549);
nand U4968 (N_4968,N_4633,N_4722);
or U4969 (N_4969,N_4524,N_4587);
nand U4970 (N_4970,N_4684,N_4701);
nand U4971 (N_4971,N_4653,N_4523);
or U4972 (N_4972,N_4581,N_4684);
and U4973 (N_4973,N_4525,N_4532);
xor U4974 (N_4974,N_4573,N_4719);
or U4975 (N_4975,N_4628,N_4740);
and U4976 (N_4976,N_4739,N_4641);
or U4977 (N_4977,N_4621,N_4604);
nor U4978 (N_4978,N_4570,N_4689);
and U4979 (N_4979,N_4698,N_4540);
and U4980 (N_4980,N_4650,N_4716);
nor U4981 (N_4981,N_4689,N_4521);
xnor U4982 (N_4982,N_4629,N_4646);
nor U4983 (N_4983,N_4571,N_4520);
nand U4984 (N_4984,N_4727,N_4710);
nand U4985 (N_4985,N_4582,N_4534);
nor U4986 (N_4986,N_4534,N_4616);
nor U4987 (N_4987,N_4605,N_4552);
nor U4988 (N_4988,N_4510,N_4597);
nand U4989 (N_4989,N_4573,N_4709);
and U4990 (N_4990,N_4664,N_4597);
nor U4991 (N_4991,N_4742,N_4614);
xnor U4992 (N_4992,N_4697,N_4511);
nand U4993 (N_4993,N_4530,N_4506);
or U4994 (N_4994,N_4611,N_4745);
and U4995 (N_4995,N_4562,N_4586);
or U4996 (N_4996,N_4602,N_4658);
and U4997 (N_4997,N_4678,N_4557);
xnor U4998 (N_4998,N_4521,N_4637);
xor U4999 (N_4999,N_4706,N_4551);
and U5000 (N_5000,N_4834,N_4825);
nor U5001 (N_5001,N_4975,N_4922);
nand U5002 (N_5002,N_4777,N_4978);
and U5003 (N_5003,N_4888,N_4788);
xnor U5004 (N_5004,N_4816,N_4915);
and U5005 (N_5005,N_4804,N_4833);
nor U5006 (N_5006,N_4895,N_4854);
or U5007 (N_5007,N_4862,N_4809);
nand U5008 (N_5008,N_4951,N_4972);
xor U5009 (N_5009,N_4892,N_4832);
nor U5010 (N_5010,N_4882,N_4756);
or U5011 (N_5011,N_4906,N_4750);
nand U5012 (N_5012,N_4931,N_4985);
nand U5013 (N_5013,N_4865,N_4878);
xor U5014 (N_5014,N_4838,N_4960);
and U5015 (N_5015,N_4797,N_4950);
nor U5016 (N_5016,N_4762,N_4904);
and U5017 (N_5017,N_4994,N_4940);
and U5018 (N_5018,N_4999,N_4856);
nor U5019 (N_5019,N_4844,N_4822);
and U5020 (N_5020,N_4925,N_4974);
or U5021 (N_5021,N_4840,N_4935);
and U5022 (N_5022,N_4875,N_4775);
xnor U5023 (N_5023,N_4963,N_4758);
nand U5024 (N_5024,N_4801,N_4981);
xnor U5025 (N_5025,N_4785,N_4824);
xor U5026 (N_5026,N_4774,N_4769);
and U5027 (N_5027,N_4843,N_4765);
xnor U5028 (N_5028,N_4884,N_4900);
and U5029 (N_5029,N_4796,N_4763);
xnor U5030 (N_5030,N_4929,N_4793);
nand U5031 (N_5031,N_4943,N_4879);
xor U5032 (N_5032,N_4913,N_4773);
nand U5033 (N_5033,N_4805,N_4992);
and U5034 (N_5034,N_4902,N_4814);
nor U5035 (N_5035,N_4799,N_4987);
nor U5036 (N_5036,N_4752,N_4941);
and U5037 (N_5037,N_4979,N_4959);
and U5038 (N_5038,N_4891,N_4909);
or U5039 (N_5039,N_4917,N_4820);
and U5040 (N_5040,N_4968,N_4971);
nor U5041 (N_5041,N_4874,N_4984);
and U5042 (N_5042,N_4962,N_4827);
nor U5043 (N_5043,N_4873,N_4764);
nor U5044 (N_5044,N_4871,N_4916);
xor U5045 (N_5045,N_4872,N_4991);
nor U5046 (N_5046,N_4953,N_4863);
xnor U5047 (N_5047,N_4828,N_4942);
and U5048 (N_5048,N_4789,N_4800);
nor U5049 (N_5049,N_4767,N_4996);
nand U5050 (N_5050,N_4795,N_4770);
and U5051 (N_5051,N_4948,N_4817);
xor U5052 (N_5052,N_4794,N_4837);
and U5053 (N_5053,N_4821,N_4926);
or U5054 (N_5054,N_4861,N_4786);
xor U5055 (N_5055,N_4835,N_4881);
xnor U5056 (N_5056,N_4957,N_4808);
and U5057 (N_5057,N_4993,N_4823);
xnor U5058 (N_5058,N_4836,N_4851);
nor U5059 (N_5059,N_4908,N_4867);
xor U5060 (N_5060,N_4815,N_4947);
or U5061 (N_5061,N_4811,N_4983);
xor U5062 (N_5062,N_4956,N_4890);
xor U5063 (N_5063,N_4829,N_4857);
or U5064 (N_5064,N_4980,N_4901);
and U5065 (N_5065,N_4858,N_4781);
or U5066 (N_5066,N_4772,N_4798);
nand U5067 (N_5067,N_4860,N_4898);
nand U5068 (N_5068,N_4806,N_4970);
nor U5069 (N_5069,N_4954,N_4792);
or U5070 (N_5070,N_4897,N_4864);
nand U5071 (N_5071,N_4899,N_4930);
nand U5072 (N_5072,N_4759,N_4761);
xor U5073 (N_5073,N_4807,N_4946);
nor U5074 (N_5074,N_4905,N_4855);
and U5075 (N_5075,N_4776,N_4880);
nor U5076 (N_5076,N_4911,N_4869);
xor U5077 (N_5077,N_4819,N_4885);
and U5078 (N_5078,N_4977,N_4768);
xor U5079 (N_5079,N_4966,N_4751);
nand U5080 (N_5080,N_4849,N_4766);
nand U5081 (N_5081,N_4883,N_4850);
nand U5082 (N_5082,N_4894,N_4967);
xor U5083 (N_5083,N_4876,N_4936);
and U5084 (N_5084,N_4877,N_4928);
and U5085 (N_5085,N_4868,N_4893);
and U5086 (N_5086,N_4784,N_4907);
and U5087 (N_5087,N_4896,N_4988);
or U5088 (N_5088,N_4755,N_4842);
or U5089 (N_5089,N_4779,N_4813);
and U5090 (N_5090,N_4754,N_4847);
and U5091 (N_5091,N_4924,N_4939);
xnor U5092 (N_5092,N_4976,N_4949);
nand U5093 (N_5093,N_4853,N_4889);
xor U5094 (N_5094,N_4790,N_4810);
xor U5095 (N_5095,N_4830,N_4919);
and U5096 (N_5096,N_4990,N_4969);
nor U5097 (N_5097,N_4927,N_4826);
nor U5098 (N_5098,N_4771,N_4886);
and U5099 (N_5099,N_4914,N_4944);
nand U5100 (N_5100,N_4903,N_4937);
nand U5101 (N_5101,N_4831,N_4812);
or U5102 (N_5102,N_4921,N_4845);
xor U5103 (N_5103,N_4802,N_4887);
nor U5104 (N_5104,N_4938,N_4920);
nor U5105 (N_5105,N_4841,N_4933);
nand U5106 (N_5106,N_4780,N_4934);
or U5107 (N_5107,N_4852,N_4848);
and U5108 (N_5108,N_4945,N_4961);
nor U5109 (N_5109,N_4753,N_4846);
nand U5110 (N_5110,N_4932,N_4859);
xnor U5111 (N_5111,N_4998,N_4866);
and U5112 (N_5112,N_4778,N_4955);
nor U5113 (N_5113,N_4918,N_4982);
or U5114 (N_5114,N_4760,N_4791);
nor U5115 (N_5115,N_4910,N_4818);
xnor U5116 (N_5116,N_4787,N_4782);
nor U5117 (N_5117,N_4965,N_4973);
xor U5118 (N_5118,N_4839,N_4986);
or U5119 (N_5119,N_4870,N_4952);
and U5120 (N_5120,N_4757,N_4997);
nand U5121 (N_5121,N_4783,N_4964);
nor U5122 (N_5122,N_4912,N_4995);
xor U5123 (N_5123,N_4803,N_4989);
xor U5124 (N_5124,N_4923,N_4958);
or U5125 (N_5125,N_4883,N_4970);
xnor U5126 (N_5126,N_4836,N_4772);
xnor U5127 (N_5127,N_4991,N_4795);
xnor U5128 (N_5128,N_4886,N_4913);
and U5129 (N_5129,N_4883,N_4900);
xnor U5130 (N_5130,N_4769,N_4938);
and U5131 (N_5131,N_4794,N_4788);
nor U5132 (N_5132,N_4916,N_4819);
and U5133 (N_5133,N_4937,N_4775);
and U5134 (N_5134,N_4802,N_4946);
nor U5135 (N_5135,N_4798,N_4918);
nand U5136 (N_5136,N_4779,N_4903);
and U5137 (N_5137,N_4988,N_4856);
nor U5138 (N_5138,N_4761,N_4794);
and U5139 (N_5139,N_4960,N_4918);
xnor U5140 (N_5140,N_4789,N_4830);
or U5141 (N_5141,N_4836,N_4792);
nor U5142 (N_5142,N_4823,N_4809);
xor U5143 (N_5143,N_4895,N_4860);
and U5144 (N_5144,N_4900,N_4988);
and U5145 (N_5145,N_4972,N_4920);
and U5146 (N_5146,N_4905,N_4859);
or U5147 (N_5147,N_4806,N_4919);
nand U5148 (N_5148,N_4789,N_4761);
nor U5149 (N_5149,N_4832,N_4755);
or U5150 (N_5150,N_4789,N_4920);
xor U5151 (N_5151,N_4800,N_4935);
xor U5152 (N_5152,N_4763,N_4791);
nor U5153 (N_5153,N_4762,N_4927);
and U5154 (N_5154,N_4999,N_4799);
nand U5155 (N_5155,N_4864,N_4837);
or U5156 (N_5156,N_4946,N_4910);
nor U5157 (N_5157,N_4881,N_4836);
xor U5158 (N_5158,N_4907,N_4800);
xnor U5159 (N_5159,N_4869,N_4887);
nor U5160 (N_5160,N_4916,N_4828);
xor U5161 (N_5161,N_4873,N_4945);
or U5162 (N_5162,N_4855,N_4932);
nand U5163 (N_5163,N_4854,N_4996);
nand U5164 (N_5164,N_4766,N_4967);
nand U5165 (N_5165,N_4872,N_4943);
nor U5166 (N_5166,N_4889,N_4905);
or U5167 (N_5167,N_4973,N_4989);
and U5168 (N_5168,N_4802,N_4940);
nor U5169 (N_5169,N_4787,N_4963);
or U5170 (N_5170,N_4885,N_4947);
nand U5171 (N_5171,N_4779,N_4956);
nand U5172 (N_5172,N_4935,N_4985);
nand U5173 (N_5173,N_4781,N_4793);
or U5174 (N_5174,N_4834,N_4817);
nand U5175 (N_5175,N_4782,N_4847);
and U5176 (N_5176,N_4819,N_4919);
nor U5177 (N_5177,N_4844,N_4986);
xnor U5178 (N_5178,N_4878,N_4978);
or U5179 (N_5179,N_4876,N_4835);
and U5180 (N_5180,N_4960,N_4928);
and U5181 (N_5181,N_4812,N_4913);
xor U5182 (N_5182,N_4801,N_4836);
or U5183 (N_5183,N_4976,N_4915);
nor U5184 (N_5184,N_4874,N_4923);
or U5185 (N_5185,N_4771,N_4898);
xnor U5186 (N_5186,N_4830,N_4925);
or U5187 (N_5187,N_4838,N_4992);
xnor U5188 (N_5188,N_4884,N_4921);
nand U5189 (N_5189,N_4921,N_4919);
or U5190 (N_5190,N_4824,N_4916);
xor U5191 (N_5191,N_4751,N_4774);
nor U5192 (N_5192,N_4808,N_4769);
or U5193 (N_5193,N_4977,N_4848);
or U5194 (N_5194,N_4910,N_4900);
or U5195 (N_5195,N_4916,N_4854);
xnor U5196 (N_5196,N_4853,N_4798);
and U5197 (N_5197,N_4883,N_4888);
xnor U5198 (N_5198,N_4848,N_4887);
and U5199 (N_5199,N_4864,N_4871);
xor U5200 (N_5200,N_4809,N_4907);
and U5201 (N_5201,N_4871,N_4949);
or U5202 (N_5202,N_4924,N_4875);
nor U5203 (N_5203,N_4885,N_4955);
nor U5204 (N_5204,N_4793,N_4770);
or U5205 (N_5205,N_4929,N_4762);
nand U5206 (N_5206,N_4964,N_4874);
and U5207 (N_5207,N_4924,N_4971);
nand U5208 (N_5208,N_4768,N_4812);
or U5209 (N_5209,N_4826,N_4925);
nor U5210 (N_5210,N_4927,N_4841);
nor U5211 (N_5211,N_4857,N_4837);
nor U5212 (N_5212,N_4791,N_4944);
and U5213 (N_5213,N_4988,N_4847);
or U5214 (N_5214,N_4874,N_4868);
xnor U5215 (N_5215,N_4777,N_4873);
nand U5216 (N_5216,N_4996,N_4883);
nand U5217 (N_5217,N_4896,N_4840);
nor U5218 (N_5218,N_4814,N_4789);
and U5219 (N_5219,N_4932,N_4881);
and U5220 (N_5220,N_4906,N_4916);
or U5221 (N_5221,N_4933,N_4984);
or U5222 (N_5222,N_4902,N_4767);
nor U5223 (N_5223,N_4966,N_4888);
nand U5224 (N_5224,N_4783,N_4958);
nand U5225 (N_5225,N_4943,N_4959);
nor U5226 (N_5226,N_4928,N_4958);
or U5227 (N_5227,N_4771,N_4952);
nand U5228 (N_5228,N_4879,N_4977);
nand U5229 (N_5229,N_4907,N_4829);
nand U5230 (N_5230,N_4786,N_4813);
xor U5231 (N_5231,N_4932,N_4994);
xor U5232 (N_5232,N_4826,N_4998);
xnor U5233 (N_5233,N_4751,N_4907);
xor U5234 (N_5234,N_4911,N_4901);
and U5235 (N_5235,N_4896,N_4775);
nor U5236 (N_5236,N_4964,N_4810);
and U5237 (N_5237,N_4871,N_4989);
nand U5238 (N_5238,N_4819,N_4880);
and U5239 (N_5239,N_4902,N_4857);
or U5240 (N_5240,N_4942,N_4763);
and U5241 (N_5241,N_4988,N_4903);
and U5242 (N_5242,N_4905,N_4880);
nor U5243 (N_5243,N_4788,N_4961);
nand U5244 (N_5244,N_4912,N_4945);
nor U5245 (N_5245,N_4936,N_4984);
nand U5246 (N_5246,N_4965,N_4846);
or U5247 (N_5247,N_4752,N_4874);
xor U5248 (N_5248,N_4942,N_4769);
or U5249 (N_5249,N_4779,N_4794);
or U5250 (N_5250,N_5057,N_5090);
nor U5251 (N_5251,N_5188,N_5089);
nor U5252 (N_5252,N_5049,N_5038);
nor U5253 (N_5253,N_5032,N_5018);
nand U5254 (N_5254,N_5026,N_5211);
and U5255 (N_5255,N_5061,N_5109);
and U5256 (N_5256,N_5149,N_5193);
and U5257 (N_5257,N_5016,N_5025);
or U5258 (N_5258,N_5230,N_5160);
or U5259 (N_5259,N_5219,N_5107);
or U5260 (N_5260,N_5248,N_5105);
xor U5261 (N_5261,N_5166,N_5088);
nor U5262 (N_5262,N_5221,N_5139);
nor U5263 (N_5263,N_5246,N_5208);
and U5264 (N_5264,N_5073,N_5147);
xor U5265 (N_5265,N_5231,N_5067);
nand U5266 (N_5266,N_5124,N_5185);
or U5267 (N_5267,N_5174,N_5177);
xor U5268 (N_5268,N_5218,N_5175);
xnor U5269 (N_5269,N_5053,N_5116);
nand U5270 (N_5270,N_5156,N_5011);
or U5271 (N_5271,N_5065,N_5228);
or U5272 (N_5272,N_5170,N_5141);
nand U5273 (N_5273,N_5191,N_5027);
and U5274 (N_5274,N_5087,N_5134);
or U5275 (N_5275,N_5126,N_5114);
or U5276 (N_5276,N_5244,N_5043);
nand U5277 (N_5277,N_5036,N_5223);
or U5278 (N_5278,N_5009,N_5146);
and U5279 (N_5279,N_5215,N_5052);
nor U5280 (N_5280,N_5080,N_5209);
nor U5281 (N_5281,N_5238,N_5072);
nor U5282 (N_5282,N_5030,N_5194);
or U5283 (N_5283,N_5119,N_5214);
or U5284 (N_5284,N_5163,N_5003);
nand U5285 (N_5285,N_5097,N_5045);
xnor U5286 (N_5286,N_5169,N_5133);
nand U5287 (N_5287,N_5148,N_5186);
and U5288 (N_5288,N_5033,N_5111);
nor U5289 (N_5289,N_5171,N_5237);
xnor U5290 (N_5290,N_5064,N_5028);
nand U5291 (N_5291,N_5137,N_5104);
nor U5292 (N_5292,N_5178,N_5142);
xnor U5293 (N_5293,N_5005,N_5180);
nor U5294 (N_5294,N_5155,N_5000);
nand U5295 (N_5295,N_5118,N_5183);
nor U5296 (N_5296,N_5200,N_5063);
nand U5297 (N_5297,N_5181,N_5096);
or U5298 (N_5298,N_5019,N_5034);
nand U5299 (N_5299,N_5070,N_5069);
nand U5300 (N_5300,N_5132,N_5010);
nand U5301 (N_5301,N_5001,N_5172);
xor U5302 (N_5302,N_5078,N_5095);
xor U5303 (N_5303,N_5161,N_5044);
xnor U5304 (N_5304,N_5024,N_5056);
or U5305 (N_5305,N_5179,N_5176);
nand U5306 (N_5306,N_5054,N_5127);
nor U5307 (N_5307,N_5076,N_5094);
and U5308 (N_5308,N_5217,N_5093);
and U5309 (N_5309,N_5182,N_5173);
nand U5310 (N_5310,N_5203,N_5234);
nand U5311 (N_5311,N_5222,N_5058);
nand U5312 (N_5312,N_5106,N_5113);
xor U5313 (N_5313,N_5190,N_5167);
nand U5314 (N_5314,N_5212,N_5079);
or U5315 (N_5315,N_5202,N_5140);
nand U5316 (N_5316,N_5224,N_5002);
or U5317 (N_5317,N_5210,N_5235);
nand U5318 (N_5318,N_5066,N_5225);
and U5319 (N_5319,N_5247,N_5195);
xnor U5320 (N_5320,N_5243,N_5216);
xor U5321 (N_5321,N_5196,N_5007);
or U5322 (N_5322,N_5062,N_5120);
nor U5323 (N_5323,N_5060,N_5039);
xnor U5324 (N_5324,N_5084,N_5187);
nor U5325 (N_5325,N_5101,N_5226);
or U5326 (N_5326,N_5136,N_5165);
nand U5327 (N_5327,N_5158,N_5037);
nand U5328 (N_5328,N_5013,N_5086);
and U5329 (N_5329,N_5242,N_5008);
nor U5330 (N_5330,N_5143,N_5152);
xor U5331 (N_5331,N_5021,N_5125);
or U5332 (N_5332,N_5122,N_5131);
nor U5333 (N_5333,N_5206,N_5110);
nand U5334 (N_5334,N_5233,N_5239);
or U5335 (N_5335,N_5098,N_5081);
and U5336 (N_5336,N_5192,N_5042);
nor U5337 (N_5337,N_5020,N_5154);
nor U5338 (N_5338,N_5041,N_5159);
xnor U5339 (N_5339,N_5074,N_5151);
nor U5340 (N_5340,N_5245,N_5071);
or U5341 (N_5341,N_5232,N_5198);
nand U5342 (N_5342,N_5117,N_5112);
or U5343 (N_5343,N_5157,N_5103);
nor U5344 (N_5344,N_5130,N_5059);
xnor U5345 (N_5345,N_5123,N_5091);
and U5346 (N_5346,N_5207,N_5035);
nand U5347 (N_5347,N_5085,N_5164);
nor U5348 (N_5348,N_5145,N_5236);
or U5349 (N_5349,N_5162,N_5050);
and U5350 (N_5350,N_5022,N_5197);
and U5351 (N_5351,N_5129,N_5153);
or U5352 (N_5352,N_5048,N_5184);
nor U5353 (N_5353,N_5040,N_5014);
nor U5354 (N_5354,N_5240,N_5083);
and U5355 (N_5355,N_5031,N_5051);
xnor U5356 (N_5356,N_5047,N_5227);
nand U5357 (N_5357,N_5138,N_5108);
or U5358 (N_5358,N_5099,N_5150);
or U5359 (N_5359,N_5029,N_5144);
and U5360 (N_5360,N_5046,N_5012);
or U5361 (N_5361,N_5055,N_5121);
nand U5362 (N_5362,N_5199,N_5023);
nor U5363 (N_5363,N_5077,N_5082);
nand U5364 (N_5364,N_5102,N_5092);
xor U5365 (N_5365,N_5100,N_5168);
xnor U5366 (N_5366,N_5229,N_5128);
nand U5367 (N_5367,N_5189,N_5220);
xor U5368 (N_5368,N_5017,N_5068);
and U5369 (N_5369,N_5204,N_5006);
xnor U5370 (N_5370,N_5004,N_5213);
nor U5371 (N_5371,N_5205,N_5115);
and U5372 (N_5372,N_5201,N_5015);
nand U5373 (N_5373,N_5135,N_5249);
xnor U5374 (N_5374,N_5241,N_5075);
and U5375 (N_5375,N_5194,N_5034);
nor U5376 (N_5376,N_5018,N_5085);
or U5377 (N_5377,N_5128,N_5045);
or U5378 (N_5378,N_5043,N_5096);
or U5379 (N_5379,N_5073,N_5165);
xor U5380 (N_5380,N_5180,N_5112);
or U5381 (N_5381,N_5143,N_5077);
nor U5382 (N_5382,N_5000,N_5083);
or U5383 (N_5383,N_5133,N_5203);
xnor U5384 (N_5384,N_5148,N_5198);
xnor U5385 (N_5385,N_5061,N_5185);
xnor U5386 (N_5386,N_5020,N_5229);
nor U5387 (N_5387,N_5028,N_5219);
or U5388 (N_5388,N_5242,N_5134);
nand U5389 (N_5389,N_5121,N_5191);
xnor U5390 (N_5390,N_5090,N_5216);
and U5391 (N_5391,N_5096,N_5056);
nand U5392 (N_5392,N_5024,N_5167);
nor U5393 (N_5393,N_5155,N_5197);
xor U5394 (N_5394,N_5120,N_5007);
or U5395 (N_5395,N_5009,N_5183);
nor U5396 (N_5396,N_5010,N_5046);
nand U5397 (N_5397,N_5200,N_5028);
xnor U5398 (N_5398,N_5095,N_5010);
or U5399 (N_5399,N_5063,N_5138);
nand U5400 (N_5400,N_5150,N_5082);
or U5401 (N_5401,N_5103,N_5244);
and U5402 (N_5402,N_5192,N_5025);
and U5403 (N_5403,N_5162,N_5161);
xor U5404 (N_5404,N_5015,N_5136);
nand U5405 (N_5405,N_5076,N_5042);
or U5406 (N_5406,N_5203,N_5069);
xor U5407 (N_5407,N_5230,N_5029);
or U5408 (N_5408,N_5137,N_5180);
nor U5409 (N_5409,N_5194,N_5161);
and U5410 (N_5410,N_5061,N_5022);
and U5411 (N_5411,N_5111,N_5082);
xnor U5412 (N_5412,N_5242,N_5175);
xnor U5413 (N_5413,N_5243,N_5068);
or U5414 (N_5414,N_5243,N_5164);
nand U5415 (N_5415,N_5084,N_5193);
nor U5416 (N_5416,N_5079,N_5084);
xor U5417 (N_5417,N_5022,N_5018);
and U5418 (N_5418,N_5186,N_5107);
nor U5419 (N_5419,N_5113,N_5155);
nor U5420 (N_5420,N_5148,N_5220);
xnor U5421 (N_5421,N_5082,N_5130);
and U5422 (N_5422,N_5241,N_5035);
nand U5423 (N_5423,N_5156,N_5061);
and U5424 (N_5424,N_5134,N_5162);
nand U5425 (N_5425,N_5031,N_5058);
nand U5426 (N_5426,N_5120,N_5071);
or U5427 (N_5427,N_5006,N_5198);
or U5428 (N_5428,N_5214,N_5240);
nor U5429 (N_5429,N_5138,N_5002);
xor U5430 (N_5430,N_5117,N_5103);
and U5431 (N_5431,N_5074,N_5165);
or U5432 (N_5432,N_5134,N_5060);
or U5433 (N_5433,N_5193,N_5232);
nand U5434 (N_5434,N_5236,N_5146);
or U5435 (N_5435,N_5067,N_5239);
nor U5436 (N_5436,N_5029,N_5238);
nor U5437 (N_5437,N_5208,N_5019);
nor U5438 (N_5438,N_5236,N_5148);
nand U5439 (N_5439,N_5007,N_5244);
nor U5440 (N_5440,N_5109,N_5165);
nor U5441 (N_5441,N_5228,N_5106);
and U5442 (N_5442,N_5233,N_5140);
or U5443 (N_5443,N_5176,N_5177);
nand U5444 (N_5444,N_5230,N_5228);
nor U5445 (N_5445,N_5113,N_5121);
and U5446 (N_5446,N_5143,N_5158);
nand U5447 (N_5447,N_5194,N_5000);
and U5448 (N_5448,N_5052,N_5072);
nor U5449 (N_5449,N_5014,N_5088);
or U5450 (N_5450,N_5183,N_5186);
nor U5451 (N_5451,N_5197,N_5085);
nand U5452 (N_5452,N_5053,N_5008);
or U5453 (N_5453,N_5043,N_5155);
nor U5454 (N_5454,N_5067,N_5089);
xor U5455 (N_5455,N_5179,N_5026);
or U5456 (N_5456,N_5102,N_5035);
xor U5457 (N_5457,N_5162,N_5120);
and U5458 (N_5458,N_5123,N_5136);
and U5459 (N_5459,N_5218,N_5074);
and U5460 (N_5460,N_5022,N_5205);
xor U5461 (N_5461,N_5030,N_5073);
and U5462 (N_5462,N_5053,N_5017);
nor U5463 (N_5463,N_5110,N_5061);
or U5464 (N_5464,N_5071,N_5198);
xor U5465 (N_5465,N_5164,N_5161);
nand U5466 (N_5466,N_5206,N_5017);
and U5467 (N_5467,N_5233,N_5021);
nand U5468 (N_5468,N_5180,N_5033);
nand U5469 (N_5469,N_5005,N_5216);
or U5470 (N_5470,N_5130,N_5004);
or U5471 (N_5471,N_5249,N_5156);
and U5472 (N_5472,N_5138,N_5223);
nand U5473 (N_5473,N_5201,N_5047);
and U5474 (N_5474,N_5148,N_5201);
or U5475 (N_5475,N_5075,N_5077);
and U5476 (N_5476,N_5031,N_5186);
nor U5477 (N_5477,N_5092,N_5236);
or U5478 (N_5478,N_5209,N_5065);
and U5479 (N_5479,N_5093,N_5242);
nand U5480 (N_5480,N_5085,N_5107);
nor U5481 (N_5481,N_5112,N_5193);
or U5482 (N_5482,N_5052,N_5240);
nand U5483 (N_5483,N_5121,N_5139);
nand U5484 (N_5484,N_5143,N_5188);
or U5485 (N_5485,N_5115,N_5055);
and U5486 (N_5486,N_5130,N_5107);
nor U5487 (N_5487,N_5062,N_5078);
nor U5488 (N_5488,N_5198,N_5107);
and U5489 (N_5489,N_5110,N_5101);
or U5490 (N_5490,N_5127,N_5118);
nor U5491 (N_5491,N_5072,N_5128);
nand U5492 (N_5492,N_5052,N_5090);
xnor U5493 (N_5493,N_5156,N_5007);
xor U5494 (N_5494,N_5249,N_5225);
and U5495 (N_5495,N_5185,N_5177);
nand U5496 (N_5496,N_5123,N_5237);
xor U5497 (N_5497,N_5043,N_5106);
nand U5498 (N_5498,N_5097,N_5039);
xor U5499 (N_5499,N_5222,N_5174);
or U5500 (N_5500,N_5411,N_5474);
and U5501 (N_5501,N_5473,N_5383);
xnor U5502 (N_5502,N_5263,N_5394);
nand U5503 (N_5503,N_5346,N_5447);
nand U5504 (N_5504,N_5461,N_5348);
xor U5505 (N_5505,N_5381,N_5262);
xor U5506 (N_5506,N_5495,N_5398);
xnor U5507 (N_5507,N_5282,N_5478);
nand U5508 (N_5508,N_5494,N_5309);
or U5509 (N_5509,N_5360,N_5337);
nor U5510 (N_5510,N_5444,N_5479);
nand U5511 (N_5511,N_5254,N_5385);
nand U5512 (N_5512,N_5256,N_5280);
nor U5513 (N_5513,N_5423,N_5438);
or U5514 (N_5514,N_5432,N_5487);
or U5515 (N_5515,N_5421,N_5267);
or U5516 (N_5516,N_5357,N_5268);
or U5517 (N_5517,N_5345,N_5260);
nor U5518 (N_5518,N_5493,N_5375);
or U5519 (N_5519,N_5320,N_5445);
nand U5520 (N_5520,N_5455,N_5472);
xor U5521 (N_5521,N_5287,N_5450);
nor U5522 (N_5522,N_5404,N_5316);
xor U5523 (N_5523,N_5436,N_5471);
or U5524 (N_5524,N_5349,N_5396);
and U5525 (N_5525,N_5433,N_5388);
xnor U5526 (N_5526,N_5257,N_5342);
and U5527 (N_5527,N_5499,N_5393);
or U5528 (N_5528,N_5326,N_5285);
and U5529 (N_5529,N_5259,N_5321);
nand U5530 (N_5530,N_5480,N_5496);
nand U5531 (N_5531,N_5469,N_5356);
nor U5532 (N_5532,N_5255,N_5422);
nor U5533 (N_5533,N_5322,N_5278);
nand U5534 (N_5534,N_5453,N_5363);
or U5535 (N_5535,N_5369,N_5352);
xor U5536 (N_5536,N_5270,N_5318);
nand U5537 (N_5537,N_5339,N_5258);
or U5538 (N_5538,N_5387,N_5372);
xor U5539 (N_5539,N_5274,N_5483);
xor U5540 (N_5540,N_5367,N_5384);
nand U5541 (N_5541,N_5334,N_5413);
and U5542 (N_5542,N_5373,N_5488);
and U5543 (N_5543,N_5490,N_5347);
xor U5544 (N_5544,N_5264,N_5415);
nor U5545 (N_5545,N_5374,N_5449);
or U5546 (N_5546,N_5359,N_5283);
nor U5547 (N_5547,N_5364,N_5498);
or U5548 (N_5548,N_5279,N_5333);
nand U5549 (N_5549,N_5301,N_5390);
nand U5550 (N_5550,N_5402,N_5335);
xnor U5551 (N_5551,N_5441,N_5417);
nor U5552 (N_5552,N_5424,N_5382);
or U5553 (N_5553,N_5416,N_5251);
or U5554 (N_5554,N_5481,N_5437);
and U5555 (N_5555,N_5492,N_5429);
xnor U5556 (N_5556,N_5440,N_5446);
nor U5557 (N_5557,N_5397,N_5408);
and U5558 (N_5558,N_5261,N_5443);
and U5559 (N_5559,N_5368,N_5484);
and U5560 (N_5560,N_5409,N_5361);
nand U5561 (N_5561,N_5330,N_5354);
xor U5562 (N_5562,N_5289,N_5298);
nor U5563 (N_5563,N_5435,N_5265);
nor U5564 (N_5564,N_5290,N_5294);
and U5565 (N_5565,N_5439,N_5366);
xnor U5566 (N_5566,N_5324,N_5344);
or U5567 (N_5567,N_5338,N_5252);
nand U5568 (N_5568,N_5253,N_5414);
or U5569 (N_5569,N_5448,N_5266);
or U5570 (N_5570,N_5271,N_5269);
and U5571 (N_5571,N_5300,N_5389);
xnor U5572 (N_5572,N_5485,N_5491);
xnor U5573 (N_5573,N_5362,N_5284);
or U5574 (N_5574,N_5426,N_5281);
nor U5575 (N_5575,N_5459,N_5482);
or U5576 (N_5576,N_5380,N_5497);
xnor U5577 (N_5577,N_5467,N_5317);
xor U5578 (N_5578,N_5371,N_5468);
nand U5579 (N_5579,N_5276,N_5305);
or U5580 (N_5580,N_5315,N_5291);
nor U5581 (N_5581,N_5272,N_5400);
or U5582 (N_5582,N_5355,N_5292);
or U5583 (N_5583,N_5406,N_5391);
nor U5584 (N_5584,N_5304,N_5419);
nand U5585 (N_5585,N_5340,N_5307);
nor U5586 (N_5586,N_5379,N_5431);
nor U5587 (N_5587,N_5475,N_5392);
xor U5588 (N_5588,N_5308,N_5299);
or U5589 (N_5589,N_5457,N_5412);
xor U5590 (N_5590,N_5465,N_5302);
or U5591 (N_5591,N_5418,N_5477);
or U5592 (N_5592,N_5350,N_5430);
and U5593 (N_5593,N_5313,N_5323);
and U5594 (N_5594,N_5319,N_5341);
nand U5595 (N_5595,N_5306,N_5442);
xnor U5596 (N_5596,N_5462,N_5310);
xnor U5597 (N_5597,N_5296,N_5297);
and U5598 (N_5598,N_5486,N_5460);
xor U5599 (N_5599,N_5456,N_5286);
xnor U5600 (N_5600,N_5476,N_5420);
xnor U5601 (N_5601,N_5288,N_5331);
xnor U5602 (N_5602,N_5376,N_5358);
nand U5603 (N_5603,N_5378,N_5403);
or U5604 (N_5604,N_5410,N_5343);
or U5605 (N_5605,N_5277,N_5451);
nor U5606 (N_5606,N_5428,N_5395);
xnor U5607 (N_5607,N_5399,N_5303);
or U5608 (N_5608,N_5489,N_5332);
nand U5609 (N_5609,N_5454,N_5405);
and U5610 (N_5610,N_5250,N_5463);
nor U5611 (N_5611,N_5325,N_5273);
or U5612 (N_5612,N_5458,N_5407);
and U5613 (N_5613,N_5311,N_5386);
nand U5614 (N_5614,N_5370,N_5329);
xor U5615 (N_5615,N_5336,N_5275);
or U5616 (N_5616,N_5351,N_5434);
nor U5617 (N_5617,N_5293,N_5470);
nand U5618 (N_5618,N_5401,N_5452);
nor U5619 (N_5619,N_5314,N_5365);
or U5620 (N_5620,N_5295,N_5466);
or U5621 (N_5621,N_5427,N_5464);
xor U5622 (N_5622,N_5377,N_5328);
and U5623 (N_5623,N_5327,N_5353);
nor U5624 (N_5624,N_5425,N_5312);
and U5625 (N_5625,N_5397,N_5250);
xnor U5626 (N_5626,N_5329,N_5419);
and U5627 (N_5627,N_5479,N_5450);
and U5628 (N_5628,N_5353,N_5492);
nand U5629 (N_5629,N_5392,N_5458);
or U5630 (N_5630,N_5278,N_5492);
or U5631 (N_5631,N_5375,N_5393);
xnor U5632 (N_5632,N_5415,N_5261);
nand U5633 (N_5633,N_5277,N_5397);
nor U5634 (N_5634,N_5438,N_5420);
nor U5635 (N_5635,N_5477,N_5258);
or U5636 (N_5636,N_5442,N_5445);
or U5637 (N_5637,N_5398,N_5273);
and U5638 (N_5638,N_5343,N_5276);
xnor U5639 (N_5639,N_5408,N_5251);
xor U5640 (N_5640,N_5499,N_5407);
nand U5641 (N_5641,N_5283,N_5255);
nand U5642 (N_5642,N_5370,N_5398);
nand U5643 (N_5643,N_5339,N_5338);
nand U5644 (N_5644,N_5418,N_5383);
or U5645 (N_5645,N_5291,N_5354);
nor U5646 (N_5646,N_5392,N_5303);
nand U5647 (N_5647,N_5430,N_5464);
and U5648 (N_5648,N_5266,N_5391);
nor U5649 (N_5649,N_5396,N_5390);
nor U5650 (N_5650,N_5436,N_5489);
nor U5651 (N_5651,N_5297,N_5486);
xor U5652 (N_5652,N_5461,N_5478);
nand U5653 (N_5653,N_5476,N_5338);
nor U5654 (N_5654,N_5493,N_5400);
nand U5655 (N_5655,N_5404,N_5276);
nor U5656 (N_5656,N_5360,N_5401);
and U5657 (N_5657,N_5481,N_5434);
and U5658 (N_5658,N_5448,N_5280);
xnor U5659 (N_5659,N_5349,N_5433);
nor U5660 (N_5660,N_5392,N_5372);
nand U5661 (N_5661,N_5459,N_5308);
nor U5662 (N_5662,N_5255,N_5373);
nor U5663 (N_5663,N_5265,N_5450);
nand U5664 (N_5664,N_5396,N_5426);
xor U5665 (N_5665,N_5272,N_5326);
or U5666 (N_5666,N_5390,N_5473);
nor U5667 (N_5667,N_5363,N_5498);
or U5668 (N_5668,N_5401,N_5364);
or U5669 (N_5669,N_5446,N_5324);
or U5670 (N_5670,N_5379,N_5395);
and U5671 (N_5671,N_5438,N_5271);
nor U5672 (N_5672,N_5306,N_5385);
nor U5673 (N_5673,N_5277,N_5316);
and U5674 (N_5674,N_5491,N_5493);
or U5675 (N_5675,N_5405,N_5275);
and U5676 (N_5676,N_5283,N_5388);
nor U5677 (N_5677,N_5425,N_5250);
nor U5678 (N_5678,N_5303,N_5430);
nor U5679 (N_5679,N_5406,N_5389);
or U5680 (N_5680,N_5299,N_5403);
nand U5681 (N_5681,N_5273,N_5280);
and U5682 (N_5682,N_5427,N_5278);
xnor U5683 (N_5683,N_5498,N_5340);
nand U5684 (N_5684,N_5468,N_5442);
nor U5685 (N_5685,N_5423,N_5313);
or U5686 (N_5686,N_5324,N_5478);
and U5687 (N_5687,N_5300,N_5388);
nor U5688 (N_5688,N_5349,N_5395);
xor U5689 (N_5689,N_5427,N_5317);
and U5690 (N_5690,N_5396,N_5470);
xor U5691 (N_5691,N_5343,N_5365);
nor U5692 (N_5692,N_5384,N_5411);
nor U5693 (N_5693,N_5278,N_5339);
and U5694 (N_5694,N_5283,N_5257);
xor U5695 (N_5695,N_5333,N_5467);
and U5696 (N_5696,N_5448,N_5316);
nor U5697 (N_5697,N_5299,N_5485);
xnor U5698 (N_5698,N_5272,N_5474);
nor U5699 (N_5699,N_5444,N_5419);
and U5700 (N_5700,N_5429,N_5476);
xor U5701 (N_5701,N_5352,N_5365);
or U5702 (N_5702,N_5250,N_5287);
nand U5703 (N_5703,N_5422,N_5404);
xnor U5704 (N_5704,N_5400,N_5365);
and U5705 (N_5705,N_5292,N_5261);
xnor U5706 (N_5706,N_5371,N_5267);
and U5707 (N_5707,N_5437,N_5337);
or U5708 (N_5708,N_5417,N_5413);
nor U5709 (N_5709,N_5417,N_5361);
xor U5710 (N_5710,N_5355,N_5468);
xnor U5711 (N_5711,N_5435,N_5376);
and U5712 (N_5712,N_5354,N_5260);
xor U5713 (N_5713,N_5340,N_5274);
nand U5714 (N_5714,N_5292,N_5266);
xnor U5715 (N_5715,N_5385,N_5383);
and U5716 (N_5716,N_5351,N_5419);
nand U5717 (N_5717,N_5300,N_5434);
or U5718 (N_5718,N_5401,N_5374);
nand U5719 (N_5719,N_5288,N_5383);
and U5720 (N_5720,N_5367,N_5470);
xnor U5721 (N_5721,N_5489,N_5449);
and U5722 (N_5722,N_5388,N_5432);
or U5723 (N_5723,N_5420,N_5465);
xnor U5724 (N_5724,N_5357,N_5295);
nor U5725 (N_5725,N_5313,N_5391);
and U5726 (N_5726,N_5381,N_5428);
nand U5727 (N_5727,N_5275,N_5417);
nor U5728 (N_5728,N_5290,N_5466);
and U5729 (N_5729,N_5341,N_5318);
and U5730 (N_5730,N_5303,N_5377);
or U5731 (N_5731,N_5368,N_5347);
and U5732 (N_5732,N_5477,N_5316);
or U5733 (N_5733,N_5344,N_5385);
and U5734 (N_5734,N_5252,N_5325);
or U5735 (N_5735,N_5440,N_5360);
xor U5736 (N_5736,N_5323,N_5451);
or U5737 (N_5737,N_5315,N_5351);
xor U5738 (N_5738,N_5275,N_5303);
nor U5739 (N_5739,N_5441,N_5431);
nand U5740 (N_5740,N_5261,N_5350);
xnor U5741 (N_5741,N_5382,N_5358);
and U5742 (N_5742,N_5472,N_5440);
and U5743 (N_5743,N_5345,N_5375);
and U5744 (N_5744,N_5451,N_5264);
nand U5745 (N_5745,N_5325,N_5401);
nand U5746 (N_5746,N_5442,N_5362);
and U5747 (N_5747,N_5324,N_5494);
and U5748 (N_5748,N_5418,N_5298);
and U5749 (N_5749,N_5284,N_5499);
xnor U5750 (N_5750,N_5559,N_5627);
or U5751 (N_5751,N_5740,N_5643);
and U5752 (N_5752,N_5557,N_5563);
nor U5753 (N_5753,N_5601,N_5529);
nand U5754 (N_5754,N_5710,N_5692);
nand U5755 (N_5755,N_5655,N_5565);
nand U5756 (N_5756,N_5743,N_5715);
and U5757 (N_5757,N_5512,N_5592);
nand U5758 (N_5758,N_5551,N_5544);
xnor U5759 (N_5759,N_5656,N_5598);
nor U5760 (N_5760,N_5675,N_5633);
xor U5761 (N_5761,N_5658,N_5620);
xnor U5762 (N_5762,N_5561,N_5687);
nor U5763 (N_5763,N_5665,N_5600);
nand U5764 (N_5764,N_5546,N_5681);
nand U5765 (N_5765,N_5732,N_5538);
nand U5766 (N_5766,N_5562,N_5713);
nor U5767 (N_5767,N_5648,N_5541);
nand U5768 (N_5768,N_5524,N_5506);
xor U5769 (N_5769,N_5688,N_5696);
and U5770 (N_5770,N_5518,N_5609);
nor U5771 (N_5771,N_5576,N_5566);
nand U5772 (N_5772,N_5618,N_5564);
xnor U5773 (N_5773,N_5735,N_5604);
nand U5774 (N_5774,N_5596,N_5702);
or U5775 (N_5775,N_5605,N_5554);
nor U5776 (N_5776,N_5626,N_5515);
nor U5777 (N_5777,N_5676,N_5575);
nand U5778 (N_5778,N_5622,N_5742);
nand U5779 (N_5779,N_5614,N_5661);
nor U5780 (N_5780,N_5582,N_5693);
nand U5781 (N_5781,N_5612,N_5660);
or U5782 (N_5782,N_5657,N_5642);
nand U5783 (N_5783,N_5654,N_5689);
xnor U5784 (N_5784,N_5581,N_5509);
xor U5785 (N_5785,N_5672,N_5542);
and U5786 (N_5786,N_5593,N_5547);
xor U5787 (N_5787,N_5703,N_5550);
nand U5788 (N_5788,N_5708,N_5639);
nor U5789 (N_5789,N_5586,N_5738);
or U5790 (N_5790,N_5719,N_5680);
or U5791 (N_5791,N_5651,N_5624);
and U5792 (N_5792,N_5523,N_5741);
nor U5793 (N_5793,N_5695,N_5500);
nor U5794 (N_5794,N_5504,N_5570);
or U5795 (N_5795,N_5638,N_5527);
and U5796 (N_5796,N_5503,N_5545);
or U5797 (N_5797,N_5646,N_5553);
nor U5798 (N_5798,N_5685,N_5629);
xnor U5799 (N_5799,N_5705,N_5528);
nand U5800 (N_5800,N_5662,N_5539);
xor U5801 (N_5801,N_5555,N_5577);
nand U5802 (N_5802,N_5595,N_5619);
nand U5803 (N_5803,N_5536,N_5694);
nor U5804 (N_5804,N_5571,N_5611);
and U5805 (N_5805,N_5625,N_5535);
or U5806 (N_5806,N_5507,N_5641);
nor U5807 (N_5807,N_5543,N_5599);
nand U5808 (N_5808,N_5591,N_5634);
or U5809 (N_5809,N_5663,N_5623);
or U5810 (N_5810,N_5522,N_5727);
xor U5811 (N_5811,N_5501,N_5587);
xor U5812 (N_5812,N_5532,N_5712);
and U5813 (N_5813,N_5690,N_5613);
and U5814 (N_5814,N_5608,N_5549);
and U5815 (N_5815,N_5736,N_5517);
nand U5816 (N_5816,N_5691,N_5704);
nor U5817 (N_5817,N_5508,N_5711);
nand U5818 (N_5818,N_5637,N_5640);
nand U5819 (N_5819,N_5537,N_5521);
xor U5820 (N_5820,N_5630,N_5516);
and U5821 (N_5821,N_5671,N_5594);
nand U5822 (N_5822,N_5664,N_5723);
nor U5823 (N_5823,N_5731,N_5686);
or U5824 (N_5824,N_5569,N_5717);
nor U5825 (N_5825,N_5653,N_5734);
xnor U5826 (N_5826,N_5628,N_5669);
xor U5827 (N_5827,N_5525,N_5631);
nor U5828 (N_5828,N_5616,N_5603);
and U5829 (N_5829,N_5739,N_5706);
or U5830 (N_5830,N_5636,N_5632);
xnor U5831 (N_5831,N_5590,N_5567);
and U5832 (N_5832,N_5645,N_5697);
xor U5833 (N_5833,N_5722,N_5585);
nand U5834 (N_5834,N_5584,N_5729);
or U5835 (N_5835,N_5677,N_5747);
nand U5836 (N_5836,N_5666,N_5745);
nor U5837 (N_5837,N_5748,N_5574);
and U5838 (N_5838,N_5698,N_5526);
xnor U5839 (N_5839,N_5511,N_5659);
xor U5840 (N_5840,N_5621,N_5530);
nor U5841 (N_5841,N_5746,N_5568);
xnor U5842 (N_5842,N_5744,N_5737);
xor U5843 (N_5843,N_5707,N_5606);
and U5844 (N_5844,N_5597,N_5579);
xnor U5845 (N_5845,N_5502,N_5725);
nor U5846 (N_5846,N_5701,N_5583);
and U5847 (N_5847,N_5647,N_5700);
nand U5848 (N_5848,N_5513,N_5602);
and U5849 (N_5849,N_5730,N_5720);
xnor U5850 (N_5850,N_5724,N_5714);
and U5851 (N_5851,N_5728,N_5589);
and U5852 (N_5852,N_5556,N_5505);
or U5853 (N_5853,N_5540,N_5519);
or U5854 (N_5854,N_5683,N_5558);
nand U5855 (N_5855,N_5635,N_5552);
and U5856 (N_5856,N_5682,N_5510);
nand U5857 (N_5857,N_5572,N_5580);
nand U5858 (N_5858,N_5749,N_5678);
and U5859 (N_5859,N_5578,N_5560);
xor U5860 (N_5860,N_5520,N_5684);
nand U5861 (N_5861,N_5644,N_5607);
or U5862 (N_5862,N_5610,N_5650);
xnor U5863 (N_5863,N_5534,N_5615);
or U5864 (N_5864,N_5709,N_5668);
or U5865 (N_5865,N_5721,N_5733);
and U5866 (N_5866,N_5726,N_5548);
nor U5867 (N_5867,N_5617,N_5667);
or U5868 (N_5868,N_5679,N_5673);
xor U5869 (N_5869,N_5674,N_5699);
xor U5870 (N_5870,N_5670,N_5533);
and U5871 (N_5871,N_5718,N_5531);
and U5872 (N_5872,N_5573,N_5649);
nor U5873 (N_5873,N_5716,N_5588);
nand U5874 (N_5874,N_5652,N_5514);
xor U5875 (N_5875,N_5503,N_5620);
nor U5876 (N_5876,N_5564,N_5720);
xnor U5877 (N_5877,N_5662,N_5557);
nand U5878 (N_5878,N_5532,N_5554);
nor U5879 (N_5879,N_5599,N_5741);
xor U5880 (N_5880,N_5547,N_5517);
nand U5881 (N_5881,N_5546,N_5623);
xnor U5882 (N_5882,N_5590,N_5538);
or U5883 (N_5883,N_5566,N_5527);
or U5884 (N_5884,N_5733,N_5591);
nor U5885 (N_5885,N_5605,N_5740);
nor U5886 (N_5886,N_5613,N_5622);
nand U5887 (N_5887,N_5587,N_5572);
nor U5888 (N_5888,N_5690,N_5607);
nand U5889 (N_5889,N_5534,N_5730);
and U5890 (N_5890,N_5565,N_5586);
or U5891 (N_5891,N_5675,N_5599);
nor U5892 (N_5892,N_5513,N_5600);
nand U5893 (N_5893,N_5623,N_5641);
and U5894 (N_5894,N_5691,N_5655);
or U5895 (N_5895,N_5602,N_5517);
and U5896 (N_5896,N_5678,N_5688);
or U5897 (N_5897,N_5578,N_5700);
or U5898 (N_5898,N_5601,N_5643);
nor U5899 (N_5899,N_5666,N_5607);
xnor U5900 (N_5900,N_5598,N_5675);
and U5901 (N_5901,N_5702,N_5592);
nand U5902 (N_5902,N_5697,N_5722);
nor U5903 (N_5903,N_5738,N_5562);
nand U5904 (N_5904,N_5703,N_5622);
xnor U5905 (N_5905,N_5644,N_5689);
xnor U5906 (N_5906,N_5737,N_5526);
xor U5907 (N_5907,N_5576,N_5605);
or U5908 (N_5908,N_5747,N_5682);
nand U5909 (N_5909,N_5500,N_5588);
xor U5910 (N_5910,N_5503,N_5506);
nand U5911 (N_5911,N_5616,N_5702);
or U5912 (N_5912,N_5665,N_5548);
and U5913 (N_5913,N_5722,N_5653);
or U5914 (N_5914,N_5724,N_5509);
xor U5915 (N_5915,N_5670,N_5672);
nand U5916 (N_5916,N_5611,N_5576);
or U5917 (N_5917,N_5563,N_5516);
or U5918 (N_5918,N_5656,N_5638);
or U5919 (N_5919,N_5711,N_5650);
nand U5920 (N_5920,N_5581,N_5526);
nand U5921 (N_5921,N_5597,N_5508);
or U5922 (N_5922,N_5656,N_5698);
xor U5923 (N_5923,N_5740,N_5719);
nand U5924 (N_5924,N_5725,N_5562);
nand U5925 (N_5925,N_5655,N_5624);
and U5926 (N_5926,N_5657,N_5561);
nand U5927 (N_5927,N_5601,N_5733);
and U5928 (N_5928,N_5685,N_5527);
nor U5929 (N_5929,N_5623,N_5537);
xnor U5930 (N_5930,N_5734,N_5666);
xnor U5931 (N_5931,N_5734,N_5565);
or U5932 (N_5932,N_5540,N_5682);
nor U5933 (N_5933,N_5701,N_5660);
xnor U5934 (N_5934,N_5700,N_5559);
or U5935 (N_5935,N_5601,N_5523);
nand U5936 (N_5936,N_5652,N_5642);
or U5937 (N_5937,N_5748,N_5681);
nor U5938 (N_5938,N_5691,N_5505);
nor U5939 (N_5939,N_5523,N_5670);
or U5940 (N_5940,N_5500,N_5613);
xnor U5941 (N_5941,N_5509,N_5678);
nand U5942 (N_5942,N_5556,N_5598);
xnor U5943 (N_5943,N_5720,N_5743);
nor U5944 (N_5944,N_5596,N_5610);
nor U5945 (N_5945,N_5708,N_5503);
xor U5946 (N_5946,N_5661,N_5735);
nor U5947 (N_5947,N_5673,N_5690);
xor U5948 (N_5948,N_5607,N_5637);
nand U5949 (N_5949,N_5732,N_5534);
nand U5950 (N_5950,N_5530,N_5708);
nand U5951 (N_5951,N_5530,N_5616);
or U5952 (N_5952,N_5647,N_5666);
or U5953 (N_5953,N_5518,N_5515);
xor U5954 (N_5954,N_5726,N_5661);
xnor U5955 (N_5955,N_5510,N_5661);
nor U5956 (N_5956,N_5559,N_5740);
xor U5957 (N_5957,N_5649,N_5615);
and U5958 (N_5958,N_5563,N_5542);
or U5959 (N_5959,N_5651,N_5617);
or U5960 (N_5960,N_5713,N_5657);
nor U5961 (N_5961,N_5631,N_5663);
nand U5962 (N_5962,N_5738,N_5684);
and U5963 (N_5963,N_5584,N_5517);
nor U5964 (N_5964,N_5527,N_5562);
and U5965 (N_5965,N_5529,N_5671);
xor U5966 (N_5966,N_5557,N_5504);
nand U5967 (N_5967,N_5731,N_5639);
and U5968 (N_5968,N_5583,N_5611);
or U5969 (N_5969,N_5584,N_5547);
or U5970 (N_5970,N_5521,N_5540);
and U5971 (N_5971,N_5571,N_5687);
nand U5972 (N_5972,N_5736,N_5612);
nand U5973 (N_5973,N_5520,N_5537);
and U5974 (N_5974,N_5518,N_5675);
xnor U5975 (N_5975,N_5537,N_5684);
nand U5976 (N_5976,N_5594,N_5675);
nor U5977 (N_5977,N_5567,N_5679);
nor U5978 (N_5978,N_5738,N_5554);
xor U5979 (N_5979,N_5667,N_5718);
xor U5980 (N_5980,N_5546,N_5647);
nor U5981 (N_5981,N_5501,N_5607);
and U5982 (N_5982,N_5626,N_5722);
or U5983 (N_5983,N_5701,N_5631);
nand U5984 (N_5984,N_5717,N_5646);
and U5985 (N_5985,N_5525,N_5732);
xor U5986 (N_5986,N_5694,N_5686);
nand U5987 (N_5987,N_5509,N_5552);
xor U5988 (N_5988,N_5711,N_5659);
or U5989 (N_5989,N_5530,N_5500);
xnor U5990 (N_5990,N_5727,N_5681);
xnor U5991 (N_5991,N_5505,N_5587);
nor U5992 (N_5992,N_5608,N_5554);
xor U5993 (N_5993,N_5591,N_5714);
and U5994 (N_5994,N_5648,N_5711);
nand U5995 (N_5995,N_5597,N_5724);
and U5996 (N_5996,N_5552,N_5550);
and U5997 (N_5997,N_5730,N_5651);
xnor U5998 (N_5998,N_5611,N_5659);
nor U5999 (N_5999,N_5719,N_5506);
and U6000 (N_6000,N_5810,N_5781);
xnor U6001 (N_6001,N_5866,N_5955);
nor U6002 (N_6002,N_5930,N_5813);
and U6003 (N_6003,N_5855,N_5932);
nor U6004 (N_6004,N_5987,N_5896);
nand U6005 (N_6005,N_5974,N_5949);
nor U6006 (N_6006,N_5939,N_5777);
xnor U6007 (N_6007,N_5938,N_5863);
and U6008 (N_6008,N_5767,N_5911);
or U6009 (N_6009,N_5837,N_5894);
nand U6010 (N_6010,N_5967,N_5796);
and U6011 (N_6011,N_5984,N_5970);
nor U6012 (N_6012,N_5768,N_5937);
nor U6013 (N_6013,N_5851,N_5758);
or U6014 (N_6014,N_5977,N_5988);
nand U6015 (N_6015,N_5785,N_5850);
nand U6016 (N_6016,N_5901,N_5854);
nor U6017 (N_6017,N_5954,N_5789);
nand U6018 (N_6018,N_5957,N_5926);
nor U6019 (N_6019,N_5834,N_5961);
or U6020 (N_6020,N_5880,N_5818);
nand U6021 (N_6021,N_5795,N_5873);
or U6022 (N_6022,N_5819,N_5890);
nand U6023 (N_6023,N_5846,N_5871);
nor U6024 (N_6024,N_5841,N_5815);
nor U6025 (N_6025,N_5919,N_5852);
or U6026 (N_6026,N_5848,N_5759);
xnor U6027 (N_6027,N_5836,N_5772);
nor U6028 (N_6028,N_5843,N_5842);
nor U6029 (N_6029,N_5760,N_5904);
nand U6030 (N_6030,N_5912,N_5933);
and U6031 (N_6031,N_5875,N_5770);
and U6032 (N_6032,N_5989,N_5874);
nor U6033 (N_6033,N_5824,N_5833);
xnor U6034 (N_6034,N_5997,N_5940);
nand U6035 (N_6035,N_5865,N_5862);
nor U6036 (N_6036,N_5787,N_5931);
nand U6037 (N_6037,N_5840,N_5895);
or U6038 (N_6038,N_5956,N_5820);
xnor U6039 (N_6039,N_5798,N_5853);
or U6040 (N_6040,N_5868,N_5838);
xnor U6041 (N_6041,N_5832,N_5946);
nor U6042 (N_6042,N_5879,N_5808);
nor U6043 (N_6043,N_5928,N_5952);
nor U6044 (N_6044,N_5971,N_5792);
xnor U6045 (N_6045,N_5965,N_5968);
or U6046 (N_6046,N_5822,N_5812);
and U6047 (N_6047,N_5753,N_5979);
nand U6048 (N_6048,N_5992,N_5814);
and U6049 (N_6049,N_5953,N_5976);
nand U6050 (N_6050,N_5856,N_5766);
and U6051 (N_6051,N_5802,N_5864);
nor U6052 (N_6052,N_5908,N_5877);
or U6053 (N_6053,N_5828,N_5751);
and U6054 (N_6054,N_5950,N_5793);
or U6055 (N_6055,N_5788,N_5907);
and U6056 (N_6056,N_5891,N_5906);
and U6057 (N_6057,N_5774,N_5993);
nand U6058 (N_6058,N_5831,N_5914);
and U6059 (N_6059,N_5804,N_5801);
and U6060 (N_6060,N_5975,N_5757);
nor U6061 (N_6061,N_5985,N_5839);
and U6062 (N_6062,N_5917,N_5948);
or U6063 (N_6063,N_5921,N_5966);
nor U6064 (N_6064,N_5927,N_5916);
or U6065 (N_6065,N_5797,N_5799);
or U6066 (N_6066,N_5978,N_5756);
xnor U6067 (N_6067,N_5805,N_5972);
and U6068 (N_6068,N_5915,N_5959);
and U6069 (N_6069,N_5951,N_5990);
nand U6070 (N_6070,N_5876,N_5821);
or U6071 (N_6071,N_5964,N_5755);
xnor U6072 (N_6072,N_5935,N_5943);
nor U6073 (N_6073,N_5769,N_5859);
nand U6074 (N_6074,N_5776,N_5924);
or U6075 (N_6075,N_5936,N_5980);
nor U6076 (N_6076,N_5860,N_5934);
nand U6077 (N_6077,N_5790,N_5897);
and U6078 (N_6078,N_5825,N_5762);
and U6079 (N_6079,N_5761,N_5765);
or U6080 (N_6080,N_5809,N_5958);
or U6081 (N_6081,N_5902,N_5807);
or U6082 (N_6082,N_5754,N_5983);
nand U6083 (N_6083,N_5986,N_5925);
and U6084 (N_6084,N_5942,N_5878);
or U6085 (N_6085,N_5991,N_5888);
and U6086 (N_6086,N_5783,N_5922);
nor U6087 (N_6087,N_5920,N_5981);
or U6088 (N_6088,N_5969,N_5889);
nand U6089 (N_6089,N_5794,N_5886);
or U6090 (N_6090,N_5918,N_5887);
nand U6091 (N_6091,N_5847,N_5867);
and U6092 (N_6092,N_5827,N_5803);
and U6093 (N_6093,N_5929,N_5913);
nor U6094 (N_6094,N_5903,N_5800);
nand U6095 (N_6095,N_5780,N_5885);
xor U6096 (N_6096,N_5923,N_5791);
and U6097 (N_6097,N_5773,N_5830);
nor U6098 (N_6098,N_5849,N_5806);
and U6099 (N_6099,N_5829,N_5899);
and U6100 (N_6100,N_5870,N_5778);
xnor U6101 (N_6101,N_5910,N_5779);
or U6102 (N_6102,N_5881,N_5905);
nand U6103 (N_6103,N_5883,N_5893);
nor U6104 (N_6104,N_5750,N_5944);
xor U6105 (N_6105,N_5900,N_5845);
nand U6106 (N_6106,N_5775,N_5996);
nor U6107 (N_6107,N_5826,N_5861);
nand U6108 (N_6108,N_5947,N_5857);
nor U6109 (N_6109,N_5869,N_5962);
xnor U6110 (N_6110,N_5817,N_5909);
or U6111 (N_6111,N_5882,N_5811);
and U6112 (N_6112,N_5982,N_5786);
or U6113 (N_6113,N_5995,N_5858);
nor U6114 (N_6114,N_5999,N_5941);
and U6115 (N_6115,N_5898,N_5960);
or U6116 (N_6116,N_5752,N_5998);
or U6117 (N_6117,N_5844,N_5763);
or U6118 (N_6118,N_5835,N_5945);
xnor U6119 (N_6119,N_5784,N_5764);
or U6120 (N_6120,N_5872,N_5823);
nand U6121 (N_6121,N_5994,N_5782);
nand U6122 (N_6122,N_5771,N_5892);
nand U6123 (N_6123,N_5973,N_5963);
and U6124 (N_6124,N_5884,N_5816);
and U6125 (N_6125,N_5941,N_5940);
and U6126 (N_6126,N_5770,N_5811);
nand U6127 (N_6127,N_5929,N_5806);
nor U6128 (N_6128,N_5808,N_5914);
nand U6129 (N_6129,N_5853,N_5831);
nor U6130 (N_6130,N_5915,N_5992);
xor U6131 (N_6131,N_5794,N_5965);
nand U6132 (N_6132,N_5961,N_5771);
and U6133 (N_6133,N_5964,N_5772);
xnor U6134 (N_6134,N_5896,N_5907);
xnor U6135 (N_6135,N_5888,N_5753);
nand U6136 (N_6136,N_5771,N_5857);
and U6137 (N_6137,N_5910,N_5887);
and U6138 (N_6138,N_5818,N_5795);
nand U6139 (N_6139,N_5938,N_5794);
nand U6140 (N_6140,N_5762,N_5874);
nor U6141 (N_6141,N_5897,N_5807);
and U6142 (N_6142,N_5881,N_5985);
nor U6143 (N_6143,N_5889,N_5776);
xnor U6144 (N_6144,N_5818,N_5754);
nor U6145 (N_6145,N_5957,N_5872);
nand U6146 (N_6146,N_5884,N_5857);
xor U6147 (N_6147,N_5845,N_5877);
xor U6148 (N_6148,N_5961,N_5977);
nand U6149 (N_6149,N_5795,N_5816);
nand U6150 (N_6150,N_5843,N_5932);
nor U6151 (N_6151,N_5807,N_5926);
and U6152 (N_6152,N_5960,N_5762);
or U6153 (N_6153,N_5930,N_5846);
nor U6154 (N_6154,N_5866,N_5885);
xnor U6155 (N_6155,N_5768,N_5771);
or U6156 (N_6156,N_5845,N_5820);
and U6157 (N_6157,N_5782,N_5788);
xor U6158 (N_6158,N_5800,N_5835);
nand U6159 (N_6159,N_5958,N_5907);
xor U6160 (N_6160,N_5892,N_5852);
nor U6161 (N_6161,N_5768,N_5778);
or U6162 (N_6162,N_5809,N_5929);
nor U6163 (N_6163,N_5798,N_5759);
xor U6164 (N_6164,N_5796,N_5837);
xor U6165 (N_6165,N_5838,N_5867);
nand U6166 (N_6166,N_5801,N_5896);
or U6167 (N_6167,N_5771,N_5844);
nor U6168 (N_6168,N_5994,N_5973);
nand U6169 (N_6169,N_5975,N_5888);
nand U6170 (N_6170,N_5882,N_5794);
xor U6171 (N_6171,N_5795,N_5826);
nor U6172 (N_6172,N_5968,N_5754);
or U6173 (N_6173,N_5962,N_5828);
nand U6174 (N_6174,N_5988,N_5817);
nor U6175 (N_6175,N_5958,N_5983);
and U6176 (N_6176,N_5845,N_5969);
nand U6177 (N_6177,N_5989,N_5792);
nor U6178 (N_6178,N_5958,N_5929);
or U6179 (N_6179,N_5925,N_5946);
xor U6180 (N_6180,N_5921,N_5886);
nor U6181 (N_6181,N_5960,N_5948);
or U6182 (N_6182,N_5772,N_5776);
nor U6183 (N_6183,N_5961,N_5804);
and U6184 (N_6184,N_5908,N_5925);
xor U6185 (N_6185,N_5903,N_5830);
or U6186 (N_6186,N_5972,N_5895);
xor U6187 (N_6187,N_5849,N_5796);
nor U6188 (N_6188,N_5812,N_5815);
or U6189 (N_6189,N_5832,N_5856);
or U6190 (N_6190,N_5818,N_5895);
nand U6191 (N_6191,N_5802,N_5775);
xnor U6192 (N_6192,N_5936,N_5810);
xor U6193 (N_6193,N_5774,N_5836);
nor U6194 (N_6194,N_5927,N_5897);
and U6195 (N_6195,N_5886,N_5939);
and U6196 (N_6196,N_5907,N_5981);
or U6197 (N_6197,N_5814,N_5990);
nor U6198 (N_6198,N_5988,N_5942);
nand U6199 (N_6199,N_5845,N_5779);
xnor U6200 (N_6200,N_5844,N_5980);
nand U6201 (N_6201,N_5811,N_5839);
or U6202 (N_6202,N_5833,N_5853);
or U6203 (N_6203,N_5786,N_5825);
xor U6204 (N_6204,N_5913,N_5810);
xor U6205 (N_6205,N_5752,N_5861);
and U6206 (N_6206,N_5827,N_5890);
or U6207 (N_6207,N_5807,N_5943);
xnor U6208 (N_6208,N_5910,N_5920);
nand U6209 (N_6209,N_5820,N_5903);
and U6210 (N_6210,N_5922,N_5851);
or U6211 (N_6211,N_5781,N_5866);
xnor U6212 (N_6212,N_5907,N_5977);
nor U6213 (N_6213,N_5991,N_5845);
nand U6214 (N_6214,N_5869,N_5978);
xor U6215 (N_6215,N_5795,N_5783);
and U6216 (N_6216,N_5937,N_5947);
and U6217 (N_6217,N_5839,N_5942);
and U6218 (N_6218,N_5917,N_5927);
nor U6219 (N_6219,N_5810,N_5825);
xor U6220 (N_6220,N_5994,N_5908);
and U6221 (N_6221,N_5874,N_5967);
nand U6222 (N_6222,N_5947,N_5910);
xor U6223 (N_6223,N_5780,N_5802);
and U6224 (N_6224,N_5955,N_5770);
nand U6225 (N_6225,N_5805,N_5776);
or U6226 (N_6226,N_5985,N_5974);
nor U6227 (N_6227,N_5938,N_5832);
nand U6228 (N_6228,N_5861,N_5885);
nand U6229 (N_6229,N_5922,N_5771);
or U6230 (N_6230,N_5889,N_5974);
nand U6231 (N_6231,N_5802,N_5897);
or U6232 (N_6232,N_5995,N_5967);
nand U6233 (N_6233,N_5925,N_5905);
and U6234 (N_6234,N_5805,N_5990);
or U6235 (N_6235,N_5824,N_5946);
xnor U6236 (N_6236,N_5968,N_5960);
or U6237 (N_6237,N_5855,N_5951);
or U6238 (N_6238,N_5925,N_5969);
nor U6239 (N_6239,N_5992,N_5904);
or U6240 (N_6240,N_5951,N_5887);
nor U6241 (N_6241,N_5851,N_5825);
nor U6242 (N_6242,N_5838,N_5986);
and U6243 (N_6243,N_5808,N_5940);
or U6244 (N_6244,N_5768,N_5786);
xnor U6245 (N_6245,N_5813,N_5974);
xor U6246 (N_6246,N_5798,N_5925);
or U6247 (N_6247,N_5818,N_5768);
and U6248 (N_6248,N_5787,N_5981);
and U6249 (N_6249,N_5957,N_5786);
or U6250 (N_6250,N_6013,N_6185);
and U6251 (N_6251,N_6181,N_6169);
and U6252 (N_6252,N_6008,N_6066);
xnor U6253 (N_6253,N_6166,N_6159);
or U6254 (N_6254,N_6041,N_6020);
or U6255 (N_6255,N_6133,N_6113);
and U6256 (N_6256,N_6165,N_6168);
xor U6257 (N_6257,N_6043,N_6059);
and U6258 (N_6258,N_6176,N_6045);
or U6259 (N_6259,N_6068,N_6147);
xor U6260 (N_6260,N_6153,N_6070);
nand U6261 (N_6261,N_6017,N_6227);
and U6262 (N_6262,N_6178,N_6237);
xnor U6263 (N_6263,N_6230,N_6211);
and U6264 (N_6264,N_6038,N_6218);
nand U6265 (N_6265,N_6145,N_6188);
nor U6266 (N_6266,N_6240,N_6057);
or U6267 (N_6267,N_6044,N_6026);
xor U6268 (N_6268,N_6174,N_6122);
and U6269 (N_6269,N_6137,N_6238);
and U6270 (N_6270,N_6042,N_6002);
xnor U6271 (N_6271,N_6035,N_6050);
and U6272 (N_6272,N_6074,N_6106);
nor U6273 (N_6273,N_6183,N_6047);
nand U6274 (N_6274,N_6032,N_6156);
and U6275 (N_6275,N_6158,N_6239);
nor U6276 (N_6276,N_6061,N_6036);
nand U6277 (N_6277,N_6062,N_6224);
xnor U6278 (N_6278,N_6099,N_6162);
xnor U6279 (N_6279,N_6234,N_6131);
nor U6280 (N_6280,N_6167,N_6023);
and U6281 (N_6281,N_6246,N_6187);
xor U6282 (N_6282,N_6228,N_6104);
or U6283 (N_6283,N_6049,N_6090);
and U6284 (N_6284,N_6076,N_6132);
nor U6285 (N_6285,N_6248,N_6190);
xnor U6286 (N_6286,N_6005,N_6103);
or U6287 (N_6287,N_6154,N_6189);
or U6288 (N_6288,N_6182,N_6112);
nand U6289 (N_6289,N_6051,N_6121);
and U6290 (N_6290,N_6069,N_6083);
nor U6291 (N_6291,N_6192,N_6216);
xor U6292 (N_6292,N_6223,N_6202);
nand U6293 (N_6293,N_6152,N_6204);
nand U6294 (N_6294,N_6033,N_6136);
or U6295 (N_6295,N_6195,N_6207);
xor U6296 (N_6296,N_6079,N_6040);
xor U6297 (N_6297,N_6086,N_6117);
nand U6298 (N_6298,N_6193,N_6191);
or U6299 (N_6299,N_6214,N_6096);
xnor U6300 (N_6300,N_6134,N_6215);
and U6301 (N_6301,N_6012,N_6179);
and U6302 (N_6302,N_6011,N_6205);
xor U6303 (N_6303,N_6072,N_6082);
nand U6304 (N_6304,N_6025,N_6243);
or U6305 (N_6305,N_6115,N_6031);
xnor U6306 (N_6306,N_6039,N_6199);
nor U6307 (N_6307,N_6063,N_6155);
and U6308 (N_6308,N_6100,N_6089);
nor U6309 (N_6309,N_6245,N_6180);
and U6310 (N_6310,N_6014,N_6004);
or U6311 (N_6311,N_6016,N_6060);
or U6312 (N_6312,N_6030,N_6077);
and U6313 (N_6313,N_6236,N_6110);
nand U6314 (N_6314,N_6128,N_6015);
nand U6315 (N_6315,N_6209,N_6226);
or U6316 (N_6316,N_6138,N_6171);
xnor U6317 (N_6317,N_6056,N_6092);
xnor U6318 (N_6318,N_6139,N_6130);
xor U6319 (N_6319,N_6151,N_6196);
and U6320 (N_6320,N_6124,N_6194);
nor U6321 (N_6321,N_6007,N_6241);
or U6322 (N_6322,N_6078,N_6127);
and U6323 (N_6323,N_6114,N_6098);
nand U6324 (N_6324,N_6225,N_6198);
or U6325 (N_6325,N_6095,N_6144);
nor U6326 (N_6326,N_6029,N_6107);
nor U6327 (N_6327,N_6231,N_6048);
and U6328 (N_6328,N_6233,N_6105);
xor U6329 (N_6329,N_6102,N_6081);
nor U6330 (N_6330,N_6173,N_6054);
xnor U6331 (N_6331,N_6009,N_6142);
and U6332 (N_6332,N_6160,N_6170);
and U6333 (N_6333,N_6071,N_6157);
xnor U6334 (N_6334,N_6203,N_6125);
nand U6335 (N_6335,N_6101,N_6242);
or U6336 (N_6336,N_6097,N_6119);
xor U6337 (N_6337,N_6212,N_6148);
and U6338 (N_6338,N_6210,N_6172);
xnor U6339 (N_6339,N_6088,N_6052);
nor U6340 (N_6340,N_6085,N_6163);
and U6341 (N_6341,N_6094,N_6164);
nor U6342 (N_6342,N_6001,N_6150);
xor U6343 (N_6343,N_6175,N_6232);
or U6344 (N_6344,N_6080,N_6000);
xnor U6345 (N_6345,N_6186,N_6037);
or U6346 (N_6346,N_6244,N_6084);
xnor U6347 (N_6347,N_6093,N_6024);
and U6348 (N_6348,N_6247,N_6221);
nor U6349 (N_6349,N_6006,N_6177);
nor U6350 (N_6350,N_6220,N_6197);
and U6351 (N_6351,N_6065,N_6208);
or U6352 (N_6352,N_6010,N_6201);
nor U6353 (N_6353,N_6141,N_6027);
xor U6354 (N_6354,N_6149,N_6058);
nor U6355 (N_6355,N_6111,N_6126);
or U6356 (N_6356,N_6200,N_6123);
nand U6357 (N_6357,N_6046,N_6022);
nor U6358 (N_6358,N_6213,N_6249);
and U6359 (N_6359,N_6073,N_6108);
and U6360 (N_6360,N_6064,N_6109);
xnor U6361 (N_6361,N_6003,N_6019);
or U6362 (N_6362,N_6140,N_6219);
and U6363 (N_6363,N_6116,N_6235);
xnor U6364 (N_6364,N_6120,N_6184);
xnor U6365 (N_6365,N_6146,N_6222);
and U6366 (N_6366,N_6028,N_6053);
nor U6367 (N_6367,N_6118,N_6217);
or U6368 (N_6368,N_6034,N_6055);
nand U6369 (N_6369,N_6229,N_6206);
and U6370 (N_6370,N_6091,N_6135);
nand U6371 (N_6371,N_6161,N_6129);
and U6372 (N_6372,N_6018,N_6087);
nand U6373 (N_6373,N_6021,N_6143);
nor U6374 (N_6374,N_6067,N_6075);
and U6375 (N_6375,N_6145,N_6036);
or U6376 (N_6376,N_6197,N_6163);
and U6377 (N_6377,N_6180,N_6201);
xor U6378 (N_6378,N_6057,N_6094);
or U6379 (N_6379,N_6077,N_6249);
or U6380 (N_6380,N_6115,N_6129);
and U6381 (N_6381,N_6021,N_6162);
or U6382 (N_6382,N_6160,N_6188);
or U6383 (N_6383,N_6069,N_6093);
xor U6384 (N_6384,N_6031,N_6162);
or U6385 (N_6385,N_6073,N_6176);
and U6386 (N_6386,N_6141,N_6080);
nor U6387 (N_6387,N_6077,N_6044);
or U6388 (N_6388,N_6006,N_6210);
and U6389 (N_6389,N_6037,N_6004);
nand U6390 (N_6390,N_6167,N_6178);
nand U6391 (N_6391,N_6160,N_6175);
xnor U6392 (N_6392,N_6083,N_6205);
xnor U6393 (N_6393,N_6014,N_6215);
or U6394 (N_6394,N_6030,N_6004);
or U6395 (N_6395,N_6096,N_6209);
and U6396 (N_6396,N_6077,N_6176);
xor U6397 (N_6397,N_6159,N_6244);
xnor U6398 (N_6398,N_6168,N_6109);
nand U6399 (N_6399,N_6193,N_6057);
nor U6400 (N_6400,N_6143,N_6152);
nor U6401 (N_6401,N_6100,N_6128);
xor U6402 (N_6402,N_6199,N_6191);
or U6403 (N_6403,N_6008,N_6020);
nor U6404 (N_6404,N_6149,N_6223);
nand U6405 (N_6405,N_6009,N_6206);
nand U6406 (N_6406,N_6160,N_6142);
nor U6407 (N_6407,N_6130,N_6090);
and U6408 (N_6408,N_6025,N_6244);
nand U6409 (N_6409,N_6157,N_6154);
and U6410 (N_6410,N_6080,N_6037);
nor U6411 (N_6411,N_6162,N_6041);
nor U6412 (N_6412,N_6242,N_6205);
nand U6413 (N_6413,N_6150,N_6232);
nor U6414 (N_6414,N_6177,N_6128);
or U6415 (N_6415,N_6144,N_6236);
nor U6416 (N_6416,N_6104,N_6223);
nand U6417 (N_6417,N_6167,N_6202);
xor U6418 (N_6418,N_6053,N_6043);
and U6419 (N_6419,N_6207,N_6010);
nor U6420 (N_6420,N_6173,N_6037);
and U6421 (N_6421,N_6234,N_6230);
or U6422 (N_6422,N_6086,N_6240);
or U6423 (N_6423,N_6247,N_6170);
or U6424 (N_6424,N_6205,N_6200);
and U6425 (N_6425,N_6203,N_6034);
or U6426 (N_6426,N_6223,N_6097);
or U6427 (N_6427,N_6213,N_6150);
nor U6428 (N_6428,N_6167,N_6206);
nor U6429 (N_6429,N_6099,N_6154);
xor U6430 (N_6430,N_6218,N_6204);
nor U6431 (N_6431,N_6196,N_6126);
or U6432 (N_6432,N_6025,N_6190);
and U6433 (N_6433,N_6012,N_6090);
nand U6434 (N_6434,N_6019,N_6069);
or U6435 (N_6435,N_6245,N_6201);
xor U6436 (N_6436,N_6125,N_6089);
and U6437 (N_6437,N_6127,N_6137);
or U6438 (N_6438,N_6229,N_6104);
xor U6439 (N_6439,N_6186,N_6174);
or U6440 (N_6440,N_6243,N_6199);
and U6441 (N_6441,N_6148,N_6129);
and U6442 (N_6442,N_6085,N_6231);
xnor U6443 (N_6443,N_6016,N_6245);
or U6444 (N_6444,N_6205,N_6220);
nor U6445 (N_6445,N_6246,N_6033);
nand U6446 (N_6446,N_6054,N_6122);
and U6447 (N_6447,N_6022,N_6005);
nor U6448 (N_6448,N_6041,N_6137);
xnor U6449 (N_6449,N_6203,N_6155);
nor U6450 (N_6450,N_6129,N_6112);
nor U6451 (N_6451,N_6080,N_6043);
nor U6452 (N_6452,N_6091,N_6147);
and U6453 (N_6453,N_6168,N_6120);
nor U6454 (N_6454,N_6097,N_6061);
and U6455 (N_6455,N_6018,N_6164);
nor U6456 (N_6456,N_6033,N_6093);
nand U6457 (N_6457,N_6196,N_6166);
nand U6458 (N_6458,N_6147,N_6100);
and U6459 (N_6459,N_6098,N_6229);
or U6460 (N_6460,N_6180,N_6050);
or U6461 (N_6461,N_6024,N_6019);
xor U6462 (N_6462,N_6045,N_6064);
nor U6463 (N_6463,N_6201,N_6177);
or U6464 (N_6464,N_6009,N_6228);
or U6465 (N_6465,N_6084,N_6153);
and U6466 (N_6466,N_6225,N_6022);
xnor U6467 (N_6467,N_6020,N_6040);
or U6468 (N_6468,N_6077,N_6199);
nor U6469 (N_6469,N_6002,N_6136);
and U6470 (N_6470,N_6052,N_6001);
and U6471 (N_6471,N_6025,N_6023);
xnor U6472 (N_6472,N_6085,N_6049);
or U6473 (N_6473,N_6114,N_6103);
and U6474 (N_6474,N_6148,N_6160);
or U6475 (N_6475,N_6240,N_6118);
or U6476 (N_6476,N_6024,N_6226);
xor U6477 (N_6477,N_6010,N_6193);
and U6478 (N_6478,N_6194,N_6140);
xnor U6479 (N_6479,N_6156,N_6172);
and U6480 (N_6480,N_6030,N_6172);
xnor U6481 (N_6481,N_6181,N_6193);
nand U6482 (N_6482,N_6159,N_6201);
and U6483 (N_6483,N_6045,N_6063);
nand U6484 (N_6484,N_6226,N_6147);
and U6485 (N_6485,N_6109,N_6234);
or U6486 (N_6486,N_6139,N_6244);
nand U6487 (N_6487,N_6090,N_6040);
and U6488 (N_6488,N_6131,N_6014);
xnor U6489 (N_6489,N_6202,N_6133);
nand U6490 (N_6490,N_6229,N_6035);
and U6491 (N_6491,N_6152,N_6075);
or U6492 (N_6492,N_6210,N_6022);
nand U6493 (N_6493,N_6240,N_6142);
nor U6494 (N_6494,N_6225,N_6185);
xor U6495 (N_6495,N_6126,N_6027);
nand U6496 (N_6496,N_6057,N_6083);
nand U6497 (N_6497,N_6204,N_6065);
nor U6498 (N_6498,N_6195,N_6075);
and U6499 (N_6499,N_6135,N_6096);
nand U6500 (N_6500,N_6340,N_6277);
nand U6501 (N_6501,N_6405,N_6300);
nand U6502 (N_6502,N_6395,N_6272);
and U6503 (N_6503,N_6275,N_6386);
nor U6504 (N_6504,N_6389,N_6298);
xnor U6505 (N_6505,N_6454,N_6486);
nand U6506 (N_6506,N_6335,N_6318);
and U6507 (N_6507,N_6338,N_6266);
or U6508 (N_6508,N_6323,N_6437);
xor U6509 (N_6509,N_6351,N_6418);
nor U6510 (N_6510,N_6406,N_6430);
nor U6511 (N_6511,N_6281,N_6285);
xnor U6512 (N_6512,N_6381,N_6439);
nand U6513 (N_6513,N_6304,N_6403);
nand U6514 (N_6514,N_6459,N_6413);
and U6515 (N_6515,N_6470,N_6344);
nand U6516 (N_6516,N_6356,N_6354);
or U6517 (N_6517,N_6267,N_6326);
nor U6518 (N_6518,N_6442,N_6489);
nor U6519 (N_6519,N_6445,N_6319);
xor U6520 (N_6520,N_6460,N_6457);
and U6521 (N_6521,N_6301,N_6481);
nand U6522 (N_6522,N_6333,N_6369);
nand U6523 (N_6523,N_6312,N_6392);
nor U6524 (N_6524,N_6342,N_6420);
or U6525 (N_6525,N_6366,N_6363);
xnor U6526 (N_6526,N_6327,N_6296);
or U6527 (N_6527,N_6265,N_6484);
and U6528 (N_6528,N_6339,N_6350);
xor U6529 (N_6529,N_6260,N_6379);
nor U6530 (N_6530,N_6295,N_6343);
nor U6531 (N_6531,N_6436,N_6331);
and U6532 (N_6532,N_6357,N_6468);
nor U6533 (N_6533,N_6269,N_6255);
nand U6534 (N_6534,N_6416,N_6314);
or U6535 (N_6535,N_6419,N_6313);
xnor U6536 (N_6536,N_6299,N_6496);
nand U6537 (N_6537,N_6359,N_6257);
nor U6538 (N_6538,N_6493,N_6310);
xnor U6539 (N_6539,N_6495,N_6407);
or U6540 (N_6540,N_6377,N_6380);
nor U6541 (N_6541,N_6293,N_6308);
xor U6542 (N_6542,N_6458,N_6303);
or U6543 (N_6543,N_6251,N_6316);
and U6544 (N_6544,N_6402,N_6353);
nand U6545 (N_6545,N_6305,N_6446);
nand U6546 (N_6546,N_6273,N_6280);
xnor U6547 (N_6547,N_6271,N_6401);
and U6548 (N_6548,N_6261,N_6375);
nor U6549 (N_6549,N_6412,N_6371);
and U6550 (N_6550,N_6411,N_6428);
nor U6551 (N_6551,N_6394,N_6367);
nor U6552 (N_6552,N_6317,N_6337);
nor U6553 (N_6553,N_6288,N_6362);
nor U6554 (N_6554,N_6347,N_6341);
or U6555 (N_6555,N_6276,N_6348);
nor U6556 (N_6556,N_6441,N_6487);
and U6557 (N_6557,N_6302,N_6452);
nand U6558 (N_6558,N_6480,N_6451);
and U6559 (N_6559,N_6398,N_6384);
nand U6560 (N_6560,N_6252,N_6315);
and U6561 (N_6561,N_6426,N_6438);
xnor U6562 (N_6562,N_6453,N_6250);
and U6563 (N_6563,N_6283,N_6393);
nor U6564 (N_6564,N_6262,N_6471);
nor U6565 (N_6565,N_6254,N_6469);
or U6566 (N_6566,N_6372,N_6455);
nand U6567 (N_6567,N_6488,N_6424);
or U6568 (N_6568,N_6473,N_6408);
nor U6569 (N_6569,N_6440,N_6490);
nor U6570 (N_6570,N_6332,N_6425);
nand U6571 (N_6571,N_6434,N_6382);
and U6572 (N_6572,N_6361,N_6387);
nor U6573 (N_6573,N_6461,N_6433);
nand U6574 (N_6574,N_6499,N_6378);
nor U6575 (N_6575,N_6328,N_6329);
and U6576 (N_6576,N_6467,N_6309);
nand U6577 (N_6577,N_6383,N_6294);
nor U6578 (N_6578,N_6306,N_6409);
xor U6579 (N_6579,N_6345,N_6476);
nand U6580 (N_6580,N_6324,N_6376);
or U6581 (N_6581,N_6368,N_6270);
nand U6582 (N_6582,N_6464,N_6259);
xnor U6583 (N_6583,N_6390,N_6292);
and U6584 (N_6584,N_6448,N_6475);
and U6585 (N_6585,N_6482,N_6494);
nor U6586 (N_6586,N_6391,N_6397);
or U6587 (N_6587,N_6360,N_6421);
nand U6588 (N_6588,N_6410,N_6497);
xnor U6589 (N_6589,N_6462,N_6365);
xor U6590 (N_6590,N_6320,N_6336);
nand U6591 (N_6591,N_6289,N_6474);
or U6592 (N_6592,N_6447,N_6492);
xnor U6593 (N_6593,N_6286,N_6290);
nand U6594 (N_6594,N_6274,N_6429);
nand U6595 (N_6595,N_6431,N_6256);
nor U6596 (N_6596,N_6472,N_6449);
nor U6597 (N_6597,N_6352,N_6491);
nand U6598 (N_6598,N_6479,N_6334);
or U6599 (N_6599,N_6435,N_6417);
xor U6600 (N_6600,N_6465,N_6355);
xor U6601 (N_6601,N_6330,N_6423);
or U6602 (N_6602,N_6385,N_6399);
xnor U6603 (N_6603,N_6263,N_6400);
or U6604 (N_6604,N_6450,N_6427);
nand U6605 (N_6605,N_6422,N_6404);
or U6606 (N_6606,N_6374,N_6443);
and U6607 (N_6607,N_6297,N_6415);
xor U6608 (N_6608,N_6485,N_6311);
xnor U6609 (N_6609,N_6456,N_6466);
xnor U6610 (N_6610,N_6349,N_6321);
nand U6611 (N_6611,N_6364,N_6370);
nand U6612 (N_6612,N_6498,N_6307);
or U6613 (N_6613,N_6325,N_6258);
xor U6614 (N_6614,N_6388,N_6432);
and U6615 (N_6615,N_6444,N_6414);
nor U6616 (N_6616,N_6291,N_6278);
nand U6617 (N_6617,N_6373,N_6358);
or U6618 (N_6618,N_6478,N_6253);
xnor U6619 (N_6619,N_6483,N_6282);
xnor U6620 (N_6620,N_6346,N_6279);
nor U6621 (N_6621,N_6322,N_6287);
nor U6622 (N_6622,N_6396,N_6264);
or U6623 (N_6623,N_6463,N_6284);
nand U6624 (N_6624,N_6477,N_6268);
nor U6625 (N_6625,N_6314,N_6347);
nor U6626 (N_6626,N_6388,N_6320);
nor U6627 (N_6627,N_6386,N_6356);
or U6628 (N_6628,N_6386,N_6362);
xor U6629 (N_6629,N_6316,N_6424);
xor U6630 (N_6630,N_6427,N_6426);
or U6631 (N_6631,N_6301,N_6267);
nand U6632 (N_6632,N_6440,N_6338);
or U6633 (N_6633,N_6437,N_6496);
or U6634 (N_6634,N_6252,N_6371);
nand U6635 (N_6635,N_6499,N_6411);
nand U6636 (N_6636,N_6485,N_6296);
xor U6637 (N_6637,N_6374,N_6345);
nor U6638 (N_6638,N_6369,N_6471);
xor U6639 (N_6639,N_6368,N_6372);
nor U6640 (N_6640,N_6389,N_6361);
and U6641 (N_6641,N_6368,N_6383);
xnor U6642 (N_6642,N_6267,N_6288);
or U6643 (N_6643,N_6434,N_6496);
and U6644 (N_6644,N_6473,N_6389);
xor U6645 (N_6645,N_6384,N_6412);
nor U6646 (N_6646,N_6361,N_6293);
nor U6647 (N_6647,N_6257,N_6479);
xnor U6648 (N_6648,N_6254,N_6432);
and U6649 (N_6649,N_6280,N_6401);
nor U6650 (N_6650,N_6266,N_6469);
xnor U6651 (N_6651,N_6342,N_6307);
nand U6652 (N_6652,N_6303,N_6429);
nand U6653 (N_6653,N_6330,N_6387);
or U6654 (N_6654,N_6287,N_6363);
nor U6655 (N_6655,N_6414,N_6484);
or U6656 (N_6656,N_6394,N_6295);
and U6657 (N_6657,N_6418,N_6461);
nor U6658 (N_6658,N_6454,N_6358);
and U6659 (N_6659,N_6326,N_6439);
or U6660 (N_6660,N_6484,N_6378);
nor U6661 (N_6661,N_6406,N_6471);
or U6662 (N_6662,N_6324,N_6360);
and U6663 (N_6663,N_6463,N_6438);
xor U6664 (N_6664,N_6433,N_6286);
nor U6665 (N_6665,N_6451,N_6392);
nor U6666 (N_6666,N_6475,N_6410);
nor U6667 (N_6667,N_6430,N_6441);
nand U6668 (N_6668,N_6324,N_6382);
nand U6669 (N_6669,N_6408,N_6257);
nor U6670 (N_6670,N_6277,N_6252);
nand U6671 (N_6671,N_6393,N_6398);
or U6672 (N_6672,N_6347,N_6455);
xnor U6673 (N_6673,N_6436,N_6288);
or U6674 (N_6674,N_6356,N_6466);
or U6675 (N_6675,N_6314,N_6385);
or U6676 (N_6676,N_6302,N_6401);
or U6677 (N_6677,N_6310,N_6439);
and U6678 (N_6678,N_6354,N_6309);
nor U6679 (N_6679,N_6349,N_6427);
nand U6680 (N_6680,N_6427,N_6294);
or U6681 (N_6681,N_6479,N_6406);
xnor U6682 (N_6682,N_6293,N_6420);
nor U6683 (N_6683,N_6355,N_6445);
nor U6684 (N_6684,N_6336,N_6278);
or U6685 (N_6685,N_6330,N_6259);
or U6686 (N_6686,N_6271,N_6301);
nand U6687 (N_6687,N_6298,N_6412);
and U6688 (N_6688,N_6481,N_6492);
nor U6689 (N_6689,N_6476,N_6263);
or U6690 (N_6690,N_6333,N_6386);
nor U6691 (N_6691,N_6468,N_6442);
nor U6692 (N_6692,N_6252,N_6401);
nand U6693 (N_6693,N_6455,N_6496);
or U6694 (N_6694,N_6469,N_6293);
nand U6695 (N_6695,N_6466,N_6335);
or U6696 (N_6696,N_6492,N_6495);
nor U6697 (N_6697,N_6309,N_6370);
nor U6698 (N_6698,N_6496,N_6447);
and U6699 (N_6699,N_6314,N_6365);
xnor U6700 (N_6700,N_6343,N_6456);
or U6701 (N_6701,N_6346,N_6283);
nor U6702 (N_6702,N_6442,N_6274);
xor U6703 (N_6703,N_6438,N_6476);
nor U6704 (N_6704,N_6297,N_6253);
or U6705 (N_6705,N_6420,N_6277);
xnor U6706 (N_6706,N_6320,N_6447);
nor U6707 (N_6707,N_6423,N_6372);
xnor U6708 (N_6708,N_6445,N_6425);
and U6709 (N_6709,N_6330,N_6322);
nand U6710 (N_6710,N_6361,N_6480);
nor U6711 (N_6711,N_6303,N_6461);
nor U6712 (N_6712,N_6435,N_6278);
nand U6713 (N_6713,N_6337,N_6397);
or U6714 (N_6714,N_6334,N_6357);
xnor U6715 (N_6715,N_6477,N_6439);
or U6716 (N_6716,N_6492,N_6332);
and U6717 (N_6717,N_6456,N_6250);
nand U6718 (N_6718,N_6456,N_6482);
nor U6719 (N_6719,N_6253,N_6359);
and U6720 (N_6720,N_6259,N_6346);
nand U6721 (N_6721,N_6413,N_6312);
xor U6722 (N_6722,N_6460,N_6311);
and U6723 (N_6723,N_6395,N_6256);
xnor U6724 (N_6724,N_6454,N_6414);
nor U6725 (N_6725,N_6384,N_6287);
and U6726 (N_6726,N_6254,N_6378);
xor U6727 (N_6727,N_6349,N_6369);
nor U6728 (N_6728,N_6281,N_6317);
or U6729 (N_6729,N_6269,N_6354);
nand U6730 (N_6730,N_6289,N_6315);
nand U6731 (N_6731,N_6337,N_6398);
or U6732 (N_6732,N_6328,N_6432);
nand U6733 (N_6733,N_6251,N_6299);
nand U6734 (N_6734,N_6486,N_6333);
or U6735 (N_6735,N_6396,N_6355);
nor U6736 (N_6736,N_6391,N_6410);
xnor U6737 (N_6737,N_6388,N_6262);
nand U6738 (N_6738,N_6430,N_6472);
nor U6739 (N_6739,N_6404,N_6453);
or U6740 (N_6740,N_6373,N_6265);
xnor U6741 (N_6741,N_6408,N_6312);
or U6742 (N_6742,N_6459,N_6326);
nor U6743 (N_6743,N_6358,N_6410);
xnor U6744 (N_6744,N_6417,N_6358);
xnor U6745 (N_6745,N_6342,N_6470);
nand U6746 (N_6746,N_6361,N_6274);
nor U6747 (N_6747,N_6277,N_6464);
or U6748 (N_6748,N_6314,N_6373);
nand U6749 (N_6749,N_6323,N_6293);
nand U6750 (N_6750,N_6518,N_6535);
xnor U6751 (N_6751,N_6714,N_6511);
xnor U6752 (N_6752,N_6633,N_6603);
and U6753 (N_6753,N_6508,N_6559);
nand U6754 (N_6754,N_6607,N_6719);
or U6755 (N_6755,N_6534,N_6734);
and U6756 (N_6756,N_6568,N_6722);
nor U6757 (N_6757,N_6537,N_6606);
xor U6758 (N_6758,N_6563,N_6707);
xor U6759 (N_6759,N_6590,N_6666);
or U6760 (N_6760,N_6713,N_6687);
xor U6761 (N_6761,N_6558,N_6622);
or U6762 (N_6762,N_6639,N_6708);
or U6763 (N_6763,N_6548,N_6598);
xor U6764 (N_6764,N_6663,N_6723);
nand U6765 (N_6765,N_6740,N_6531);
nor U6766 (N_6766,N_6655,N_6553);
xnor U6767 (N_6767,N_6576,N_6582);
nand U6768 (N_6768,N_6571,N_6503);
nor U6769 (N_6769,N_6521,N_6502);
and U6770 (N_6770,N_6745,N_6549);
xnor U6771 (N_6771,N_6680,N_6579);
or U6772 (N_6772,N_6523,N_6599);
or U6773 (N_6773,N_6570,N_6584);
nand U6774 (N_6774,N_6660,N_6676);
or U6775 (N_6775,N_6540,N_6684);
or U6776 (N_6776,N_6519,N_6536);
xor U6777 (N_6777,N_6645,N_6657);
nand U6778 (N_6778,N_6569,N_6730);
and U6779 (N_6779,N_6644,N_6669);
nand U6780 (N_6780,N_6642,N_6573);
nand U6781 (N_6781,N_6661,N_6529);
or U6782 (N_6782,N_6544,N_6501);
and U6783 (N_6783,N_6715,N_6585);
or U6784 (N_6784,N_6630,N_6705);
xor U6785 (N_6785,N_6512,N_6637);
nor U6786 (N_6786,N_6577,N_6741);
and U6787 (N_6787,N_6706,N_6641);
or U6788 (N_6788,N_6728,N_6675);
or U6789 (N_6789,N_6618,N_6547);
xor U6790 (N_6790,N_6651,N_6506);
xnor U6791 (N_6791,N_6703,N_6698);
nand U6792 (N_6792,N_6556,N_6593);
and U6793 (N_6793,N_6673,N_6597);
and U6794 (N_6794,N_6737,N_6688);
nor U6795 (N_6795,N_6566,N_6628);
and U6796 (N_6796,N_6574,N_6662);
xor U6797 (N_6797,N_6646,N_6691);
nor U6798 (N_6798,N_6643,N_6612);
nor U6799 (N_6799,N_6500,N_6635);
nand U6800 (N_6800,N_6677,N_6561);
nand U6801 (N_6801,N_6654,N_6700);
nor U6802 (N_6802,N_6681,N_6736);
or U6803 (N_6803,N_6743,N_6526);
or U6804 (N_6804,N_6514,N_6564);
and U6805 (N_6805,N_6659,N_6664);
and U6806 (N_6806,N_6626,N_6504);
nand U6807 (N_6807,N_6554,N_6527);
and U6808 (N_6808,N_6693,N_6739);
and U6809 (N_6809,N_6742,N_6710);
and U6810 (N_6810,N_6682,N_6636);
or U6811 (N_6811,N_6711,N_6701);
and U6812 (N_6812,N_6516,N_6727);
nor U6813 (N_6813,N_6510,N_6704);
xnor U6814 (N_6814,N_6671,N_6505);
nor U6815 (N_6815,N_6557,N_6726);
and U6816 (N_6816,N_6692,N_6620);
or U6817 (N_6817,N_6670,N_6609);
or U6818 (N_6818,N_6539,N_6513);
xnor U6819 (N_6819,N_6572,N_6621);
nor U6820 (N_6820,N_6749,N_6578);
or U6821 (N_6821,N_6591,N_6594);
nor U6822 (N_6822,N_6595,N_6614);
nor U6823 (N_6823,N_6545,N_6507);
xor U6824 (N_6824,N_6672,N_6530);
or U6825 (N_6825,N_6602,N_6533);
or U6826 (N_6826,N_6588,N_6515);
or U6827 (N_6827,N_6592,N_6709);
nand U6828 (N_6828,N_6640,N_6697);
and U6829 (N_6829,N_6565,N_6532);
nor U6830 (N_6830,N_6702,N_6520);
xor U6831 (N_6831,N_6611,N_6509);
xnor U6832 (N_6832,N_6648,N_6668);
nand U6833 (N_6833,N_6667,N_6616);
xnor U6834 (N_6834,N_6522,N_6586);
xor U6835 (N_6835,N_6623,N_6689);
or U6836 (N_6836,N_6721,N_6580);
or U6837 (N_6837,N_6731,N_6674);
and U6838 (N_6838,N_6625,N_6542);
nand U6839 (N_6839,N_6634,N_6617);
and U6840 (N_6840,N_6696,N_6744);
and U6841 (N_6841,N_6613,N_6624);
nor U6842 (N_6842,N_6658,N_6665);
and U6843 (N_6843,N_6543,N_6524);
nand U6844 (N_6844,N_6699,N_6647);
nor U6845 (N_6845,N_6567,N_6608);
nand U6846 (N_6846,N_6656,N_6733);
xor U6847 (N_6847,N_6695,N_6528);
and U6848 (N_6848,N_6629,N_6725);
nand U6849 (N_6849,N_6729,N_6627);
nor U6850 (N_6850,N_6638,N_6583);
and U6851 (N_6851,N_6690,N_6738);
nand U6852 (N_6852,N_6604,N_6678);
xnor U6853 (N_6853,N_6685,N_6746);
nor U6854 (N_6854,N_6748,N_6747);
nor U6855 (N_6855,N_6525,N_6716);
and U6856 (N_6856,N_6652,N_6610);
or U6857 (N_6857,N_6615,N_6650);
nor U6858 (N_6858,N_6517,N_6619);
or U6859 (N_6859,N_6601,N_6605);
and U6860 (N_6860,N_6589,N_6649);
xor U6861 (N_6861,N_6560,N_6653);
xor U6862 (N_6862,N_6631,N_6551);
and U6863 (N_6863,N_6575,N_6550);
nor U6864 (N_6864,N_6724,N_6683);
xnor U6865 (N_6865,N_6732,N_6720);
or U6866 (N_6866,N_6679,N_6587);
nor U6867 (N_6867,N_6686,N_6562);
nand U6868 (N_6868,N_6718,N_6552);
xnor U6869 (N_6869,N_6555,N_6581);
xnor U6870 (N_6870,N_6541,N_6694);
nand U6871 (N_6871,N_6712,N_6735);
and U6872 (N_6872,N_6596,N_6600);
nand U6873 (N_6873,N_6632,N_6538);
and U6874 (N_6874,N_6717,N_6546);
and U6875 (N_6875,N_6540,N_6721);
xnor U6876 (N_6876,N_6609,N_6710);
and U6877 (N_6877,N_6550,N_6652);
and U6878 (N_6878,N_6728,N_6673);
nor U6879 (N_6879,N_6715,N_6654);
and U6880 (N_6880,N_6625,N_6577);
xnor U6881 (N_6881,N_6660,N_6524);
nor U6882 (N_6882,N_6670,N_6714);
xnor U6883 (N_6883,N_6592,N_6703);
and U6884 (N_6884,N_6633,N_6694);
or U6885 (N_6885,N_6593,N_6575);
or U6886 (N_6886,N_6592,N_6690);
and U6887 (N_6887,N_6663,N_6695);
xor U6888 (N_6888,N_6561,N_6579);
and U6889 (N_6889,N_6562,N_6704);
nand U6890 (N_6890,N_6694,N_6580);
and U6891 (N_6891,N_6593,N_6599);
and U6892 (N_6892,N_6638,N_6737);
xnor U6893 (N_6893,N_6538,N_6595);
and U6894 (N_6894,N_6723,N_6646);
nand U6895 (N_6895,N_6605,N_6671);
xor U6896 (N_6896,N_6732,N_6607);
or U6897 (N_6897,N_6568,N_6645);
xor U6898 (N_6898,N_6715,N_6684);
nand U6899 (N_6899,N_6564,N_6607);
nor U6900 (N_6900,N_6632,N_6550);
xnor U6901 (N_6901,N_6635,N_6533);
xnor U6902 (N_6902,N_6542,N_6690);
nor U6903 (N_6903,N_6577,N_6678);
xnor U6904 (N_6904,N_6575,N_6609);
nand U6905 (N_6905,N_6703,N_6542);
or U6906 (N_6906,N_6634,N_6613);
xnor U6907 (N_6907,N_6571,N_6708);
and U6908 (N_6908,N_6608,N_6553);
or U6909 (N_6909,N_6583,N_6516);
nand U6910 (N_6910,N_6570,N_6637);
and U6911 (N_6911,N_6505,N_6577);
and U6912 (N_6912,N_6656,N_6540);
nor U6913 (N_6913,N_6509,N_6599);
nor U6914 (N_6914,N_6634,N_6567);
and U6915 (N_6915,N_6544,N_6588);
and U6916 (N_6916,N_6744,N_6603);
or U6917 (N_6917,N_6675,N_6737);
and U6918 (N_6918,N_6529,N_6516);
nor U6919 (N_6919,N_6687,N_6609);
nand U6920 (N_6920,N_6703,N_6602);
xnor U6921 (N_6921,N_6521,N_6654);
nor U6922 (N_6922,N_6659,N_6541);
nand U6923 (N_6923,N_6520,N_6581);
nand U6924 (N_6924,N_6646,N_6641);
nor U6925 (N_6925,N_6506,N_6566);
and U6926 (N_6926,N_6633,N_6636);
nand U6927 (N_6927,N_6695,N_6540);
or U6928 (N_6928,N_6663,N_6510);
nand U6929 (N_6929,N_6612,N_6500);
and U6930 (N_6930,N_6507,N_6586);
and U6931 (N_6931,N_6517,N_6562);
or U6932 (N_6932,N_6637,N_6539);
nand U6933 (N_6933,N_6538,N_6582);
nand U6934 (N_6934,N_6623,N_6710);
nor U6935 (N_6935,N_6527,N_6639);
nor U6936 (N_6936,N_6651,N_6556);
nor U6937 (N_6937,N_6520,N_6555);
nand U6938 (N_6938,N_6530,N_6677);
or U6939 (N_6939,N_6744,N_6654);
or U6940 (N_6940,N_6584,N_6523);
nand U6941 (N_6941,N_6735,N_6682);
and U6942 (N_6942,N_6603,N_6505);
or U6943 (N_6943,N_6620,N_6593);
xor U6944 (N_6944,N_6627,N_6686);
nor U6945 (N_6945,N_6684,N_6588);
xor U6946 (N_6946,N_6591,N_6711);
nor U6947 (N_6947,N_6535,N_6585);
nand U6948 (N_6948,N_6549,N_6570);
nor U6949 (N_6949,N_6696,N_6652);
and U6950 (N_6950,N_6505,N_6742);
nand U6951 (N_6951,N_6694,N_6511);
or U6952 (N_6952,N_6638,N_6710);
or U6953 (N_6953,N_6725,N_6568);
nor U6954 (N_6954,N_6598,N_6549);
or U6955 (N_6955,N_6593,N_6699);
and U6956 (N_6956,N_6633,N_6700);
nand U6957 (N_6957,N_6548,N_6661);
nor U6958 (N_6958,N_6671,N_6585);
xnor U6959 (N_6959,N_6556,N_6618);
or U6960 (N_6960,N_6664,N_6522);
nand U6961 (N_6961,N_6717,N_6597);
or U6962 (N_6962,N_6747,N_6570);
or U6963 (N_6963,N_6698,N_6536);
nand U6964 (N_6964,N_6643,N_6737);
xnor U6965 (N_6965,N_6732,N_6599);
xor U6966 (N_6966,N_6540,N_6700);
and U6967 (N_6967,N_6551,N_6716);
or U6968 (N_6968,N_6702,N_6735);
nand U6969 (N_6969,N_6657,N_6731);
nor U6970 (N_6970,N_6508,N_6717);
nor U6971 (N_6971,N_6641,N_6501);
or U6972 (N_6972,N_6570,N_6650);
and U6973 (N_6973,N_6734,N_6610);
and U6974 (N_6974,N_6503,N_6520);
or U6975 (N_6975,N_6623,N_6673);
nor U6976 (N_6976,N_6663,N_6710);
and U6977 (N_6977,N_6698,N_6576);
nor U6978 (N_6978,N_6581,N_6662);
nor U6979 (N_6979,N_6535,N_6524);
nand U6980 (N_6980,N_6505,N_6653);
or U6981 (N_6981,N_6652,N_6744);
or U6982 (N_6982,N_6529,N_6655);
and U6983 (N_6983,N_6609,N_6734);
nand U6984 (N_6984,N_6696,N_6571);
and U6985 (N_6985,N_6559,N_6552);
xnor U6986 (N_6986,N_6692,N_6635);
or U6987 (N_6987,N_6692,N_6723);
xnor U6988 (N_6988,N_6702,N_6747);
xnor U6989 (N_6989,N_6570,N_6689);
or U6990 (N_6990,N_6585,N_6621);
and U6991 (N_6991,N_6553,N_6582);
xor U6992 (N_6992,N_6504,N_6642);
nand U6993 (N_6993,N_6556,N_6573);
or U6994 (N_6994,N_6623,N_6741);
and U6995 (N_6995,N_6524,N_6743);
and U6996 (N_6996,N_6702,N_6586);
nor U6997 (N_6997,N_6575,N_6673);
and U6998 (N_6998,N_6501,N_6592);
nor U6999 (N_6999,N_6733,N_6696);
nor U7000 (N_7000,N_6885,N_6882);
or U7001 (N_7001,N_6946,N_6891);
xnor U7002 (N_7002,N_6792,N_6789);
xnor U7003 (N_7003,N_6832,N_6790);
and U7004 (N_7004,N_6788,N_6984);
nand U7005 (N_7005,N_6861,N_6835);
nor U7006 (N_7006,N_6991,N_6897);
xor U7007 (N_7007,N_6869,N_6932);
and U7008 (N_7008,N_6921,N_6973);
nand U7009 (N_7009,N_6983,N_6848);
and U7010 (N_7010,N_6878,N_6987);
nor U7011 (N_7011,N_6990,N_6913);
nand U7012 (N_7012,N_6845,N_6962);
and U7013 (N_7013,N_6884,N_6802);
and U7014 (N_7014,N_6778,N_6819);
nand U7015 (N_7015,N_6931,N_6756);
and U7016 (N_7016,N_6957,N_6886);
or U7017 (N_7017,N_6902,N_6982);
nor U7018 (N_7018,N_6895,N_6814);
nor U7019 (N_7019,N_6879,N_6944);
and U7020 (N_7020,N_6883,N_6951);
or U7021 (N_7021,N_6852,N_6785);
and U7022 (N_7022,N_6784,N_6866);
and U7023 (N_7023,N_6933,N_6764);
nand U7024 (N_7024,N_6971,N_6812);
and U7025 (N_7025,N_6782,N_6820);
nor U7026 (N_7026,N_6755,N_6928);
nor U7027 (N_7027,N_6965,N_6894);
or U7028 (N_7028,N_6841,N_6837);
xnor U7029 (N_7029,N_6994,N_6849);
nor U7030 (N_7030,N_6808,N_6753);
nand U7031 (N_7031,N_6876,N_6858);
or U7032 (N_7032,N_6949,N_6801);
nand U7033 (N_7033,N_6769,N_6762);
or U7034 (N_7034,N_6956,N_6900);
or U7035 (N_7035,N_6935,N_6803);
nor U7036 (N_7036,N_6945,N_6823);
nand U7037 (N_7037,N_6775,N_6793);
xor U7038 (N_7038,N_6818,N_6972);
nor U7039 (N_7039,N_6875,N_6824);
nand U7040 (N_7040,N_6822,N_6761);
and U7041 (N_7041,N_6865,N_6815);
nand U7042 (N_7042,N_6988,N_6846);
nor U7043 (N_7043,N_6927,N_6859);
xor U7044 (N_7044,N_6805,N_6963);
nor U7045 (N_7045,N_6766,N_6840);
nand U7046 (N_7046,N_6947,N_6877);
or U7047 (N_7047,N_6918,N_6839);
nand U7048 (N_7048,N_6804,N_6938);
nor U7049 (N_7049,N_6958,N_6850);
nor U7050 (N_7050,N_6833,N_6758);
and U7051 (N_7051,N_6888,N_6893);
nor U7052 (N_7052,N_6796,N_6989);
or U7053 (N_7053,N_6903,N_6843);
xor U7054 (N_7054,N_6996,N_6862);
nor U7055 (N_7055,N_6797,N_6867);
nor U7056 (N_7056,N_6809,N_6922);
and U7057 (N_7057,N_6826,N_6967);
or U7058 (N_7058,N_6774,N_6970);
xnor U7059 (N_7059,N_6977,N_6794);
xor U7060 (N_7060,N_6889,N_6836);
xnor U7061 (N_7061,N_6979,N_6847);
xor U7062 (N_7062,N_6941,N_6993);
and U7063 (N_7063,N_6914,N_6874);
nand U7064 (N_7064,N_6871,N_6856);
nor U7065 (N_7065,N_6919,N_6810);
nand U7066 (N_7066,N_6910,N_6887);
xor U7067 (N_7067,N_6817,N_6939);
xor U7068 (N_7068,N_6806,N_6770);
or U7069 (N_7069,N_6923,N_6924);
nand U7070 (N_7070,N_6901,N_6828);
or U7071 (N_7071,N_6767,N_6930);
xnor U7072 (N_7072,N_6853,N_6995);
nor U7073 (N_7073,N_6976,N_6777);
and U7074 (N_7074,N_6783,N_6953);
nor U7075 (N_7075,N_6969,N_6892);
or U7076 (N_7076,N_6773,N_6798);
nand U7077 (N_7077,N_6915,N_6752);
nor U7078 (N_7078,N_6934,N_6807);
or U7079 (N_7079,N_6959,N_6964);
xnor U7080 (N_7080,N_6760,N_6978);
nor U7081 (N_7081,N_6940,N_6872);
xor U7082 (N_7082,N_6912,N_6907);
xor U7083 (N_7083,N_6998,N_6920);
and U7084 (N_7084,N_6911,N_6825);
nor U7085 (N_7085,N_6816,N_6800);
and U7086 (N_7086,N_6992,N_6829);
and U7087 (N_7087,N_6870,N_6986);
nand U7088 (N_7088,N_6779,N_6855);
or U7089 (N_7089,N_6772,N_6961);
nor U7090 (N_7090,N_6942,N_6966);
nand U7091 (N_7091,N_6950,N_6880);
nor U7092 (N_7092,N_6868,N_6881);
and U7093 (N_7093,N_6759,N_6751);
nor U7094 (N_7094,N_6771,N_6838);
and U7095 (N_7095,N_6926,N_6864);
xnor U7096 (N_7096,N_6763,N_6765);
xnor U7097 (N_7097,N_6795,N_6860);
xor U7098 (N_7098,N_6821,N_6842);
nand U7099 (N_7099,N_6943,N_6898);
xnor U7100 (N_7100,N_6811,N_6936);
or U7101 (N_7101,N_6960,N_6948);
nand U7102 (N_7102,N_6916,N_6905);
xor U7103 (N_7103,N_6974,N_6981);
xnor U7104 (N_7104,N_6997,N_6937);
xnor U7105 (N_7105,N_6851,N_6791);
and U7106 (N_7106,N_6863,N_6929);
or U7107 (N_7107,N_6830,N_6909);
nor U7108 (N_7108,N_6857,N_6768);
or U7109 (N_7109,N_6954,N_6754);
and U7110 (N_7110,N_6985,N_6757);
nor U7111 (N_7111,N_6904,N_6813);
xor U7112 (N_7112,N_6799,N_6750);
nor U7113 (N_7113,N_6827,N_6831);
nand U7114 (N_7114,N_6786,N_6908);
nand U7115 (N_7115,N_6873,N_6980);
or U7116 (N_7116,N_6854,N_6896);
and U7117 (N_7117,N_6780,N_6844);
xnor U7118 (N_7118,N_6925,N_6899);
nand U7119 (N_7119,N_6975,N_6834);
or U7120 (N_7120,N_6781,N_6999);
nor U7121 (N_7121,N_6787,N_6906);
and U7122 (N_7122,N_6955,N_6968);
xnor U7123 (N_7123,N_6952,N_6776);
and U7124 (N_7124,N_6890,N_6917);
or U7125 (N_7125,N_6995,N_6864);
nor U7126 (N_7126,N_6982,N_6976);
or U7127 (N_7127,N_6855,N_6987);
nand U7128 (N_7128,N_6858,N_6994);
xor U7129 (N_7129,N_6953,N_6917);
and U7130 (N_7130,N_6877,N_6909);
nor U7131 (N_7131,N_6759,N_6913);
nor U7132 (N_7132,N_6986,N_6820);
or U7133 (N_7133,N_6906,N_6752);
nand U7134 (N_7134,N_6931,N_6868);
or U7135 (N_7135,N_6951,N_6966);
or U7136 (N_7136,N_6971,N_6965);
xor U7137 (N_7137,N_6941,N_6871);
and U7138 (N_7138,N_6826,N_6936);
nor U7139 (N_7139,N_6961,N_6934);
xor U7140 (N_7140,N_6855,N_6893);
xor U7141 (N_7141,N_6774,N_6858);
nand U7142 (N_7142,N_6773,N_6776);
or U7143 (N_7143,N_6761,N_6875);
and U7144 (N_7144,N_6761,N_6879);
nand U7145 (N_7145,N_6855,N_6950);
or U7146 (N_7146,N_6776,N_6806);
or U7147 (N_7147,N_6835,N_6832);
and U7148 (N_7148,N_6819,N_6927);
and U7149 (N_7149,N_6974,N_6792);
or U7150 (N_7150,N_6893,N_6976);
and U7151 (N_7151,N_6773,N_6861);
or U7152 (N_7152,N_6993,N_6905);
and U7153 (N_7153,N_6876,N_6965);
xor U7154 (N_7154,N_6962,N_6815);
and U7155 (N_7155,N_6829,N_6846);
nand U7156 (N_7156,N_6851,N_6973);
nor U7157 (N_7157,N_6918,N_6848);
xnor U7158 (N_7158,N_6789,N_6964);
nor U7159 (N_7159,N_6950,N_6944);
nor U7160 (N_7160,N_6991,N_6778);
nand U7161 (N_7161,N_6835,N_6854);
xor U7162 (N_7162,N_6906,N_6769);
or U7163 (N_7163,N_6779,N_6885);
nor U7164 (N_7164,N_6805,N_6862);
and U7165 (N_7165,N_6805,N_6941);
or U7166 (N_7166,N_6786,N_6833);
xor U7167 (N_7167,N_6855,N_6877);
nor U7168 (N_7168,N_6909,N_6851);
or U7169 (N_7169,N_6954,N_6784);
nand U7170 (N_7170,N_6945,N_6757);
nand U7171 (N_7171,N_6857,N_6790);
and U7172 (N_7172,N_6938,N_6771);
nand U7173 (N_7173,N_6942,N_6880);
nand U7174 (N_7174,N_6809,N_6781);
xor U7175 (N_7175,N_6775,N_6921);
and U7176 (N_7176,N_6928,N_6906);
nor U7177 (N_7177,N_6820,N_6902);
nor U7178 (N_7178,N_6771,N_6996);
xor U7179 (N_7179,N_6791,N_6823);
xnor U7180 (N_7180,N_6966,N_6962);
or U7181 (N_7181,N_6770,N_6852);
or U7182 (N_7182,N_6854,N_6768);
nor U7183 (N_7183,N_6866,N_6966);
nand U7184 (N_7184,N_6988,N_6773);
xnor U7185 (N_7185,N_6827,N_6935);
xor U7186 (N_7186,N_6787,N_6962);
nand U7187 (N_7187,N_6965,N_6990);
nor U7188 (N_7188,N_6784,N_6802);
and U7189 (N_7189,N_6976,N_6887);
and U7190 (N_7190,N_6889,N_6901);
nand U7191 (N_7191,N_6795,N_6947);
and U7192 (N_7192,N_6790,N_6824);
nor U7193 (N_7193,N_6886,N_6823);
nor U7194 (N_7194,N_6893,N_6842);
and U7195 (N_7195,N_6873,N_6957);
and U7196 (N_7196,N_6987,N_6982);
and U7197 (N_7197,N_6883,N_6835);
and U7198 (N_7198,N_6972,N_6999);
xor U7199 (N_7199,N_6941,N_6987);
or U7200 (N_7200,N_6898,N_6779);
nor U7201 (N_7201,N_6908,N_6883);
and U7202 (N_7202,N_6889,N_6981);
and U7203 (N_7203,N_6982,N_6895);
or U7204 (N_7204,N_6768,N_6885);
nand U7205 (N_7205,N_6777,N_6806);
nand U7206 (N_7206,N_6756,N_6840);
and U7207 (N_7207,N_6824,N_6972);
or U7208 (N_7208,N_6771,N_6860);
or U7209 (N_7209,N_6812,N_6942);
and U7210 (N_7210,N_6968,N_6801);
or U7211 (N_7211,N_6830,N_6844);
xnor U7212 (N_7212,N_6853,N_6810);
nor U7213 (N_7213,N_6999,N_6834);
nor U7214 (N_7214,N_6910,N_6779);
xor U7215 (N_7215,N_6753,N_6834);
or U7216 (N_7216,N_6775,N_6836);
nor U7217 (N_7217,N_6916,N_6949);
nor U7218 (N_7218,N_6805,N_6884);
or U7219 (N_7219,N_6962,N_6821);
or U7220 (N_7220,N_6948,N_6834);
or U7221 (N_7221,N_6865,N_6930);
xnor U7222 (N_7222,N_6835,N_6947);
or U7223 (N_7223,N_6986,N_6943);
nand U7224 (N_7224,N_6776,N_6834);
xnor U7225 (N_7225,N_6764,N_6918);
nand U7226 (N_7226,N_6985,N_6927);
xor U7227 (N_7227,N_6979,N_6794);
and U7228 (N_7228,N_6913,N_6963);
nor U7229 (N_7229,N_6936,N_6759);
xor U7230 (N_7230,N_6796,N_6905);
nand U7231 (N_7231,N_6797,N_6832);
nand U7232 (N_7232,N_6980,N_6755);
nor U7233 (N_7233,N_6782,N_6830);
xor U7234 (N_7234,N_6773,N_6843);
or U7235 (N_7235,N_6990,N_6854);
nor U7236 (N_7236,N_6762,N_6869);
or U7237 (N_7237,N_6956,N_6940);
nor U7238 (N_7238,N_6970,N_6849);
and U7239 (N_7239,N_6846,N_6850);
xor U7240 (N_7240,N_6977,N_6789);
nor U7241 (N_7241,N_6829,N_6825);
xor U7242 (N_7242,N_6883,N_6757);
nand U7243 (N_7243,N_6856,N_6874);
xnor U7244 (N_7244,N_6769,N_6910);
or U7245 (N_7245,N_6805,N_6791);
nor U7246 (N_7246,N_6857,N_6893);
xnor U7247 (N_7247,N_6938,N_6912);
xnor U7248 (N_7248,N_6821,N_6808);
or U7249 (N_7249,N_6758,N_6917);
and U7250 (N_7250,N_7047,N_7152);
xor U7251 (N_7251,N_7124,N_7054);
xor U7252 (N_7252,N_7131,N_7053);
nand U7253 (N_7253,N_7127,N_7189);
nand U7254 (N_7254,N_7090,N_7030);
nor U7255 (N_7255,N_7082,N_7093);
or U7256 (N_7256,N_7242,N_7027);
nand U7257 (N_7257,N_7138,N_7241);
xnor U7258 (N_7258,N_7011,N_7033);
or U7259 (N_7259,N_7227,N_7007);
and U7260 (N_7260,N_7078,N_7118);
or U7261 (N_7261,N_7052,N_7029);
and U7262 (N_7262,N_7101,N_7248);
xnor U7263 (N_7263,N_7038,N_7154);
nand U7264 (N_7264,N_7020,N_7133);
nand U7265 (N_7265,N_7235,N_7068);
nor U7266 (N_7266,N_7085,N_7086);
and U7267 (N_7267,N_7119,N_7141);
and U7268 (N_7268,N_7039,N_7192);
or U7269 (N_7269,N_7217,N_7087);
xnor U7270 (N_7270,N_7043,N_7112);
xor U7271 (N_7271,N_7204,N_7057);
nor U7272 (N_7272,N_7048,N_7153);
xor U7273 (N_7273,N_7002,N_7171);
nand U7274 (N_7274,N_7003,N_7247);
nand U7275 (N_7275,N_7240,N_7223);
nand U7276 (N_7276,N_7182,N_7088);
or U7277 (N_7277,N_7063,N_7005);
or U7278 (N_7278,N_7009,N_7099);
nor U7279 (N_7279,N_7215,N_7169);
and U7280 (N_7280,N_7246,N_7165);
nand U7281 (N_7281,N_7208,N_7113);
nand U7282 (N_7282,N_7091,N_7032);
nand U7283 (N_7283,N_7128,N_7092);
or U7284 (N_7284,N_7156,N_7239);
nand U7285 (N_7285,N_7103,N_7185);
xnor U7286 (N_7286,N_7183,N_7230);
and U7287 (N_7287,N_7200,N_7193);
nor U7288 (N_7288,N_7015,N_7197);
nor U7289 (N_7289,N_7137,N_7140);
nand U7290 (N_7290,N_7037,N_7058);
or U7291 (N_7291,N_7213,N_7019);
nand U7292 (N_7292,N_7237,N_7205);
nand U7293 (N_7293,N_7238,N_7022);
nand U7294 (N_7294,N_7123,N_7014);
nor U7295 (N_7295,N_7172,N_7198);
or U7296 (N_7296,N_7122,N_7083);
nor U7297 (N_7297,N_7195,N_7041);
or U7298 (N_7298,N_7219,N_7233);
and U7299 (N_7299,N_7164,N_7143);
nand U7300 (N_7300,N_7186,N_7142);
nand U7301 (N_7301,N_7162,N_7207);
and U7302 (N_7302,N_7146,N_7206);
xor U7303 (N_7303,N_7034,N_7025);
and U7304 (N_7304,N_7049,N_7046);
nor U7305 (N_7305,N_7071,N_7216);
xnor U7306 (N_7306,N_7144,N_7024);
or U7307 (N_7307,N_7076,N_7159);
nand U7308 (N_7308,N_7060,N_7023);
or U7309 (N_7309,N_7132,N_7218);
or U7310 (N_7310,N_7098,N_7021);
or U7311 (N_7311,N_7097,N_7036);
nand U7312 (N_7312,N_7061,N_7191);
xnor U7313 (N_7313,N_7167,N_7194);
or U7314 (N_7314,N_7106,N_7069);
nor U7315 (N_7315,N_7120,N_7070);
and U7316 (N_7316,N_7175,N_7190);
nor U7317 (N_7317,N_7042,N_7160);
and U7318 (N_7318,N_7028,N_7055);
nand U7319 (N_7319,N_7109,N_7136);
or U7320 (N_7320,N_7077,N_7229);
nand U7321 (N_7321,N_7126,N_7107);
nor U7322 (N_7322,N_7170,N_7040);
and U7323 (N_7323,N_7199,N_7050);
nand U7324 (N_7324,N_7187,N_7010);
and U7325 (N_7325,N_7125,N_7111);
xnor U7326 (N_7326,N_7100,N_7114);
and U7327 (N_7327,N_7031,N_7157);
nand U7328 (N_7328,N_7177,N_7224);
nand U7329 (N_7329,N_7081,N_7004);
xnor U7330 (N_7330,N_7129,N_7145);
and U7331 (N_7331,N_7176,N_7108);
nand U7332 (N_7332,N_7209,N_7075);
and U7333 (N_7333,N_7163,N_7135);
nor U7334 (N_7334,N_7151,N_7155);
or U7335 (N_7335,N_7196,N_7105);
nor U7336 (N_7336,N_7096,N_7116);
xor U7337 (N_7337,N_7202,N_7212);
and U7338 (N_7338,N_7188,N_7161);
or U7339 (N_7339,N_7073,N_7067);
or U7340 (N_7340,N_7228,N_7117);
nand U7341 (N_7341,N_7220,N_7211);
xnor U7342 (N_7342,N_7089,N_7221);
nor U7343 (N_7343,N_7035,N_7179);
xnor U7344 (N_7344,N_7173,N_7222);
and U7345 (N_7345,N_7018,N_7184);
xor U7346 (N_7346,N_7074,N_7168);
nor U7347 (N_7347,N_7079,N_7017);
and U7348 (N_7348,N_7044,N_7006);
nand U7349 (N_7349,N_7016,N_7121);
nand U7350 (N_7350,N_7178,N_7226);
nor U7351 (N_7351,N_7059,N_7214);
nand U7352 (N_7352,N_7115,N_7243);
xor U7353 (N_7353,N_7001,N_7064);
nand U7354 (N_7354,N_7062,N_7150);
and U7355 (N_7355,N_7056,N_7210);
nor U7356 (N_7356,N_7072,N_7139);
nor U7357 (N_7357,N_7249,N_7134);
nand U7358 (N_7358,N_7166,N_7244);
and U7359 (N_7359,N_7065,N_7094);
nand U7360 (N_7360,N_7013,N_7201);
or U7361 (N_7361,N_7203,N_7012);
and U7362 (N_7362,N_7095,N_7234);
nand U7363 (N_7363,N_7000,N_7236);
nor U7364 (N_7364,N_7008,N_7066);
nor U7365 (N_7365,N_7051,N_7225);
xor U7366 (N_7366,N_7110,N_7232);
nand U7367 (N_7367,N_7102,N_7180);
or U7368 (N_7368,N_7245,N_7181);
and U7369 (N_7369,N_7149,N_7080);
and U7370 (N_7370,N_7147,N_7174);
or U7371 (N_7371,N_7158,N_7084);
nand U7372 (N_7372,N_7130,N_7104);
nand U7373 (N_7373,N_7148,N_7045);
and U7374 (N_7374,N_7231,N_7026);
and U7375 (N_7375,N_7121,N_7018);
nand U7376 (N_7376,N_7123,N_7241);
nand U7377 (N_7377,N_7107,N_7097);
or U7378 (N_7378,N_7046,N_7230);
and U7379 (N_7379,N_7134,N_7055);
and U7380 (N_7380,N_7147,N_7066);
or U7381 (N_7381,N_7003,N_7021);
xor U7382 (N_7382,N_7188,N_7081);
xnor U7383 (N_7383,N_7026,N_7006);
nor U7384 (N_7384,N_7119,N_7005);
or U7385 (N_7385,N_7124,N_7065);
or U7386 (N_7386,N_7099,N_7027);
nand U7387 (N_7387,N_7140,N_7187);
and U7388 (N_7388,N_7099,N_7134);
xnor U7389 (N_7389,N_7208,N_7106);
xor U7390 (N_7390,N_7235,N_7155);
and U7391 (N_7391,N_7078,N_7184);
nor U7392 (N_7392,N_7121,N_7087);
and U7393 (N_7393,N_7188,N_7127);
and U7394 (N_7394,N_7227,N_7186);
xnor U7395 (N_7395,N_7165,N_7128);
or U7396 (N_7396,N_7051,N_7119);
xnor U7397 (N_7397,N_7003,N_7176);
nor U7398 (N_7398,N_7029,N_7132);
nand U7399 (N_7399,N_7218,N_7117);
nand U7400 (N_7400,N_7162,N_7027);
or U7401 (N_7401,N_7227,N_7235);
or U7402 (N_7402,N_7135,N_7016);
nor U7403 (N_7403,N_7184,N_7216);
or U7404 (N_7404,N_7117,N_7048);
xnor U7405 (N_7405,N_7132,N_7142);
or U7406 (N_7406,N_7246,N_7220);
or U7407 (N_7407,N_7221,N_7108);
nor U7408 (N_7408,N_7213,N_7205);
nor U7409 (N_7409,N_7223,N_7206);
or U7410 (N_7410,N_7174,N_7203);
or U7411 (N_7411,N_7140,N_7018);
or U7412 (N_7412,N_7120,N_7027);
nand U7413 (N_7413,N_7133,N_7145);
nand U7414 (N_7414,N_7125,N_7171);
and U7415 (N_7415,N_7104,N_7239);
or U7416 (N_7416,N_7208,N_7225);
nor U7417 (N_7417,N_7119,N_7165);
or U7418 (N_7418,N_7040,N_7065);
or U7419 (N_7419,N_7112,N_7178);
or U7420 (N_7420,N_7184,N_7208);
or U7421 (N_7421,N_7188,N_7141);
nand U7422 (N_7422,N_7167,N_7214);
or U7423 (N_7423,N_7230,N_7216);
or U7424 (N_7424,N_7196,N_7052);
xor U7425 (N_7425,N_7210,N_7138);
and U7426 (N_7426,N_7214,N_7130);
xnor U7427 (N_7427,N_7021,N_7176);
and U7428 (N_7428,N_7177,N_7211);
nand U7429 (N_7429,N_7240,N_7179);
nand U7430 (N_7430,N_7038,N_7083);
or U7431 (N_7431,N_7225,N_7227);
or U7432 (N_7432,N_7230,N_7040);
nor U7433 (N_7433,N_7014,N_7122);
or U7434 (N_7434,N_7162,N_7173);
xor U7435 (N_7435,N_7237,N_7181);
or U7436 (N_7436,N_7042,N_7082);
and U7437 (N_7437,N_7185,N_7051);
xor U7438 (N_7438,N_7074,N_7203);
and U7439 (N_7439,N_7164,N_7173);
or U7440 (N_7440,N_7040,N_7152);
and U7441 (N_7441,N_7154,N_7235);
or U7442 (N_7442,N_7193,N_7093);
and U7443 (N_7443,N_7145,N_7231);
xor U7444 (N_7444,N_7107,N_7004);
nor U7445 (N_7445,N_7094,N_7172);
xnor U7446 (N_7446,N_7100,N_7168);
nand U7447 (N_7447,N_7120,N_7090);
nor U7448 (N_7448,N_7061,N_7150);
nand U7449 (N_7449,N_7019,N_7207);
or U7450 (N_7450,N_7144,N_7026);
and U7451 (N_7451,N_7213,N_7094);
nand U7452 (N_7452,N_7100,N_7189);
nand U7453 (N_7453,N_7100,N_7092);
nand U7454 (N_7454,N_7042,N_7115);
nor U7455 (N_7455,N_7079,N_7176);
xor U7456 (N_7456,N_7042,N_7119);
nor U7457 (N_7457,N_7243,N_7083);
nor U7458 (N_7458,N_7127,N_7115);
or U7459 (N_7459,N_7233,N_7182);
and U7460 (N_7460,N_7094,N_7032);
xor U7461 (N_7461,N_7009,N_7061);
xor U7462 (N_7462,N_7246,N_7168);
xor U7463 (N_7463,N_7129,N_7041);
and U7464 (N_7464,N_7233,N_7168);
and U7465 (N_7465,N_7210,N_7156);
xor U7466 (N_7466,N_7224,N_7245);
nand U7467 (N_7467,N_7237,N_7136);
and U7468 (N_7468,N_7062,N_7026);
nor U7469 (N_7469,N_7112,N_7187);
or U7470 (N_7470,N_7148,N_7239);
and U7471 (N_7471,N_7127,N_7146);
xnor U7472 (N_7472,N_7115,N_7180);
nand U7473 (N_7473,N_7081,N_7116);
nand U7474 (N_7474,N_7232,N_7152);
and U7475 (N_7475,N_7212,N_7227);
or U7476 (N_7476,N_7051,N_7067);
or U7477 (N_7477,N_7111,N_7121);
or U7478 (N_7478,N_7222,N_7238);
or U7479 (N_7479,N_7241,N_7092);
or U7480 (N_7480,N_7227,N_7034);
or U7481 (N_7481,N_7064,N_7208);
nor U7482 (N_7482,N_7145,N_7096);
or U7483 (N_7483,N_7201,N_7217);
nor U7484 (N_7484,N_7234,N_7149);
xnor U7485 (N_7485,N_7146,N_7145);
xor U7486 (N_7486,N_7054,N_7037);
nor U7487 (N_7487,N_7223,N_7242);
nand U7488 (N_7488,N_7189,N_7040);
and U7489 (N_7489,N_7245,N_7128);
nand U7490 (N_7490,N_7032,N_7097);
nand U7491 (N_7491,N_7240,N_7117);
nor U7492 (N_7492,N_7149,N_7017);
xnor U7493 (N_7493,N_7051,N_7022);
nand U7494 (N_7494,N_7041,N_7111);
nor U7495 (N_7495,N_7129,N_7112);
and U7496 (N_7496,N_7036,N_7148);
nor U7497 (N_7497,N_7082,N_7097);
or U7498 (N_7498,N_7042,N_7158);
or U7499 (N_7499,N_7107,N_7170);
or U7500 (N_7500,N_7284,N_7256);
and U7501 (N_7501,N_7322,N_7462);
and U7502 (N_7502,N_7382,N_7427);
xnor U7503 (N_7503,N_7344,N_7375);
or U7504 (N_7504,N_7254,N_7476);
nand U7505 (N_7505,N_7474,N_7315);
nor U7506 (N_7506,N_7250,N_7394);
nor U7507 (N_7507,N_7434,N_7361);
and U7508 (N_7508,N_7417,N_7346);
or U7509 (N_7509,N_7477,N_7333);
or U7510 (N_7510,N_7472,N_7255);
and U7511 (N_7511,N_7395,N_7410);
nor U7512 (N_7512,N_7279,N_7483);
and U7513 (N_7513,N_7331,N_7321);
nand U7514 (N_7514,N_7492,N_7459);
xor U7515 (N_7515,N_7314,N_7305);
xnor U7516 (N_7516,N_7251,N_7493);
or U7517 (N_7517,N_7408,N_7264);
xnor U7518 (N_7518,N_7450,N_7429);
nand U7519 (N_7519,N_7411,N_7336);
or U7520 (N_7520,N_7262,N_7350);
nor U7521 (N_7521,N_7405,N_7392);
nand U7522 (N_7522,N_7400,N_7376);
and U7523 (N_7523,N_7357,N_7292);
xor U7524 (N_7524,N_7290,N_7340);
and U7525 (N_7525,N_7478,N_7372);
or U7526 (N_7526,N_7311,N_7325);
and U7527 (N_7527,N_7317,N_7277);
nor U7528 (N_7528,N_7287,N_7419);
xor U7529 (N_7529,N_7380,N_7454);
xnor U7530 (N_7530,N_7275,N_7297);
nor U7531 (N_7531,N_7300,N_7289);
nand U7532 (N_7532,N_7258,N_7366);
and U7533 (N_7533,N_7466,N_7433);
xnor U7534 (N_7534,N_7413,N_7443);
or U7535 (N_7535,N_7378,N_7332);
nor U7536 (N_7536,N_7278,N_7288);
nor U7537 (N_7537,N_7407,N_7269);
and U7538 (N_7538,N_7482,N_7316);
xor U7539 (N_7539,N_7460,N_7402);
and U7540 (N_7540,N_7456,N_7270);
nor U7541 (N_7541,N_7498,N_7267);
or U7542 (N_7542,N_7319,N_7324);
or U7543 (N_7543,N_7370,N_7312);
or U7544 (N_7544,N_7309,N_7307);
nor U7545 (N_7545,N_7449,N_7391);
or U7546 (N_7546,N_7455,N_7488);
xor U7547 (N_7547,N_7355,N_7435);
nor U7548 (N_7548,N_7441,N_7379);
xor U7549 (N_7549,N_7327,N_7383);
xnor U7550 (N_7550,N_7257,N_7403);
nand U7551 (N_7551,N_7369,N_7389);
and U7552 (N_7552,N_7368,N_7387);
xor U7553 (N_7553,N_7323,N_7363);
or U7554 (N_7554,N_7479,N_7373);
and U7555 (N_7555,N_7426,N_7320);
and U7556 (N_7556,N_7351,N_7281);
xnor U7557 (N_7557,N_7365,N_7499);
nand U7558 (N_7558,N_7438,N_7416);
nor U7559 (N_7559,N_7458,N_7354);
nor U7560 (N_7560,N_7345,N_7381);
or U7561 (N_7561,N_7339,N_7457);
xnor U7562 (N_7562,N_7259,N_7385);
xnor U7563 (N_7563,N_7306,N_7406);
nor U7564 (N_7564,N_7296,N_7442);
nor U7565 (N_7565,N_7489,N_7304);
and U7566 (N_7566,N_7447,N_7283);
nand U7567 (N_7567,N_7465,N_7253);
nand U7568 (N_7568,N_7282,N_7390);
and U7569 (N_7569,N_7470,N_7495);
nand U7570 (N_7570,N_7347,N_7341);
and U7571 (N_7571,N_7342,N_7485);
and U7572 (N_7572,N_7494,N_7431);
nand U7573 (N_7573,N_7446,N_7348);
or U7574 (N_7574,N_7261,N_7352);
xor U7575 (N_7575,N_7263,N_7418);
and U7576 (N_7576,N_7440,N_7334);
or U7577 (N_7577,N_7404,N_7424);
and U7578 (N_7578,N_7299,N_7266);
nor U7579 (N_7579,N_7329,N_7497);
nor U7580 (N_7580,N_7415,N_7445);
or U7581 (N_7581,N_7401,N_7409);
and U7582 (N_7582,N_7298,N_7393);
nor U7583 (N_7583,N_7448,N_7285);
or U7584 (N_7584,N_7353,N_7301);
xor U7585 (N_7585,N_7265,N_7484);
or U7586 (N_7586,N_7295,N_7496);
xor U7587 (N_7587,N_7422,N_7293);
nand U7588 (N_7588,N_7471,N_7469);
nor U7589 (N_7589,N_7313,N_7272);
xor U7590 (N_7590,N_7308,N_7467);
nor U7591 (N_7591,N_7388,N_7384);
xnor U7592 (N_7592,N_7421,N_7252);
nand U7593 (N_7593,N_7359,N_7364);
nor U7594 (N_7594,N_7420,N_7291);
or U7595 (N_7595,N_7439,N_7428);
xor U7596 (N_7596,N_7463,N_7374);
or U7597 (N_7597,N_7343,N_7260);
xor U7598 (N_7598,N_7453,N_7280);
and U7599 (N_7599,N_7432,N_7436);
nand U7600 (N_7600,N_7475,N_7437);
or U7601 (N_7601,N_7386,N_7464);
xor U7602 (N_7602,N_7358,N_7414);
xnor U7603 (N_7603,N_7362,N_7360);
nand U7604 (N_7604,N_7326,N_7480);
xor U7605 (N_7605,N_7423,N_7330);
xor U7606 (N_7606,N_7398,N_7349);
xor U7607 (N_7607,N_7273,N_7444);
nor U7608 (N_7608,N_7268,N_7490);
or U7609 (N_7609,N_7452,N_7396);
and U7610 (N_7610,N_7377,N_7271);
nand U7611 (N_7611,N_7294,N_7371);
nand U7612 (N_7612,N_7487,N_7274);
nor U7613 (N_7613,N_7481,N_7399);
nand U7614 (N_7614,N_7473,N_7412);
xnor U7615 (N_7615,N_7302,N_7356);
xor U7616 (N_7616,N_7430,N_7335);
xnor U7617 (N_7617,N_7318,N_7491);
and U7618 (N_7618,N_7461,N_7303);
nand U7619 (N_7619,N_7486,N_7310);
nand U7620 (N_7620,N_7468,N_7451);
or U7621 (N_7621,N_7338,N_7397);
and U7622 (N_7622,N_7328,N_7337);
and U7623 (N_7623,N_7286,N_7276);
nor U7624 (N_7624,N_7367,N_7425);
xor U7625 (N_7625,N_7352,N_7298);
nor U7626 (N_7626,N_7367,N_7445);
nand U7627 (N_7627,N_7492,N_7340);
and U7628 (N_7628,N_7422,N_7264);
nand U7629 (N_7629,N_7281,N_7288);
or U7630 (N_7630,N_7436,N_7433);
or U7631 (N_7631,N_7267,N_7279);
and U7632 (N_7632,N_7466,N_7467);
xor U7633 (N_7633,N_7437,N_7418);
nor U7634 (N_7634,N_7289,N_7385);
and U7635 (N_7635,N_7342,N_7436);
nor U7636 (N_7636,N_7333,N_7418);
xor U7637 (N_7637,N_7457,N_7259);
nand U7638 (N_7638,N_7302,N_7430);
nand U7639 (N_7639,N_7270,N_7497);
and U7640 (N_7640,N_7482,N_7277);
nor U7641 (N_7641,N_7472,N_7257);
nand U7642 (N_7642,N_7422,N_7333);
or U7643 (N_7643,N_7376,N_7426);
or U7644 (N_7644,N_7331,N_7286);
or U7645 (N_7645,N_7348,N_7337);
nand U7646 (N_7646,N_7492,N_7489);
xor U7647 (N_7647,N_7352,N_7468);
or U7648 (N_7648,N_7412,N_7339);
nor U7649 (N_7649,N_7286,N_7259);
xnor U7650 (N_7650,N_7352,N_7318);
nor U7651 (N_7651,N_7323,N_7264);
nor U7652 (N_7652,N_7284,N_7305);
nand U7653 (N_7653,N_7498,N_7284);
nor U7654 (N_7654,N_7482,N_7468);
or U7655 (N_7655,N_7395,N_7305);
or U7656 (N_7656,N_7312,N_7491);
and U7657 (N_7657,N_7486,N_7364);
nor U7658 (N_7658,N_7394,N_7384);
and U7659 (N_7659,N_7287,N_7318);
xor U7660 (N_7660,N_7250,N_7426);
nor U7661 (N_7661,N_7295,N_7461);
and U7662 (N_7662,N_7398,N_7357);
nand U7663 (N_7663,N_7364,N_7269);
nand U7664 (N_7664,N_7339,N_7397);
nor U7665 (N_7665,N_7422,N_7376);
nor U7666 (N_7666,N_7399,N_7295);
xor U7667 (N_7667,N_7302,N_7416);
and U7668 (N_7668,N_7337,N_7262);
nor U7669 (N_7669,N_7375,N_7473);
and U7670 (N_7670,N_7391,N_7304);
xor U7671 (N_7671,N_7369,N_7378);
xor U7672 (N_7672,N_7307,N_7283);
nor U7673 (N_7673,N_7440,N_7401);
and U7674 (N_7674,N_7490,N_7426);
and U7675 (N_7675,N_7367,N_7459);
or U7676 (N_7676,N_7447,N_7363);
nand U7677 (N_7677,N_7396,N_7425);
nand U7678 (N_7678,N_7301,N_7351);
nand U7679 (N_7679,N_7410,N_7327);
or U7680 (N_7680,N_7474,N_7408);
nor U7681 (N_7681,N_7272,N_7464);
xor U7682 (N_7682,N_7258,N_7344);
or U7683 (N_7683,N_7324,N_7356);
nand U7684 (N_7684,N_7386,N_7329);
or U7685 (N_7685,N_7476,N_7438);
xor U7686 (N_7686,N_7426,N_7287);
and U7687 (N_7687,N_7481,N_7292);
nand U7688 (N_7688,N_7312,N_7290);
nand U7689 (N_7689,N_7420,N_7322);
and U7690 (N_7690,N_7475,N_7320);
nand U7691 (N_7691,N_7272,N_7264);
nor U7692 (N_7692,N_7445,N_7406);
xnor U7693 (N_7693,N_7352,N_7265);
or U7694 (N_7694,N_7419,N_7361);
nand U7695 (N_7695,N_7335,N_7393);
xnor U7696 (N_7696,N_7408,N_7274);
and U7697 (N_7697,N_7319,N_7409);
nand U7698 (N_7698,N_7369,N_7269);
nand U7699 (N_7699,N_7312,N_7414);
nor U7700 (N_7700,N_7256,N_7439);
nor U7701 (N_7701,N_7417,N_7321);
xor U7702 (N_7702,N_7446,N_7497);
or U7703 (N_7703,N_7437,N_7327);
nand U7704 (N_7704,N_7377,N_7465);
xnor U7705 (N_7705,N_7252,N_7351);
and U7706 (N_7706,N_7366,N_7375);
nand U7707 (N_7707,N_7410,N_7253);
and U7708 (N_7708,N_7369,N_7467);
or U7709 (N_7709,N_7499,N_7254);
nand U7710 (N_7710,N_7352,N_7359);
xor U7711 (N_7711,N_7499,N_7466);
and U7712 (N_7712,N_7277,N_7374);
and U7713 (N_7713,N_7331,N_7289);
nor U7714 (N_7714,N_7376,N_7438);
xor U7715 (N_7715,N_7499,N_7356);
nand U7716 (N_7716,N_7333,N_7314);
and U7717 (N_7717,N_7492,N_7281);
nand U7718 (N_7718,N_7356,N_7386);
or U7719 (N_7719,N_7305,N_7430);
nand U7720 (N_7720,N_7286,N_7250);
nor U7721 (N_7721,N_7491,N_7370);
nor U7722 (N_7722,N_7429,N_7283);
xnor U7723 (N_7723,N_7280,N_7497);
and U7724 (N_7724,N_7309,N_7301);
nand U7725 (N_7725,N_7296,N_7259);
xnor U7726 (N_7726,N_7343,N_7461);
and U7727 (N_7727,N_7423,N_7371);
nor U7728 (N_7728,N_7339,N_7293);
and U7729 (N_7729,N_7417,N_7267);
nand U7730 (N_7730,N_7265,N_7467);
or U7731 (N_7731,N_7403,N_7385);
nor U7732 (N_7732,N_7387,N_7477);
xnor U7733 (N_7733,N_7466,N_7419);
and U7734 (N_7734,N_7454,N_7372);
nor U7735 (N_7735,N_7476,N_7282);
xnor U7736 (N_7736,N_7258,N_7451);
and U7737 (N_7737,N_7332,N_7363);
nand U7738 (N_7738,N_7394,N_7386);
nand U7739 (N_7739,N_7419,N_7426);
or U7740 (N_7740,N_7384,N_7312);
nand U7741 (N_7741,N_7319,N_7482);
nor U7742 (N_7742,N_7455,N_7492);
and U7743 (N_7743,N_7255,N_7312);
or U7744 (N_7744,N_7369,N_7280);
and U7745 (N_7745,N_7301,N_7314);
xnor U7746 (N_7746,N_7364,N_7296);
and U7747 (N_7747,N_7356,N_7423);
and U7748 (N_7748,N_7414,N_7428);
or U7749 (N_7749,N_7403,N_7448);
nand U7750 (N_7750,N_7598,N_7630);
and U7751 (N_7751,N_7726,N_7657);
or U7752 (N_7752,N_7645,N_7700);
or U7753 (N_7753,N_7651,N_7658);
or U7754 (N_7754,N_7639,N_7673);
xor U7755 (N_7755,N_7519,N_7669);
nand U7756 (N_7756,N_7563,N_7614);
nand U7757 (N_7757,N_7525,N_7650);
nor U7758 (N_7758,N_7637,N_7540);
and U7759 (N_7759,N_7594,N_7617);
or U7760 (N_7760,N_7547,N_7682);
nand U7761 (N_7761,N_7578,N_7719);
nand U7762 (N_7762,N_7609,N_7735);
xnor U7763 (N_7763,N_7572,N_7557);
or U7764 (N_7764,N_7672,N_7646);
and U7765 (N_7765,N_7661,N_7693);
nor U7766 (N_7766,N_7718,N_7686);
xnor U7767 (N_7767,N_7517,N_7599);
or U7768 (N_7768,N_7558,N_7644);
nand U7769 (N_7769,N_7605,N_7505);
or U7770 (N_7770,N_7641,N_7706);
nand U7771 (N_7771,N_7668,N_7539);
or U7772 (N_7772,N_7627,N_7511);
nand U7773 (N_7773,N_7733,N_7723);
or U7774 (N_7774,N_7732,N_7537);
or U7775 (N_7775,N_7656,N_7667);
and U7776 (N_7776,N_7549,N_7579);
nand U7777 (N_7777,N_7591,N_7555);
xor U7778 (N_7778,N_7683,N_7606);
and U7779 (N_7779,N_7602,N_7701);
xor U7780 (N_7780,N_7649,N_7575);
or U7781 (N_7781,N_7721,N_7541);
nand U7782 (N_7782,N_7642,N_7516);
or U7783 (N_7783,N_7622,N_7526);
nand U7784 (N_7784,N_7713,N_7708);
nand U7785 (N_7785,N_7648,N_7633);
nand U7786 (N_7786,N_7694,N_7687);
or U7787 (N_7787,N_7666,N_7534);
nand U7788 (N_7788,N_7556,N_7738);
xor U7789 (N_7789,N_7520,N_7685);
xnor U7790 (N_7790,N_7565,N_7542);
or U7791 (N_7791,N_7566,N_7709);
or U7792 (N_7792,N_7613,N_7634);
nor U7793 (N_7793,N_7736,N_7740);
and U7794 (N_7794,N_7731,N_7724);
xnor U7795 (N_7795,N_7524,N_7628);
or U7796 (N_7796,N_7638,N_7521);
or U7797 (N_7797,N_7576,N_7569);
nand U7798 (N_7798,N_7715,N_7678);
nor U7799 (N_7799,N_7507,N_7523);
nand U7800 (N_7800,N_7528,N_7500);
and U7801 (N_7801,N_7664,N_7704);
nor U7802 (N_7802,N_7546,N_7691);
xnor U7803 (N_7803,N_7562,N_7508);
nand U7804 (N_7804,N_7545,N_7655);
nand U7805 (N_7805,N_7714,N_7616);
or U7806 (N_7806,N_7544,N_7699);
xnor U7807 (N_7807,N_7611,N_7564);
nor U7808 (N_7808,N_7727,N_7696);
or U7809 (N_7809,N_7502,N_7527);
nor U7810 (N_7810,N_7745,N_7529);
nor U7811 (N_7811,N_7515,N_7554);
nor U7812 (N_7812,N_7747,N_7601);
nor U7813 (N_7813,N_7741,N_7550);
nor U7814 (N_7814,N_7621,N_7504);
xnor U7815 (N_7815,N_7739,N_7584);
nand U7816 (N_7816,N_7671,N_7513);
or U7817 (N_7817,N_7670,N_7543);
nor U7818 (N_7818,N_7625,N_7593);
nand U7819 (N_7819,N_7716,N_7619);
nand U7820 (N_7820,N_7618,N_7744);
or U7821 (N_7821,N_7580,N_7624);
xor U7822 (N_7822,N_7567,N_7577);
and U7823 (N_7823,N_7743,N_7503);
nand U7824 (N_7824,N_7588,N_7612);
nand U7825 (N_7825,N_7560,N_7742);
or U7826 (N_7826,N_7688,N_7623);
nand U7827 (N_7827,N_7573,N_7610);
xnor U7828 (N_7828,N_7674,N_7695);
nand U7829 (N_7829,N_7553,N_7631);
xnor U7830 (N_7830,N_7681,N_7662);
and U7831 (N_7831,N_7707,N_7582);
nand U7832 (N_7832,N_7589,N_7665);
nand U7833 (N_7833,N_7531,N_7568);
or U7834 (N_7834,N_7533,N_7587);
nor U7835 (N_7835,N_7675,N_7561);
or U7836 (N_7836,N_7679,N_7538);
or U7837 (N_7837,N_7663,N_7676);
nand U7838 (N_7838,N_7603,N_7720);
or U7839 (N_7839,N_7703,N_7729);
or U7840 (N_7840,N_7640,N_7710);
nand U7841 (N_7841,N_7725,N_7607);
nand U7842 (N_7842,N_7643,N_7570);
or U7843 (N_7843,N_7711,N_7522);
nand U7844 (N_7844,N_7514,N_7501);
nor U7845 (N_7845,N_7660,N_7530);
nor U7846 (N_7846,N_7548,N_7712);
nor U7847 (N_7847,N_7728,N_7652);
nor U7848 (N_7848,N_7592,N_7597);
and U7849 (N_7849,N_7559,N_7532);
nand U7850 (N_7850,N_7659,N_7722);
nor U7851 (N_7851,N_7692,N_7680);
or U7852 (N_7852,N_7626,N_7535);
nand U7853 (N_7853,N_7734,N_7629);
and U7854 (N_7854,N_7596,N_7571);
and U7855 (N_7855,N_7509,N_7653);
or U7856 (N_7856,N_7512,N_7581);
nand U7857 (N_7857,N_7510,N_7590);
xor U7858 (N_7858,N_7737,N_7551);
xor U7859 (N_7859,N_7574,N_7749);
and U7860 (N_7860,N_7615,N_7698);
or U7861 (N_7861,N_7697,N_7552);
and U7862 (N_7862,N_7717,N_7595);
or U7863 (N_7863,N_7604,N_7635);
and U7864 (N_7864,N_7690,N_7702);
and U7865 (N_7865,N_7684,N_7632);
nand U7866 (N_7866,N_7586,N_7705);
nor U7867 (N_7867,N_7506,N_7600);
and U7868 (N_7868,N_7730,N_7636);
nand U7869 (N_7869,N_7585,N_7647);
nand U7870 (N_7870,N_7746,N_7536);
or U7871 (N_7871,N_7620,N_7518);
or U7872 (N_7872,N_7748,N_7583);
nand U7873 (N_7873,N_7677,N_7689);
xnor U7874 (N_7874,N_7654,N_7608);
xor U7875 (N_7875,N_7507,N_7524);
and U7876 (N_7876,N_7625,N_7694);
nand U7877 (N_7877,N_7519,N_7553);
and U7878 (N_7878,N_7589,N_7570);
or U7879 (N_7879,N_7653,N_7507);
or U7880 (N_7880,N_7527,N_7707);
and U7881 (N_7881,N_7614,N_7702);
nor U7882 (N_7882,N_7700,N_7586);
nand U7883 (N_7883,N_7562,N_7529);
and U7884 (N_7884,N_7503,N_7736);
nor U7885 (N_7885,N_7690,N_7526);
or U7886 (N_7886,N_7560,N_7670);
xnor U7887 (N_7887,N_7678,N_7604);
or U7888 (N_7888,N_7662,N_7628);
nand U7889 (N_7889,N_7552,N_7728);
and U7890 (N_7890,N_7619,N_7709);
nand U7891 (N_7891,N_7607,N_7599);
xor U7892 (N_7892,N_7515,N_7575);
nor U7893 (N_7893,N_7650,N_7684);
or U7894 (N_7894,N_7641,N_7591);
nand U7895 (N_7895,N_7667,N_7553);
nand U7896 (N_7896,N_7744,N_7630);
xor U7897 (N_7897,N_7625,N_7623);
and U7898 (N_7898,N_7739,N_7668);
and U7899 (N_7899,N_7724,N_7603);
nand U7900 (N_7900,N_7500,N_7681);
xor U7901 (N_7901,N_7597,N_7694);
xor U7902 (N_7902,N_7641,N_7701);
and U7903 (N_7903,N_7523,N_7545);
and U7904 (N_7904,N_7644,N_7646);
nor U7905 (N_7905,N_7707,N_7535);
xor U7906 (N_7906,N_7703,N_7632);
or U7907 (N_7907,N_7680,N_7644);
or U7908 (N_7908,N_7574,N_7696);
xor U7909 (N_7909,N_7653,N_7613);
and U7910 (N_7910,N_7533,N_7579);
nor U7911 (N_7911,N_7646,N_7507);
xnor U7912 (N_7912,N_7511,N_7618);
and U7913 (N_7913,N_7557,N_7532);
or U7914 (N_7914,N_7569,N_7648);
or U7915 (N_7915,N_7657,N_7555);
xnor U7916 (N_7916,N_7655,N_7653);
xnor U7917 (N_7917,N_7641,N_7660);
xor U7918 (N_7918,N_7559,N_7561);
or U7919 (N_7919,N_7507,N_7568);
and U7920 (N_7920,N_7605,N_7717);
nor U7921 (N_7921,N_7689,N_7583);
and U7922 (N_7922,N_7575,N_7502);
nand U7923 (N_7923,N_7524,N_7600);
nor U7924 (N_7924,N_7742,N_7507);
nand U7925 (N_7925,N_7526,N_7582);
xor U7926 (N_7926,N_7676,N_7621);
or U7927 (N_7927,N_7633,N_7661);
xnor U7928 (N_7928,N_7701,N_7654);
xnor U7929 (N_7929,N_7590,N_7558);
nand U7930 (N_7930,N_7674,N_7620);
nor U7931 (N_7931,N_7696,N_7718);
nand U7932 (N_7932,N_7642,N_7601);
and U7933 (N_7933,N_7611,N_7666);
xnor U7934 (N_7934,N_7743,N_7598);
and U7935 (N_7935,N_7708,N_7640);
or U7936 (N_7936,N_7552,N_7677);
and U7937 (N_7937,N_7748,N_7728);
or U7938 (N_7938,N_7671,N_7599);
and U7939 (N_7939,N_7616,N_7709);
and U7940 (N_7940,N_7655,N_7693);
and U7941 (N_7941,N_7582,N_7626);
or U7942 (N_7942,N_7568,N_7610);
nor U7943 (N_7943,N_7712,N_7624);
nor U7944 (N_7944,N_7683,N_7707);
nand U7945 (N_7945,N_7646,N_7668);
or U7946 (N_7946,N_7640,N_7518);
or U7947 (N_7947,N_7591,N_7513);
xor U7948 (N_7948,N_7651,N_7741);
or U7949 (N_7949,N_7630,N_7517);
or U7950 (N_7950,N_7565,N_7691);
nand U7951 (N_7951,N_7572,N_7619);
nor U7952 (N_7952,N_7671,N_7740);
and U7953 (N_7953,N_7737,N_7673);
and U7954 (N_7954,N_7727,N_7640);
nand U7955 (N_7955,N_7733,N_7643);
or U7956 (N_7956,N_7712,N_7502);
and U7957 (N_7957,N_7603,N_7606);
and U7958 (N_7958,N_7551,N_7693);
nand U7959 (N_7959,N_7556,N_7656);
xnor U7960 (N_7960,N_7647,N_7576);
and U7961 (N_7961,N_7540,N_7728);
xnor U7962 (N_7962,N_7561,N_7564);
and U7963 (N_7963,N_7689,N_7525);
nand U7964 (N_7964,N_7729,N_7582);
nor U7965 (N_7965,N_7515,N_7658);
nor U7966 (N_7966,N_7523,N_7661);
and U7967 (N_7967,N_7542,N_7609);
xnor U7968 (N_7968,N_7533,N_7738);
nand U7969 (N_7969,N_7620,N_7683);
nor U7970 (N_7970,N_7747,N_7620);
xor U7971 (N_7971,N_7653,N_7514);
and U7972 (N_7972,N_7634,N_7697);
and U7973 (N_7973,N_7574,N_7590);
nand U7974 (N_7974,N_7737,N_7677);
xnor U7975 (N_7975,N_7511,N_7516);
nand U7976 (N_7976,N_7707,N_7612);
or U7977 (N_7977,N_7593,N_7728);
nand U7978 (N_7978,N_7626,N_7638);
and U7979 (N_7979,N_7668,N_7564);
or U7980 (N_7980,N_7581,N_7556);
nand U7981 (N_7981,N_7674,N_7505);
nor U7982 (N_7982,N_7618,N_7626);
xnor U7983 (N_7983,N_7549,N_7695);
and U7984 (N_7984,N_7538,N_7618);
and U7985 (N_7985,N_7736,N_7716);
nor U7986 (N_7986,N_7573,N_7710);
and U7987 (N_7987,N_7695,N_7507);
nand U7988 (N_7988,N_7539,N_7720);
xor U7989 (N_7989,N_7511,N_7745);
xor U7990 (N_7990,N_7731,N_7627);
nor U7991 (N_7991,N_7649,N_7546);
or U7992 (N_7992,N_7745,N_7615);
or U7993 (N_7993,N_7611,N_7677);
or U7994 (N_7994,N_7587,N_7620);
or U7995 (N_7995,N_7616,N_7707);
nor U7996 (N_7996,N_7602,N_7690);
nor U7997 (N_7997,N_7505,N_7696);
xor U7998 (N_7998,N_7692,N_7678);
and U7999 (N_7999,N_7574,N_7512);
nor U8000 (N_8000,N_7751,N_7871);
nand U8001 (N_8001,N_7813,N_7977);
and U8002 (N_8002,N_7825,N_7865);
or U8003 (N_8003,N_7873,N_7788);
nand U8004 (N_8004,N_7759,N_7796);
nand U8005 (N_8005,N_7911,N_7899);
or U8006 (N_8006,N_7864,N_7889);
and U8007 (N_8007,N_7815,N_7845);
nand U8008 (N_8008,N_7883,N_7920);
or U8009 (N_8009,N_7757,N_7786);
nor U8010 (N_8010,N_7863,N_7988);
nand U8011 (N_8011,N_7772,N_7769);
and U8012 (N_8012,N_7995,N_7999);
and U8013 (N_8013,N_7805,N_7846);
and U8014 (N_8014,N_7997,N_7758);
or U8015 (N_8015,N_7798,N_7937);
or U8016 (N_8016,N_7902,N_7755);
and U8017 (N_8017,N_7934,N_7910);
nor U8018 (N_8018,N_7963,N_7784);
nor U8019 (N_8019,N_7985,N_7981);
xor U8020 (N_8020,N_7917,N_7840);
nor U8021 (N_8021,N_7993,N_7848);
nor U8022 (N_8022,N_7967,N_7909);
nor U8023 (N_8023,N_7955,N_7959);
nand U8024 (N_8024,N_7996,N_7836);
nor U8025 (N_8025,N_7881,N_7927);
and U8026 (N_8026,N_7768,N_7913);
and U8027 (N_8027,N_7794,N_7940);
nor U8028 (N_8028,N_7898,N_7832);
xnor U8029 (N_8029,N_7808,N_7849);
xor U8030 (N_8030,N_7842,N_7753);
nand U8031 (N_8031,N_7953,N_7931);
and U8032 (N_8032,N_7976,N_7847);
xor U8033 (N_8033,N_7994,N_7947);
xnor U8034 (N_8034,N_7965,N_7879);
or U8035 (N_8035,N_7990,N_7904);
nor U8036 (N_8036,N_7775,N_7973);
or U8037 (N_8037,N_7754,N_7799);
nand U8038 (N_8038,N_7958,N_7801);
or U8039 (N_8039,N_7893,N_7980);
and U8040 (N_8040,N_7935,N_7966);
and U8041 (N_8041,N_7826,N_7960);
or U8042 (N_8042,N_7766,N_7945);
or U8043 (N_8043,N_7835,N_7892);
or U8044 (N_8044,N_7928,N_7764);
nor U8045 (N_8045,N_7860,N_7903);
xnor U8046 (N_8046,N_7831,N_7918);
xor U8047 (N_8047,N_7936,N_7867);
nand U8048 (N_8048,N_7854,N_7880);
nand U8049 (N_8049,N_7908,N_7861);
nor U8050 (N_8050,N_7816,N_7779);
nand U8051 (N_8051,N_7807,N_7773);
or U8052 (N_8052,N_7986,N_7791);
nor U8053 (N_8053,N_7789,N_7915);
and U8054 (N_8054,N_7774,N_7933);
xnor U8055 (N_8055,N_7824,N_7767);
and U8056 (N_8056,N_7869,N_7752);
xor U8057 (N_8057,N_7841,N_7888);
xor U8058 (N_8058,N_7763,N_7961);
and U8059 (N_8059,N_7803,N_7851);
nor U8060 (N_8060,N_7852,N_7942);
or U8061 (N_8061,N_7761,N_7785);
nand U8062 (N_8062,N_7930,N_7975);
nor U8063 (N_8063,N_7837,N_7951);
and U8064 (N_8064,N_7897,N_7964);
nor U8065 (N_8065,N_7885,N_7790);
xor U8066 (N_8066,N_7810,N_7797);
xnor U8067 (N_8067,N_7954,N_7868);
nand U8068 (N_8068,N_7820,N_7912);
nor U8069 (N_8069,N_7962,N_7821);
and U8070 (N_8070,N_7957,N_7890);
xor U8071 (N_8071,N_7787,N_7968);
and U8072 (N_8072,N_7882,N_7819);
xor U8073 (N_8073,N_7877,N_7900);
xor U8074 (N_8074,N_7828,N_7924);
and U8075 (N_8075,N_7943,N_7853);
nor U8076 (N_8076,N_7916,N_7983);
nor U8077 (N_8077,N_7950,N_7843);
and U8078 (N_8078,N_7829,N_7974);
and U8079 (N_8079,N_7891,N_7948);
nand U8080 (N_8080,N_7765,N_7907);
xor U8081 (N_8081,N_7858,N_7781);
or U8082 (N_8082,N_7972,N_7795);
xnor U8083 (N_8083,N_7834,N_7938);
xor U8084 (N_8084,N_7875,N_7992);
and U8085 (N_8085,N_7776,N_7770);
nor U8086 (N_8086,N_7894,N_7982);
nand U8087 (N_8087,N_7946,N_7809);
nand U8088 (N_8088,N_7830,N_7896);
or U8089 (N_8089,N_7949,N_7923);
nor U8090 (N_8090,N_7922,N_7804);
nand U8091 (N_8091,N_7901,N_7906);
and U8092 (N_8092,N_7921,N_7970);
xnor U8093 (N_8093,N_7792,N_7811);
xor U8094 (N_8094,N_7929,N_7783);
and U8095 (N_8095,N_7862,N_7979);
or U8096 (N_8096,N_7812,N_7823);
nor U8097 (N_8097,N_7822,N_7800);
xnor U8098 (N_8098,N_7956,N_7844);
nor U8099 (N_8099,N_7866,N_7857);
xor U8100 (N_8100,N_7760,N_7941);
nand U8101 (N_8101,N_7778,N_7878);
nand U8102 (N_8102,N_7838,N_7814);
nor U8103 (N_8103,N_7850,N_7855);
nand U8104 (N_8104,N_7756,N_7969);
xor U8105 (N_8105,N_7919,N_7872);
xor U8106 (N_8106,N_7839,N_7905);
xnor U8107 (N_8107,N_7827,N_7884);
nand U8108 (N_8108,N_7793,N_7818);
nor U8109 (N_8109,N_7802,N_7887);
nand U8110 (N_8110,N_7856,N_7870);
or U8111 (N_8111,N_7750,N_7952);
and U8112 (N_8112,N_7925,N_7989);
or U8113 (N_8113,N_7971,N_7874);
xor U8114 (N_8114,N_7984,N_7895);
xnor U8115 (N_8115,N_7932,N_7978);
nand U8116 (N_8116,N_7833,N_7886);
nand U8117 (N_8117,N_7817,N_7998);
or U8118 (N_8118,N_7806,N_7859);
nand U8119 (N_8119,N_7771,N_7926);
and U8120 (N_8120,N_7780,N_7939);
xnor U8121 (N_8121,N_7782,N_7777);
nor U8122 (N_8122,N_7762,N_7876);
nor U8123 (N_8123,N_7944,N_7991);
nand U8124 (N_8124,N_7914,N_7987);
xnor U8125 (N_8125,N_7874,N_7949);
nand U8126 (N_8126,N_7815,N_7997);
and U8127 (N_8127,N_7926,N_7778);
nand U8128 (N_8128,N_7891,N_7811);
xnor U8129 (N_8129,N_7894,N_7881);
xor U8130 (N_8130,N_7889,N_7999);
xnor U8131 (N_8131,N_7802,N_7833);
and U8132 (N_8132,N_7793,N_7974);
nor U8133 (N_8133,N_7892,N_7908);
xnor U8134 (N_8134,N_7938,N_7777);
nor U8135 (N_8135,N_7979,N_7831);
nand U8136 (N_8136,N_7844,N_7829);
or U8137 (N_8137,N_7918,N_7895);
nor U8138 (N_8138,N_7979,N_7776);
and U8139 (N_8139,N_7835,N_7837);
nor U8140 (N_8140,N_7807,N_7800);
nor U8141 (N_8141,N_7800,N_7836);
nand U8142 (N_8142,N_7839,N_7922);
or U8143 (N_8143,N_7915,N_7866);
nand U8144 (N_8144,N_7893,N_7996);
xnor U8145 (N_8145,N_7839,N_7847);
or U8146 (N_8146,N_7839,N_7849);
nor U8147 (N_8147,N_7947,N_7973);
and U8148 (N_8148,N_7760,N_7906);
nand U8149 (N_8149,N_7927,N_7813);
or U8150 (N_8150,N_7819,N_7927);
xnor U8151 (N_8151,N_7762,N_7954);
xnor U8152 (N_8152,N_7878,N_7819);
nand U8153 (N_8153,N_7887,N_7783);
or U8154 (N_8154,N_7918,N_7854);
and U8155 (N_8155,N_7774,N_7922);
nor U8156 (N_8156,N_7755,N_7800);
nand U8157 (N_8157,N_7894,N_7916);
nor U8158 (N_8158,N_7879,N_7828);
nor U8159 (N_8159,N_7900,N_7755);
nor U8160 (N_8160,N_7921,N_7828);
or U8161 (N_8161,N_7963,N_7981);
nand U8162 (N_8162,N_7904,N_7929);
and U8163 (N_8163,N_7946,N_7772);
or U8164 (N_8164,N_7890,N_7819);
or U8165 (N_8165,N_7939,N_7876);
or U8166 (N_8166,N_7958,N_7813);
and U8167 (N_8167,N_7805,N_7818);
nor U8168 (N_8168,N_7788,N_7776);
and U8169 (N_8169,N_7751,N_7775);
or U8170 (N_8170,N_7968,N_7809);
nand U8171 (N_8171,N_7876,N_7977);
xnor U8172 (N_8172,N_7800,N_7898);
or U8173 (N_8173,N_7896,N_7751);
or U8174 (N_8174,N_7914,N_7949);
and U8175 (N_8175,N_7907,N_7933);
nand U8176 (N_8176,N_7765,N_7876);
and U8177 (N_8177,N_7945,N_7982);
and U8178 (N_8178,N_7987,N_7755);
nand U8179 (N_8179,N_7762,N_7798);
or U8180 (N_8180,N_7920,N_7926);
nand U8181 (N_8181,N_7926,N_7987);
or U8182 (N_8182,N_7755,N_7886);
nor U8183 (N_8183,N_7796,N_7828);
or U8184 (N_8184,N_7811,N_7941);
xnor U8185 (N_8185,N_7986,N_7753);
xor U8186 (N_8186,N_7855,N_7974);
nor U8187 (N_8187,N_7825,N_7773);
nor U8188 (N_8188,N_7903,N_7886);
xnor U8189 (N_8189,N_7839,N_7846);
or U8190 (N_8190,N_7753,N_7838);
nor U8191 (N_8191,N_7961,N_7983);
or U8192 (N_8192,N_7829,N_7751);
xor U8193 (N_8193,N_7779,N_7894);
xor U8194 (N_8194,N_7804,N_7906);
and U8195 (N_8195,N_7860,N_7919);
or U8196 (N_8196,N_7854,N_7983);
or U8197 (N_8197,N_7994,N_7903);
and U8198 (N_8198,N_7993,N_7911);
nor U8199 (N_8199,N_7971,N_7941);
or U8200 (N_8200,N_7825,N_7815);
xor U8201 (N_8201,N_7864,N_7814);
nor U8202 (N_8202,N_7853,N_7820);
and U8203 (N_8203,N_7938,N_7903);
nor U8204 (N_8204,N_7930,N_7923);
and U8205 (N_8205,N_7752,N_7863);
and U8206 (N_8206,N_7771,N_7862);
nor U8207 (N_8207,N_7837,N_7997);
and U8208 (N_8208,N_7845,N_7836);
nor U8209 (N_8209,N_7976,N_7780);
nand U8210 (N_8210,N_7898,N_7915);
nand U8211 (N_8211,N_7952,N_7766);
or U8212 (N_8212,N_7986,N_7879);
or U8213 (N_8213,N_7840,N_7898);
and U8214 (N_8214,N_7787,N_7839);
and U8215 (N_8215,N_7926,N_7790);
or U8216 (N_8216,N_7758,N_7764);
nand U8217 (N_8217,N_7882,N_7931);
or U8218 (N_8218,N_7884,N_7875);
nor U8219 (N_8219,N_7874,N_7970);
nand U8220 (N_8220,N_7813,N_7951);
or U8221 (N_8221,N_7970,N_7976);
and U8222 (N_8222,N_7887,N_7943);
xnor U8223 (N_8223,N_7783,N_7960);
nor U8224 (N_8224,N_7894,N_7990);
xnor U8225 (N_8225,N_7923,N_7802);
or U8226 (N_8226,N_7914,N_7957);
nor U8227 (N_8227,N_7792,N_7801);
or U8228 (N_8228,N_7931,N_7930);
nor U8229 (N_8229,N_7946,N_7842);
nand U8230 (N_8230,N_7860,N_7833);
nand U8231 (N_8231,N_7780,N_7935);
nand U8232 (N_8232,N_7763,N_7810);
nor U8233 (N_8233,N_7929,N_7806);
xor U8234 (N_8234,N_7936,N_7792);
nand U8235 (N_8235,N_7971,N_7758);
nor U8236 (N_8236,N_7966,N_7978);
or U8237 (N_8237,N_7950,N_7858);
and U8238 (N_8238,N_7977,N_7782);
and U8239 (N_8239,N_7934,N_7755);
xor U8240 (N_8240,N_7774,N_7770);
xnor U8241 (N_8241,N_7906,N_7931);
or U8242 (N_8242,N_7873,N_7945);
nor U8243 (N_8243,N_7989,N_7933);
and U8244 (N_8244,N_7870,N_7781);
nor U8245 (N_8245,N_7795,N_7803);
and U8246 (N_8246,N_7985,N_7927);
xnor U8247 (N_8247,N_7760,N_7773);
xor U8248 (N_8248,N_7781,N_7903);
nor U8249 (N_8249,N_7940,N_7766);
xnor U8250 (N_8250,N_8002,N_8074);
nand U8251 (N_8251,N_8070,N_8038);
xor U8252 (N_8252,N_8129,N_8235);
xnor U8253 (N_8253,N_8149,N_8046);
nor U8254 (N_8254,N_8131,N_8023);
and U8255 (N_8255,N_8158,N_8113);
nor U8256 (N_8256,N_8160,N_8075);
xor U8257 (N_8257,N_8213,N_8217);
nor U8258 (N_8258,N_8206,N_8030);
nand U8259 (N_8259,N_8226,N_8190);
and U8260 (N_8260,N_8133,N_8114);
or U8261 (N_8261,N_8056,N_8007);
nand U8262 (N_8262,N_8045,N_8001);
and U8263 (N_8263,N_8037,N_8130);
xor U8264 (N_8264,N_8016,N_8197);
or U8265 (N_8265,N_8135,N_8151);
xnor U8266 (N_8266,N_8044,N_8048);
or U8267 (N_8267,N_8145,N_8193);
or U8268 (N_8268,N_8186,N_8202);
or U8269 (N_8269,N_8050,N_8214);
and U8270 (N_8270,N_8146,N_8248);
nor U8271 (N_8271,N_8153,N_8087);
xor U8272 (N_8272,N_8054,N_8142);
xor U8273 (N_8273,N_8010,N_8168);
xnor U8274 (N_8274,N_8165,N_8052);
or U8275 (N_8275,N_8116,N_8127);
or U8276 (N_8276,N_8065,N_8161);
and U8277 (N_8277,N_8000,N_8204);
and U8278 (N_8278,N_8096,N_8148);
nand U8279 (N_8279,N_8195,N_8123);
xnor U8280 (N_8280,N_8015,N_8067);
nor U8281 (N_8281,N_8072,N_8024);
or U8282 (N_8282,N_8141,N_8107);
xor U8283 (N_8283,N_8063,N_8053);
and U8284 (N_8284,N_8109,N_8042);
or U8285 (N_8285,N_8021,N_8064);
nand U8286 (N_8286,N_8079,N_8180);
xnor U8287 (N_8287,N_8220,N_8118);
nand U8288 (N_8288,N_8208,N_8147);
xnor U8289 (N_8289,N_8237,N_8035);
or U8290 (N_8290,N_8081,N_8150);
nand U8291 (N_8291,N_8101,N_8051);
and U8292 (N_8292,N_8122,N_8120);
xnor U8293 (N_8293,N_8209,N_8012);
nor U8294 (N_8294,N_8084,N_8091);
xor U8295 (N_8295,N_8144,N_8232);
and U8296 (N_8296,N_8152,N_8013);
or U8297 (N_8297,N_8031,N_8178);
xor U8298 (N_8298,N_8156,N_8032);
nand U8299 (N_8299,N_8225,N_8242);
nor U8300 (N_8300,N_8028,N_8134);
nand U8301 (N_8301,N_8119,N_8216);
or U8302 (N_8302,N_8092,N_8103);
or U8303 (N_8303,N_8177,N_8246);
nand U8304 (N_8304,N_8061,N_8174);
or U8305 (N_8305,N_8157,N_8179);
nand U8306 (N_8306,N_8059,N_8243);
and U8307 (N_8307,N_8229,N_8058);
nand U8308 (N_8308,N_8020,N_8117);
xnor U8309 (N_8309,N_8078,N_8018);
nand U8310 (N_8310,N_8201,N_8019);
xor U8311 (N_8311,N_8223,N_8100);
or U8312 (N_8312,N_8139,N_8191);
or U8313 (N_8313,N_8060,N_8200);
and U8314 (N_8314,N_8004,N_8138);
or U8315 (N_8315,N_8094,N_8057);
or U8316 (N_8316,N_8073,N_8184);
xor U8317 (N_8317,N_8227,N_8047);
and U8318 (N_8318,N_8108,N_8083);
xor U8319 (N_8319,N_8222,N_8187);
nor U8320 (N_8320,N_8086,N_8155);
and U8321 (N_8321,N_8173,N_8231);
or U8322 (N_8322,N_8136,N_8090);
and U8323 (N_8323,N_8125,N_8106);
xnor U8324 (N_8324,N_8185,N_8172);
nand U8325 (N_8325,N_8115,N_8234);
nor U8326 (N_8326,N_8163,N_8039);
xnor U8327 (N_8327,N_8011,N_8068);
or U8328 (N_8328,N_8128,N_8017);
and U8329 (N_8329,N_8183,N_8049);
nor U8330 (N_8330,N_8203,N_8236);
nand U8331 (N_8331,N_8169,N_8027);
nand U8332 (N_8332,N_8082,N_8196);
and U8333 (N_8333,N_8080,N_8009);
or U8334 (N_8334,N_8062,N_8167);
xor U8335 (N_8335,N_8181,N_8110);
xor U8336 (N_8336,N_8102,N_8014);
nand U8337 (N_8337,N_8249,N_8228);
nor U8338 (N_8338,N_8171,N_8224);
nand U8339 (N_8339,N_8126,N_8245);
nor U8340 (N_8340,N_8071,N_8112);
and U8341 (N_8341,N_8198,N_8188);
nor U8342 (N_8342,N_8003,N_8239);
xnor U8343 (N_8343,N_8170,N_8137);
nand U8344 (N_8344,N_8212,N_8207);
xnor U8345 (N_8345,N_8033,N_8066);
or U8346 (N_8346,N_8069,N_8192);
and U8347 (N_8347,N_8182,N_8132);
nor U8348 (N_8348,N_8041,N_8055);
and U8349 (N_8349,N_8205,N_8247);
or U8350 (N_8350,N_8029,N_8240);
nor U8351 (N_8351,N_8238,N_8219);
nor U8352 (N_8352,N_8194,N_8221);
xor U8353 (N_8353,N_8043,N_8121);
nor U8354 (N_8354,N_8124,N_8233);
nor U8355 (N_8355,N_8005,N_8025);
xor U8356 (N_8356,N_8006,N_8143);
nand U8357 (N_8357,N_8022,N_8077);
xor U8358 (N_8358,N_8230,N_8085);
and U8359 (N_8359,N_8154,N_8199);
nand U8360 (N_8360,N_8215,N_8176);
and U8361 (N_8361,N_8099,N_8036);
nor U8362 (N_8362,N_8162,N_8097);
xor U8363 (N_8363,N_8140,N_8093);
nand U8364 (N_8364,N_8210,N_8111);
nor U8365 (N_8365,N_8189,N_8088);
xnor U8366 (N_8366,N_8089,N_8076);
and U8367 (N_8367,N_8026,N_8008);
nor U8368 (N_8368,N_8244,N_8105);
or U8369 (N_8369,N_8159,N_8095);
xnor U8370 (N_8370,N_8040,N_8218);
and U8371 (N_8371,N_8211,N_8164);
and U8372 (N_8372,N_8166,N_8034);
and U8373 (N_8373,N_8241,N_8098);
nor U8374 (N_8374,N_8104,N_8175);
nand U8375 (N_8375,N_8137,N_8025);
nor U8376 (N_8376,N_8168,N_8190);
or U8377 (N_8377,N_8096,N_8185);
nand U8378 (N_8378,N_8064,N_8177);
or U8379 (N_8379,N_8179,N_8015);
and U8380 (N_8380,N_8169,N_8069);
nor U8381 (N_8381,N_8228,N_8019);
xnor U8382 (N_8382,N_8193,N_8056);
and U8383 (N_8383,N_8098,N_8057);
and U8384 (N_8384,N_8010,N_8103);
and U8385 (N_8385,N_8141,N_8046);
nor U8386 (N_8386,N_8009,N_8135);
xor U8387 (N_8387,N_8205,N_8103);
nor U8388 (N_8388,N_8003,N_8231);
xor U8389 (N_8389,N_8181,N_8050);
nor U8390 (N_8390,N_8144,N_8191);
nand U8391 (N_8391,N_8151,N_8105);
and U8392 (N_8392,N_8129,N_8031);
and U8393 (N_8393,N_8003,N_8009);
and U8394 (N_8394,N_8121,N_8202);
nor U8395 (N_8395,N_8063,N_8047);
and U8396 (N_8396,N_8199,N_8183);
nand U8397 (N_8397,N_8004,N_8077);
or U8398 (N_8398,N_8054,N_8122);
nand U8399 (N_8399,N_8199,N_8064);
xnor U8400 (N_8400,N_8047,N_8178);
or U8401 (N_8401,N_8064,N_8186);
xnor U8402 (N_8402,N_8167,N_8133);
nand U8403 (N_8403,N_8096,N_8169);
xnor U8404 (N_8404,N_8132,N_8063);
nand U8405 (N_8405,N_8017,N_8066);
or U8406 (N_8406,N_8095,N_8016);
nand U8407 (N_8407,N_8143,N_8137);
xnor U8408 (N_8408,N_8133,N_8168);
and U8409 (N_8409,N_8204,N_8202);
nand U8410 (N_8410,N_8036,N_8222);
xor U8411 (N_8411,N_8108,N_8032);
nand U8412 (N_8412,N_8101,N_8156);
nor U8413 (N_8413,N_8129,N_8155);
xnor U8414 (N_8414,N_8210,N_8047);
or U8415 (N_8415,N_8026,N_8088);
nor U8416 (N_8416,N_8111,N_8154);
xnor U8417 (N_8417,N_8227,N_8237);
xnor U8418 (N_8418,N_8079,N_8166);
xor U8419 (N_8419,N_8090,N_8203);
nor U8420 (N_8420,N_8166,N_8189);
and U8421 (N_8421,N_8224,N_8010);
nor U8422 (N_8422,N_8133,N_8072);
nor U8423 (N_8423,N_8090,N_8165);
nor U8424 (N_8424,N_8206,N_8200);
nor U8425 (N_8425,N_8028,N_8152);
nand U8426 (N_8426,N_8075,N_8098);
nand U8427 (N_8427,N_8196,N_8025);
or U8428 (N_8428,N_8219,N_8046);
or U8429 (N_8429,N_8193,N_8158);
nand U8430 (N_8430,N_8235,N_8161);
nor U8431 (N_8431,N_8034,N_8030);
or U8432 (N_8432,N_8239,N_8180);
or U8433 (N_8433,N_8058,N_8225);
or U8434 (N_8434,N_8065,N_8194);
nor U8435 (N_8435,N_8100,N_8027);
nor U8436 (N_8436,N_8154,N_8180);
or U8437 (N_8437,N_8213,N_8206);
nor U8438 (N_8438,N_8148,N_8204);
nor U8439 (N_8439,N_8062,N_8031);
nand U8440 (N_8440,N_8161,N_8114);
nand U8441 (N_8441,N_8097,N_8017);
xor U8442 (N_8442,N_8220,N_8215);
nor U8443 (N_8443,N_8172,N_8131);
and U8444 (N_8444,N_8044,N_8099);
nor U8445 (N_8445,N_8198,N_8124);
xnor U8446 (N_8446,N_8001,N_8216);
and U8447 (N_8447,N_8212,N_8200);
or U8448 (N_8448,N_8114,N_8149);
nor U8449 (N_8449,N_8239,N_8006);
or U8450 (N_8450,N_8196,N_8042);
nand U8451 (N_8451,N_8181,N_8216);
xnor U8452 (N_8452,N_8053,N_8030);
and U8453 (N_8453,N_8079,N_8164);
nand U8454 (N_8454,N_8028,N_8195);
or U8455 (N_8455,N_8164,N_8012);
and U8456 (N_8456,N_8155,N_8173);
or U8457 (N_8457,N_8046,N_8022);
or U8458 (N_8458,N_8018,N_8086);
or U8459 (N_8459,N_8137,N_8053);
xor U8460 (N_8460,N_8058,N_8050);
and U8461 (N_8461,N_8144,N_8075);
xnor U8462 (N_8462,N_8186,N_8021);
nand U8463 (N_8463,N_8045,N_8130);
and U8464 (N_8464,N_8046,N_8021);
nand U8465 (N_8465,N_8090,N_8053);
or U8466 (N_8466,N_8065,N_8090);
xnor U8467 (N_8467,N_8189,N_8012);
xor U8468 (N_8468,N_8062,N_8037);
or U8469 (N_8469,N_8040,N_8069);
nand U8470 (N_8470,N_8164,N_8043);
nand U8471 (N_8471,N_8056,N_8167);
xor U8472 (N_8472,N_8135,N_8187);
nor U8473 (N_8473,N_8112,N_8166);
and U8474 (N_8474,N_8227,N_8185);
nor U8475 (N_8475,N_8017,N_8161);
xor U8476 (N_8476,N_8005,N_8020);
xnor U8477 (N_8477,N_8071,N_8223);
and U8478 (N_8478,N_8213,N_8185);
and U8479 (N_8479,N_8180,N_8139);
nor U8480 (N_8480,N_8242,N_8021);
nand U8481 (N_8481,N_8233,N_8165);
nor U8482 (N_8482,N_8146,N_8066);
xor U8483 (N_8483,N_8079,N_8002);
nand U8484 (N_8484,N_8104,N_8155);
nor U8485 (N_8485,N_8151,N_8166);
and U8486 (N_8486,N_8015,N_8111);
and U8487 (N_8487,N_8092,N_8016);
nand U8488 (N_8488,N_8234,N_8101);
nor U8489 (N_8489,N_8000,N_8081);
and U8490 (N_8490,N_8095,N_8085);
nand U8491 (N_8491,N_8094,N_8065);
or U8492 (N_8492,N_8033,N_8003);
and U8493 (N_8493,N_8079,N_8019);
or U8494 (N_8494,N_8138,N_8058);
nand U8495 (N_8495,N_8214,N_8148);
xnor U8496 (N_8496,N_8055,N_8218);
and U8497 (N_8497,N_8078,N_8032);
or U8498 (N_8498,N_8016,N_8045);
and U8499 (N_8499,N_8123,N_8235);
nor U8500 (N_8500,N_8267,N_8467);
and U8501 (N_8501,N_8383,N_8262);
nand U8502 (N_8502,N_8310,N_8324);
xnor U8503 (N_8503,N_8285,N_8353);
nor U8504 (N_8504,N_8462,N_8389);
xnor U8505 (N_8505,N_8459,N_8322);
nor U8506 (N_8506,N_8306,N_8347);
or U8507 (N_8507,N_8356,N_8369);
xnor U8508 (N_8508,N_8361,N_8295);
xnor U8509 (N_8509,N_8445,N_8435);
or U8510 (N_8510,N_8354,N_8349);
xor U8511 (N_8511,N_8357,N_8482);
nand U8512 (N_8512,N_8301,N_8374);
nand U8513 (N_8513,N_8478,N_8392);
or U8514 (N_8514,N_8496,N_8279);
xnor U8515 (N_8515,N_8486,N_8377);
and U8516 (N_8516,N_8391,N_8469);
and U8517 (N_8517,N_8373,N_8323);
nand U8518 (N_8518,N_8280,N_8408);
nand U8519 (N_8519,N_8390,N_8458);
or U8520 (N_8520,N_8457,N_8316);
xnor U8521 (N_8521,N_8474,N_8471);
nor U8522 (N_8522,N_8343,N_8406);
xnor U8523 (N_8523,N_8437,N_8481);
or U8524 (N_8524,N_8433,N_8276);
nand U8525 (N_8525,N_8363,N_8325);
and U8526 (N_8526,N_8410,N_8272);
xnor U8527 (N_8527,N_8455,N_8485);
nand U8528 (N_8528,N_8450,N_8460);
or U8529 (N_8529,N_8387,N_8345);
and U8530 (N_8530,N_8335,N_8362);
and U8531 (N_8531,N_8344,N_8275);
nor U8532 (N_8532,N_8328,N_8380);
or U8533 (N_8533,N_8261,N_8329);
nand U8534 (N_8534,N_8398,N_8254);
xor U8535 (N_8535,N_8400,N_8307);
xnor U8536 (N_8536,N_8304,N_8427);
and U8537 (N_8537,N_8303,N_8465);
and U8538 (N_8538,N_8309,N_8271);
nand U8539 (N_8539,N_8340,N_8250);
or U8540 (N_8540,N_8413,N_8265);
nor U8541 (N_8541,N_8479,N_8281);
nand U8542 (N_8542,N_8430,N_8404);
or U8543 (N_8543,N_8268,N_8299);
and U8544 (N_8544,N_8424,N_8302);
or U8545 (N_8545,N_8346,N_8257);
and U8546 (N_8546,N_8263,N_8417);
xnor U8547 (N_8547,N_8376,N_8282);
xnor U8548 (N_8548,N_8290,N_8399);
or U8549 (N_8549,N_8422,N_8348);
and U8550 (N_8550,N_8315,N_8423);
and U8551 (N_8551,N_8494,N_8456);
xnor U8552 (N_8552,N_8296,N_8498);
nand U8553 (N_8553,N_8490,N_8350);
nor U8554 (N_8554,N_8468,N_8421);
and U8555 (N_8555,N_8414,N_8431);
and U8556 (N_8556,N_8405,N_8330);
nand U8557 (N_8557,N_8293,N_8397);
and U8558 (N_8558,N_8440,N_8446);
and U8559 (N_8559,N_8360,N_8379);
xor U8560 (N_8560,N_8388,N_8256);
nor U8561 (N_8561,N_8463,N_8341);
xor U8562 (N_8562,N_8278,N_8451);
nand U8563 (N_8563,N_8407,N_8333);
and U8564 (N_8564,N_8251,N_8339);
or U8565 (N_8565,N_8365,N_8375);
and U8566 (N_8566,N_8452,N_8402);
and U8567 (N_8567,N_8447,N_8409);
or U8568 (N_8568,N_8491,N_8338);
nor U8569 (N_8569,N_8286,N_8370);
or U8570 (N_8570,N_8252,N_8497);
or U8571 (N_8571,N_8300,N_8264);
and U8572 (N_8572,N_8411,N_8274);
and U8573 (N_8573,N_8284,N_8288);
and U8574 (N_8574,N_8326,N_8308);
nand U8575 (N_8575,N_8493,N_8294);
xnor U8576 (N_8576,N_8342,N_8253);
and U8577 (N_8577,N_8287,N_8386);
and U8578 (N_8578,N_8311,N_8283);
or U8579 (N_8579,N_8359,N_8475);
nand U8580 (N_8580,N_8327,N_8461);
and U8581 (N_8581,N_8378,N_8260);
or U8582 (N_8582,N_8319,N_8438);
and U8583 (N_8583,N_8298,N_8443);
nand U8584 (N_8584,N_8434,N_8368);
xnor U8585 (N_8585,N_8403,N_8499);
nor U8586 (N_8586,N_8332,N_8255);
and U8587 (N_8587,N_8489,N_8289);
nor U8588 (N_8588,N_8305,N_8381);
xnor U8589 (N_8589,N_8367,N_8384);
xnor U8590 (N_8590,N_8396,N_8395);
nand U8591 (N_8591,N_8312,N_8416);
or U8592 (N_8592,N_8259,N_8321);
nand U8593 (N_8593,N_8415,N_8320);
nor U8594 (N_8594,N_8436,N_8495);
xor U8595 (N_8595,N_8426,N_8382);
xnor U8596 (N_8596,N_8472,N_8292);
xnor U8597 (N_8597,N_8476,N_8366);
nand U8598 (N_8598,N_8466,N_8355);
and U8599 (N_8599,N_8492,N_8394);
or U8600 (N_8600,N_8334,N_8331);
and U8601 (N_8601,N_8444,N_8258);
nand U8602 (N_8602,N_8266,N_8483);
nor U8603 (N_8603,N_8432,N_8439);
xnor U8604 (N_8604,N_8425,N_8297);
xnor U8605 (N_8605,N_8270,N_8358);
or U8606 (N_8606,N_8372,N_8449);
or U8607 (N_8607,N_8441,N_8420);
nor U8608 (N_8608,N_8336,N_8453);
and U8609 (N_8609,N_8412,N_8454);
or U8610 (N_8610,N_8273,N_8269);
and U8611 (N_8611,N_8442,N_8488);
nand U8612 (N_8612,N_8371,N_8364);
nor U8613 (N_8613,N_8464,N_8480);
and U8614 (N_8614,N_8448,N_8313);
or U8615 (N_8615,N_8393,N_8418);
xor U8616 (N_8616,N_8352,N_8351);
nand U8617 (N_8617,N_8337,N_8385);
or U8618 (N_8618,N_8317,N_8291);
or U8619 (N_8619,N_8428,N_8473);
and U8620 (N_8620,N_8401,N_8477);
xor U8621 (N_8621,N_8419,N_8314);
and U8622 (N_8622,N_8484,N_8318);
and U8623 (N_8623,N_8277,N_8429);
nor U8624 (N_8624,N_8470,N_8487);
or U8625 (N_8625,N_8445,N_8293);
and U8626 (N_8626,N_8471,N_8264);
xor U8627 (N_8627,N_8431,N_8380);
nor U8628 (N_8628,N_8416,N_8335);
or U8629 (N_8629,N_8331,N_8303);
nor U8630 (N_8630,N_8314,N_8258);
xor U8631 (N_8631,N_8439,N_8312);
xnor U8632 (N_8632,N_8476,N_8376);
xnor U8633 (N_8633,N_8480,N_8308);
and U8634 (N_8634,N_8375,N_8296);
or U8635 (N_8635,N_8461,N_8443);
xor U8636 (N_8636,N_8492,N_8250);
and U8637 (N_8637,N_8447,N_8434);
nand U8638 (N_8638,N_8399,N_8440);
nor U8639 (N_8639,N_8356,N_8321);
nor U8640 (N_8640,N_8257,N_8472);
and U8641 (N_8641,N_8381,N_8300);
xor U8642 (N_8642,N_8362,N_8319);
nor U8643 (N_8643,N_8496,N_8282);
xnor U8644 (N_8644,N_8308,N_8438);
and U8645 (N_8645,N_8425,N_8466);
or U8646 (N_8646,N_8276,N_8457);
xor U8647 (N_8647,N_8419,N_8345);
nand U8648 (N_8648,N_8322,N_8282);
or U8649 (N_8649,N_8347,N_8363);
nor U8650 (N_8650,N_8271,N_8299);
nand U8651 (N_8651,N_8457,N_8283);
nand U8652 (N_8652,N_8250,N_8408);
and U8653 (N_8653,N_8329,N_8356);
nand U8654 (N_8654,N_8341,N_8258);
nand U8655 (N_8655,N_8310,N_8449);
nand U8656 (N_8656,N_8280,N_8267);
nor U8657 (N_8657,N_8400,N_8387);
and U8658 (N_8658,N_8470,N_8381);
or U8659 (N_8659,N_8256,N_8489);
or U8660 (N_8660,N_8317,N_8496);
nand U8661 (N_8661,N_8315,N_8365);
nand U8662 (N_8662,N_8294,N_8464);
xor U8663 (N_8663,N_8350,N_8437);
and U8664 (N_8664,N_8343,N_8399);
or U8665 (N_8665,N_8386,N_8379);
nand U8666 (N_8666,N_8326,N_8415);
nand U8667 (N_8667,N_8273,N_8404);
xor U8668 (N_8668,N_8409,N_8450);
nand U8669 (N_8669,N_8255,N_8399);
nand U8670 (N_8670,N_8344,N_8414);
nor U8671 (N_8671,N_8460,N_8252);
or U8672 (N_8672,N_8464,N_8276);
nor U8673 (N_8673,N_8259,N_8436);
nor U8674 (N_8674,N_8313,N_8270);
and U8675 (N_8675,N_8423,N_8416);
and U8676 (N_8676,N_8433,N_8345);
and U8677 (N_8677,N_8479,N_8374);
and U8678 (N_8678,N_8277,N_8347);
nor U8679 (N_8679,N_8345,N_8280);
nor U8680 (N_8680,N_8373,N_8308);
or U8681 (N_8681,N_8484,N_8488);
xnor U8682 (N_8682,N_8376,N_8357);
nand U8683 (N_8683,N_8448,N_8401);
xnor U8684 (N_8684,N_8375,N_8347);
nor U8685 (N_8685,N_8403,N_8498);
nand U8686 (N_8686,N_8436,N_8362);
xnor U8687 (N_8687,N_8301,N_8273);
nor U8688 (N_8688,N_8430,N_8332);
nor U8689 (N_8689,N_8369,N_8287);
or U8690 (N_8690,N_8418,N_8326);
and U8691 (N_8691,N_8299,N_8432);
nor U8692 (N_8692,N_8444,N_8488);
and U8693 (N_8693,N_8392,N_8283);
and U8694 (N_8694,N_8326,N_8306);
nand U8695 (N_8695,N_8495,N_8473);
and U8696 (N_8696,N_8333,N_8285);
or U8697 (N_8697,N_8300,N_8337);
or U8698 (N_8698,N_8262,N_8459);
nand U8699 (N_8699,N_8441,N_8320);
nor U8700 (N_8700,N_8494,N_8394);
xnor U8701 (N_8701,N_8288,N_8388);
or U8702 (N_8702,N_8497,N_8305);
xor U8703 (N_8703,N_8393,N_8498);
or U8704 (N_8704,N_8342,N_8454);
nor U8705 (N_8705,N_8327,N_8407);
nor U8706 (N_8706,N_8300,N_8484);
xnor U8707 (N_8707,N_8364,N_8328);
and U8708 (N_8708,N_8375,N_8440);
nor U8709 (N_8709,N_8427,N_8389);
and U8710 (N_8710,N_8296,N_8388);
nor U8711 (N_8711,N_8409,N_8426);
or U8712 (N_8712,N_8274,N_8298);
xor U8713 (N_8713,N_8268,N_8450);
xnor U8714 (N_8714,N_8274,N_8427);
and U8715 (N_8715,N_8265,N_8276);
nor U8716 (N_8716,N_8305,N_8464);
and U8717 (N_8717,N_8345,N_8489);
xnor U8718 (N_8718,N_8435,N_8262);
or U8719 (N_8719,N_8327,N_8455);
or U8720 (N_8720,N_8480,N_8409);
or U8721 (N_8721,N_8252,N_8487);
nor U8722 (N_8722,N_8457,N_8272);
xor U8723 (N_8723,N_8482,N_8282);
nand U8724 (N_8724,N_8270,N_8347);
and U8725 (N_8725,N_8421,N_8458);
and U8726 (N_8726,N_8434,N_8264);
nand U8727 (N_8727,N_8353,N_8487);
or U8728 (N_8728,N_8306,N_8458);
nand U8729 (N_8729,N_8458,N_8462);
nor U8730 (N_8730,N_8296,N_8319);
xor U8731 (N_8731,N_8408,N_8344);
nand U8732 (N_8732,N_8326,N_8358);
nand U8733 (N_8733,N_8433,N_8327);
xor U8734 (N_8734,N_8286,N_8272);
nor U8735 (N_8735,N_8378,N_8393);
or U8736 (N_8736,N_8424,N_8364);
and U8737 (N_8737,N_8272,N_8344);
and U8738 (N_8738,N_8380,N_8295);
nor U8739 (N_8739,N_8289,N_8390);
xor U8740 (N_8740,N_8272,N_8255);
nor U8741 (N_8741,N_8310,N_8412);
or U8742 (N_8742,N_8325,N_8434);
or U8743 (N_8743,N_8341,N_8486);
nor U8744 (N_8744,N_8260,N_8488);
xor U8745 (N_8745,N_8458,N_8378);
or U8746 (N_8746,N_8297,N_8453);
or U8747 (N_8747,N_8465,N_8367);
nand U8748 (N_8748,N_8310,N_8430);
and U8749 (N_8749,N_8364,N_8354);
and U8750 (N_8750,N_8698,N_8638);
nand U8751 (N_8751,N_8648,N_8603);
or U8752 (N_8752,N_8609,N_8588);
or U8753 (N_8753,N_8580,N_8735);
or U8754 (N_8754,N_8724,N_8667);
nor U8755 (N_8755,N_8688,N_8645);
nor U8756 (N_8756,N_8662,N_8519);
xor U8757 (N_8757,N_8591,N_8517);
nand U8758 (N_8758,N_8722,N_8652);
or U8759 (N_8759,N_8614,N_8738);
nor U8760 (N_8760,N_8598,N_8727);
nor U8761 (N_8761,N_8681,N_8550);
nor U8762 (N_8762,N_8547,N_8716);
nand U8763 (N_8763,N_8587,N_8546);
or U8764 (N_8764,N_8538,N_8739);
xor U8765 (N_8765,N_8533,N_8705);
nor U8766 (N_8766,N_8637,N_8683);
nand U8767 (N_8767,N_8695,N_8567);
or U8768 (N_8768,N_8551,N_8701);
nand U8769 (N_8769,N_8711,N_8647);
nand U8770 (N_8770,N_8685,N_8513);
nor U8771 (N_8771,N_8526,N_8624);
nor U8772 (N_8772,N_8694,N_8534);
nor U8773 (N_8773,N_8635,N_8561);
and U8774 (N_8774,N_8541,N_8634);
nand U8775 (N_8775,N_8682,N_8617);
or U8776 (N_8776,N_8602,N_8625);
nor U8777 (N_8777,N_8516,N_8610);
and U8778 (N_8778,N_8572,N_8560);
or U8779 (N_8779,N_8657,N_8573);
and U8780 (N_8780,N_8743,N_8696);
and U8781 (N_8781,N_8619,N_8578);
nor U8782 (N_8782,N_8510,N_8712);
nor U8783 (N_8783,N_8726,N_8502);
or U8784 (N_8784,N_8514,N_8639);
xor U8785 (N_8785,N_8655,N_8713);
xnor U8786 (N_8786,N_8564,N_8720);
or U8787 (N_8787,N_8706,N_8545);
xnor U8788 (N_8788,N_8595,N_8656);
or U8789 (N_8789,N_8605,N_8626);
and U8790 (N_8790,N_8693,N_8710);
and U8791 (N_8791,N_8697,N_8521);
xnor U8792 (N_8792,N_8568,N_8554);
nor U8793 (N_8793,N_8737,N_8660);
and U8794 (N_8794,N_8615,N_8601);
or U8795 (N_8795,N_8552,N_8562);
or U8796 (N_8796,N_8632,N_8718);
nand U8797 (N_8797,N_8542,N_8641);
nand U8798 (N_8798,N_8576,N_8671);
or U8799 (N_8799,N_8721,N_8649);
and U8800 (N_8800,N_8748,N_8673);
and U8801 (N_8801,N_8644,N_8725);
and U8802 (N_8802,N_8708,N_8537);
nand U8803 (N_8803,N_8563,N_8640);
nand U8804 (N_8804,N_8627,N_8575);
nand U8805 (N_8805,N_8666,N_8599);
xor U8806 (N_8806,N_8663,N_8672);
nor U8807 (N_8807,N_8523,N_8642);
nor U8808 (N_8808,N_8529,N_8643);
nand U8809 (N_8809,N_8679,N_8636);
xnor U8810 (N_8810,N_8553,N_8584);
nand U8811 (N_8811,N_8661,N_8525);
nand U8812 (N_8812,N_8539,N_8717);
xnor U8813 (N_8813,N_8675,N_8629);
nand U8814 (N_8814,N_8507,N_8571);
xnor U8815 (N_8815,N_8594,N_8628);
xnor U8816 (N_8816,N_8719,N_8596);
xnor U8817 (N_8817,N_8749,N_8506);
nand U8818 (N_8818,N_8549,N_8618);
xnor U8819 (N_8819,N_8590,N_8616);
or U8820 (N_8820,N_8728,N_8723);
and U8821 (N_8821,N_8565,N_8503);
or U8822 (N_8822,N_8544,N_8518);
xor U8823 (N_8823,N_8597,N_8703);
and U8824 (N_8824,N_8524,N_8742);
nand U8825 (N_8825,N_8585,N_8579);
and U8826 (N_8826,N_8633,N_8511);
xnor U8827 (N_8827,N_8670,N_8566);
and U8828 (N_8828,N_8620,N_8592);
or U8829 (N_8829,N_8669,N_8570);
xnor U8830 (N_8830,N_8500,N_8650);
nand U8831 (N_8831,N_8715,N_8678);
or U8832 (N_8832,N_8622,N_8582);
and U8833 (N_8833,N_8548,N_8687);
nand U8834 (N_8834,N_8532,N_8508);
and U8835 (N_8835,N_8677,N_8606);
or U8836 (N_8836,N_8556,N_8736);
and U8837 (N_8837,N_8714,N_8522);
xnor U8838 (N_8838,N_8630,N_8680);
nand U8839 (N_8839,N_8691,N_8515);
nor U8840 (N_8840,N_8528,N_8654);
xnor U8841 (N_8841,N_8540,N_8668);
and U8842 (N_8842,N_8690,N_8707);
xor U8843 (N_8843,N_8505,N_8658);
xor U8844 (N_8844,N_8709,N_8689);
and U8845 (N_8845,N_8729,N_8699);
nand U8846 (N_8846,N_8745,N_8593);
nor U8847 (N_8847,N_8577,N_8744);
and U8848 (N_8848,N_8520,N_8730);
nor U8849 (N_8849,N_8686,N_8608);
xnor U8850 (N_8850,N_8530,N_8734);
nor U8851 (N_8851,N_8581,N_8527);
and U8852 (N_8852,N_8574,N_8512);
or U8853 (N_8853,N_8557,N_8704);
or U8854 (N_8854,N_8611,N_8676);
nand U8855 (N_8855,N_8535,N_8731);
xor U8856 (N_8856,N_8674,N_8558);
nor U8857 (N_8857,N_8586,N_8659);
and U8858 (N_8858,N_8631,N_8589);
nand U8859 (N_8859,N_8733,N_8607);
or U8860 (N_8860,N_8653,N_8600);
nand U8861 (N_8861,N_8536,N_8741);
and U8862 (N_8862,N_8555,N_8700);
xnor U8863 (N_8863,N_8651,N_8665);
or U8864 (N_8864,N_8684,N_8702);
nor U8865 (N_8865,N_8531,N_8732);
or U8866 (N_8866,N_8692,N_8746);
and U8867 (N_8867,N_8543,N_8740);
or U8868 (N_8868,N_8509,N_8646);
nor U8869 (N_8869,N_8621,N_8559);
and U8870 (N_8870,N_8747,N_8613);
nand U8871 (N_8871,N_8612,N_8623);
or U8872 (N_8872,N_8504,N_8664);
or U8873 (N_8873,N_8583,N_8569);
or U8874 (N_8874,N_8604,N_8501);
nand U8875 (N_8875,N_8500,N_8656);
xor U8876 (N_8876,N_8540,N_8544);
nand U8877 (N_8877,N_8728,N_8680);
xnor U8878 (N_8878,N_8615,N_8530);
nor U8879 (N_8879,N_8703,N_8606);
and U8880 (N_8880,N_8581,N_8588);
nand U8881 (N_8881,N_8610,N_8714);
nand U8882 (N_8882,N_8577,N_8641);
nor U8883 (N_8883,N_8629,N_8748);
and U8884 (N_8884,N_8689,N_8738);
or U8885 (N_8885,N_8725,N_8555);
nor U8886 (N_8886,N_8549,N_8520);
xor U8887 (N_8887,N_8717,N_8719);
or U8888 (N_8888,N_8724,N_8577);
nor U8889 (N_8889,N_8741,N_8684);
or U8890 (N_8890,N_8590,N_8703);
nand U8891 (N_8891,N_8665,N_8682);
xor U8892 (N_8892,N_8639,N_8572);
and U8893 (N_8893,N_8613,N_8542);
and U8894 (N_8894,N_8612,N_8748);
xor U8895 (N_8895,N_8535,N_8563);
nor U8896 (N_8896,N_8647,N_8539);
nor U8897 (N_8897,N_8707,N_8702);
nand U8898 (N_8898,N_8671,N_8610);
or U8899 (N_8899,N_8555,N_8593);
nand U8900 (N_8900,N_8728,N_8671);
or U8901 (N_8901,N_8681,N_8590);
nand U8902 (N_8902,N_8597,N_8515);
nand U8903 (N_8903,N_8624,N_8674);
xnor U8904 (N_8904,N_8672,N_8520);
or U8905 (N_8905,N_8503,N_8625);
xor U8906 (N_8906,N_8724,N_8545);
nand U8907 (N_8907,N_8515,N_8679);
or U8908 (N_8908,N_8624,N_8616);
nand U8909 (N_8909,N_8507,N_8623);
or U8910 (N_8910,N_8558,N_8603);
xnor U8911 (N_8911,N_8678,N_8503);
nand U8912 (N_8912,N_8542,N_8722);
xor U8913 (N_8913,N_8678,N_8567);
and U8914 (N_8914,N_8655,N_8656);
nor U8915 (N_8915,N_8549,N_8604);
and U8916 (N_8916,N_8552,N_8654);
and U8917 (N_8917,N_8745,N_8660);
and U8918 (N_8918,N_8718,N_8732);
xnor U8919 (N_8919,N_8589,N_8747);
or U8920 (N_8920,N_8676,N_8589);
xnor U8921 (N_8921,N_8571,N_8688);
xnor U8922 (N_8922,N_8733,N_8549);
nor U8923 (N_8923,N_8663,N_8701);
and U8924 (N_8924,N_8621,N_8640);
or U8925 (N_8925,N_8739,N_8653);
or U8926 (N_8926,N_8670,N_8568);
nand U8927 (N_8927,N_8538,N_8622);
nand U8928 (N_8928,N_8643,N_8718);
nor U8929 (N_8929,N_8737,N_8595);
and U8930 (N_8930,N_8528,N_8522);
and U8931 (N_8931,N_8698,N_8740);
and U8932 (N_8932,N_8665,N_8674);
nor U8933 (N_8933,N_8695,N_8706);
nor U8934 (N_8934,N_8544,N_8743);
nor U8935 (N_8935,N_8509,N_8545);
xnor U8936 (N_8936,N_8699,N_8686);
xor U8937 (N_8937,N_8692,N_8624);
xor U8938 (N_8938,N_8526,N_8521);
nor U8939 (N_8939,N_8526,N_8621);
nor U8940 (N_8940,N_8654,N_8725);
nor U8941 (N_8941,N_8708,N_8723);
nand U8942 (N_8942,N_8544,N_8708);
nand U8943 (N_8943,N_8706,N_8668);
xnor U8944 (N_8944,N_8510,N_8664);
or U8945 (N_8945,N_8709,N_8746);
nand U8946 (N_8946,N_8665,N_8695);
or U8947 (N_8947,N_8524,N_8622);
nand U8948 (N_8948,N_8530,N_8623);
nand U8949 (N_8949,N_8672,N_8535);
nand U8950 (N_8950,N_8555,N_8690);
or U8951 (N_8951,N_8556,N_8535);
xor U8952 (N_8952,N_8595,N_8630);
nand U8953 (N_8953,N_8538,N_8537);
and U8954 (N_8954,N_8523,N_8697);
xnor U8955 (N_8955,N_8653,N_8501);
nor U8956 (N_8956,N_8547,N_8619);
or U8957 (N_8957,N_8648,N_8643);
xnor U8958 (N_8958,N_8667,N_8704);
and U8959 (N_8959,N_8735,N_8720);
xnor U8960 (N_8960,N_8659,N_8748);
nand U8961 (N_8961,N_8515,N_8556);
xor U8962 (N_8962,N_8606,N_8660);
xor U8963 (N_8963,N_8712,N_8574);
or U8964 (N_8964,N_8659,N_8713);
nand U8965 (N_8965,N_8611,N_8626);
nand U8966 (N_8966,N_8719,N_8672);
or U8967 (N_8967,N_8745,N_8557);
nand U8968 (N_8968,N_8646,N_8555);
nor U8969 (N_8969,N_8742,N_8565);
nand U8970 (N_8970,N_8592,N_8577);
nor U8971 (N_8971,N_8558,N_8628);
nor U8972 (N_8972,N_8653,N_8737);
nor U8973 (N_8973,N_8695,N_8531);
and U8974 (N_8974,N_8513,N_8544);
nand U8975 (N_8975,N_8647,N_8740);
and U8976 (N_8976,N_8656,N_8616);
xnor U8977 (N_8977,N_8600,N_8694);
or U8978 (N_8978,N_8529,N_8543);
xor U8979 (N_8979,N_8566,N_8548);
xor U8980 (N_8980,N_8546,N_8601);
and U8981 (N_8981,N_8711,N_8527);
nand U8982 (N_8982,N_8591,N_8735);
nand U8983 (N_8983,N_8673,N_8694);
nand U8984 (N_8984,N_8718,N_8609);
nand U8985 (N_8985,N_8675,N_8573);
nand U8986 (N_8986,N_8729,N_8621);
nor U8987 (N_8987,N_8732,N_8641);
nand U8988 (N_8988,N_8641,N_8510);
nand U8989 (N_8989,N_8725,N_8590);
or U8990 (N_8990,N_8712,N_8728);
nand U8991 (N_8991,N_8710,N_8593);
or U8992 (N_8992,N_8518,N_8680);
xor U8993 (N_8993,N_8749,N_8541);
nor U8994 (N_8994,N_8696,N_8731);
nand U8995 (N_8995,N_8637,N_8737);
nor U8996 (N_8996,N_8731,N_8525);
nor U8997 (N_8997,N_8546,N_8612);
nand U8998 (N_8998,N_8700,N_8738);
nor U8999 (N_8999,N_8522,N_8716);
xor U9000 (N_9000,N_8953,N_8955);
xnor U9001 (N_9001,N_8789,N_8946);
nor U9002 (N_9002,N_8945,N_8813);
nand U9003 (N_9003,N_8897,N_8923);
or U9004 (N_9004,N_8832,N_8862);
xor U9005 (N_9005,N_8792,N_8755);
and U9006 (N_9006,N_8770,N_8973);
or U9007 (N_9007,N_8938,N_8825);
nand U9008 (N_9008,N_8970,N_8849);
xor U9009 (N_9009,N_8799,N_8936);
xor U9010 (N_9010,N_8848,N_8925);
nand U9011 (N_9011,N_8888,N_8989);
nand U9012 (N_9012,N_8758,N_8983);
xor U9013 (N_9013,N_8981,N_8948);
nand U9014 (N_9014,N_8884,N_8878);
xnor U9015 (N_9015,N_8778,N_8918);
and U9016 (N_9016,N_8971,N_8992);
or U9017 (N_9017,N_8837,N_8867);
nand U9018 (N_9018,N_8975,N_8805);
nand U9019 (N_9019,N_8829,N_8851);
xor U9020 (N_9020,N_8899,N_8987);
xnor U9021 (N_9021,N_8920,N_8937);
nand U9022 (N_9022,N_8869,N_8822);
nor U9023 (N_9023,N_8819,N_8927);
nand U9024 (N_9024,N_8828,N_8783);
and U9025 (N_9025,N_8787,N_8754);
nor U9026 (N_9026,N_8874,N_8919);
nor U9027 (N_9027,N_8908,N_8934);
xor U9028 (N_9028,N_8810,N_8785);
or U9029 (N_9029,N_8842,N_8904);
nand U9030 (N_9030,N_8894,N_8876);
nand U9031 (N_9031,N_8891,N_8944);
nor U9032 (N_9032,N_8980,N_8809);
or U9033 (N_9033,N_8976,N_8871);
nor U9034 (N_9034,N_8866,N_8863);
or U9035 (N_9035,N_8969,N_8850);
and U9036 (N_9036,N_8839,N_8759);
nor U9037 (N_9037,N_8926,N_8782);
nor U9038 (N_9038,N_8930,N_8966);
and U9039 (N_9039,N_8812,N_8830);
xor U9040 (N_9040,N_8816,N_8793);
xnor U9041 (N_9041,N_8988,N_8776);
nand U9042 (N_9042,N_8898,N_8803);
or U9043 (N_9043,N_8796,N_8751);
or U9044 (N_9044,N_8882,N_8913);
nand U9045 (N_9045,N_8996,N_8870);
and U9046 (N_9046,N_8774,N_8999);
or U9047 (N_9047,N_8942,N_8932);
or U9048 (N_9048,N_8772,N_8761);
xor U9049 (N_9049,N_8947,N_8967);
and U9050 (N_9050,N_8858,N_8826);
or U9051 (N_9051,N_8846,N_8784);
and U9052 (N_9052,N_8771,N_8833);
and U9053 (N_9053,N_8977,N_8814);
or U9054 (N_9054,N_8795,N_8941);
nand U9055 (N_9055,N_8963,N_8887);
and U9056 (N_9056,N_8997,N_8979);
nand U9057 (N_9057,N_8998,N_8921);
nand U9058 (N_9058,N_8857,N_8961);
nor U9059 (N_9059,N_8804,N_8959);
xnor U9060 (N_9060,N_8929,N_8956);
nand U9061 (N_9061,N_8911,N_8794);
nand U9062 (N_9062,N_8815,N_8924);
and U9063 (N_9063,N_8914,N_8843);
nand U9064 (N_9064,N_8905,N_8893);
or U9065 (N_9065,N_8972,N_8958);
nand U9066 (N_9066,N_8852,N_8982);
xnor U9067 (N_9067,N_8768,N_8917);
xnor U9068 (N_9068,N_8864,N_8800);
nand U9069 (N_9069,N_8844,N_8993);
and U9070 (N_9070,N_8957,N_8949);
nor U9071 (N_9071,N_8841,N_8818);
xnor U9072 (N_9072,N_8881,N_8964);
nor U9073 (N_9073,N_8877,N_8909);
nand U9074 (N_9074,N_8885,N_8788);
nand U9075 (N_9075,N_8994,N_8984);
xnor U9076 (N_9076,N_8817,N_8798);
xnor U9077 (N_9077,N_8875,N_8883);
or U9078 (N_9078,N_8950,N_8939);
and U9079 (N_9079,N_8859,N_8775);
or U9080 (N_9080,N_8797,N_8889);
and U9081 (N_9081,N_8780,N_8901);
nand U9082 (N_9082,N_8890,N_8868);
or U9083 (N_9083,N_8880,N_8808);
nor U9084 (N_9084,N_8892,N_8847);
and U9085 (N_9085,N_8886,N_8995);
xnor U9086 (N_9086,N_8763,N_8990);
or U9087 (N_9087,N_8786,N_8827);
nor U9088 (N_9088,N_8824,N_8991);
and U9089 (N_9089,N_8960,N_8855);
nor U9090 (N_9090,N_8757,N_8836);
nor U9091 (N_9091,N_8912,N_8802);
nor U9092 (N_9092,N_8974,N_8767);
nor U9093 (N_9093,N_8806,N_8766);
and U9094 (N_9094,N_8861,N_8952);
and U9095 (N_9095,N_8838,N_8860);
and U9096 (N_9096,N_8915,N_8845);
nand U9097 (N_9097,N_8962,N_8895);
or U9098 (N_9098,N_8965,N_8943);
nand U9099 (N_9099,N_8773,N_8823);
nand U9100 (N_9100,N_8873,N_8900);
and U9101 (N_9101,N_8807,N_8954);
or U9102 (N_9102,N_8896,N_8762);
or U9103 (N_9103,N_8801,N_8779);
and U9104 (N_9104,N_8986,N_8916);
nand U9105 (N_9105,N_8933,N_8907);
and U9106 (N_9106,N_8978,N_8854);
nor U9107 (N_9107,N_8811,N_8791);
nor U9108 (N_9108,N_8935,N_8750);
xnor U9109 (N_9109,N_8752,N_8902);
and U9110 (N_9110,N_8853,N_8756);
nor U9111 (N_9111,N_8831,N_8985);
or U9112 (N_9112,N_8760,N_8951);
or U9113 (N_9113,N_8856,N_8903);
and U9114 (N_9114,N_8821,N_8765);
or U9115 (N_9115,N_8835,N_8872);
nor U9116 (N_9116,N_8820,N_8840);
and U9117 (N_9117,N_8906,N_8910);
or U9118 (N_9118,N_8865,N_8931);
xnor U9119 (N_9119,N_8764,N_8834);
or U9120 (N_9120,N_8769,N_8928);
xnor U9121 (N_9121,N_8968,N_8879);
and U9122 (N_9122,N_8790,N_8922);
xnor U9123 (N_9123,N_8940,N_8777);
nand U9124 (N_9124,N_8781,N_8753);
and U9125 (N_9125,N_8931,N_8897);
nand U9126 (N_9126,N_8760,N_8922);
or U9127 (N_9127,N_8760,N_8782);
nor U9128 (N_9128,N_8829,N_8809);
nor U9129 (N_9129,N_8880,N_8782);
xor U9130 (N_9130,N_8907,N_8837);
xnor U9131 (N_9131,N_8833,N_8943);
xnor U9132 (N_9132,N_8825,N_8843);
nor U9133 (N_9133,N_8827,N_8763);
nor U9134 (N_9134,N_8979,N_8809);
and U9135 (N_9135,N_8786,N_8857);
nand U9136 (N_9136,N_8875,N_8852);
and U9137 (N_9137,N_8819,N_8788);
nand U9138 (N_9138,N_8771,N_8751);
nand U9139 (N_9139,N_8992,N_8809);
and U9140 (N_9140,N_8770,N_8870);
or U9141 (N_9141,N_8866,N_8893);
and U9142 (N_9142,N_8896,N_8993);
xor U9143 (N_9143,N_8932,N_8986);
and U9144 (N_9144,N_8996,N_8941);
or U9145 (N_9145,N_8937,N_8854);
nor U9146 (N_9146,N_8884,N_8902);
nand U9147 (N_9147,N_8890,N_8777);
xnor U9148 (N_9148,N_8936,N_8984);
nor U9149 (N_9149,N_8915,N_8806);
nor U9150 (N_9150,N_8956,N_8836);
nor U9151 (N_9151,N_8817,N_8884);
xor U9152 (N_9152,N_8824,N_8994);
xor U9153 (N_9153,N_8769,N_8964);
nor U9154 (N_9154,N_8865,N_8792);
xor U9155 (N_9155,N_8884,N_8932);
or U9156 (N_9156,N_8826,N_8913);
xor U9157 (N_9157,N_8799,N_8823);
or U9158 (N_9158,N_8949,N_8781);
xor U9159 (N_9159,N_8835,N_8888);
and U9160 (N_9160,N_8909,N_8967);
or U9161 (N_9161,N_8848,N_8999);
and U9162 (N_9162,N_8890,N_8983);
xnor U9163 (N_9163,N_8750,N_8888);
and U9164 (N_9164,N_8808,N_8806);
nand U9165 (N_9165,N_8869,N_8831);
and U9166 (N_9166,N_8864,N_8986);
xnor U9167 (N_9167,N_8838,N_8894);
xor U9168 (N_9168,N_8945,N_8929);
xor U9169 (N_9169,N_8997,N_8788);
nand U9170 (N_9170,N_8859,N_8951);
nand U9171 (N_9171,N_8979,N_8792);
xnor U9172 (N_9172,N_8965,N_8803);
or U9173 (N_9173,N_8870,N_8968);
xor U9174 (N_9174,N_8938,N_8787);
xnor U9175 (N_9175,N_8955,N_8922);
nor U9176 (N_9176,N_8876,N_8801);
xnor U9177 (N_9177,N_8792,N_8776);
xnor U9178 (N_9178,N_8954,N_8876);
xor U9179 (N_9179,N_8775,N_8999);
or U9180 (N_9180,N_8922,N_8985);
or U9181 (N_9181,N_8834,N_8938);
xnor U9182 (N_9182,N_8783,N_8762);
nor U9183 (N_9183,N_8883,N_8904);
xnor U9184 (N_9184,N_8989,N_8803);
nand U9185 (N_9185,N_8948,N_8755);
and U9186 (N_9186,N_8870,N_8956);
nand U9187 (N_9187,N_8889,N_8781);
or U9188 (N_9188,N_8766,N_8870);
or U9189 (N_9189,N_8849,N_8986);
xnor U9190 (N_9190,N_8884,N_8863);
nor U9191 (N_9191,N_8791,N_8774);
nand U9192 (N_9192,N_8778,N_8878);
and U9193 (N_9193,N_8941,N_8952);
nor U9194 (N_9194,N_8837,N_8899);
or U9195 (N_9195,N_8907,N_8883);
nor U9196 (N_9196,N_8983,N_8946);
or U9197 (N_9197,N_8903,N_8964);
xor U9198 (N_9198,N_8918,N_8827);
xor U9199 (N_9199,N_8834,N_8868);
or U9200 (N_9200,N_8843,N_8803);
xnor U9201 (N_9201,N_8789,N_8928);
nand U9202 (N_9202,N_8921,N_8969);
and U9203 (N_9203,N_8863,N_8869);
nand U9204 (N_9204,N_8998,N_8873);
and U9205 (N_9205,N_8829,N_8915);
or U9206 (N_9206,N_8950,N_8865);
xor U9207 (N_9207,N_8974,N_8933);
or U9208 (N_9208,N_8876,N_8870);
nand U9209 (N_9209,N_8882,N_8942);
xor U9210 (N_9210,N_8985,N_8767);
or U9211 (N_9211,N_8767,N_8950);
nor U9212 (N_9212,N_8853,N_8880);
xor U9213 (N_9213,N_8774,N_8866);
nand U9214 (N_9214,N_8845,N_8903);
nand U9215 (N_9215,N_8830,N_8834);
xor U9216 (N_9216,N_8984,N_8771);
and U9217 (N_9217,N_8856,N_8851);
or U9218 (N_9218,N_8769,N_8987);
or U9219 (N_9219,N_8782,N_8856);
nand U9220 (N_9220,N_8935,N_8964);
and U9221 (N_9221,N_8975,N_8790);
or U9222 (N_9222,N_8801,N_8822);
nor U9223 (N_9223,N_8847,N_8837);
nand U9224 (N_9224,N_8808,N_8774);
nand U9225 (N_9225,N_8754,N_8757);
or U9226 (N_9226,N_8762,N_8900);
xor U9227 (N_9227,N_8845,N_8764);
nand U9228 (N_9228,N_8980,N_8757);
nand U9229 (N_9229,N_8808,N_8895);
nand U9230 (N_9230,N_8923,N_8970);
nand U9231 (N_9231,N_8792,N_8808);
and U9232 (N_9232,N_8949,N_8761);
xor U9233 (N_9233,N_8824,N_8803);
or U9234 (N_9234,N_8947,N_8883);
xor U9235 (N_9235,N_8978,N_8866);
nand U9236 (N_9236,N_8845,N_8829);
xnor U9237 (N_9237,N_8927,N_8864);
and U9238 (N_9238,N_8973,N_8800);
and U9239 (N_9239,N_8852,N_8800);
nor U9240 (N_9240,N_8892,N_8787);
nor U9241 (N_9241,N_8778,N_8861);
and U9242 (N_9242,N_8821,N_8833);
or U9243 (N_9243,N_8954,N_8983);
xnor U9244 (N_9244,N_8918,N_8975);
or U9245 (N_9245,N_8984,N_8781);
nor U9246 (N_9246,N_8979,N_8782);
nor U9247 (N_9247,N_8925,N_8830);
nand U9248 (N_9248,N_8906,N_8914);
or U9249 (N_9249,N_8872,N_8830);
nand U9250 (N_9250,N_9024,N_9005);
or U9251 (N_9251,N_9177,N_9208);
nor U9252 (N_9252,N_9142,N_9109);
nand U9253 (N_9253,N_9118,N_9135);
nand U9254 (N_9254,N_9078,N_9096);
and U9255 (N_9255,N_9237,N_9000);
nor U9256 (N_9256,N_9161,N_9119);
nor U9257 (N_9257,N_9199,N_9094);
nand U9258 (N_9258,N_9011,N_9105);
or U9259 (N_9259,N_9056,N_9144);
and U9260 (N_9260,N_9092,N_9063);
and U9261 (N_9261,N_9107,N_9110);
and U9262 (N_9262,N_9185,N_9182);
nor U9263 (N_9263,N_9216,N_9245);
nand U9264 (N_9264,N_9085,N_9190);
nand U9265 (N_9265,N_9246,N_9018);
xnor U9266 (N_9266,N_9002,N_9089);
or U9267 (N_9267,N_9053,N_9115);
xor U9268 (N_9268,N_9202,N_9090);
nor U9269 (N_9269,N_9134,N_9131);
or U9270 (N_9270,N_9243,N_9223);
and U9271 (N_9271,N_9108,N_9219);
nand U9272 (N_9272,N_9066,N_9213);
and U9273 (N_9273,N_9062,N_9009);
xor U9274 (N_9274,N_9129,N_9174);
nand U9275 (N_9275,N_9151,N_9195);
xnor U9276 (N_9276,N_9097,N_9086);
xnor U9277 (N_9277,N_9212,N_9095);
or U9278 (N_9278,N_9079,N_9081);
or U9279 (N_9279,N_9031,N_9065);
nor U9280 (N_9280,N_9111,N_9075);
and U9281 (N_9281,N_9116,N_9047);
nor U9282 (N_9282,N_9167,N_9023);
xor U9283 (N_9283,N_9132,N_9193);
xor U9284 (N_9284,N_9046,N_9071);
or U9285 (N_9285,N_9013,N_9049);
and U9286 (N_9286,N_9206,N_9221);
xnor U9287 (N_9287,N_9186,N_9055);
and U9288 (N_9288,N_9020,N_9137);
nor U9289 (N_9289,N_9165,N_9088);
nand U9290 (N_9290,N_9189,N_9231);
or U9291 (N_9291,N_9001,N_9048);
and U9292 (N_9292,N_9117,N_9150);
nand U9293 (N_9293,N_9217,N_9042);
and U9294 (N_9294,N_9082,N_9247);
xnor U9295 (N_9295,N_9229,N_9008);
xnor U9296 (N_9296,N_9074,N_9010);
nand U9297 (N_9297,N_9139,N_9122);
nor U9298 (N_9298,N_9197,N_9239);
or U9299 (N_9299,N_9044,N_9033);
and U9300 (N_9300,N_9068,N_9136);
xor U9301 (N_9301,N_9210,N_9163);
nor U9302 (N_9302,N_9228,N_9224);
and U9303 (N_9303,N_9158,N_9032);
and U9304 (N_9304,N_9160,N_9077);
and U9305 (N_9305,N_9026,N_9232);
nor U9306 (N_9306,N_9021,N_9192);
and U9307 (N_9307,N_9125,N_9244);
nor U9308 (N_9308,N_9249,N_9155);
xor U9309 (N_9309,N_9015,N_9181);
nand U9310 (N_9310,N_9169,N_9054);
or U9311 (N_9311,N_9133,N_9104);
nand U9312 (N_9312,N_9146,N_9016);
nand U9313 (N_9313,N_9162,N_9043);
or U9314 (N_9314,N_9130,N_9183);
or U9315 (N_9315,N_9187,N_9112);
or U9316 (N_9316,N_9236,N_9200);
nand U9317 (N_9317,N_9178,N_9076);
xor U9318 (N_9318,N_9204,N_9027);
nand U9319 (N_9319,N_9087,N_9203);
nor U9320 (N_9320,N_9149,N_9173);
and U9321 (N_9321,N_9205,N_9194);
nor U9322 (N_9322,N_9198,N_9050);
nand U9323 (N_9323,N_9113,N_9060);
and U9324 (N_9324,N_9017,N_9226);
and U9325 (N_9325,N_9099,N_9179);
nand U9326 (N_9326,N_9022,N_9093);
or U9327 (N_9327,N_9128,N_9240);
or U9328 (N_9328,N_9038,N_9220);
and U9329 (N_9329,N_9123,N_9138);
nand U9330 (N_9330,N_9171,N_9126);
nand U9331 (N_9331,N_9103,N_9188);
or U9332 (N_9332,N_9045,N_9121);
nand U9333 (N_9333,N_9234,N_9170);
xnor U9334 (N_9334,N_9004,N_9242);
nand U9335 (N_9335,N_9176,N_9153);
or U9336 (N_9336,N_9030,N_9083);
xnor U9337 (N_9337,N_9148,N_9012);
nor U9338 (N_9338,N_9057,N_9218);
nor U9339 (N_9339,N_9145,N_9070);
and U9340 (N_9340,N_9003,N_9102);
nand U9341 (N_9341,N_9191,N_9230);
nor U9342 (N_9342,N_9064,N_9124);
nor U9343 (N_9343,N_9114,N_9152);
xor U9344 (N_9344,N_9052,N_9209);
nand U9345 (N_9345,N_9073,N_9039);
nand U9346 (N_9346,N_9215,N_9147);
xor U9347 (N_9347,N_9225,N_9059);
nor U9348 (N_9348,N_9007,N_9157);
nor U9349 (N_9349,N_9248,N_9069);
and U9350 (N_9350,N_9154,N_9025);
nand U9351 (N_9351,N_9241,N_9091);
and U9352 (N_9352,N_9201,N_9072);
nor U9353 (N_9353,N_9006,N_9040);
xnor U9354 (N_9354,N_9196,N_9159);
and U9355 (N_9355,N_9061,N_9214);
nor U9356 (N_9356,N_9175,N_9166);
nor U9357 (N_9357,N_9227,N_9235);
and U9358 (N_9358,N_9098,N_9051);
and U9359 (N_9359,N_9067,N_9164);
or U9360 (N_9360,N_9041,N_9035);
and U9361 (N_9361,N_9034,N_9233);
or U9362 (N_9362,N_9084,N_9222);
nand U9363 (N_9363,N_9036,N_9211);
nor U9364 (N_9364,N_9058,N_9037);
and U9365 (N_9365,N_9080,N_9156);
nand U9366 (N_9366,N_9029,N_9238);
and U9367 (N_9367,N_9014,N_9207);
or U9368 (N_9368,N_9120,N_9141);
xnor U9369 (N_9369,N_9172,N_9101);
nor U9370 (N_9370,N_9180,N_9168);
nand U9371 (N_9371,N_9019,N_9140);
or U9372 (N_9372,N_9106,N_9143);
and U9373 (N_9373,N_9127,N_9100);
and U9374 (N_9374,N_9028,N_9184);
nand U9375 (N_9375,N_9058,N_9170);
nor U9376 (N_9376,N_9246,N_9085);
nand U9377 (N_9377,N_9198,N_9243);
nor U9378 (N_9378,N_9186,N_9172);
xor U9379 (N_9379,N_9247,N_9132);
and U9380 (N_9380,N_9211,N_9106);
nor U9381 (N_9381,N_9114,N_9086);
or U9382 (N_9382,N_9004,N_9164);
and U9383 (N_9383,N_9147,N_9036);
nand U9384 (N_9384,N_9117,N_9201);
nor U9385 (N_9385,N_9192,N_9120);
xor U9386 (N_9386,N_9182,N_9136);
nor U9387 (N_9387,N_9170,N_9150);
and U9388 (N_9388,N_9094,N_9151);
or U9389 (N_9389,N_9119,N_9136);
and U9390 (N_9390,N_9141,N_9031);
or U9391 (N_9391,N_9085,N_9220);
nor U9392 (N_9392,N_9217,N_9027);
nor U9393 (N_9393,N_9242,N_9117);
xor U9394 (N_9394,N_9187,N_9199);
nor U9395 (N_9395,N_9164,N_9175);
nor U9396 (N_9396,N_9054,N_9151);
nor U9397 (N_9397,N_9046,N_9154);
and U9398 (N_9398,N_9046,N_9211);
xor U9399 (N_9399,N_9083,N_9191);
nor U9400 (N_9400,N_9084,N_9064);
nand U9401 (N_9401,N_9001,N_9173);
xnor U9402 (N_9402,N_9188,N_9161);
nor U9403 (N_9403,N_9176,N_9220);
xor U9404 (N_9404,N_9237,N_9002);
xnor U9405 (N_9405,N_9167,N_9085);
nand U9406 (N_9406,N_9111,N_9201);
nand U9407 (N_9407,N_9161,N_9089);
and U9408 (N_9408,N_9027,N_9041);
or U9409 (N_9409,N_9182,N_9042);
nand U9410 (N_9410,N_9036,N_9175);
nor U9411 (N_9411,N_9129,N_9218);
nor U9412 (N_9412,N_9246,N_9135);
xnor U9413 (N_9413,N_9154,N_9115);
and U9414 (N_9414,N_9181,N_9109);
nand U9415 (N_9415,N_9063,N_9122);
nor U9416 (N_9416,N_9185,N_9067);
nor U9417 (N_9417,N_9015,N_9222);
nor U9418 (N_9418,N_9234,N_9185);
nor U9419 (N_9419,N_9031,N_9056);
and U9420 (N_9420,N_9128,N_9107);
nor U9421 (N_9421,N_9248,N_9053);
or U9422 (N_9422,N_9118,N_9143);
and U9423 (N_9423,N_9138,N_9019);
nand U9424 (N_9424,N_9178,N_9148);
nand U9425 (N_9425,N_9000,N_9112);
nor U9426 (N_9426,N_9142,N_9223);
or U9427 (N_9427,N_9172,N_9056);
and U9428 (N_9428,N_9152,N_9190);
nor U9429 (N_9429,N_9028,N_9062);
xor U9430 (N_9430,N_9224,N_9065);
or U9431 (N_9431,N_9050,N_9060);
xnor U9432 (N_9432,N_9087,N_9120);
nand U9433 (N_9433,N_9008,N_9219);
and U9434 (N_9434,N_9138,N_9107);
xnor U9435 (N_9435,N_9084,N_9121);
nand U9436 (N_9436,N_9185,N_9055);
or U9437 (N_9437,N_9223,N_9047);
and U9438 (N_9438,N_9215,N_9003);
nand U9439 (N_9439,N_9108,N_9202);
and U9440 (N_9440,N_9155,N_9058);
xnor U9441 (N_9441,N_9122,N_9196);
xnor U9442 (N_9442,N_9101,N_9116);
nor U9443 (N_9443,N_9028,N_9010);
or U9444 (N_9444,N_9135,N_9117);
and U9445 (N_9445,N_9088,N_9119);
nor U9446 (N_9446,N_9139,N_9064);
xor U9447 (N_9447,N_9026,N_9066);
xnor U9448 (N_9448,N_9163,N_9048);
or U9449 (N_9449,N_9151,N_9249);
nor U9450 (N_9450,N_9179,N_9248);
nor U9451 (N_9451,N_9244,N_9013);
or U9452 (N_9452,N_9196,N_9029);
or U9453 (N_9453,N_9246,N_9205);
nand U9454 (N_9454,N_9161,N_9021);
nand U9455 (N_9455,N_9179,N_9050);
and U9456 (N_9456,N_9228,N_9149);
xor U9457 (N_9457,N_9051,N_9010);
and U9458 (N_9458,N_9117,N_9070);
nor U9459 (N_9459,N_9094,N_9177);
xor U9460 (N_9460,N_9109,N_9212);
or U9461 (N_9461,N_9072,N_9191);
or U9462 (N_9462,N_9206,N_9145);
xor U9463 (N_9463,N_9070,N_9009);
and U9464 (N_9464,N_9133,N_9213);
xor U9465 (N_9465,N_9086,N_9048);
nand U9466 (N_9466,N_9133,N_9175);
nor U9467 (N_9467,N_9107,N_9017);
xor U9468 (N_9468,N_9111,N_9016);
and U9469 (N_9469,N_9042,N_9192);
nor U9470 (N_9470,N_9239,N_9133);
or U9471 (N_9471,N_9072,N_9079);
and U9472 (N_9472,N_9222,N_9149);
nand U9473 (N_9473,N_9026,N_9141);
xnor U9474 (N_9474,N_9146,N_9086);
or U9475 (N_9475,N_9129,N_9064);
or U9476 (N_9476,N_9205,N_9207);
nand U9477 (N_9477,N_9158,N_9065);
xnor U9478 (N_9478,N_9146,N_9066);
nand U9479 (N_9479,N_9107,N_9160);
xor U9480 (N_9480,N_9144,N_9214);
or U9481 (N_9481,N_9202,N_9235);
nand U9482 (N_9482,N_9242,N_9134);
nor U9483 (N_9483,N_9078,N_9188);
nor U9484 (N_9484,N_9156,N_9032);
xor U9485 (N_9485,N_9137,N_9088);
nor U9486 (N_9486,N_9097,N_9126);
and U9487 (N_9487,N_9059,N_9088);
or U9488 (N_9488,N_9245,N_9069);
or U9489 (N_9489,N_9176,N_9196);
and U9490 (N_9490,N_9135,N_9245);
and U9491 (N_9491,N_9141,N_9103);
and U9492 (N_9492,N_9202,N_9077);
nor U9493 (N_9493,N_9060,N_9109);
xor U9494 (N_9494,N_9204,N_9008);
xnor U9495 (N_9495,N_9219,N_9207);
xnor U9496 (N_9496,N_9006,N_9106);
and U9497 (N_9497,N_9244,N_9015);
and U9498 (N_9498,N_9105,N_9179);
nor U9499 (N_9499,N_9034,N_9176);
xor U9500 (N_9500,N_9313,N_9375);
nor U9501 (N_9501,N_9455,N_9438);
nand U9502 (N_9502,N_9323,N_9333);
nor U9503 (N_9503,N_9339,N_9409);
or U9504 (N_9504,N_9273,N_9349);
nand U9505 (N_9505,N_9487,N_9454);
nand U9506 (N_9506,N_9382,N_9472);
nor U9507 (N_9507,N_9256,N_9496);
and U9508 (N_9508,N_9378,N_9254);
and U9509 (N_9509,N_9396,N_9327);
or U9510 (N_9510,N_9316,N_9367);
nor U9511 (N_9511,N_9253,N_9473);
and U9512 (N_9512,N_9440,N_9425);
or U9513 (N_9513,N_9419,N_9450);
nor U9514 (N_9514,N_9366,N_9486);
nand U9515 (N_9515,N_9309,N_9312);
xnor U9516 (N_9516,N_9481,N_9439);
and U9517 (N_9517,N_9457,N_9497);
and U9518 (N_9518,N_9337,N_9255);
nor U9519 (N_9519,N_9281,N_9494);
and U9520 (N_9520,N_9374,N_9342);
xor U9521 (N_9521,N_9403,N_9401);
and U9522 (N_9522,N_9356,N_9263);
nor U9523 (N_9523,N_9391,N_9357);
or U9524 (N_9524,N_9354,N_9371);
or U9525 (N_9525,N_9428,N_9365);
xor U9526 (N_9526,N_9474,N_9379);
nor U9527 (N_9527,N_9271,N_9402);
nand U9528 (N_9528,N_9362,N_9293);
or U9529 (N_9529,N_9329,N_9251);
and U9530 (N_9530,N_9288,N_9390);
xnor U9531 (N_9531,N_9338,N_9261);
nand U9532 (N_9532,N_9360,N_9277);
or U9533 (N_9533,N_9319,N_9389);
and U9534 (N_9534,N_9314,N_9465);
nor U9535 (N_9535,N_9305,N_9344);
or U9536 (N_9536,N_9355,N_9431);
nand U9537 (N_9537,N_9284,N_9377);
nor U9538 (N_9538,N_9274,N_9317);
or U9539 (N_9539,N_9423,N_9266);
or U9540 (N_9540,N_9296,N_9446);
nor U9541 (N_9541,N_9257,N_9410);
nor U9542 (N_9542,N_9348,N_9321);
nand U9543 (N_9543,N_9453,N_9491);
and U9544 (N_9544,N_9399,N_9262);
xor U9545 (N_9545,N_9426,N_9299);
nor U9546 (N_9546,N_9372,N_9370);
or U9547 (N_9547,N_9435,N_9437);
nor U9548 (N_9548,N_9275,N_9413);
and U9549 (N_9549,N_9298,N_9373);
xnor U9550 (N_9550,N_9482,N_9480);
and U9551 (N_9551,N_9477,N_9363);
nand U9552 (N_9552,N_9458,N_9405);
nor U9553 (N_9553,N_9272,N_9325);
xor U9554 (N_9554,N_9304,N_9485);
nor U9555 (N_9555,N_9394,N_9442);
xor U9556 (N_9556,N_9259,N_9301);
and U9557 (N_9557,N_9387,N_9369);
nor U9558 (N_9558,N_9295,N_9290);
nor U9559 (N_9559,N_9286,N_9311);
nand U9560 (N_9560,N_9269,N_9483);
nor U9561 (N_9561,N_9397,N_9398);
xnor U9562 (N_9562,N_9408,N_9278);
nand U9563 (N_9563,N_9383,N_9441);
nand U9564 (N_9564,N_9350,N_9459);
xor U9565 (N_9565,N_9452,N_9386);
nand U9566 (N_9566,N_9451,N_9420);
nor U9567 (N_9567,N_9490,N_9267);
nor U9568 (N_9568,N_9411,N_9404);
nand U9569 (N_9569,N_9447,N_9292);
or U9570 (N_9570,N_9385,N_9331);
or U9571 (N_9571,N_9388,N_9334);
or U9572 (N_9572,N_9471,N_9318);
nand U9573 (N_9573,N_9466,N_9392);
xor U9574 (N_9574,N_9358,N_9421);
nand U9575 (N_9575,N_9467,N_9484);
nand U9576 (N_9576,N_9489,N_9340);
xor U9577 (N_9577,N_9282,N_9265);
or U9578 (N_9578,N_9315,N_9361);
xor U9579 (N_9579,N_9499,N_9456);
nand U9580 (N_9580,N_9332,N_9308);
xor U9581 (N_9581,N_9444,N_9406);
xnor U9582 (N_9582,N_9297,N_9343);
and U9583 (N_9583,N_9488,N_9280);
or U9584 (N_9584,N_9407,N_9336);
and U9585 (N_9585,N_9364,N_9498);
nor U9586 (N_9586,N_9307,N_9368);
nor U9587 (N_9587,N_9463,N_9433);
or U9588 (N_9588,N_9470,N_9341);
nor U9589 (N_9589,N_9283,N_9449);
or U9590 (N_9590,N_9434,N_9381);
xor U9591 (N_9591,N_9264,N_9351);
or U9592 (N_9592,N_9276,N_9335);
nand U9593 (N_9593,N_9279,N_9306);
xnor U9594 (N_9594,N_9395,N_9476);
nand U9595 (N_9595,N_9414,N_9352);
nor U9596 (N_9596,N_9478,N_9424);
nand U9597 (N_9597,N_9422,N_9287);
xnor U9598 (N_9598,N_9479,N_9427);
or U9599 (N_9599,N_9436,N_9418);
nor U9600 (N_9600,N_9291,N_9464);
nand U9601 (N_9601,N_9400,N_9416);
nor U9602 (N_9602,N_9322,N_9324);
xnor U9603 (N_9603,N_9330,N_9300);
xnor U9604 (N_9604,N_9415,N_9493);
and U9605 (N_9605,N_9492,N_9495);
xor U9606 (N_9606,N_9268,N_9320);
or U9607 (N_9607,N_9468,N_9285);
nand U9608 (N_9608,N_9376,N_9302);
xnor U9609 (N_9609,N_9475,N_9260);
and U9610 (N_9610,N_9443,N_9384);
xnor U9611 (N_9611,N_9310,N_9294);
or U9612 (N_9612,N_9252,N_9412);
or U9613 (N_9613,N_9347,N_9462);
xor U9614 (N_9614,N_9432,N_9417);
nor U9615 (N_9615,N_9469,N_9445);
and U9616 (N_9616,N_9353,N_9289);
and U9617 (N_9617,N_9448,N_9380);
or U9618 (N_9618,N_9303,N_9430);
nor U9619 (N_9619,N_9429,N_9460);
nand U9620 (N_9620,N_9326,N_9328);
xnor U9621 (N_9621,N_9258,N_9359);
and U9622 (N_9622,N_9250,N_9270);
and U9623 (N_9623,N_9345,N_9393);
xor U9624 (N_9624,N_9461,N_9346);
or U9625 (N_9625,N_9326,N_9300);
or U9626 (N_9626,N_9276,N_9359);
or U9627 (N_9627,N_9421,N_9495);
and U9628 (N_9628,N_9352,N_9293);
nor U9629 (N_9629,N_9258,N_9364);
and U9630 (N_9630,N_9409,N_9393);
and U9631 (N_9631,N_9388,N_9259);
nor U9632 (N_9632,N_9442,N_9365);
xnor U9633 (N_9633,N_9378,N_9337);
nand U9634 (N_9634,N_9296,N_9434);
nor U9635 (N_9635,N_9272,N_9469);
and U9636 (N_9636,N_9410,N_9255);
or U9637 (N_9637,N_9322,N_9424);
and U9638 (N_9638,N_9367,N_9477);
nor U9639 (N_9639,N_9307,N_9277);
nor U9640 (N_9640,N_9373,N_9350);
xor U9641 (N_9641,N_9436,N_9467);
nor U9642 (N_9642,N_9412,N_9369);
and U9643 (N_9643,N_9411,N_9373);
xnor U9644 (N_9644,N_9267,N_9252);
nor U9645 (N_9645,N_9462,N_9455);
nand U9646 (N_9646,N_9408,N_9391);
nor U9647 (N_9647,N_9449,N_9466);
nor U9648 (N_9648,N_9252,N_9288);
nand U9649 (N_9649,N_9432,N_9478);
xnor U9650 (N_9650,N_9389,N_9342);
xnor U9651 (N_9651,N_9263,N_9467);
nor U9652 (N_9652,N_9253,N_9316);
nand U9653 (N_9653,N_9496,N_9264);
xor U9654 (N_9654,N_9444,N_9458);
or U9655 (N_9655,N_9262,N_9459);
xnor U9656 (N_9656,N_9453,N_9338);
nand U9657 (N_9657,N_9284,N_9426);
or U9658 (N_9658,N_9372,N_9307);
nor U9659 (N_9659,N_9276,N_9319);
xor U9660 (N_9660,N_9316,N_9353);
or U9661 (N_9661,N_9346,N_9359);
nand U9662 (N_9662,N_9466,N_9379);
and U9663 (N_9663,N_9384,N_9379);
or U9664 (N_9664,N_9261,N_9440);
nand U9665 (N_9665,N_9445,N_9479);
and U9666 (N_9666,N_9285,N_9387);
and U9667 (N_9667,N_9415,N_9323);
nor U9668 (N_9668,N_9349,N_9329);
xnor U9669 (N_9669,N_9280,N_9406);
nor U9670 (N_9670,N_9321,N_9334);
or U9671 (N_9671,N_9354,N_9471);
nand U9672 (N_9672,N_9370,N_9400);
or U9673 (N_9673,N_9358,N_9363);
xnor U9674 (N_9674,N_9459,N_9411);
xnor U9675 (N_9675,N_9350,N_9337);
nand U9676 (N_9676,N_9439,N_9295);
xnor U9677 (N_9677,N_9381,N_9302);
and U9678 (N_9678,N_9397,N_9442);
and U9679 (N_9679,N_9335,N_9449);
and U9680 (N_9680,N_9334,N_9418);
and U9681 (N_9681,N_9476,N_9313);
nand U9682 (N_9682,N_9313,N_9278);
or U9683 (N_9683,N_9258,N_9316);
nand U9684 (N_9684,N_9473,N_9427);
or U9685 (N_9685,N_9405,N_9417);
or U9686 (N_9686,N_9360,N_9274);
or U9687 (N_9687,N_9446,N_9455);
nor U9688 (N_9688,N_9493,N_9354);
nor U9689 (N_9689,N_9291,N_9340);
nor U9690 (N_9690,N_9416,N_9277);
nor U9691 (N_9691,N_9344,N_9343);
and U9692 (N_9692,N_9293,N_9375);
xnor U9693 (N_9693,N_9487,N_9273);
nor U9694 (N_9694,N_9352,N_9436);
or U9695 (N_9695,N_9340,N_9313);
and U9696 (N_9696,N_9423,N_9441);
nand U9697 (N_9697,N_9309,N_9466);
nand U9698 (N_9698,N_9344,N_9378);
or U9699 (N_9699,N_9476,N_9255);
nor U9700 (N_9700,N_9447,N_9493);
and U9701 (N_9701,N_9267,N_9464);
xnor U9702 (N_9702,N_9325,N_9311);
and U9703 (N_9703,N_9450,N_9411);
xnor U9704 (N_9704,N_9498,N_9297);
nor U9705 (N_9705,N_9484,N_9387);
nand U9706 (N_9706,N_9455,N_9449);
nand U9707 (N_9707,N_9297,N_9272);
nand U9708 (N_9708,N_9250,N_9417);
and U9709 (N_9709,N_9306,N_9392);
nor U9710 (N_9710,N_9404,N_9492);
xnor U9711 (N_9711,N_9476,N_9388);
or U9712 (N_9712,N_9261,N_9466);
or U9713 (N_9713,N_9467,N_9424);
nand U9714 (N_9714,N_9280,N_9443);
nor U9715 (N_9715,N_9469,N_9396);
nor U9716 (N_9716,N_9348,N_9487);
nor U9717 (N_9717,N_9313,N_9321);
or U9718 (N_9718,N_9291,N_9351);
nor U9719 (N_9719,N_9349,N_9482);
xor U9720 (N_9720,N_9485,N_9268);
nand U9721 (N_9721,N_9265,N_9340);
or U9722 (N_9722,N_9444,N_9466);
xor U9723 (N_9723,N_9385,N_9369);
and U9724 (N_9724,N_9491,N_9314);
or U9725 (N_9725,N_9393,N_9334);
xor U9726 (N_9726,N_9367,N_9360);
nor U9727 (N_9727,N_9497,N_9292);
nand U9728 (N_9728,N_9341,N_9396);
xor U9729 (N_9729,N_9252,N_9369);
or U9730 (N_9730,N_9420,N_9496);
or U9731 (N_9731,N_9411,N_9318);
or U9732 (N_9732,N_9403,N_9347);
nand U9733 (N_9733,N_9380,N_9278);
and U9734 (N_9734,N_9477,N_9300);
nand U9735 (N_9735,N_9408,N_9479);
nand U9736 (N_9736,N_9331,N_9267);
xor U9737 (N_9737,N_9380,N_9459);
and U9738 (N_9738,N_9345,N_9480);
nor U9739 (N_9739,N_9269,N_9352);
nor U9740 (N_9740,N_9277,N_9427);
nor U9741 (N_9741,N_9333,N_9376);
and U9742 (N_9742,N_9382,N_9431);
or U9743 (N_9743,N_9489,N_9445);
and U9744 (N_9744,N_9490,N_9270);
or U9745 (N_9745,N_9381,N_9478);
nor U9746 (N_9746,N_9492,N_9354);
or U9747 (N_9747,N_9422,N_9274);
nand U9748 (N_9748,N_9426,N_9371);
nor U9749 (N_9749,N_9411,N_9417);
nor U9750 (N_9750,N_9728,N_9546);
nand U9751 (N_9751,N_9740,N_9540);
and U9752 (N_9752,N_9696,N_9517);
or U9753 (N_9753,N_9605,N_9744);
xor U9754 (N_9754,N_9746,N_9619);
and U9755 (N_9755,N_9661,N_9691);
nor U9756 (N_9756,N_9622,N_9577);
nor U9757 (N_9757,N_9646,N_9555);
nor U9758 (N_9758,N_9738,N_9736);
and U9759 (N_9759,N_9557,N_9719);
and U9760 (N_9760,N_9668,N_9552);
or U9761 (N_9761,N_9588,N_9548);
nor U9762 (N_9762,N_9521,N_9582);
nand U9763 (N_9763,N_9504,N_9604);
xor U9764 (N_9764,N_9595,N_9730);
or U9765 (N_9765,N_9729,N_9589);
or U9766 (N_9766,N_9702,N_9614);
nor U9767 (N_9767,N_9524,N_9710);
and U9768 (N_9768,N_9683,N_9623);
or U9769 (N_9769,N_9749,N_9655);
nor U9770 (N_9770,N_9695,N_9525);
nand U9771 (N_9771,N_9535,N_9585);
or U9772 (N_9772,N_9732,N_9628);
or U9773 (N_9773,N_9648,N_9579);
and U9774 (N_9774,N_9505,N_9583);
xor U9775 (N_9775,N_9694,N_9603);
nor U9776 (N_9776,N_9624,N_9539);
nor U9777 (N_9777,N_9608,N_9671);
nor U9778 (N_9778,N_9503,N_9739);
nor U9779 (N_9779,N_9592,N_9533);
or U9780 (N_9780,N_9613,N_9530);
nand U9781 (N_9781,N_9742,N_9572);
or U9782 (N_9782,N_9641,N_9669);
nand U9783 (N_9783,N_9692,N_9645);
and U9784 (N_9784,N_9593,N_9637);
nand U9785 (N_9785,N_9570,N_9534);
nor U9786 (N_9786,N_9680,N_9610);
xor U9787 (N_9787,N_9629,N_9647);
nor U9788 (N_9788,N_9515,N_9650);
nand U9789 (N_9789,N_9700,N_9649);
or U9790 (N_9790,N_9586,N_9529);
nand U9791 (N_9791,N_9507,N_9576);
nor U9792 (N_9792,N_9639,N_9725);
xnor U9793 (N_9793,N_9541,N_9707);
xor U9794 (N_9794,N_9676,N_9634);
and U9795 (N_9795,N_9745,N_9667);
nor U9796 (N_9796,N_9544,N_9545);
or U9797 (N_9797,N_9554,N_9712);
or U9798 (N_9798,N_9558,N_9727);
and U9799 (N_9799,N_9550,N_9704);
nor U9800 (N_9800,N_9563,N_9510);
nor U9801 (N_9801,N_9713,N_9711);
and U9802 (N_9802,N_9726,N_9620);
and U9803 (N_9803,N_9717,N_9596);
and U9804 (N_9804,N_9573,N_9528);
nor U9805 (N_9805,N_9615,N_9748);
xnor U9806 (N_9806,N_9594,N_9574);
nand U9807 (N_9807,N_9684,N_9735);
nand U9808 (N_9808,N_9658,N_9724);
or U9809 (N_9809,N_9666,N_9512);
xor U9810 (N_9810,N_9643,N_9502);
or U9811 (N_9811,N_9743,N_9638);
or U9812 (N_9812,N_9537,N_9686);
or U9813 (N_9813,N_9568,N_9723);
nand U9814 (N_9814,N_9578,N_9602);
xor U9815 (N_9815,N_9531,N_9630);
xor U9816 (N_9816,N_9697,N_9714);
xor U9817 (N_9817,N_9690,N_9653);
nor U9818 (N_9818,N_9681,N_9564);
nor U9819 (N_9819,N_9560,N_9642);
nand U9820 (N_9820,N_9553,N_9705);
xnor U9821 (N_9821,N_9543,N_9616);
and U9822 (N_9822,N_9556,N_9571);
or U9823 (N_9823,N_9536,N_9685);
and U9824 (N_9824,N_9565,N_9514);
or U9825 (N_9825,N_9532,N_9654);
or U9826 (N_9826,N_9609,N_9513);
nand U9827 (N_9827,N_9689,N_9584);
xnor U9828 (N_9828,N_9509,N_9741);
nand U9829 (N_9829,N_9617,N_9734);
and U9830 (N_9830,N_9567,N_9551);
or U9831 (N_9831,N_9611,N_9698);
or U9832 (N_9832,N_9511,N_9597);
nand U9833 (N_9833,N_9652,N_9670);
nand U9834 (N_9834,N_9518,N_9591);
nand U9835 (N_9835,N_9651,N_9635);
and U9836 (N_9836,N_9660,N_9720);
xnor U9837 (N_9837,N_9612,N_9519);
and U9838 (N_9838,N_9547,N_9715);
and U9839 (N_9839,N_9674,N_9506);
nand U9840 (N_9840,N_9699,N_9598);
and U9841 (N_9841,N_9662,N_9632);
and U9842 (N_9842,N_9644,N_9500);
or U9843 (N_9843,N_9561,N_9527);
or U9844 (N_9844,N_9562,N_9523);
nand U9845 (N_9845,N_9747,N_9657);
or U9846 (N_9846,N_9587,N_9633);
nand U9847 (N_9847,N_9607,N_9520);
xnor U9848 (N_9848,N_9678,N_9542);
xor U9849 (N_9849,N_9627,N_9693);
nand U9850 (N_9850,N_9731,N_9631);
or U9851 (N_9851,N_9709,N_9590);
and U9852 (N_9852,N_9675,N_9664);
nand U9853 (N_9853,N_9640,N_9508);
or U9854 (N_9854,N_9737,N_9716);
and U9855 (N_9855,N_9621,N_9625);
nand U9856 (N_9856,N_9501,N_9663);
nand U9857 (N_9857,N_9687,N_9706);
and U9858 (N_9858,N_9703,N_9600);
or U9859 (N_9859,N_9626,N_9559);
nor U9860 (N_9860,N_9708,N_9718);
or U9861 (N_9861,N_9580,N_9526);
nand U9862 (N_9862,N_9516,N_9722);
nand U9863 (N_9863,N_9701,N_9659);
xor U9864 (N_9864,N_9656,N_9679);
and U9865 (N_9865,N_9601,N_9538);
nand U9866 (N_9866,N_9549,N_9682);
nor U9867 (N_9867,N_9688,N_9733);
nor U9868 (N_9868,N_9581,N_9599);
nor U9869 (N_9869,N_9665,N_9575);
or U9870 (N_9870,N_9522,N_9606);
nand U9871 (N_9871,N_9721,N_9569);
or U9872 (N_9872,N_9677,N_9618);
nand U9873 (N_9873,N_9636,N_9672);
and U9874 (N_9874,N_9566,N_9673);
and U9875 (N_9875,N_9697,N_9568);
nand U9876 (N_9876,N_9609,N_9706);
nand U9877 (N_9877,N_9741,N_9645);
nor U9878 (N_9878,N_9744,N_9535);
or U9879 (N_9879,N_9553,N_9573);
and U9880 (N_9880,N_9520,N_9703);
xor U9881 (N_9881,N_9579,N_9635);
and U9882 (N_9882,N_9719,N_9682);
xnor U9883 (N_9883,N_9524,N_9684);
nand U9884 (N_9884,N_9617,N_9607);
xnor U9885 (N_9885,N_9691,N_9610);
nor U9886 (N_9886,N_9629,N_9543);
or U9887 (N_9887,N_9564,N_9650);
and U9888 (N_9888,N_9565,N_9595);
nand U9889 (N_9889,N_9518,N_9744);
nand U9890 (N_9890,N_9609,N_9543);
xnor U9891 (N_9891,N_9519,N_9614);
and U9892 (N_9892,N_9650,N_9605);
nor U9893 (N_9893,N_9710,N_9501);
xor U9894 (N_9894,N_9615,N_9504);
or U9895 (N_9895,N_9598,N_9734);
or U9896 (N_9896,N_9642,N_9635);
xor U9897 (N_9897,N_9505,N_9563);
and U9898 (N_9898,N_9740,N_9601);
nor U9899 (N_9899,N_9504,N_9742);
and U9900 (N_9900,N_9738,N_9530);
nor U9901 (N_9901,N_9705,N_9509);
or U9902 (N_9902,N_9646,N_9585);
nand U9903 (N_9903,N_9744,N_9712);
or U9904 (N_9904,N_9639,N_9593);
xnor U9905 (N_9905,N_9677,N_9543);
nand U9906 (N_9906,N_9580,N_9715);
and U9907 (N_9907,N_9573,N_9739);
and U9908 (N_9908,N_9659,N_9575);
nand U9909 (N_9909,N_9508,N_9746);
and U9910 (N_9910,N_9530,N_9742);
nand U9911 (N_9911,N_9710,N_9669);
or U9912 (N_9912,N_9612,N_9642);
nand U9913 (N_9913,N_9511,N_9725);
nor U9914 (N_9914,N_9540,N_9562);
nand U9915 (N_9915,N_9550,N_9635);
nand U9916 (N_9916,N_9564,N_9600);
nor U9917 (N_9917,N_9524,N_9676);
nor U9918 (N_9918,N_9593,N_9592);
and U9919 (N_9919,N_9683,N_9588);
xnor U9920 (N_9920,N_9646,N_9651);
nor U9921 (N_9921,N_9670,N_9598);
nor U9922 (N_9922,N_9504,N_9548);
and U9923 (N_9923,N_9518,N_9708);
and U9924 (N_9924,N_9652,N_9679);
and U9925 (N_9925,N_9523,N_9689);
and U9926 (N_9926,N_9656,N_9579);
nor U9927 (N_9927,N_9542,N_9535);
xnor U9928 (N_9928,N_9702,N_9707);
or U9929 (N_9929,N_9585,N_9507);
xor U9930 (N_9930,N_9712,N_9708);
xnor U9931 (N_9931,N_9599,N_9505);
nor U9932 (N_9932,N_9583,N_9745);
xor U9933 (N_9933,N_9662,N_9613);
nand U9934 (N_9934,N_9699,N_9666);
xor U9935 (N_9935,N_9629,N_9705);
xor U9936 (N_9936,N_9721,N_9602);
xnor U9937 (N_9937,N_9592,N_9610);
xnor U9938 (N_9938,N_9711,N_9568);
nor U9939 (N_9939,N_9573,N_9602);
nand U9940 (N_9940,N_9566,N_9734);
nor U9941 (N_9941,N_9524,N_9530);
nand U9942 (N_9942,N_9593,N_9719);
xnor U9943 (N_9943,N_9601,N_9579);
xor U9944 (N_9944,N_9687,N_9644);
nor U9945 (N_9945,N_9593,N_9741);
nor U9946 (N_9946,N_9702,N_9626);
and U9947 (N_9947,N_9715,N_9636);
nor U9948 (N_9948,N_9531,N_9707);
or U9949 (N_9949,N_9633,N_9575);
and U9950 (N_9950,N_9577,N_9714);
or U9951 (N_9951,N_9511,N_9685);
or U9952 (N_9952,N_9617,N_9582);
and U9953 (N_9953,N_9530,N_9582);
and U9954 (N_9954,N_9500,N_9535);
nor U9955 (N_9955,N_9503,N_9749);
nand U9956 (N_9956,N_9560,N_9688);
nor U9957 (N_9957,N_9626,N_9690);
nor U9958 (N_9958,N_9561,N_9707);
nor U9959 (N_9959,N_9725,N_9507);
nand U9960 (N_9960,N_9692,N_9640);
or U9961 (N_9961,N_9514,N_9578);
nand U9962 (N_9962,N_9659,N_9571);
xnor U9963 (N_9963,N_9598,N_9550);
or U9964 (N_9964,N_9729,N_9736);
xor U9965 (N_9965,N_9734,N_9690);
and U9966 (N_9966,N_9611,N_9505);
xnor U9967 (N_9967,N_9547,N_9530);
and U9968 (N_9968,N_9557,N_9549);
nor U9969 (N_9969,N_9546,N_9509);
and U9970 (N_9970,N_9517,N_9707);
xor U9971 (N_9971,N_9727,N_9711);
nor U9972 (N_9972,N_9616,N_9601);
nor U9973 (N_9973,N_9573,N_9586);
nand U9974 (N_9974,N_9715,N_9639);
nand U9975 (N_9975,N_9561,N_9722);
xnor U9976 (N_9976,N_9561,N_9540);
nand U9977 (N_9977,N_9569,N_9633);
and U9978 (N_9978,N_9658,N_9565);
xor U9979 (N_9979,N_9542,N_9537);
or U9980 (N_9980,N_9553,N_9690);
xor U9981 (N_9981,N_9722,N_9642);
nand U9982 (N_9982,N_9716,N_9504);
xor U9983 (N_9983,N_9656,N_9676);
or U9984 (N_9984,N_9742,N_9637);
and U9985 (N_9985,N_9556,N_9513);
xor U9986 (N_9986,N_9519,N_9651);
or U9987 (N_9987,N_9691,N_9722);
or U9988 (N_9988,N_9685,N_9634);
nor U9989 (N_9989,N_9609,N_9643);
or U9990 (N_9990,N_9552,N_9648);
and U9991 (N_9991,N_9747,N_9614);
xnor U9992 (N_9992,N_9535,N_9583);
xor U9993 (N_9993,N_9641,N_9715);
or U9994 (N_9994,N_9711,N_9731);
nand U9995 (N_9995,N_9656,N_9733);
nor U9996 (N_9996,N_9710,N_9519);
nor U9997 (N_9997,N_9690,N_9715);
and U9998 (N_9998,N_9588,N_9616);
or U9999 (N_9999,N_9621,N_9670);
xor U10000 (N_10000,N_9804,N_9838);
nand U10001 (N_10001,N_9905,N_9952);
xnor U10002 (N_10002,N_9778,N_9876);
and U10003 (N_10003,N_9877,N_9767);
xor U10004 (N_10004,N_9947,N_9812);
nand U10005 (N_10005,N_9752,N_9816);
and U10006 (N_10006,N_9854,N_9865);
or U10007 (N_10007,N_9789,N_9795);
and U10008 (N_10008,N_9924,N_9824);
or U10009 (N_10009,N_9867,N_9935);
and U10010 (N_10010,N_9933,N_9794);
nor U10011 (N_10011,N_9834,N_9982);
nor U10012 (N_10012,N_9820,N_9988);
nor U10013 (N_10013,N_9870,N_9873);
nand U10014 (N_10014,N_9814,N_9875);
and U10015 (N_10015,N_9949,N_9826);
and U10016 (N_10016,N_9861,N_9929);
and U10017 (N_10017,N_9844,N_9950);
xor U10018 (N_10018,N_9993,N_9991);
and U10019 (N_10019,N_9997,N_9846);
nand U10020 (N_10020,N_9848,N_9827);
and U10021 (N_10021,N_9966,N_9998);
nor U10022 (N_10022,N_9766,N_9866);
or U10023 (N_10023,N_9891,N_9774);
nor U10024 (N_10024,N_9822,N_9967);
xor U10025 (N_10025,N_9979,N_9823);
nand U10026 (N_10026,N_9970,N_9953);
nor U10027 (N_10027,N_9761,N_9811);
nor U10028 (N_10028,N_9995,N_9780);
nand U10029 (N_10029,N_9828,N_9971);
or U10030 (N_10030,N_9863,N_9959);
nand U10031 (N_10031,N_9840,N_9962);
nand U10032 (N_10032,N_9808,N_9839);
xnor U10033 (N_10033,N_9939,N_9888);
nand U10034 (N_10034,N_9978,N_9882);
nand U10035 (N_10035,N_9917,N_9769);
nand U10036 (N_10036,N_9755,N_9800);
or U10037 (N_10037,N_9897,N_9868);
nand U10038 (N_10038,N_9750,N_9777);
and U10039 (N_10039,N_9799,N_9954);
nand U10040 (N_10040,N_9773,N_9832);
xnor U10041 (N_10041,N_9847,N_9910);
nand U10042 (N_10042,N_9806,N_9909);
and U10043 (N_10043,N_9906,N_9898);
nand U10044 (N_10044,N_9759,N_9860);
nor U10045 (N_10045,N_9754,N_9790);
xnor U10046 (N_10046,N_9992,N_9829);
nand U10047 (N_10047,N_9874,N_9864);
and U10048 (N_10048,N_9879,N_9785);
xnor U10049 (N_10049,N_9851,N_9931);
or U10050 (N_10050,N_9983,N_9934);
and U10051 (N_10051,N_9768,N_9810);
or U10052 (N_10052,N_9922,N_9842);
and U10053 (N_10053,N_9833,N_9821);
nor U10054 (N_10054,N_9914,N_9764);
nand U10055 (N_10055,N_9858,N_9932);
xnor U10056 (N_10056,N_9765,N_9825);
xnor U10057 (N_10057,N_9943,N_9835);
nor U10058 (N_10058,N_9757,N_9880);
nand U10059 (N_10059,N_9969,N_9802);
or U10060 (N_10060,N_9902,N_9981);
or U10061 (N_10061,N_9787,N_9855);
xnor U10062 (N_10062,N_9984,N_9915);
or U10063 (N_10063,N_9972,N_9771);
nor U10064 (N_10064,N_9907,N_9890);
or U10065 (N_10065,N_9895,N_9964);
and U10066 (N_10066,N_9941,N_9976);
or U10067 (N_10067,N_9975,N_9869);
xnor U10068 (N_10068,N_9920,N_9892);
nor U10069 (N_10069,N_9996,N_9786);
xor U10070 (N_10070,N_9883,N_9796);
nand U10071 (N_10071,N_9776,N_9887);
and U10072 (N_10072,N_9999,N_9942);
nor U10073 (N_10073,N_9884,N_9893);
nor U10074 (N_10074,N_9760,N_9817);
xnor U10075 (N_10075,N_9797,N_9770);
xor U10076 (N_10076,N_9805,N_9801);
or U10077 (N_10077,N_9836,N_9936);
or U10078 (N_10078,N_9901,N_9974);
xor U10079 (N_10079,N_9803,N_9798);
xnor U10080 (N_10080,N_9753,N_9762);
xor U10081 (N_10081,N_9818,N_9779);
and U10082 (N_10082,N_9807,N_9782);
and U10083 (N_10083,N_9894,N_9763);
nor U10084 (N_10084,N_9788,N_9921);
nand U10085 (N_10085,N_9948,N_9815);
xnor U10086 (N_10086,N_9913,N_9783);
xor U10087 (N_10087,N_9850,N_9925);
nand U10088 (N_10088,N_9857,N_9899);
and U10089 (N_10089,N_9945,N_9937);
nand U10090 (N_10090,N_9963,N_9955);
or U10091 (N_10091,N_9878,N_9756);
and U10092 (N_10092,N_9830,N_9852);
xor U10093 (N_10093,N_9940,N_9841);
and U10094 (N_10094,N_9911,N_9946);
and U10095 (N_10095,N_9791,N_9986);
nor U10096 (N_10096,N_9896,N_9813);
nand U10097 (N_10097,N_9938,N_9928);
and U10098 (N_10098,N_9886,N_9793);
nand U10099 (N_10099,N_9961,N_9926);
nor U10100 (N_10100,N_9784,N_9927);
and U10101 (N_10101,N_9977,N_9916);
and U10102 (N_10102,N_9871,N_9985);
nand U10103 (N_10103,N_9859,N_9900);
or U10104 (N_10104,N_9994,N_9965);
nor U10105 (N_10105,N_9987,N_9957);
nor U10106 (N_10106,N_9872,N_9968);
and U10107 (N_10107,N_9849,N_9845);
xnor U10108 (N_10108,N_9973,N_9958);
and U10109 (N_10109,N_9881,N_9912);
nand U10110 (N_10110,N_9758,N_9944);
or U10111 (N_10111,N_9889,N_9792);
or U10112 (N_10112,N_9919,N_9951);
or U10113 (N_10113,N_9918,N_9781);
and U10114 (N_10114,N_9819,N_9775);
or U10115 (N_10115,N_9831,N_9980);
and U10116 (N_10116,N_9809,N_9908);
or U10117 (N_10117,N_9772,N_9751);
nor U10118 (N_10118,N_9956,N_9837);
nand U10119 (N_10119,N_9853,N_9843);
xor U10120 (N_10120,N_9862,N_9885);
or U10121 (N_10121,N_9990,N_9960);
and U10122 (N_10122,N_9989,N_9903);
nor U10123 (N_10123,N_9856,N_9930);
and U10124 (N_10124,N_9904,N_9923);
nor U10125 (N_10125,N_9777,N_9917);
nor U10126 (N_10126,N_9889,N_9856);
and U10127 (N_10127,N_9958,N_9856);
and U10128 (N_10128,N_9885,N_9947);
xor U10129 (N_10129,N_9799,N_9761);
nand U10130 (N_10130,N_9928,N_9915);
and U10131 (N_10131,N_9856,N_9872);
or U10132 (N_10132,N_9879,N_9779);
nor U10133 (N_10133,N_9772,N_9756);
xor U10134 (N_10134,N_9900,N_9964);
or U10135 (N_10135,N_9891,N_9848);
xor U10136 (N_10136,N_9813,N_9979);
and U10137 (N_10137,N_9931,N_9751);
nor U10138 (N_10138,N_9784,N_9768);
nor U10139 (N_10139,N_9930,N_9957);
and U10140 (N_10140,N_9936,N_9872);
nand U10141 (N_10141,N_9938,N_9877);
or U10142 (N_10142,N_9775,N_9861);
nor U10143 (N_10143,N_9997,N_9959);
xnor U10144 (N_10144,N_9809,N_9939);
or U10145 (N_10145,N_9764,N_9815);
nor U10146 (N_10146,N_9837,N_9906);
xnor U10147 (N_10147,N_9886,N_9943);
nand U10148 (N_10148,N_9909,N_9962);
and U10149 (N_10149,N_9980,N_9760);
nor U10150 (N_10150,N_9780,N_9884);
xor U10151 (N_10151,N_9831,N_9860);
xor U10152 (N_10152,N_9930,N_9836);
and U10153 (N_10153,N_9773,N_9869);
nor U10154 (N_10154,N_9988,N_9757);
nor U10155 (N_10155,N_9899,N_9889);
nor U10156 (N_10156,N_9854,N_9804);
nand U10157 (N_10157,N_9999,N_9931);
nor U10158 (N_10158,N_9839,N_9873);
nor U10159 (N_10159,N_9936,N_9887);
or U10160 (N_10160,N_9967,N_9895);
or U10161 (N_10161,N_9889,N_9844);
or U10162 (N_10162,N_9768,N_9782);
xnor U10163 (N_10163,N_9855,N_9912);
or U10164 (N_10164,N_9909,N_9815);
nor U10165 (N_10165,N_9954,N_9839);
nor U10166 (N_10166,N_9869,N_9798);
xnor U10167 (N_10167,N_9899,N_9805);
nor U10168 (N_10168,N_9972,N_9760);
nor U10169 (N_10169,N_9940,N_9900);
or U10170 (N_10170,N_9908,N_9889);
and U10171 (N_10171,N_9883,N_9905);
xor U10172 (N_10172,N_9763,N_9956);
nor U10173 (N_10173,N_9804,N_9757);
or U10174 (N_10174,N_9866,N_9810);
xor U10175 (N_10175,N_9823,N_9861);
xnor U10176 (N_10176,N_9769,N_9970);
nand U10177 (N_10177,N_9877,N_9880);
or U10178 (N_10178,N_9760,N_9768);
or U10179 (N_10179,N_9774,N_9877);
xnor U10180 (N_10180,N_9915,N_9869);
nand U10181 (N_10181,N_9932,N_9822);
nand U10182 (N_10182,N_9764,N_9917);
or U10183 (N_10183,N_9864,N_9848);
and U10184 (N_10184,N_9864,N_9850);
or U10185 (N_10185,N_9906,N_9822);
nor U10186 (N_10186,N_9974,N_9949);
and U10187 (N_10187,N_9846,N_9877);
nor U10188 (N_10188,N_9902,N_9936);
and U10189 (N_10189,N_9796,N_9814);
xnor U10190 (N_10190,N_9981,N_9876);
nor U10191 (N_10191,N_9872,N_9773);
or U10192 (N_10192,N_9867,N_9982);
or U10193 (N_10193,N_9755,N_9783);
and U10194 (N_10194,N_9925,N_9867);
and U10195 (N_10195,N_9868,N_9755);
and U10196 (N_10196,N_9925,N_9881);
nor U10197 (N_10197,N_9891,N_9785);
nor U10198 (N_10198,N_9920,N_9934);
nand U10199 (N_10199,N_9958,N_9807);
xnor U10200 (N_10200,N_9809,N_9844);
or U10201 (N_10201,N_9872,N_9904);
or U10202 (N_10202,N_9789,N_9782);
and U10203 (N_10203,N_9789,N_9924);
nor U10204 (N_10204,N_9873,N_9827);
nor U10205 (N_10205,N_9935,N_9987);
xor U10206 (N_10206,N_9929,N_9907);
or U10207 (N_10207,N_9761,N_9937);
nor U10208 (N_10208,N_9869,N_9858);
or U10209 (N_10209,N_9982,N_9993);
nand U10210 (N_10210,N_9891,N_9887);
xor U10211 (N_10211,N_9794,N_9964);
nor U10212 (N_10212,N_9761,N_9780);
xnor U10213 (N_10213,N_9876,N_9804);
nor U10214 (N_10214,N_9865,N_9967);
nor U10215 (N_10215,N_9780,N_9849);
nand U10216 (N_10216,N_9879,N_9880);
or U10217 (N_10217,N_9906,N_9802);
nor U10218 (N_10218,N_9783,N_9785);
xnor U10219 (N_10219,N_9826,N_9838);
or U10220 (N_10220,N_9823,N_9928);
nand U10221 (N_10221,N_9895,N_9829);
or U10222 (N_10222,N_9916,N_9883);
and U10223 (N_10223,N_9938,N_9868);
nor U10224 (N_10224,N_9760,N_9845);
or U10225 (N_10225,N_9752,N_9880);
xor U10226 (N_10226,N_9962,N_9966);
nand U10227 (N_10227,N_9883,N_9824);
nor U10228 (N_10228,N_9944,N_9845);
nand U10229 (N_10229,N_9866,N_9919);
nand U10230 (N_10230,N_9915,N_9764);
and U10231 (N_10231,N_9906,N_9931);
nor U10232 (N_10232,N_9816,N_9945);
nand U10233 (N_10233,N_9871,N_9909);
nand U10234 (N_10234,N_9759,N_9767);
xor U10235 (N_10235,N_9855,N_9756);
or U10236 (N_10236,N_9934,N_9947);
nor U10237 (N_10237,N_9751,N_9992);
xor U10238 (N_10238,N_9895,N_9831);
nor U10239 (N_10239,N_9946,N_9910);
and U10240 (N_10240,N_9815,N_9786);
nor U10241 (N_10241,N_9802,N_9970);
xor U10242 (N_10242,N_9947,N_9820);
and U10243 (N_10243,N_9801,N_9910);
or U10244 (N_10244,N_9955,N_9769);
nand U10245 (N_10245,N_9799,N_9937);
nand U10246 (N_10246,N_9908,N_9885);
nor U10247 (N_10247,N_9896,N_9761);
nor U10248 (N_10248,N_9780,N_9858);
xnor U10249 (N_10249,N_9797,N_9791);
nand U10250 (N_10250,N_10086,N_10113);
and U10251 (N_10251,N_10065,N_10052);
and U10252 (N_10252,N_10159,N_10219);
nor U10253 (N_10253,N_10078,N_10116);
nor U10254 (N_10254,N_10018,N_10148);
xnor U10255 (N_10255,N_10202,N_10079);
or U10256 (N_10256,N_10197,N_10004);
nor U10257 (N_10257,N_10165,N_10147);
nand U10258 (N_10258,N_10076,N_10184);
nand U10259 (N_10259,N_10029,N_10097);
nor U10260 (N_10260,N_10226,N_10246);
xnor U10261 (N_10261,N_10046,N_10214);
nand U10262 (N_10262,N_10200,N_10245);
nor U10263 (N_10263,N_10217,N_10024);
nor U10264 (N_10264,N_10223,N_10111);
or U10265 (N_10265,N_10005,N_10106);
nor U10266 (N_10266,N_10025,N_10092);
nor U10267 (N_10267,N_10208,N_10166);
or U10268 (N_10268,N_10198,N_10068);
and U10269 (N_10269,N_10152,N_10093);
xnor U10270 (N_10270,N_10058,N_10021);
nand U10271 (N_10271,N_10187,N_10191);
or U10272 (N_10272,N_10061,N_10201);
and U10273 (N_10273,N_10178,N_10188);
and U10274 (N_10274,N_10149,N_10129);
nor U10275 (N_10275,N_10209,N_10088);
nor U10276 (N_10276,N_10141,N_10199);
and U10277 (N_10277,N_10080,N_10062);
nor U10278 (N_10278,N_10193,N_10205);
or U10279 (N_10279,N_10185,N_10011);
or U10280 (N_10280,N_10027,N_10244);
nor U10281 (N_10281,N_10035,N_10161);
xnor U10282 (N_10282,N_10098,N_10054);
or U10283 (N_10283,N_10233,N_10010);
xor U10284 (N_10284,N_10006,N_10108);
xor U10285 (N_10285,N_10134,N_10124);
or U10286 (N_10286,N_10123,N_10069);
and U10287 (N_10287,N_10121,N_10213);
xnor U10288 (N_10288,N_10229,N_10158);
nor U10289 (N_10289,N_10037,N_10231);
nand U10290 (N_10290,N_10167,N_10090);
and U10291 (N_10291,N_10089,N_10127);
nor U10292 (N_10292,N_10162,N_10125);
xnor U10293 (N_10293,N_10059,N_10212);
or U10294 (N_10294,N_10242,N_10072);
nand U10295 (N_10295,N_10221,N_10057);
or U10296 (N_10296,N_10241,N_10215);
nor U10297 (N_10297,N_10102,N_10204);
and U10298 (N_10298,N_10074,N_10136);
or U10299 (N_10299,N_10033,N_10218);
or U10300 (N_10300,N_10032,N_10207);
nor U10301 (N_10301,N_10138,N_10145);
nor U10302 (N_10302,N_10118,N_10120);
nor U10303 (N_10303,N_10016,N_10066);
nand U10304 (N_10304,N_10169,N_10195);
xor U10305 (N_10305,N_10186,N_10060);
or U10306 (N_10306,N_10103,N_10132);
or U10307 (N_10307,N_10085,N_10154);
nand U10308 (N_10308,N_10012,N_10084);
or U10309 (N_10309,N_10056,N_10101);
or U10310 (N_10310,N_10164,N_10156);
nor U10311 (N_10311,N_10104,N_10181);
xor U10312 (N_10312,N_10177,N_10237);
and U10313 (N_10313,N_10003,N_10105);
nand U10314 (N_10314,N_10155,N_10007);
xnor U10315 (N_10315,N_10063,N_10210);
or U10316 (N_10316,N_10216,N_10232);
or U10317 (N_10317,N_10023,N_10110);
nand U10318 (N_10318,N_10128,N_10153);
or U10319 (N_10319,N_10131,N_10049);
nor U10320 (N_10320,N_10094,N_10031);
and U10321 (N_10321,N_10075,N_10115);
or U10322 (N_10322,N_10206,N_10170);
xnor U10323 (N_10323,N_10100,N_10034);
xnor U10324 (N_10324,N_10107,N_10014);
xnor U10325 (N_10325,N_10183,N_10042);
nand U10326 (N_10326,N_10143,N_10236);
xor U10327 (N_10327,N_10122,N_10142);
nor U10328 (N_10328,N_10082,N_10000);
nor U10329 (N_10329,N_10146,N_10243);
xnor U10330 (N_10330,N_10020,N_10126);
nor U10331 (N_10331,N_10220,N_10176);
nand U10332 (N_10332,N_10119,N_10081);
nor U10333 (N_10333,N_10174,N_10070);
nand U10334 (N_10334,N_10077,N_10117);
nor U10335 (N_10335,N_10248,N_10045);
and U10336 (N_10336,N_10190,N_10180);
nor U10337 (N_10337,N_10038,N_10175);
nor U10338 (N_10338,N_10151,N_10234);
or U10339 (N_10339,N_10225,N_10172);
or U10340 (N_10340,N_10048,N_10073);
nand U10341 (N_10341,N_10247,N_10071);
nand U10342 (N_10342,N_10150,N_10022);
and U10343 (N_10343,N_10194,N_10019);
nand U10344 (N_10344,N_10168,N_10224);
xnor U10345 (N_10345,N_10053,N_10095);
nor U10346 (N_10346,N_10140,N_10087);
xor U10347 (N_10347,N_10083,N_10055);
nand U10348 (N_10348,N_10238,N_10064);
and U10349 (N_10349,N_10051,N_10114);
nor U10350 (N_10350,N_10192,N_10239);
or U10351 (N_10351,N_10189,N_10235);
or U10352 (N_10352,N_10028,N_10015);
xnor U10353 (N_10353,N_10171,N_10026);
or U10354 (N_10354,N_10139,N_10009);
and U10355 (N_10355,N_10179,N_10017);
and U10356 (N_10356,N_10112,N_10203);
xor U10357 (N_10357,N_10091,N_10144);
nand U10358 (N_10358,N_10249,N_10030);
or U10359 (N_10359,N_10109,N_10002);
nand U10360 (N_10360,N_10096,N_10039);
or U10361 (N_10361,N_10163,N_10040);
nor U10362 (N_10362,N_10130,N_10157);
and U10363 (N_10363,N_10211,N_10067);
or U10364 (N_10364,N_10173,N_10044);
and U10365 (N_10365,N_10182,N_10008);
nor U10366 (N_10366,N_10228,N_10041);
and U10367 (N_10367,N_10240,N_10160);
or U10368 (N_10368,N_10043,N_10001);
or U10369 (N_10369,N_10013,N_10036);
xor U10370 (N_10370,N_10227,N_10196);
and U10371 (N_10371,N_10222,N_10230);
or U10372 (N_10372,N_10135,N_10137);
nand U10373 (N_10373,N_10047,N_10099);
xor U10374 (N_10374,N_10133,N_10050);
xor U10375 (N_10375,N_10191,N_10100);
xnor U10376 (N_10376,N_10023,N_10145);
and U10377 (N_10377,N_10188,N_10172);
xnor U10378 (N_10378,N_10211,N_10060);
xnor U10379 (N_10379,N_10221,N_10021);
nand U10380 (N_10380,N_10088,N_10092);
nand U10381 (N_10381,N_10007,N_10193);
xnor U10382 (N_10382,N_10161,N_10151);
xnor U10383 (N_10383,N_10039,N_10044);
xor U10384 (N_10384,N_10188,N_10238);
xnor U10385 (N_10385,N_10164,N_10011);
or U10386 (N_10386,N_10041,N_10154);
and U10387 (N_10387,N_10086,N_10067);
nor U10388 (N_10388,N_10013,N_10072);
nand U10389 (N_10389,N_10104,N_10183);
and U10390 (N_10390,N_10168,N_10171);
or U10391 (N_10391,N_10161,N_10070);
and U10392 (N_10392,N_10226,N_10147);
nand U10393 (N_10393,N_10139,N_10034);
nand U10394 (N_10394,N_10139,N_10228);
or U10395 (N_10395,N_10135,N_10091);
nand U10396 (N_10396,N_10130,N_10087);
or U10397 (N_10397,N_10151,N_10222);
nor U10398 (N_10398,N_10214,N_10230);
and U10399 (N_10399,N_10231,N_10017);
xor U10400 (N_10400,N_10034,N_10078);
or U10401 (N_10401,N_10152,N_10187);
or U10402 (N_10402,N_10015,N_10228);
nand U10403 (N_10403,N_10029,N_10025);
nor U10404 (N_10404,N_10135,N_10193);
nor U10405 (N_10405,N_10218,N_10243);
xor U10406 (N_10406,N_10238,N_10167);
nand U10407 (N_10407,N_10129,N_10177);
or U10408 (N_10408,N_10043,N_10109);
xor U10409 (N_10409,N_10089,N_10164);
or U10410 (N_10410,N_10033,N_10173);
nor U10411 (N_10411,N_10020,N_10042);
and U10412 (N_10412,N_10157,N_10006);
xnor U10413 (N_10413,N_10236,N_10162);
and U10414 (N_10414,N_10170,N_10066);
xor U10415 (N_10415,N_10092,N_10215);
or U10416 (N_10416,N_10090,N_10242);
and U10417 (N_10417,N_10195,N_10047);
nand U10418 (N_10418,N_10075,N_10192);
or U10419 (N_10419,N_10103,N_10211);
nand U10420 (N_10420,N_10111,N_10031);
xnor U10421 (N_10421,N_10108,N_10185);
nand U10422 (N_10422,N_10130,N_10109);
and U10423 (N_10423,N_10183,N_10084);
nor U10424 (N_10424,N_10120,N_10002);
or U10425 (N_10425,N_10034,N_10165);
nand U10426 (N_10426,N_10248,N_10194);
or U10427 (N_10427,N_10053,N_10224);
nor U10428 (N_10428,N_10109,N_10114);
xnor U10429 (N_10429,N_10222,N_10092);
nand U10430 (N_10430,N_10130,N_10100);
nand U10431 (N_10431,N_10014,N_10118);
nor U10432 (N_10432,N_10129,N_10123);
or U10433 (N_10433,N_10027,N_10043);
xnor U10434 (N_10434,N_10217,N_10243);
and U10435 (N_10435,N_10055,N_10004);
or U10436 (N_10436,N_10096,N_10061);
or U10437 (N_10437,N_10208,N_10217);
xor U10438 (N_10438,N_10097,N_10162);
nand U10439 (N_10439,N_10126,N_10075);
or U10440 (N_10440,N_10049,N_10164);
xnor U10441 (N_10441,N_10013,N_10098);
and U10442 (N_10442,N_10185,N_10208);
nand U10443 (N_10443,N_10192,N_10244);
nor U10444 (N_10444,N_10231,N_10170);
nor U10445 (N_10445,N_10224,N_10207);
and U10446 (N_10446,N_10210,N_10021);
and U10447 (N_10447,N_10198,N_10216);
and U10448 (N_10448,N_10204,N_10026);
xnor U10449 (N_10449,N_10068,N_10128);
nor U10450 (N_10450,N_10156,N_10000);
nand U10451 (N_10451,N_10037,N_10116);
xnor U10452 (N_10452,N_10176,N_10003);
and U10453 (N_10453,N_10029,N_10022);
or U10454 (N_10454,N_10112,N_10075);
nor U10455 (N_10455,N_10228,N_10106);
nor U10456 (N_10456,N_10057,N_10249);
nor U10457 (N_10457,N_10137,N_10002);
nand U10458 (N_10458,N_10159,N_10015);
nor U10459 (N_10459,N_10090,N_10154);
and U10460 (N_10460,N_10146,N_10010);
nand U10461 (N_10461,N_10001,N_10137);
xnor U10462 (N_10462,N_10068,N_10056);
or U10463 (N_10463,N_10028,N_10230);
and U10464 (N_10464,N_10248,N_10200);
or U10465 (N_10465,N_10086,N_10111);
and U10466 (N_10466,N_10126,N_10067);
nand U10467 (N_10467,N_10019,N_10078);
and U10468 (N_10468,N_10232,N_10095);
or U10469 (N_10469,N_10136,N_10033);
nand U10470 (N_10470,N_10055,N_10072);
xnor U10471 (N_10471,N_10131,N_10106);
xnor U10472 (N_10472,N_10160,N_10067);
xnor U10473 (N_10473,N_10108,N_10127);
nor U10474 (N_10474,N_10011,N_10043);
and U10475 (N_10475,N_10205,N_10200);
nor U10476 (N_10476,N_10152,N_10066);
xnor U10477 (N_10477,N_10065,N_10224);
nor U10478 (N_10478,N_10143,N_10152);
or U10479 (N_10479,N_10228,N_10108);
xnor U10480 (N_10480,N_10211,N_10038);
xnor U10481 (N_10481,N_10190,N_10085);
or U10482 (N_10482,N_10051,N_10200);
xnor U10483 (N_10483,N_10114,N_10184);
or U10484 (N_10484,N_10180,N_10172);
xor U10485 (N_10485,N_10079,N_10120);
and U10486 (N_10486,N_10034,N_10085);
or U10487 (N_10487,N_10134,N_10020);
nor U10488 (N_10488,N_10123,N_10108);
and U10489 (N_10489,N_10233,N_10000);
and U10490 (N_10490,N_10088,N_10181);
nor U10491 (N_10491,N_10218,N_10028);
nor U10492 (N_10492,N_10114,N_10032);
and U10493 (N_10493,N_10074,N_10115);
or U10494 (N_10494,N_10016,N_10080);
xor U10495 (N_10495,N_10189,N_10023);
nor U10496 (N_10496,N_10119,N_10049);
nand U10497 (N_10497,N_10163,N_10244);
xor U10498 (N_10498,N_10129,N_10178);
or U10499 (N_10499,N_10207,N_10085);
nor U10500 (N_10500,N_10382,N_10487);
nand U10501 (N_10501,N_10320,N_10464);
or U10502 (N_10502,N_10287,N_10356);
nor U10503 (N_10503,N_10353,N_10313);
or U10504 (N_10504,N_10404,N_10298);
nor U10505 (N_10505,N_10316,N_10424);
nand U10506 (N_10506,N_10486,N_10453);
and U10507 (N_10507,N_10395,N_10273);
and U10508 (N_10508,N_10389,N_10458);
xor U10509 (N_10509,N_10375,N_10303);
and U10510 (N_10510,N_10300,N_10488);
and U10511 (N_10511,N_10272,N_10335);
xnor U10512 (N_10512,N_10454,N_10333);
xor U10513 (N_10513,N_10388,N_10429);
nand U10514 (N_10514,N_10283,N_10430);
nor U10515 (N_10515,N_10485,N_10324);
and U10516 (N_10516,N_10436,N_10263);
nor U10517 (N_10517,N_10416,N_10269);
xor U10518 (N_10518,N_10460,N_10426);
xnor U10519 (N_10519,N_10299,N_10425);
nand U10520 (N_10520,N_10367,N_10337);
nand U10521 (N_10521,N_10448,N_10476);
nand U10522 (N_10522,N_10258,N_10341);
and U10523 (N_10523,N_10312,N_10332);
xor U10524 (N_10524,N_10260,N_10346);
xnor U10525 (N_10525,N_10253,N_10366);
xnor U10526 (N_10526,N_10469,N_10363);
nor U10527 (N_10527,N_10493,N_10403);
or U10528 (N_10528,N_10280,N_10307);
xnor U10529 (N_10529,N_10317,N_10481);
nor U10530 (N_10530,N_10314,N_10496);
and U10531 (N_10531,N_10490,N_10265);
and U10532 (N_10532,N_10284,N_10465);
and U10533 (N_10533,N_10431,N_10259);
xnor U10534 (N_10534,N_10277,N_10295);
nor U10535 (N_10535,N_10463,N_10378);
or U10536 (N_10536,N_10359,N_10380);
and U10537 (N_10537,N_10438,N_10405);
xor U10538 (N_10538,N_10472,N_10264);
nor U10539 (N_10539,N_10385,N_10386);
nor U10540 (N_10540,N_10445,N_10310);
xor U10541 (N_10541,N_10330,N_10348);
nor U10542 (N_10542,N_10250,N_10281);
or U10543 (N_10543,N_10285,N_10440);
nor U10544 (N_10544,N_10398,N_10396);
or U10545 (N_10545,N_10446,N_10443);
nand U10546 (N_10546,N_10336,N_10468);
and U10547 (N_10547,N_10351,N_10489);
nor U10548 (N_10548,N_10302,N_10370);
or U10549 (N_10549,N_10392,N_10291);
or U10550 (N_10550,N_10399,N_10288);
nand U10551 (N_10551,N_10467,N_10305);
xnor U10552 (N_10552,N_10301,N_10358);
xor U10553 (N_10553,N_10421,N_10318);
nand U10554 (N_10554,N_10270,N_10406);
nor U10555 (N_10555,N_10345,N_10296);
and U10556 (N_10556,N_10274,N_10457);
nand U10557 (N_10557,N_10290,N_10322);
nand U10558 (N_10558,N_10402,N_10384);
and U10559 (N_10559,N_10364,N_10474);
and U10560 (N_10560,N_10254,N_10420);
nor U10561 (N_10561,N_10338,N_10462);
nand U10562 (N_10562,N_10441,N_10297);
and U10563 (N_10563,N_10444,N_10365);
or U10564 (N_10564,N_10482,N_10374);
nor U10565 (N_10565,N_10412,N_10319);
and U10566 (N_10566,N_10452,N_10450);
or U10567 (N_10567,N_10262,N_10439);
xor U10568 (N_10568,N_10306,N_10347);
xnor U10569 (N_10569,N_10355,N_10331);
nor U10570 (N_10570,N_10471,N_10477);
xnor U10571 (N_10571,N_10393,N_10286);
xor U10572 (N_10572,N_10315,N_10499);
nor U10573 (N_10573,N_10266,N_10282);
xor U10574 (N_10574,N_10276,N_10304);
nand U10575 (N_10575,N_10350,N_10261);
nor U10576 (N_10576,N_10255,N_10410);
xnor U10577 (N_10577,N_10328,N_10362);
nand U10578 (N_10578,N_10326,N_10417);
xnor U10579 (N_10579,N_10478,N_10294);
xnor U10580 (N_10580,N_10434,N_10354);
or U10581 (N_10581,N_10271,N_10433);
or U10582 (N_10582,N_10484,N_10432);
xor U10583 (N_10583,N_10407,N_10437);
xnor U10584 (N_10584,N_10372,N_10479);
xor U10585 (N_10585,N_10498,N_10394);
nor U10586 (N_10586,N_10414,N_10279);
nand U10587 (N_10587,N_10377,N_10428);
nor U10588 (N_10588,N_10495,N_10267);
and U10589 (N_10589,N_10352,N_10413);
or U10590 (N_10590,N_10342,N_10309);
nor U10591 (N_10591,N_10383,N_10268);
nor U10592 (N_10592,N_10449,N_10387);
nor U10593 (N_10593,N_10423,N_10349);
nor U10594 (N_10594,N_10409,N_10289);
xor U10595 (N_10595,N_10397,N_10418);
and U10596 (N_10596,N_10376,N_10390);
xnor U10597 (N_10597,N_10334,N_10292);
or U10598 (N_10598,N_10340,N_10325);
xnor U10599 (N_10599,N_10293,N_10422);
nand U10600 (N_10600,N_10427,N_10494);
xnor U10601 (N_10601,N_10483,N_10357);
nor U10602 (N_10602,N_10329,N_10461);
or U10603 (N_10603,N_10278,N_10360);
nor U10604 (N_10604,N_10497,N_10442);
nand U10605 (N_10605,N_10339,N_10419);
nor U10606 (N_10606,N_10408,N_10411);
xnor U10607 (N_10607,N_10368,N_10492);
nor U10608 (N_10608,N_10308,N_10275);
nand U10609 (N_10609,N_10379,N_10451);
nor U10610 (N_10610,N_10373,N_10473);
nor U10611 (N_10611,N_10470,N_10251);
nand U10612 (N_10612,N_10491,N_10257);
nor U10613 (N_10613,N_10455,N_10311);
nor U10614 (N_10614,N_10447,N_10435);
xor U10615 (N_10615,N_10381,N_10371);
nand U10616 (N_10616,N_10400,N_10327);
nor U10617 (N_10617,N_10401,N_10252);
and U10618 (N_10618,N_10344,N_10475);
and U10619 (N_10619,N_10480,N_10323);
xnor U10620 (N_10620,N_10369,N_10466);
nand U10621 (N_10621,N_10415,N_10459);
nor U10622 (N_10622,N_10343,N_10456);
nor U10623 (N_10623,N_10256,N_10321);
or U10624 (N_10624,N_10361,N_10391);
or U10625 (N_10625,N_10424,N_10402);
and U10626 (N_10626,N_10384,N_10281);
and U10627 (N_10627,N_10487,N_10345);
and U10628 (N_10628,N_10295,N_10406);
nand U10629 (N_10629,N_10477,N_10480);
nor U10630 (N_10630,N_10421,N_10410);
and U10631 (N_10631,N_10429,N_10311);
nand U10632 (N_10632,N_10334,N_10308);
nor U10633 (N_10633,N_10497,N_10416);
or U10634 (N_10634,N_10378,N_10494);
nand U10635 (N_10635,N_10290,N_10414);
xor U10636 (N_10636,N_10399,N_10271);
or U10637 (N_10637,N_10251,N_10343);
and U10638 (N_10638,N_10455,N_10369);
and U10639 (N_10639,N_10359,N_10353);
nor U10640 (N_10640,N_10287,N_10274);
nor U10641 (N_10641,N_10466,N_10486);
nor U10642 (N_10642,N_10327,N_10304);
nand U10643 (N_10643,N_10486,N_10250);
or U10644 (N_10644,N_10475,N_10358);
nor U10645 (N_10645,N_10340,N_10335);
nand U10646 (N_10646,N_10253,N_10423);
nor U10647 (N_10647,N_10254,N_10415);
xor U10648 (N_10648,N_10400,N_10343);
nor U10649 (N_10649,N_10332,N_10456);
and U10650 (N_10650,N_10266,N_10289);
nor U10651 (N_10651,N_10403,N_10362);
xor U10652 (N_10652,N_10290,N_10453);
or U10653 (N_10653,N_10437,N_10482);
or U10654 (N_10654,N_10382,N_10473);
xnor U10655 (N_10655,N_10358,N_10483);
nand U10656 (N_10656,N_10278,N_10481);
nor U10657 (N_10657,N_10285,N_10309);
nor U10658 (N_10658,N_10471,N_10377);
or U10659 (N_10659,N_10423,N_10300);
and U10660 (N_10660,N_10468,N_10277);
nor U10661 (N_10661,N_10416,N_10473);
or U10662 (N_10662,N_10388,N_10441);
nor U10663 (N_10663,N_10318,N_10365);
nand U10664 (N_10664,N_10340,N_10327);
or U10665 (N_10665,N_10316,N_10408);
and U10666 (N_10666,N_10453,N_10282);
and U10667 (N_10667,N_10446,N_10496);
xor U10668 (N_10668,N_10425,N_10345);
and U10669 (N_10669,N_10452,N_10451);
and U10670 (N_10670,N_10312,N_10368);
nand U10671 (N_10671,N_10438,N_10472);
nand U10672 (N_10672,N_10399,N_10361);
or U10673 (N_10673,N_10476,N_10420);
nand U10674 (N_10674,N_10404,N_10285);
nor U10675 (N_10675,N_10411,N_10278);
xnor U10676 (N_10676,N_10283,N_10391);
xnor U10677 (N_10677,N_10499,N_10418);
xor U10678 (N_10678,N_10378,N_10318);
or U10679 (N_10679,N_10252,N_10286);
or U10680 (N_10680,N_10265,N_10327);
or U10681 (N_10681,N_10396,N_10437);
and U10682 (N_10682,N_10492,N_10447);
or U10683 (N_10683,N_10473,N_10440);
nand U10684 (N_10684,N_10423,N_10366);
and U10685 (N_10685,N_10382,N_10370);
and U10686 (N_10686,N_10390,N_10268);
and U10687 (N_10687,N_10339,N_10285);
and U10688 (N_10688,N_10274,N_10401);
nor U10689 (N_10689,N_10493,N_10400);
xor U10690 (N_10690,N_10370,N_10366);
nand U10691 (N_10691,N_10273,N_10252);
or U10692 (N_10692,N_10410,N_10449);
and U10693 (N_10693,N_10439,N_10402);
and U10694 (N_10694,N_10314,N_10293);
nand U10695 (N_10695,N_10412,N_10356);
nor U10696 (N_10696,N_10457,N_10411);
or U10697 (N_10697,N_10375,N_10487);
xor U10698 (N_10698,N_10314,N_10292);
and U10699 (N_10699,N_10405,N_10351);
xnor U10700 (N_10700,N_10279,N_10268);
nor U10701 (N_10701,N_10448,N_10263);
and U10702 (N_10702,N_10278,N_10378);
or U10703 (N_10703,N_10263,N_10353);
and U10704 (N_10704,N_10368,N_10285);
or U10705 (N_10705,N_10474,N_10398);
xnor U10706 (N_10706,N_10485,N_10304);
nand U10707 (N_10707,N_10458,N_10305);
nor U10708 (N_10708,N_10342,N_10446);
nor U10709 (N_10709,N_10400,N_10410);
xor U10710 (N_10710,N_10438,N_10254);
nand U10711 (N_10711,N_10340,N_10477);
nand U10712 (N_10712,N_10281,N_10280);
nor U10713 (N_10713,N_10402,N_10489);
and U10714 (N_10714,N_10425,N_10400);
and U10715 (N_10715,N_10379,N_10353);
and U10716 (N_10716,N_10256,N_10407);
xor U10717 (N_10717,N_10402,N_10256);
or U10718 (N_10718,N_10427,N_10285);
or U10719 (N_10719,N_10321,N_10449);
nand U10720 (N_10720,N_10490,N_10254);
and U10721 (N_10721,N_10321,N_10427);
nor U10722 (N_10722,N_10311,N_10460);
and U10723 (N_10723,N_10336,N_10470);
xor U10724 (N_10724,N_10283,N_10438);
nand U10725 (N_10725,N_10407,N_10263);
xnor U10726 (N_10726,N_10346,N_10478);
or U10727 (N_10727,N_10470,N_10253);
nand U10728 (N_10728,N_10335,N_10495);
or U10729 (N_10729,N_10282,N_10250);
nor U10730 (N_10730,N_10312,N_10303);
nor U10731 (N_10731,N_10473,N_10496);
and U10732 (N_10732,N_10497,N_10460);
nand U10733 (N_10733,N_10403,N_10296);
xor U10734 (N_10734,N_10327,N_10317);
and U10735 (N_10735,N_10474,N_10491);
nand U10736 (N_10736,N_10279,N_10280);
or U10737 (N_10737,N_10358,N_10383);
xnor U10738 (N_10738,N_10456,N_10259);
nor U10739 (N_10739,N_10311,N_10491);
and U10740 (N_10740,N_10330,N_10351);
nor U10741 (N_10741,N_10420,N_10392);
or U10742 (N_10742,N_10484,N_10320);
nand U10743 (N_10743,N_10396,N_10322);
and U10744 (N_10744,N_10441,N_10452);
or U10745 (N_10745,N_10416,N_10418);
xnor U10746 (N_10746,N_10368,N_10258);
and U10747 (N_10747,N_10461,N_10334);
or U10748 (N_10748,N_10358,N_10416);
nor U10749 (N_10749,N_10430,N_10412);
or U10750 (N_10750,N_10577,N_10658);
xor U10751 (N_10751,N_10598,N_10745);
nor U10752 (N_10752,N_10503,N_10548);
or U10753 (N_10753,N_10669,N_10648);
and U10754 (N_10754,N_10667,N_10518);
and U10755 (N_10755,N_10511,N_10689);
xor U10756 (N_10756,N_10501,N_10706);
nand U10757 (N_10757,N_10715,N_10678);
nor U10758 (N_10758,N_10543,N_10684);
nor U10759 (N_10759,N_10728,N_10544);
nand U10760 (N_10760,N_10614,N_10569);
and U10761 (N_10761,N_10583,N_10610);
nand U10762 (N_10762,N_10531,N_10609);
and U10763 (N_10763,N_10585,N_10714);
nor U10764 (N_10764,N_10661,N_10733);
xor U10765 (N_10765,N_10612,N_10718);
xnor U10766 (N_10766,N_10565,N_10743);
and U10767 (N_10767,N_10551,N_10505);
and U10768 (N_10768,N_10542,N_10742);
or U10769 (N_10769,N_10692,N_10712);
xnor U10770 (N_10770,N_10557,N_10508);
nor U10771 (N_10771,N_10560,N_10704);
and U10772 (N_10772,N_10504,N_10665);
or U10773 (N_10773,N_10520,N_10666);
and U10774 (N_10774,N_10663,N_10611);
nand U10775 (N_10775,N_10682,N_10516);
or U10776 (N_10776,N_10578,N_10748);
nor U10777 (N_10777,N_10563,N_10527);
or U10778 (N_10778,N_10693,N_10581);
and U10779 (N_10779,N_10539,N_10670);
nand U10780 (N_10780,N_10618,N_10708);
nand U10781 (N_10781,N_10677,N_10650);
nand U10782 (N_10782,N_10555,N_10685);
or U10783 (N_10783,N_10546,N_10559);
or U10784 (N_10784,N_10644,N_10696);
nand U10785 (N_10785,N_10637,N_10703);
nand U10786 (N_10786,N_10575,N_10639);
and U10787 (N_10787,N_10633,N_10587);
or U10788 (N_10788,N_10690,N_10683);
nor U10789 (N_10789,N_10720,N_10737);
xnor U10790 (N_10790,N_10605,N_10675);
and U10791 (N_10791,N_10584,N_10625);
and U10792 (N_10792,N_10564,N_10595);
or U10793 (N_10793,N_10739,N_10607);
xor U10794 (N_10794,N_10654,N_10573);
xnor U10795 (N_10795,N_10632,N_10635);
or U10796 (N_10796,N_10579,N_10619);
nor U10797 (N_10797,N_10655,N_10589);
nor U10798 (N_10798,N_10602,N_10710);
or U10799 (N_10799,N_10686,N_10738);
xor U10800 (N_10800,N_10652,N_10558);
xnor U10801 (N_10801,N_10588,N_10620);
xnor U10802 (N_10802,N_10731,N_10671);
xor U10803 (N_10803,N_10734,N_10532);
nor U10804 (N_10804,N_10594,N_10590);
and U10805 (N_10805,N_10681,N_10621);
and U10806 (N_10806,N_10561,N_10608);
or U10807 (N_10807,N_10550,N_10746);
nor U10808 (N_10808,N_10672,N_10736);
nor U10809 (N_10809,N_10660,N_10638);
nand U10810 (N_10810,N_10536,N_10626);
xnor U10811 (N_10811,N_10657,N_10599);
and U10812 (N_10812,N_10547,N_10524);
or U10813 (N_10813,N_10730,N_10519);
nand U10814 (N_10814,N_10534,N_10656);
nor U10815 (N_10815,N_10662,N_10735);
nor U10816 (N_10816,N_10562,N_10593);
nand U10817 (N_10817,N_10597,N_10641);
and U10818 (N_10818,N_10615,N_10568);
xor U10819 (N_10819,N_10721,N_10673);
and U10820 (N_10820,N_10507,N_10537);
and U10821 (N_10821,N_10512,N_10647);
nand U10822 (N_10822,N_10576,N_10687);
nand U10823 (N_10823,N_10521,N_10553);
and U10824 (N_10824,N_10727,N_10556);
xor U10825 (N_10825,N_10526,N_10749);
nand U10826 (N_10826,N_10740,N_10674);
nand U10827 (N_10827,N_10522,N_10566);
nand U10828 (N_10828,N_10567,N_10688);
nor U10829 (N_10829,N_10651,N_10523);
or U10830 (N_10830,N_10592,N_10645);
nand U10831 (N_10831,N_10617,N_10517);
and U10832 (N_10832,N_10747,N_10668);
nor U10833 (N_10833,N_10552,N_10634);
nand U10834 (N_10834,N_10525,N_10676);
xnor U10835 (N_10835,N_10659,N_10723);
nand U10836 (N_10836,N_10500,N_10741);
and U10837 (N_10837,N_10636,N_10570);
xnor U10838 (N_10838,N_10700,N_10699);
xor U10839 (N_10839,N_10646,N_10724);
and U10840 (N_10840,N_10535,N_10628);
nand U10841 (N_10841,N_10716,N_10515);
xor U10842 (N_10842,N_10600,N_10729);
and U10843 (N_10843,N_10580,N_10514);
nor U10844 (N_10844,N_10616,N_10627);
and U10845 (N_10845,N_10623,N_10719);
or U10846 (N_10846,N_10640,N_10586);
or U10847 (N_10847,N_10702,N_10722);
and U10848 (N_10848,N_10613,N_10606);
xor U10849 (N_10849,N_10506,N_10698);
nand U10850 (N_10850,N_10538,N_10691);
or U10851 (N_10851,N_10653,N_10629);
and U10852 (N_10852,N_10709,N_10631);
xor U10853 (N_10853,N_10622,N_10554);
nand U10854 (N_10854,N_10694,N_10697);
nand U10855 (N_10855,N_10717,N_10502);
or U10856 (N_10856,N_10574,N_10744);
xnor U10857 (N_10857,N_10732,N_10711);
nand U10858 (N_10858,N_10530,N_10571);
or U10859 (N_10859,N_10603,N_10649);
nor U10860 (N_10860,N_10713,N_10642);
and U10861 (N_10861,N_10510,N_10601);
and U10862 (N_10862,N_10705,N_10591);
and U10863 (N_10863,N_10549,N_10695);
nor U10864 (N_10864,N_10664,N_10726);
and U10865 (N_10865,N_10529,N_10509);
and U10866 (N_10866,N_10604,N_10596);
nor U10867 (N_10867,N_10679,N_10533);
and U10868 (N_10868,N_10680,N_10572);
nand U10869 (N_10869,N_10513,N_10528);
nand U10870 (N_10870,N_10624,N_10541);
xor U10871 (N_10871,N_10540,N_10582);
nor U10872 (N_10872,N_10701,N_10630);
nand U10873 (N_10873,N_10545,N_10725);
and U10874 (N_10874,N_10707,N_10643);
nor U10875 (N_10875,N_10595,N_10707);
or U10876 (N_10876,N_10632,N_10500);
nor U10877 (N_10877,N_10578,N_10661);
nand U10878 (N_10878,N_10660,N_10608);
nand U10879 (N_10879,N_10630,N_10716);
nor U10880 (N_10880,N_10539,N_10737);
xor U10881 (N_10881,N_10737,N_10596);
nor U10882 (N_10882,N_10577,N_10725);
nand U10883 (N_10883,N_10733,N_10557);
xor U10884 (N_10884,N_10612,N_10551);
nand U10885 (N_10885,N_10558,N_10677);
xnor U10886 (N_10886,N_10654,N_10663);
or U10887 (N_10887,N_10638,N_10564);
nand U10888 (N_10888,N_10655,N_10500);
nor U10889 (N_10889,N_10646,N_10637);
or U10890 (N_10890,N_10630,N_10535);
or U10891 (N_10891,N_10642,N_10521);
nand U10892 (N_10892,N_10648,N_10663);
and U10893 (N_10893,N_10635,N_10741);
or U10894 (N_10894,N_10605,N_10641);
or U10895 (N_10895,N_10641,N_10539);
or U10896 (N_10896,N_10512,N_10578);
or U10897 (N_10897,N_10580,N_10613);
nor U10898 (N_10898,N_10692,N_10662);
nand U10899 (N_10899,N_10528,N_10592);
xnor U10900 (N_10900,N_10667,N_10598);
nor U10901 (N_10901,N_10601,N_10693);
and U10902 (N_10902,N_10565,N_10580);
or U10903 (N_10903,N_10695,N_10689);
nor U10904 (N_10904,N_10506,N_10666);
nand U10905 (N_10905,N_10560,N_10631);
and U10906 (N_10906,N_10594,N_10691);
and U10907 (N_10907,N_10536,N_10628);
nor U10908 (N_10908,N_10636,N_10674);
nand U10909 (N_10909,N_10622,N_10658);
and U10910 (N_10910,N_10684,N_10731);
or U10911 (N_10911,N_10716,N_10601);
nand U10912 (N_10912,N_10736,N_10710);
nand U10913 (N_10913,N_10717,N_10623);
nor U10914 (N_10914,N_10530,N_10627);
and U10915 (N_10915,N_10542,N_10605);
or U10916 (N_10916,N_10690,N_10718);
and U10917 (N_10917,N_10701,N_10558);
nor U10918 (N_10918,N_10608,N_10569);
nor U10919 (N_10919,N_10535,N_10668);
or U10920 (N_10920,N_10699,N_10728);
nand U10921 (N_10921,N_10510,N_10676);
nand U10922 (N_10922,N_10691,N_10703);
and U10923 (N_10923,N_10513,N_10714);
xor U10924 (N_10924,N_10559,N_10507);
or U10925 (N_10925,N_10530,N_10589);
nor U10926 (N_10926,N_10736,N_10631);
nand U10927 (N_10927,N_10622,N_10643);
or U10928 (N_10928,N_10515,N_10633);
or U10929 (N_10929,N_10576,N_10645);
xnor U10930 (N_10930,N_10661,N_10675);
nand U10931 (N_10931,N_10580,N_10590);
nor U10932 (N_10932,N_10713,N_10614);
nand U10933 (N_10933,N_10598,N_10540);
nand U10934 (N_10934,N_10668,N_10745);
nor U10935 (N_10935,N_10724,N_10507);
nand U10936 (N_10936,N_10586,N_10712);
and U10937 (N_10937,N_10591,N_10638);
xnor U10938 (N_10938,N_10692,N_10554);
nor U10939 (N_10939,N_10697,N_10743);
and U10940 (N_10940,N_10539,N_10648);
xor U10941 (N_10941,N_10546,N_10715);
and U10942 (N_10942,N_10646,N_10657);
and U10943 (N_10943,N_10662,N_10541);
nand U10944 (N_10944,N_10560,N_10613);
xnor U10945 (N_10945,N_10508,N_10740);
xnor U10946 (N_10946,N_10596,N_10683);
xor U10947 (N_10947,N_10580,N_10673);
and U10948 (N_10948,N_10749,N_10624);
nor U10949 (N_10949,N_10576,N_10551);
and U10950 (N_10950,N_10670,N_10678);
nand U10951 (N_10951,N_10685,N_10500);
nor U10952 (N_10952,N_10573,N_10644);
xnor U10953 (N_10953,N_10705,N_10694);
nor U10954 (N_10954,N_10609,N_10535);
xor U10955 (N_10955,N_10742,N_10532);
nand U10956 (N_10956,N_10531,N_10697);
xor U10957 (N_10957,N_10556,N_10559);
or U10958 (N_10958,N_10654,N_10657);
nor U10959 (N_10959,N_10635,N_10515);
nand U10960 (N_10960,N_10649,N_10699);
nor U10961 (N_10961,N_10714,N_10592);
nand U10962 (N_10962,N_10639,N_10644);
nor U10963 (N_10963,N_10529,N_10576);
or U10964 (N_10964,N_10678,N_10608);
and U10965 (N_10965,N_10670,N_10542);
and U10966 (N_10966,N_10685,N_10560);
and U10967 (N_10967,N_10629,N_10656);
or U10968 (N_10968,N_10509,N_10559);
nand U10969 (N_10969,N_10665,N_10722);
or U10970 (N_10970,N_10534,N_10727);
or U10971 (N_10971,N_10645,N_10607);
xor U10972 (N_10972,N_10713,N_10674);
nand U10973 (N_10973,N_10509,N_10573);
xor U10974 (N_10974,N_10637,N_10649);
nand U10975 (N_10975,N_10603,N_10627);
and U10976 (N_10976,N_10688,N_10583);
and U10977 (N_10977,N_10608,N_10537);
nor U10978 (N_10978,N_10669,N_10744);
and U10979 (N_10979,N_10619,N_10608);
nor U10980 (N_10980,N_10622,N_10601);
xor U10981 (N_10981,N_10690,N_10624);
xor U10982 (N_10982,N_10655,N_10638);
nor U10983 (N_10983,N_10604,N_10526);
xnor U10984 (N_10984,N_10619,N_10749);
nand U10985 (N_10985,N_10692,N_10626);
and U10986 (N_10986,N_10507,N_10667);
nor U10987 (N_10987,N_10648,N_10692);
xor U10988 (N_10988,N_10616,N_10661);
or U10989 (N_10989,N_10563,N_10619);
or U10990 (N_10990,N_10744,N_10555);
or U10991 (N_10991,N_10621,N_10574);
nor U10992 (N_10992,N_10534,N_10583);
nand U10993 (N_10993,N_10641,N_10719);
xnor U10994 (N_10994,N_10645,N_10677);
and U10995 (N_10995,N_10538,N_10581);
nand U10996 (N_10996,N_10681,N_10533);
and U10997 (N_10997,N_10710,N_10720);
and U10998 (N_10998,N_10524,N_10540);
and U10999 (N_10999,N_10501,N_10679);
and U11000 (N_11000,N_10983,N_10917);
and U11001 (N_11001,N_10839,N_10848);
or U11002 (N_11002,N_10794,N_10928);
and U11003 (N_11003,N_10845,N_10957);
and U11004 (N_11004,N_10932,N_10945);
nand U11005 (N_11005,N_10900,N_10851);
nand U11006 (N_11006,N_10757,N_10925);
nand U11007 (N_11007,N_10986,N_10806);
and U11008 (N_11008,N_10860,N_10823);
and U11009 (N_11009,N_10956,N_10800);
xnor U11010 (N_11010,N_10871,N_10922);
and U11011 (N_11011,N_10758,N_10979);
xor U11012 (N_11012,N_10958,N_10993);
or U11013 (N_11013,N_10831,N_10943);
or U11014 (N_11014,N_10804,N_10942);
nand U11015 (N_11015,N_10841,N_10878);
nor U11016 (N_11016,N_10793,N_10809);
nand U11017 (N_11017,N_10760,N_10777);
or U11018 (N_11018,N_10852,N_10931);
nand U11019 (N_11019,N_10994,N_10797);
nor U11020 (N_11020,N_10818,N_10939);
or U11021 (N_11021,N_10781,N_10791);
nor U11022 (N_11022,N_10962,N_10888);
xor U11023 (N_11023,N_10837,N_10899);
and U11024 (N_11024,N_10768,N_10889);
xnor U11025 (N_11025,N_10886,N_10955);
and U11026 (N_11026,N_10775,N_10981);
xnor U11027 (N_11027,N_10952,N_10906);
nor U11028 (N_11028,N_10842,N_10798);
nor U11029 (N_11029,N_10950,N_10903);
or U11030 (N_11030,N_10897,N_10976);
or U11031 (N_11031,N_10905,N_10951);
and U11032 (N_11032,N_10868,N_10808);
xnor U11033 (N_11033,N_10918,N_10773);
and U11034 (N_11034,N_10762,N_10884);
nand U11035 (N_11035,N_10829,N_10991);
xnor U11036 (N_11036,N_10916,N_10980);
and U11037 (N_11037,N_10990,N_10813);
or U11038 (N_11038,N_10850,N_10894);
nor U11039 (N_11039,N_10778,N_10985);
xnor U11040 (N_11040,N_10834,N_10914);
xnor U11041 (N_11041,N_10796,N_10862);
or U11042 (N_11042,N_10828,N_10946);
nand U11043 (N_11043,N_10998,N_10859);
xor U11044 (N_11044,N_10812,N_10966);
and U11045 (N_11045,N_10814,N_10937);
xor U11046 (N_11046,N_10774,N_10959);
nand U11047 (N_11047,N_10915,N_10953);
or U11048 (N_11048,N_10861,N_10787);
or U11049 (N_11049,N_10938,N_10934);
nor U11050 (N_11050,N_10904,N_10987);
nor U11051 (N_11051,N_10876,N_10854);
and U11052 (N_11052,N_10929,N_10896);
or U11053 (N_11053,N_10795,N_10927);
xor U11054 (N_11054,N_10961,N_10909);
or U11055 (N_11055,N_10867,N_10750);
or U11056 (N_11056,N_10954,N_10844);
xnor U11057 (N_11057,N_10965,N_10941);
xor U11058 (N_11058,N_10963,N_10754);
and U11059 (N_11059,N_10866,N_10835);
and U11060 (N_11060,N_10920,N_10996);
and U11061 (N_11061,N_10790,N_10995);
xnor U11062 (N_11062,N_10870,N_10944);
nor U11063 (N_11063,N_10857,N_10856);
nor U11064 (N_11064,N_10902,N_10765);
and U11065 (N_11065,N_10817,N_10924);
nand U11066 (N_11066,N_10849,N_10752);
nor U11067 (N_11067,N_10893,N_10891);
or U11068 (N_11068,N_10820,N_10973);
xor U11069 (N_11069,N_10877,N_10913);
nor U11070 (N_11070,N_10982,N_10788);
and U11071 (N_11071,N_10949,N_10799);
nor U11072 (N_11072,N_10948,N_10780);
and U11073 (N_11073,N_10971,N_10826);
nor U11074 (N_11074,N_10838,N_10833);
nand U11075 (N_11075,N_10978,N_10907);
xnor U11076 (N_11076,N_10970,N_10771);
xnor U11077 (N_11077,N_10853,N_10974);
xor U11078 (N_11078,N_10881,N_10759);
xor U11079 (N_11079,N_10807,N_10989);
nand U11080 (N_11080,N_10769,N_10821);
nor U11081 (N_11081,N_10782,N_10910);
or U11082 (N_11082,N_10975,N_10824);
or U11083 (N_11083,N_10764,N_10885);
nor U11084 (N_11084,N_10873,N_10936);
nand U11085 (N_11085,N_10882,N_10865);
nand U11086 (N_11086,N_10783,N_10815);
or U11087 (N_11087,N_10977,N_10776);
nor U11088 (N_11088,N_10840,N_10912);
xor U11089 (N_11089,N_10761,N_10969);
or U11090 (N_11090,N_10803,N_10858);
or U11091 (N_11091,N_10830,N_10811);
nor U11092 (N_11092,N_10827,N_10947);
nor U11093 (N_11093,N_10935,N_10872);
xnor U11094 (N_11094,N_10836,N_10772);
or U11095 (N_11095,N_10864,N_10802);
nor U11096 (N_11096,N_10846,N_10869);
nand U11097 (N_11097,N_10874,N_10786);
xor U11098 (N_11098,N_10898,N_10919);
or U11099 (N_11099,N_10960,N_10847);
or U11100 (N_11100,N_10789,N_10940);
and U11101 (N_11101,N_10766,N_10972);
or U11102 (N_11102,N_10816,N_10887);
and U11103 (N_11103,N_10855,N_10923);
nor U11104 (N_11104,N_10753,N_10892);
and U11105 (N_11105,N_10968,N_10895);
nor U11106 (N_11106,N_10801,N_10911);
nand U11107 (N_11107,N_10984,N_10767);
and U11108 (N_11108,N_10810,N_10832);
nand U11109 (N_11109,N_10779,N_10926);
xnor U11110 (N_11110,N_10921,N_10822);
nand U11111 (N_11111,N_10908,N_10825);
xor U11112 (N_11112,N_10784,N_10863);
nand U11113 (N_11113,N_10964,N_10879);
or U11114 (N_11114,N_10819,N_10843);
nand U11115 (N_11115,N_10875,N_10763);
xor U11116 (N_11116,N_10933,N_10792);
xor U11117 (N_11117,N_10999,N_10756);
or U11118 (N_11118,N_10930,N_10883);
and U11119 (N_11119,N_10997,N_10901);
and U11120 (N_11120,N_10992,N_10890);
or U11121 (N_11121,N_10770,N_10751);
nand U11122 (N_11122,N_10880,N_10805);
or U11123 (N_11123,N_10967,N_10785);
nand U11124 (N_11124,N_10755,N_10988);
and U11125 (N_11125,N_10785,N_10784);
and U11126 (N_11126,N_10917,N_10877);
or U11127 (N_11127,N_10942,N_10956);
xor U11128 (N_11128,N_10872,N_10986);
and U11129 (N_11129,N_10874,N_10892);
xnor U11130 (N_11130,N_10985,N_10974);
and U11131 (N_11131,N_10855,N_10904);
xnor U11132 (N_11132,N_10819,N_10902);
and U11133 (N_11133,N_10829,N_10893);
nand U11134 (N_11134,N_10825,N_10946);
or U11135 (N_11135,N_10948,N_10754);
and U11136 (N_11136,N_10813,N_10982);
xnor U11137 (N_11137,N_10962,N_10801);
or U11138 (N_11138,N_10782,N_10945);
and U11139 (N_11139,N_10891,N_10998);
xnor U11140 (N_11140,N_10934,N_10854);
or U11141 (N_11141,N_10819,N_10895);
nor U11142 (N_11142,N_10886,N_10938);
nand U11143 (N_11143,N_10884,N_10768);
or U11144 (N_11144,N_10993,N_10961);
and U11145 (N_11145,N_10877,N_10850);
or U11146 (N_11146,N_10921,N_10928);
nand U11147 (N_11147,N_10998,N_10830);
xnor U11148 (N_11148,N_10790,N_10869);
nor U11149 (N_11149,N_10999,N_10853);
xor U11150 (N_11150,N_10791,N_10895);
nand U11151 (N_11151,N_10873,N_10920);
nand U11152 (N_11152,N_10830,N_10789);
or U11153 (N_11153,N_10892,N_10952);
nand U11154 (N_11154,N_10839,N_10963);
xnor U11155 (N_11155,N_10787,N_10945);
or U11156 (N_11156,N_10988,N_10817);
nor U11157 (N_11157,N_10836,N_10804);
nor U11158 (N_11158,N_10947,N_10934);
or U11159 (N_11159,N_10889,N_10814);
or U11160 (N_11160,N_10813,N_10752);
nor U11161 (N_11161,N_10753,N_10927);
and U11162 (N_11162,N_10903,N_10949);
nor U11163 (N_11163,N_10841,N_10799);
xnor U11164 (N_11164,N_10772,N_10901);
nand U11165 (N_11165,N_10805,N_10915);
and U11166 (N_11166,N_10760,N_10996);
nor U11167 (N_11167,N_10758,N_10796);
xnor U11168 (N_11168,N_10921,N_10824);
nand U11169 (N_11169,N_10995,N_10872);
xnor U11170 (N_11170,N_10811,N_10769);
nor U11171 (N_11171,N_10938,N_10829);
and U11172 (N_11172,N_10991,N_10885);
nand U11173 (N_11173,N_10969,N_10889);
xor U11174 (N_11174,N_10770,N_10965);
nor U11175 (N_11175,N_10976,N_10783);
or U11176 (N_11176,N_10956,N_10782);
or U11177 (N_11177,N_10931,N_10813);
xor U11178 (N_11178,N_10824,N_10907);
nor U11179 (N_11179,N_10978,N_10910);
nor U11180 (N_11180,N_10971,N_10806);
xnor U11181 (N_11181,N_10757,N_10955);
nand U11182 (N_11182,N_10977,N_10886);
xor U11183 (N_11183,N_10762,N_10901);
nor U11184 (N_11184,N_10888,N_10925);
nor U11185 (N_11185,N_10950,N_10901);
and U11186 (N_11186,N_10844,N_10895);
or U11187 (N_11187,N_10996,N_10879);
nor U11188 (N_11188,N_10783,N_10839);
nor U11189 (N_11189,N_10775,N_10794);
nor U11190 (N_11190,N_10938,N_10968);
and U11191 (N_11191,N_10932,N_10786);
xor U11192 (N_11192,N_10764,N_10910);
or U11193 (N_11193,N_10977,N_10842);
or U11194 (N_11194,N_10776,N_10823);
and U11195 (N_11195,N_10861,N_10939);
or U11196 (N_11196,N_10803,N_10761);
or U11197 (N_11197,N_10876,N_10799);
nand U11198 (N_11198,N_10852,N_10770);
nor U11199 (N_11199,N_10857,N_10984);
nand U11200 (N_11200,N_10974,N_10886);
nor U11201 (N_11201,N_10935,N_10877);
nand U11202 (N_11202,N_10955,N_10937);
xnor U11203 (N_11203,N_10932,N_10878);
xor U11204 (N_11204,N_10816,N_10753);
nor U11205 (N_11205,N_10772,N_10916);
or U11206 (N_11206,N_10938,N_10952);
nand U11207 (N_11207,N_10808,N_10975);
nand U11208 (N_11208,N_10925,N_10879);
nor U11209 (N_11209,N_10840,N_10985);
nor U11210 (N_11210,N_10757,N_10831);
or U11211 (N_11211,N_10822,N_10823);
and U11212 (N_11212,N_10926,N_10956);
xor U11213 (N_11213,N_10984,N_10975);
xor U11214 (N_11214,N_10783,N_10789);
xor U11215 (N_11215,N_10896,N_10846);
xor U11216 (N_11216,N_10756,N_10947);
xnor U11217 (N_11217,N_10882,N_10919);
and U11218 (N_11218,N_10926,N_10984);
nand U11219 (N_11219,N_10965,N_10848);
or U11220 (N_11220,N_10978,N_10817);
xnor U11221 (N_11221,N_10756,N_10803);
xor U11222 (N_11222,N_10798,N_10759);
nor U11223 (N_11223,N_10874,N_10875);
xor U11224 (N_11224,N_10923,N_10862);
and U11225 (N_11225,N_10845,N_10956);
nor U11226 (N_11226,N_10793,N_10919);
and U11227 (N_11227,N_10888,N_10804);
nor U11228 (N_11228,N_10866,N_10990);
and U11229 (N_11229,N_10968,N_10866);
or U11230 (N_11230,N_10783,N_10872);
nand U11231 (N_11231,N_10814,N_10807);
nand U11232 (N_11232,N_10890,N_10940);
nand U11233 (N_11233,N_10874,N_10850);
and U11234 (N_11234,N_10915,N_10851);
nand U11235 (N_11235,N_10783,N_10952);
nor U11236 (N_11236,N_10901,N_10929);
and U11237 (N_11237,N_10850,N_10820);
nor U11238 (N_11238,N_10836,N_10997);
and U11239 (N_11239,N_10832,N_10938);
or U11240 (N_11240,N_10777,N_10926);
or U11241 (N_11241,N_10821,N_10954);
and U11242 (N_11242,N_10994,N_10939);
xnor U11243 (N_11243,N_10809,N_10846);
and U11244 (N_11244,N_10752,N_10967);
xor U11245 (N_11245,N_10978,N_10820);
nor U11246 (N_11246,N_10943,N_10974);
and U11247 (N_11247,N_10965,N_10759);
nor U11248 (N_11248,N_10865,N_10813);
nor U11249 (N_11249,N_10830,N_10941);
nand U11250 (N_11250,N_11035,N_11186);
nand U11251 (N_11251,N_11234,N_11166);
or U11252 (N_11252,N_11167,N_11165);
nand U11253 (N_11253,N_11066,N_11136);
nand U11254 (N_11254,N_11081,N_11156);
and U11255 (N_11255,N_11192,N_11087);
nand U11256 (N_11256,N_11162,N_11021);
xor U11257 (N_11257,N_11005,N_11086);
or U11258 (N_11258,N_11188,N_11172);
or U11259 (N_11259,N_11152,N_11109);
or U11260 (N_11260,N_11230,N_11213);
and U11261 (N_11261,N_11033,N_11044);
nand U11262 (N_11262,N_11198,N_11052);
nand U11263 (N_11263,N_11204,N_11113);
or U11264 (N_11264,N_11106,N_11013);
or U11265 (N_11265,N_11110,N_11229);
nand U11266 (N_11266,N_11088,N_11043);
nand U11267 (N_11267,N_11148,N_11080);
or U11268 (N_11268,N_11182,N_11134);
and U11269 (N_11269,N_11037,N_11050);
or U11270 (N_11270,N_11190,N_11155);
nand U11271 (N_11271,N_11111,N_11246);
or U11272 (N_11272,N_11040,N_11057);
xnor U11273 (N_11273,N_11239,N_11144);
and U11274 (N_11274,N_11116,N_11107);
nor U11275 (N_11275,N_11158,N_11220);
and U11276 (N_11276,N_11170,N_11130);
xnor U11277 (N_11277,N_11059,N_11224);
nand U11278 (N_11278,N_11211,N_11024);
or U11279 (N_11279,N_11048,N_11245);
xnor U11280 (N_11280,N_11221,N_11233);
nor U11281 (N_11281,N_11053,N_11014);
xnor U11282 (N_11282,N_11092,N_11058);
nor U11283 (N_11283,N_11120,N_11199);
xnor U11284 (N_11284,N_11098,N_11159);
or U11285 (N_11285,N_11191,N_11184);
xnor U11286 (N_11286,N_11138,N_11197);
or U11287 (N_11287,N_11002,N_11225);
xor U11288 (N_11288,N_11029,N_11232);
xor U11289 (N_11289,N_11183,N_11179);
nor U11290 (N_11290,N_11085,N_11164);
nand U11291 (N_11291,N_11031,N_11222);
or U11292 (N_11292,N_11101,N_11026);
nand U11293 (N_11293,N_11163,N_11124);
xnor U11294 (N_11294,N_11215,N_11042);
xor U11295 (N_11295,N_11147,N_11151);
xor U11296 (N_11296,N_11032,N_11030);
nor U11297 (N_11297,N_11028,N_11169);
and U11298 (N_11298,N_11209,N_11056);
and U11299 (N_11299,N_11006,N_11160);
nor U11300 (N_11300,N_11034,N_11196);
nor U11301 (N_11301,N_11011,N_11063);
nand U11302 (N_11302,N_11016,N_11076);
and U11303 (N_11303,N_11047,N_11001);
nor U11304 (N_11304,N_11149,N_11214);
xor U11305 (N_11305,N_11127,N_11126);
and U11306 (N_11306,N_11150,N_11062);
or U11307 (N_11307,N_11038,N_11089);
and U11308 (N_11308,N_11157,N_11025);
nor U11309 (N_11309,N_11242,N_11114);
nand U11310 (N_11310,N_11175,N_11228);
nor U11311 (N_11311,N_11119,N_11243);
nor U11312 (N_11312,N_11096,N_11223);
xor U11313 (N_11313,N_11212,N_11015);
xor U11314 (N_11314,N_11105,N_11200);
nand U11315 (N_11315,N_11174,N_11065);
nor U11316 (N_11316,N_11054,N_11100);
nor U11317 (N_11317,N_11128,N_11210);
and U11318 (N_11318,N_11168,N_11181);
nand U11319 (N_11319,N_11131,N_11073);
or U11320 (N_11320,N_11041,N_11123);
nor U11321 (N_11321,N_11061,N_11208);
and U11322 (N_11322,N_11241,N_11143);
or U11323 (N_11323,N_11115,N_11012);
nand U11324 (N_11324,N_11187,N_11008);
nor U11325 (N_11325,N_11132,N_11248);
xnor U11326 (N_11326,N_11046,N_11146);
nor U11327 (N_11327,N_11231,N_11099);
xor U11328 (N_11328,N_11064,N_11010);
nand U11329 (N_11329,N_11205,N_11071);
and U11330 (N_11330,N_11083,N_11102);
and U11331 (N_11331,N_11129,N_11216);
nor U11332 (N_11332,N_11218,N_11009);
nand U11333 (N_11333,N_11000,N_11018);
and U11334 (N_11334,N_11017,N_11079);
or U11335 (N_11335,N_11074,N_11090);
nand U11336 (N_11336,N_11135,N_11139);
and U11337 (N_11337,N_11121,N_11173);
or U11338 (N_11338,N_11118,N_11019);
xor U11339 (N_11339,N_11133,N_11180);
and U11340 (N_11340,N_11206,N_11078);
nor U11341 (N_11341,N_11249,N_11070);
nor U11342 (N_11342,N_11226,N_11091);
nand U11343 (N_11343,N_11072,N_11171);
and U11344 (N_11344,N_11244,N_11176);
nor U11345 (N_11345,N_11145,N_11161);
nand U11346 (N_11346,N_11003,N_11084);
xnor U11347 (N_11347,N_11142,N_11240);
xor U11348 (N_11348,N_11140,N_11238);
xnor U11349 (N_11349,N_11108,N_11022);
nand U11350 (N_11350,N_11051,N_11117);
or U11351 (N_11351,N_11045,N_11219);
or U11352 (N_11352,N_11194,N_11068);
nor U11353 (N_11353,N_11039,N_11077);
or U11354 (N_11354,N_11247,N_11082);
nor U11355 (N_11355,N_11201,N_11235);
xnor U11356 (N_11356,N_11023,N_11097);
xor U11357 (N_11357,N_11075,N_11178);
or U11358 (N_11358,N_11153,N_11203);
nor U11359 (N_11359,N_11236,N_11193);
xnor U11360 (N_11360,N_11217,N_11237);
nand U11361 (N_11361,N_11122,N_11195);
nor U11362 (N_11362,N_11004,N_11137);
nand U11363 (N_11363,N_11036,N_11125);
xnor U11364 (N_11364,N_11007,N_11093);
nor U11365 (N_11365,N_11227,N_11177);
or U11366 (N_11366,N_11067,N_11095);
xnor U11367 (N_11367,N_11094,N_11189);
nor U11368 (N_11368,N_11141,N_11049);
nor U11369 (N_11369,N_11202,N_11185);
nand U11370 (N_11370,N_11069,N_11103);
nor U11371 (N_11371,N_11020,N_11027);
xor U11372 (N_11372,N_11154,N_11207);
nand U11373 (N_11373,N_11104,N_11055);
xnor U11374 (N_11374,N_11060,N_11112);
and U11375 (N_11375,N_11218,N_11021);
or U11376 (N_11376,N_11130,N_11212);
and U11377 (N_11377,N_11094,N_11074);
nand U11378 (N_11378,N_11104,N_11205);
or U11379 (N_11379,N_11232,N_11229);
nor U11380 (N_11380,N_11140,N_11059);
or U11381 (N_11381,N_11236,N_11042);
xor U11382 (N_11382,N_11069,N_11175);
xor U11383 (N_11383,N_11012,N_11041);
or U11384 (N_11384,N_11244,N_11017);
and U11385 (N_11385,N_11201,N_11011);
xor U11386 (N_11386,N_11054,N_11101);
nand U11387 (N_11387,N_11014,N_11077);
or U11388 (N_11388,N_11117,N_11193);
xor U11389 (N_11389,N_11004,N_11009);
or U11390 (N_11390,N_11228,N_11212);
nand U11391 (N_11391,N_11225,N_11027);
and U11392 (N_11392,N_11026,N_11247);
and U11393 (N_11393,N_11021,N_11070);
nand U11394 (N_11394,N_11032,N_11119);
and U11395 (N_11395,N_11123,N_11097);
nor U11396 (N_11396,N_11004,N_11057);
nand U11397 (N_11397,N_11056,N_11170);
and U11398 (N_11398,N_11227,N_11044);
nand U11399 (N_11399,N_11220,N_11069);
nor U11400 (N_11400,N_11049,N_11004);
nor U11401 (N_11401,N_11171,N_11110);
nor U11402 (N_11402,N_11227,N_11214);
nor U11403 (N_11403,N_11109,N_11209);
and U11404 (N_11404,N_11000,N_11052);
and U11405 (N_11405,N_11139,N_11171);
and U11406 (N_11406,N_11044,N_11050);
or U11407 (N_11407,N_11103,N_11106);
and U11408 (N_11408,N_11016,N_11144);
nor U11409 (N_11409,N_11026,N_11200);
and U11410 (N_11410,N_11140,N_11013);
xor U11411 (N_11411,N_11231,N_11235);
or U11412 (N_11412,N_11168,N_11093);
xor U11413 (N_11413,N_11203,N_11021);
or U11414 (N_11414,N_11204,N_11082);
and U11415 (N_11415,N_11124,N_11207);
or U11416 (N_11416,N_11027,N_11006);
xor U11417 (N_11417,N_11045,N_11074);
or U11418 (N_11418,N_11221,N_11042);
xor U11419 (N_11419,N_11039,N_11199);
or U11420 (N_11420,N_11148,N_11179);
nor U11421 (N_11421,N_11041,N_11224);
or U11422 (N_11422,N_11243,N_11174);
or U11423 (N_11423,N_11173,N_11183);
nand U11424 (N_11424,N_11210,N_11228);
nand U11425 (N_11425,N_11098,N_11105);
xnor U11426 (N_11426,N_11099,N_11235);
and U11427 (N_11427,N_11132,N_11025);
and U11428 (N_11428,N_11131,N_11097);
and U11429 (N_11429,N_11163,N_11179);
xor U11430 (N_11430,N_11181,N_11215);
nand U11431 (N_11431,N_11034,N_11112);
nand U11432 (N_11432,N_11153,N_11212);
or U11433 (N_11433,N_11211,N_11121);
or U11434 (N_11434,N_11007,N_11186);
nor U11435 (N_11435,N_11070,N_11024);
xor U11436 (N_11436,N_11024,N_11025);
xor U11437 (N_11437,N_11068,N_11190);
nand U11438 (N_11438,N_11060,N_11017);
or U11439 (N_11439,N_11122,N_11212);
nor U11440 (N_11440,N_11141,N_11067);
or U11441 (N_11441,N_11050,N_11234);
and U11442 (N_11442,N_11212,N_11211);
and U11443 (N_11443,N_11187,N_11117);
nand U11444 (N_11444,N_11027,N_11217);
or U11445 (N_11445,N_11215,N_11045);
or U11446 (N_11446,N_11172,N_11040);
or U11447 (N_11447,N_11185,N_11165);
and U11448 (N_11448,N_11028,N_11098);
or U11449 (N_11449,N_11198,N_11214);
nor U11450 (N_11450,N_11179,N_11171);
nor U11451 (N_11451,N_11039,N_11204);
and U11452 (N_11452,N_11023,N_11148);
nor U11453 (N_11453,N_11064,N_11142);
nor U11454 (N_11454,N_11246,N_11123);
nand U11455 (N_11455,N_11132,N_11181);
and U11456 (N_11456,N_11041,N_11223);
nor U11457 (N_11457,N_11040,N_11232);
nand U11458 (N_11458,N_11158,N_11058);
and U11459 (N_11459,N_11060,N_11124);
nor U11460 (N_11460,N_11102,N_11118);
xnor U11461 (N_11461,N_11217,N_11185);
nand U11462 (N_11462,N_11049,N_11187);
or U11463 (N_11463,N_11094,N_11192);
or U11464 (N_11464,N_11184,N_11211);
or U11465 (N_11465,N_11102,N_11214);
nand U11466 (N_11466,N_11104,N_11046);
xor U11467 (N_11467,N_11032,N_11182);
and U11468 (N_11468,N_11011,N_11077);
xnor U11469 (N_11469,N_11130,N_11109);
nand U11470 (N_11470,N_11062,N_11201);
xnor U11471 (N_11471,N_11112,N_11063);
nand U11472 (N_11472,N_11101,N_11177);
xor U11473 (N_11473,N_11014,N_11046);
or U11474 (N_11474,N_11109,N_11017);
nand U11475 (N_11475,N_11025,N_11126);
nor U11476 (N_11476,N_11099,N_11200);
xor U11477 (N_11477,N_11223,N_11216);
or U11478 (N_11478,N_11087,N_11171);
and U11479 (N_11479,N_11197,N_11117);
nand U11480 (N_11480,N_11109,N_11095);
nand U11481 (N_11481,N_11069,N_11222);
and U11482 (N_11482,N_11094,N_11118);
nand U11483 (N_11483,N_11000,N_11234);
nand U11484 (N_11484,N_11035,N_11005);
and U11485 (N_11485,N_11145,N_11046);
nand U11486 (N_11486,N_11161,N_11159);
and U11487 (N_11487,N_11142,N_11068);
xnor U11488 (N_11488,N_11147,N_11243);
and U11489 (N_11489,N_11079,N_11131);
or U11490 (N_11490,N_11089,N_11166);
xor U11491 (N_11491,N_11045,N_11085);
nor U11492 (N_11492,N_11090,N_11133);
xor U11493 (N_11493,N_11049,N_11203);
or U11494 (N_11494,N_11124,N_11023);
and U11495 (N_11495,N_11241,N_11166);
and U11496 (N_11496,N_11091,N_11220);
xnor U11497 (N_11497,N_11086,N_11062);
and U11498 (N_11498,N_11226,N_11184);
xnor U11499 (N_11499,N_11068,N_11111);
nand U11500 (N_11500,N_11316,N_11466);
xor U11501 (N_11501,N_11490,N_11359);
and U11502 (N_11502,N_11312,N_11492);
nand U11503 (N_11503,N_11433,N_11300);
xor U11504 (N_11504,N_11352,N_11351);
or U11505 (N_11505,N_11487,N_11313);
or U11506 (N_11506,N_11323,N_11317);
and U11507 (N_11507,N_11315,N_11325);
nor U11508 (N_11508,N_11346,N_11419);
xor U11509 (N_11509,N_11395,N_11473);
xor U11510 (N_11510,N_11496,N_11471);
nor U11511 (N_11511,N_11498,N_11398);
and U11512 (N_11512,N_11274,N_11371);
nor U11513 (N_11513,N_11399,N_11376);
or U11514 (N_11514,N_11286,N_11299);
xor U11515 (N_11515,N_11354,N_11463);
and U11516 (N_11516,N_11361,N_11397);
xnor U11517 (N_11517,N_11423,N_11430);
or U11518 (N_11518,N_11409,N_11307);
xnor U11519 (N_11519,N_11332,N_11362);
nor U11520 (N_11520,N_11318,N_11445);
or U11521 (N_11521,N_11436,N_11497);
xor U11522 (N_11522,N_11278,N_11385);
and U11523 (N_11523,N_11277,N_11266);
nand U11524 (N_11524,N_11309,N_11339);
or U11525 (N_11525,N_11365,N_11413);
or U11526 (N_11526,N_11292,N_11418);
or U11527 (N_11527,N_11306,N_11401);
nor U11528 (N_11528,N_11368,N_11464);
nand U11529 (N_11529,N_11402,N_11459);
nor U11530 (N_11530,N_11265,N_11333);
or U11531 (N_11531,N_11404,N_11453);
or U11532 (N_11532,N_11485,N_11457);
or U11533 (N_11533,N_11448,N_11355);
and U11534 (N_11534,N_11383,N_11481);
nand U11535 (N_11535,N_11322,N_11386);
nor U11536 (N_11536,N_11415,N_11373);
nand U11537 (N_11537,N_11469,N_11435);
and U11538 (N_11538,N_11343,N_11293);
and U11539 (N_11539,N_11282,N_11304);
nand U11540 (N_11540,N_11478,N_11456);
and U11541 (N_11541,N_11375,N_11405);
nor U11542 (N_11542,N_11480,N_11314);
or U11543 (N_11543,N_11328,N_11334);
xnor U11544 (N_11544,N_11428,N_11283);
or U11545 (N_11545,N_11431,N_11414);
or U11546 (N_11546,N_11421,N_11252);
or U11547 (N_11547,N_11380,N_11408);
nand U11548 (N_11548,N_11310,N_11336);
or U11549 (N_11549,N_11285,N_11444);
or U11550 (N_11550,N_11337,N_11482);
nor U11551 (N_11551,N_11451,N_11450);
nand U11552 (N_11552,N_11389,N_11489);
nand U11553 (N_11553,N_11484,N_11429);
nand U11554 (N_11554,N_11446,N_11297);
and U11555 (N_11555,N_11449,N_11454);
and U11556 (N_11556,N_11338,N_11363);
and U11557 (N_11557,N_11356,N_11372);
or U11558 (N_11558,N_11335,N_11384);
nor U11559 (N_11559,N_11342,N_11479);
or U11560 (N_11560,N_11390,N_11488);
xor U11561 (N_11561,N_11493,N_11253);
or U11562 (N_11562,N_11281,N_11358);
and U11563 (N_11563,N_11269,N_11483);
nor U11564 (N_11564,N_11440,N_11259);
nor U11565 (N_11565,N_11442,N_11258);
nand U11566 (N_11566,N_11319,N_11261);
or U11567 (N_11567,N_11329,N_11400);
xor U11568 (N_11568,N_11324,N_11374);
and U11569 (N_11569,N_11452,N_11290);
and U11570 (N_11570,N_11308,N_11460);
and U11571 (N_11571,N_11364,N_11289);
xnor U11572 (N_11572,N_11391,N_11382);
and U11573 (N_11573,N_11294,N_11251);
and U11574 (N_11574,N_11296,N_11331);
nand U11575 (N_11575,N_11416,N_11392);
or U11576 (N_11576,N_11393,N_11465);
nor U11577 (N_11577,N_11271,N_11321);
and U11578 (N_11578,N_11369,N_11284);
nand U11579 (N_11579,N_11438,N_11461);
and U11580 (N_11580,N_11260,N_11357);
xnor U11581 (N_11581,N_11275,N_11437);
nor U11582 (N_11582,N_11467,N_11475);
xor U11583 (N_11583,N_11345,N_11494);
and U11584 (N_11584,N_11256,N_11360);
xnor U11585 (N_11585,N_11458,N_11311);
and U11586 (N_11586,N_11353,N_11447);
nor U11587 (N_11587,N_11476,N_11491);
nand U11588 (N_11588,N_11341,N_11381);
xor U11589 (N_11589,N_11303,N_11254);
and U11590 (N_11590,N_11330,N_11427);
nor U11591 (N_11591,N_11347,N_11406);
nand U11592 (N_11592,N_11417,N_11267);
nand U11593 (N_11593,N_11366,N_11407);
nor U11594 (N_11594,N_11378,N_11302);
xor U11595 (N_11595,N_11326,N_11268);
nand U11596 (N_11596,N_11441,N_11250);
nor U11597 (N_11597,N_11411,N_11387);
xnor U11598 (N_11598,N_11377,N_11474);
and U11599 (N_11599,N_11305,N_11470);
and U11600 (N_11600,N_11379,N_11495);
or U11601 (N_11601,N_11410,N_11396);
nor U11602 (N_11602,N_11301,N_11426);
nor U11603 (N_11603,N_11486,N_11298);
xnor U11604 (N_11604,N_11462,N_11349);
nand U11605 (N_11605,N_11270,N_11272);
xor U11606 (N_11606,N_11422,N_11412);
nand U11607 (N_11607,N_11499,N_11420);
nor U11608 (N_11608,N_11287,N_11273);
nor U11609 (N_11609,N_11472,N_11344);
nor U11610 (N_11610,N_11348,N_11327);
xnor U11611 (N_11611,N_11477,N_11280);
xor U11612 (N_11612,N_11455,N_11394);
or U11613 (N_11613,N_11424,N_11425);
or U11614 (N_11614,N_11295,N_11255);
or U11615 (N_11615,N_11276,N_11403);
nor U11616 (N_11616,N_11443,N_11370);
nand U11617 (N_11617,N_11291,N_11388);
nand U11618 (N_11618,N_11263,N_11468);
and U11619 (N_11619,N_11432,N_11320);
and U11620 (N_11620,N_11288,N_11262);
nand U11621 (N_11621,N_11279,N_11257);
and U11622 (N_11622,N_11439,N_11340);
nor U11623 (N_11623,N_11350,N_11434);
and U11624 (N_11624,N_11367,N_11264);
nor U11625 (N_11625,N_11401,N_11389);
nor U11626 (N_11626,N_11477,N_11273);
xor U11627 (N_11627,N_11483,N_11389);
or U11628 (N_11628,N_11369,N_11458);
nor U11629 (N_11629,N_11276,N_11349);
nor U11630 (N_11630,N_11491,N_11403);
nor U11631 (N_11631,N_11295,N_11332);
nor U11632 (N_11632,N_11331,N_11493);
and U11633 (N_11633,N_11337,N_11335);
xor U11634 (N_11634,N_11430,N_11252);
nand U11635 (N_11635,N_11439,N_11357);
nor U11636 (N_11636,N_11390,N_11418);
or U11637 (N_11637,N_11344,N_11358);
or U11638 (N_11638,N_11440,N_11469);
xor U11639 (N_11639,N_11305,N_11345);
nor U11640 (N_11640,N_11451,N_11318);
or U11641 (N_11641,N_11310,N_11369);
or U11642 (N_11642,N_11419,N_11305);
xor U11643 (N_11643,N_11278,N_11496);
or U11644 (N_11644,N_11469,N_11495);
nor U11645 (N_11645,N_11311,N_11359);
nor U11646 (N_11646,N_11423,N_11344);
nor U11647 (N_11647,N_11277,N_11355);
xnor U11648 (N_11648,N_11379,N_11474);
xnor U11649 (N_11649,N_11463,N_11406);
and U11650 (N_11650,N_11416,N_11321);
and U11651 (N_11651,N_11342,N_11333);
nor U11652 (N_11652,N_11497,N_11261);
xnor U11653 (N_11653,N_11443,N_11321);
nand U11654 (N_11654,N_11427,N_11402);
xor U11655 (N_11655,N_11351,N_11425);
or U11656 (N_11656,N_11253,N_11431);
xnor U11657 (N_11657,N_11260,N_11261);
nor U11658 (N_11658,N_11405,N_11388);
and U11659 (N_11659,N_11395,N_11270);
xnor U11660 (N_11660,N_11356,N_11476);
or U11661 (N_11661,N_11371,N_11361);
nand U11662 (N_11662,N_11318,N_11447);
nand U11663 (N_11663,N_11269,N_11287);
or U11664 (N_11664,N_11359,N_11279);
and U11665 (N_11665,N_11450,N_11374);
nand U11666 (N_11666,N_11352,N_11296);
nand U11667 (N_11667,N_11458,N_11471);
and U11668 (N_11668,N_11316,N_11309);
xor U11669 (N_11669,N_11308,N_11477);
and U11670 (N_11670,N_11460,N_11333);
nand U11671 (N_11671,N_11492,N_11319);
or U11672 (N_11672,N_11422,N_11298);
xnor U11673 (N_11673,N_11468,N_11398);
nand U11674 (N_11674,N_11401,N_11469);
and U11675 (N_11675,N_11291,N_11380);
nand U11676 (N_11676,N_11433,N_11338);
nor U11677 (N_11677,N_11481,N_11392);
nor U11678 (N_11678,N_11327,N_11295);
nor U11679 (N_11679,N_11314,N_11458);
nand U11680 (N_11680,N_11295,N_11497);
or U11681 (N_11681,N_11369,N_11427);
xor U11682 (N_11682,N_11471,N_11490);
nor U11683 (N_11683,N_11352,N_11420);
xnor U11684 (N_11684,N_11259,N_11373);
xnor U11685 (N_11685,N_11318,N_11418);
nand U11686 (N_11686,N_11386,N_11444);
or U11687 (N_11687,N_11410,N_11491);
and U11688 (N_11688,N_11474,N_11273);
and U11689 (N_11689,N_11352,N_11329);
and U11690 (N_11690,N_11260,N_11332);
and U11691 (N_11691,N_11281,N_11465);
xor U11692 (N_11692,N_11484,N_11268);
xor U11693 (N_11693,N_11477,N_11326);
xnor U11694 (N_11694,N_11335,N_11386);
nor U11695 (N_11695,N_11371,N_11427);
nand U11696 (N_11696,N_11469,N_11423);
nand U11697 (N_11697,N_11446,N_11385);
and U11698 (N_11698,N_11361,N_11320);
or U11699 (N_11699,N_11307,N_11300);
nor U11700 (N_11700,N_11338,N_11405);
nand U11701 (N_11701,N_11295,N_11265);
or U11702 (N_11702,N_11418,N_11473);
or U11703 (N_11703,N_11253,N_11311);
or U11704 (N_11704,N_11471,N_11327);
and U11705 (N_11705,N_11457,N_11466);
nand U11706 (N_11706,N_11346,N_11325);
nand U11707 (N_11707,N_11468,N_11412);
xnor U11708 (N_11708,N_11481,N_11302);
xnor U11709 (N_11709,N_11415,N_11263);
nor U11710 (N_11710,N_11475,N_11308);
or U11711 (N_11711,N_11344,N_11293);
xnor U11712 (N_11712,N_11351,N_11370);
and U11713 (N_11713,N_11484,N_11272);
xor U11714 (N_11714,N_11481,N_11443);
nor U11715 (N_11715,N_11405,N_11420);
xnor U11716 (N_11716,N_11374,N_11462);
nor U11717 (N_11717,N_11314,N_11360);
nor U11718 (N_11718,N_11336,N_11330);
xnor U11719 (N_11719,N_11458,N_11327);
nand U11720 (N_11720,N_11447,N_11346);
xnor U11721 (N_11721,N_11333,N_11310);
or U11722 (N_11722,N_11361,N_11253);
or U11723 (N_11723,N_11418,N_11342);
or U11724 (N_11724,N_11366,N_11420);
or U11725 (N_11725,N_11470,N_11330);
xnor U11726 (N_11726,N_11431,N_11376);
or U11727 (N_11727,N_11299,N_11259);
xor U11728 (N_11728,N_11403,N_11429);
xor U11729 (N_11729,N_11262,N_11351);
nand U11730 (N_11730,N_11435,N_11437);
nor U11731 (N_11731,N_11480,N_11350);
or U11732 (N_11732,N_11419,N_11298);
nand U11733 (N_11733,N_11250,N_11447);
or U11734 (N_11734,N_11492,N_11264);
nor U11735 (N_11735,N_11373,N_11442);
nor U11736 (N_11736,N_11260,N_11339);
nand U11737 (N_11737,N_11312,N_11389);
xor U11738 (N_11738,N_11433,N_11381);
nand U11739 (N_11739,N_11343,N_11302);
xor U11740 (N_11740,N_11268,N_11264);
nand U11741 (N_11741,N_11381,N_11387);
or U11742 (N_11742,N_11359,N_11402);
and U11743 (N_11743,N_11262,N_11356);
nor U11744 (N_11744,N_11459,N_11349);
and U11745 (N_11745,N_11467,N_11417);
nand U11746 (N_11746,N_11342,N_11313);
nor U11747 (N_11747,N_11270,N_11302);
or U11748 (N_11748,N_11465,N_11412);
xnor U11749 (N_11749,N_11362,N_11347);
nor U11750 (N_11750,N_11532,N_11571);
nor U11751 (N_11751,N_11624,N_11573);
xnor U11752 (N_11752,N_11697,N_11583);
nand U11753 (N_11753,N_11601,N_11568);
nor U11754 (N_11754,N_11739,N_11678);
and U11755 (N_11755,N_11691,N_11591);
nor U11756 (N_11756,N_11710,N_11588);
or U11757 (N_11757,N_11673,N_11689);
or U11758 (N_11758,N_11577,N_11633);
and U11759 (N_11759,N_11546,N_11749);
or U11760 (N_11760,N_11562,N_11623);
nor U11761 (N_11761,N_11614,N_11617);
xnor U11762 (N_11762,N_11555,N_11664);
or U11763 (N_11763,N_11535,N_11662);
and U11764 (N_11764,N_11629,N_11669);
nor U11765 (N_11765,N_11722,N_11742);
and U11766 (N_11766,N_11730,N_11626);
xor U11767 (N_11767,N_11675,N_11533);
or U11768 (N_11768,N_11637,N_11732);
xnor U11769 (N_11769,N_11728,N_11696);
and U11770 (N_11770,N_11744,N_11699);
or U11771 (N_11771,N_11642,N_11709);
xnor U11772 (N_11772,N_11738,N_11582);
or U11773 (N_11773,N_11719,N_11702);
and U11774 (N_11774,N_11656,N_11580);
nand U11775 (N_11775,N_11594,N_11708);
or U11776 (N_11776,N_11565,N_11586);
or U11777 (N_11777,N_11654,N_11745);
xor U11778 (N_11778,N_11505,N_11578);
nor U11779 (N_11779,N_11639,N_11552);
xor U11780 (N_11780,N_11590,N_11646);
and U11781 (N_11781,N_11519,N_11541);
or U11782 (N_11782,N_11747,N_11530);
nand U11783 (N_11783,N_11721,N_11714);
xnor U11784 (N_11784,N_11641,N_11701);
nand U11785 (N_11785,N_11706,N_11598);
nor U11786 (N_11786,N_11581,N_11584);
nor U11787 (N_11787,N_11660,N_11631);
nand U11788 (N_11788,N_11680,N_11523);
nand U11789 (N_11789,N_11632,N_11608);
nor U11790 (N_11790,N_11525,N_11677);
and U11791 (N_11791,N_11652,N_11516);
xnor U11792 (N_11792,N_11687,N_11544);
and U11793 (N_11793,N_11585,N_11645);
or U11794 (N_11794,N_11558,N_11727);
nand U11795 (N_11795,N_11597,N_11566);
nor U11796 (N_11796,N_11574,N_11653);
xor U11797 (N_11797,N_11550,N_11606);
nor U11798 (N_11798,N_11686,N_11703);
or U11799 (N_11799,N_11647,N_11735);
and U11800 (N_11800,N_11715,N_11743);
nand U11801 (N_11801,N_11640,N_11746);
or U11802 (N_11802,N_11683,N_11644);
nor U11803 (N_11803,N_11684,N_11511);
nand U11804 (N_11804,N_11643,N_11713);
and U11805 (N_11805,N_11723,N_11539);
nor U11806 (N_11806,N_11542,N_11502);
nand U11807 (N_11807,N_11726,N_11627);
and U11808 (N_11808,N_11634,N_11599);
nand U11809 (N_11809,N_11508,N_11720);
and U11810 (N_11810,N_11693,N_11668);
nor U11811 (N_11811,N_11538,N_11649);
xnor U11812 (N_11812,N_11567,N_11572);
nor U11813 (N_11813,N_11672,N_11579);
nand U11814 (N_11814,N_11587,N_11717);
xnor U11815 (N_11815,N_11712,N_11504);
nand U11816 (N_11816,N_11651,N_11724);
and U11817 (N_11817,N_11524,N_11589);
or U11818 (N_11818,N_11537,N_11635);
xnor U11819 (N_11819,N_11681,N_11501);
xnor U11820 (N_11820,N_11540,N_11548);
and U11821 (N_11821,N_11700,N_11618);
nand U11822 (N_11822,N_11671,N_11619);
nor U11823 (N_11823,N_11718,N_11625);
or U11824 (N_11824,N_11564,N_11575);
nand U11825 (N_11825,N_11518,N_11685);
nor U11826 (N_11826,N_11513,N_11650);
and U11827 (N_11827,N_11622,N_11613);
nor U11828 (N_11828,N_11688,N_11522);
nand U11829 (N_11829,N_11521,N_11596);
or U11830 (N_11830,N_11570,N_11615);
or U11831 (N_11831,N_11545,N_11657);
nor U11832 (N_11832,N_11725,N_11698);
and U11833 (N_11833,N_11682,N_11534);
nand U11834 (N_11834,N_11741,N_11512);
and U11835 (N_11835,N_11733,N_11520);
or U11836 (N_11836,N_11704,N_11561);
nand U11837 (N_11837,N_11729,N_11648);
and U11838 (N_11838,N_11517,N_11569);
or U11839 (N_11839,N_11500,N_11616);
nand U11840 (N_11840,N_11557,N_11705);
nor U11841 (N_11841,N_11554,N_11665);
xor U11842 (N_11842,N_11560,N_11630);
or U11843 (N_11843,N_11576,N_11551);
nor U11844 (N_11844,N_11663,N_11559);
xor U11845 (N_11845,N_11731,N_11628);
or U11846 (N_11846,N_11604,N_11603);
nor U11847 (N_11847,N_11612,N_11531);
nand U11848 (N_11848,N_11607,N_11610);
nor U11849 (N_11849,N_11602,N_11593);
nand U11850 (N_11850,N_11667,N_11611);
and U11851 (N_11851,N_11692,N_11621);
and U11852 (N_11852,N_11670,N_11507);
and U11853 (N_11853,N_11658,N_11528);
xnor U11854 (N_11854,N_11716,N_11514);
or U11855 (N_11855,N_11506,N_11636);
nand U11856 (N_11856,N_11620,N_11543);
and U11857 (N_11857,N_11515,N_11736);
nor U11858 (N_11858,N_11674,N_11659);
or U11859 (N_11859,N_11536,N_11609);
nand U11860 (N_11860,N_11695,N_11592);
or U11861 (N_11861,N_11509,N_11600);
nand U11862 (N_11862,N_11638,N_11679);
nor U11863 (N_11863,N_11547,N_11553);
nand U11864 (N_11864,N_11655,N_11737);
xor U11865 (N_11865,N_11595,N_11503);
and U11866 (N_11866,N_11527,N_11690);
xor U11867 (N_11867,N_11605,N_11661);
nand U11868 (N_11868,N_11748,N_11707);
nand U11869 (N_11869,N_11666,N_11556);
nand U11870 (N_11870,N_11711,N_11529);
nor U11871 (N_11871,N_11676,N_11510);
or U11872 (N_11872,N_11563,N_11549);
nand U11873 (N_11873,N_11526,N_11694);
or U11874 (N_11874,N_11740,N_11734);
and U11875 (N_11875,N_11612,N_11623);
nor U11876 (N_11876,N_11588,N_11693);
or U11877 (N_11877,N_11719,N_11562);
nor U11878 (N_11878,N_11700,N_11650);
xnor U11879 (N_11879,N_11561,N_11596);
nand U11880 (N_11880,N_11700,N_11722);
and U11881 (N_11881,N_11628,N_11551);
nor U11882 (N_11882,N_11688,N_11649);
nand U11883 (N_11883,N_11635,N_11678);
or U11884 (N_11884,N_11691,N_11510);
or U11885 (N_11885,N_11714,N_11588);
or U11886 (N_11886,N_11555,N_11578);
nor U11887 (N_11887,N_11721,N_11712);
nand U11888 (N_11888,N_11696,N_11522);
nor U11889 (N_11889,N_11645,N_11745);
nand U11890 (N_11890,N_11704,N_11668);
xnor U11891 (N_11891,N_11639,N_11572);
nor U11892 (N_11892,N_11676,N_11627);
and U11893 (N_11893,N_11598,N_11654);
xor U11894 (N_11894,N_11523,N_11629);
xnor U11895 (N_11895,N_11540,N_11693);
or U11896 (N_11896,N_11509,N_11622);
nand U11897 (N_11897,N_11603,N_11707);
nor U11898 (N_11898,N_11530,N_11679);
xnor U11899 (N_11899,N_11717,N_11500);
or U11900 (N_11900,N_11628,N_11525);
nor U11901 (N_11901,N_11596,N_11688);
nand U11902 (N_11902,N_11721,N_11677);
nand U11903 (N_11903,N_11526,N_11665);
or U11904 (N_11904,N_11522,N_11732);
or U11905 (N_11905,N_11701,N_11637);
nand U11906 (N_11906,N_11736,N_11627);
and U11907 (N_11907,N_11550,N_11705);
nand U11908 (N_11908,N_11675,N_11680);
or U11909 (N_11909,N_11662,N_11537);
nor U11910 (N_11910,N_11618,N_11698);
nand U11911 (N_11911,N_11730,N_11648);
nand U11912 (N_11912,N_11516,N_11631);
nor U11913 (N_11913,N_11545,N_11644);
nor U11914 (N_11914,N_11511,N_11527);
and U11915 (N_11915,N_11726,N_11569);
nand U11916 (N_11916,N_11599,N_11566);
xnor U11917 (N_11917,N_11516,N_11640);
and U11918 (N_11918,N_11744,N_11729);
and U11919 (N_11919,N_11528,N_11672);
xor U11920 (N_11920,N_11526,N_11707);
or U11921 (N_11921,N_11584,N_11748);
nor U11922 (N_11922,N_11600,N_11664);
xnor U11923 (N_11923,N_11578,N_11607);
or U11924 (N_11924,N_11647,N_11533);
xor U11925 (N_11925,N_11702,N_11628);
or U11926 (N_11926,N_11538,N_11527);
xor U11927 (N_11927,N_11508,N_11645);
or U11928 (N_11928,N_11508,N_11620);
nor U11929 (N_11929,N_11568,N_11583);
or U11930 (N_11930,N_11675,N_11711);
xor U11931 (N_11931,N_11568,N_11728);
or U11932 (N_11932,N_11701,N_11523);
and U11933 (N_11933,N_11748,N_11736);
nand U11934 (N_11934,N_11694,N_11622);
and U11935 (N_11935,N_11610,N_11743);
nor U11936 (N_11936,N_11721,N_11651);
xor U11937 (N_11937,N_11551,N_11746);
nor U11938 (N_11938,N_11542,N_11603);
nand U11939 (N_11939,N_11665,N_11620);
or U11940 (N_11940,N_11538,N_11563);
nand U11941 (N_11941,N_11675,N_11710);
or U11942 (N_11942,N_11679,N_11534);
or U11943 (N_11943,N_11527,N_11643);
nor U11944 (N_11944,N_11731,N_11676);
xor U11945 (N_11945,N_11514,N_11510);
nor U11946 (N_11946,N_11634,N_11693);
xor U11947 (N_11947,N_11612,N_11572);
xor U11948 (N_11948,N_11614,N_11615);
xor U11949 (N_11949,N_11721,N_11681);
or U11950 (N_11950,N_11599,N_11742);
xnor U11951 (N_11951,N_11592,N_11677);
or U11952 (N_11952,N_11647,N_11634);
or U11953 (N_11953,N_11517,N_11718);
or U11954 (N_11954,N_11632,N_11527);
or U11955 (N_11955,N_11684,N_11729);
or U11956 (N_11956,N_11725,N_11531);
nor U11957 (N_11957,N_11594,N_11592);
nor U11958 (N_11958,N_11522,N_11667);
or U11959 (N_11959,N_11629,N_11655);
xor U11960 (N_11960,N_11748,N_11659);
or U11961 (N_11961,N_11516,N_11698);
xnor U11962 (N_11962,N_11663,N_11719);
nor U11963 (N_11963,N_11737,N_11675);
nand U11964 (N_11964,N_11577,N_11524);
xnor U11965 (N_11965,N_11665,N_11643);
or U11966 (N_11966,N_11706,N_11687);
or U11967 (N_11967,N_11664,N_11554);
xnor U11968 (N_11968,N_11606,N_11694);
nand U11969 (N_11969,N_11664,N_11696);
xnor U11970 (N_11970,N_11708,N_11635);
nor U11971 (N_11971,N_11734,N_11534);
xor U11972 (N_11972,N_11721,N_11615);
nor U11973 (N_11973,N_11660,N_11732);
or U11974 (N_11974,N_11577,N_11727);
nand U11975 (N_11975,N_11702,N_11505);
xnor U11976 (N_11976,N_11655,N_11735);
xor U11977 (N_11977,N_11607,N_11723);
nand U11978 (N_11978,N_11679,N_11736);
nand U11979 (N_11979,N_11516,N_11685);
xnor U11980 (N_11980,N_11593,N_11677);
nor U11981 (N_11981,N_11556,N_11520);
xnor U11982 (N_11982,N_11718,N_11558);
nor U11983 (N_11983,N_11684,N_11664);
nor U11984 (N_11984,N_11609,N_11735);
or U11985 (N_11985,N_11610,N_11565);
xnor U11986 (N_11986,N_11697,N_11520);
nor U11987 (N_11987,N_11704,N_11555);
and U11988 (N_11988,N_11626,N_11549);
xor U11989 (N_11989,N_11670,N_11721);
or U11990 (N_11990,N_11677,N_11507);
xor U11991 (N_11991,N_11714,N_11587);
nand U11992 (N_11992,N_11626,N_11661);
nand U11993 (N_11993,N_11650,N_11693);
nor U11994 (N_11994,N_11648,N_11662);
or U11995 (N_11995,N_11539,N_11685);
xnor U11996 (N_11996,N_11555,N_11613);
nand U11997 (N_11997,N_11524,N_11739);
xnor U11998 (N_11998,N_11631,N_11566);
nor U11999 (N_11999,N_11652,N_11570);
xnor U12000 (N_12000,N_11887,N_11865);
nor U12001 (N_12001,N_11871,N_11774);
nor U12002 (N_12002,N_11772,N_11898);
or U12003 (N_12003,N_11799,N_11927);
or U12004 (N_12004,N_11833,N_11994);
or U12005 (N_12005,N_11852,N_11775);
xor U12006 (N_12006,N_11832,N_11998);
nor U12007 (N_12007,N_11925,N_11924);
or U12008 (N_12008,N_11753,N_11883);
or U12009 (N_12009,N_11837,N_11913);
nand U12010 (N_12010,N_11860,N_11894);
nand U12011 (N_12011,N_11769,N_11829);
nor U12012 (N_12012,N_11768,N_11945);
xor U12013 (N_12013,N_11784,N_11970);
and U12014 (N_12014,N_11979,N_11773);
xor U12015 (N_12015,N_11943,N_11877);
xor U12016 (N_12016,N_11941,N_11848);
xnor U12017 (N_12017,N_11880,N_11912);
nand U12018 (N_12018,N_11940,N_11757);
and U12019 (N_12019,N_11891,N_11870);
nor U12020 (N_12020,N_11752,N_11878);
xnor U12021 (N_12021,N_11886,N_11964);
nor U12022 (N_12022,N_11845,N_11782);
nand U12023 (N_12023,N_11750,N_11934);
nor U12024 (N_12024,N_11914,N_11817);
nand U12025 (N_12025,N_11956,N_11786);
and U12026 (N_12026,N_11758,N_11858);
or U12027 (N_12027,N_11787,N_11791);
and U12028 (N_12028,N_11826,N_11864);
or U12029 (N_12029,N_11897,N_11806);
nand U12030 (N_12030,N_11900,N_11946);
nor U12031 (N_12031,N_11893,N_11770);
or U12032 (N_12032,N_11780,N_11819);
xor U12033 (N_12033,N_11882,N_11908);
nand U12034 (N_12034,N_11969,N_11831);
nand U12035 (N_12035,N_11954,N_11890);
xor U12036 (N_12036,N_11944,N_11947);
or U12037 (N_12037,N_11781,N_11844);
nand U12038 (N_12038,N_11932,N_11960);
and U12039 (N_12039,N_11821,N_11754);
xor U12040 (N_12040,N_11955,N_11997);
or U12041 (N_12041,N_11972,N_11926);
xor U12042 (N_12042,N_11804,N_11899);
nand U12043 (N_12043,N_11763,N_11910);
and U12044 (N_12044,N_11834,N_11884);
or U12045 (N_12045,N_11835,N_11915);
xor U12046 (N_12046,N_11885,N_11974);
nor U12047 (N_12047,N_11823,N_11902);
xor U12048 (N_12048,N_11958,N_11755);
xnor U12049 (N_12049,N_11987,N_11777);
and U12050 (N_12050,N_11963,N_11760);
or U12051 (N_12051,N_11983,N_11857);
or U12052 (N_12052,N_11901,N_11856);
and U12053 (N_12053,N_11982,N_11978);
or U12054 (N_12054,N_11935,N_11850);
or U12055 (N_12055,N_11805,N_11977);
xor U12056 (N_12056,N_11921,N_11948);
nand U12057 (N_12057,N_11779,N_11793);
nand U12058 (N_12058,N_11869,N_11996);
nor U12059 (N_12059,N_11896,N_11989);
or U12060 (N_12060,N_11965,N_11991);
xor U12061 (N_12061,N_11942,N_11846);
and U12062 (N_12062,N_11807,N_11797);
or U12063 (N_12063,N_11872,N_11930);
and U12064 (N_12064,N_11881,N_11811);
xnor U12065 (N_12065,N_11933,N_11973);
nand U12066 (N_12066,N_11790,N_11875);
xor U12067 (N_12067,N_11962,N_11971);
or U12068 (N_12068,N_11892,N_11756);
nand U12069 (N_12069,N_11838,N_11929);
nand U12070 (N_12070,N_11868,N_11928);
nor U12071 (N_12071,N_11854,N_11789);
nor U12072 (N_12072,N_11859,N_11767);
nor U12073 (N_12073,N_11820,N_11938);
and U12074 (N_12074,N_11889,N_11866);
nand U12075 (N_12075,N_11939,N_11751);
nor U12076 (N_12076,N_11847,N_11808);
or U12077 (N_12077,N_11761,N_11814);
xnor U12078 (N_12078,N_11810,N_11861);
and U12079 (N_12079,N_11839,N_11909);
nand U12080 (N_12080,N_11794,N_11950);
xor U12081 (N_12081,N_11825,N_11798);
nand U12082 (N_12082,N_11931,N_11764);
or U12083 (N_12083,N_11842,N_11917);
nor U12084 (N_12084,N_11813,N_11984);
nor U12085 (N_12085,N_11959,N_11952);
or U12086 (N_12086,N_11995,N_11968);
nand U12087 (N_12087,N_11936,N_11836);
and U12088 (N_12088,N_11796,N_11803);
or U12089 (N_12089,N_11762,N_11822);
nand U12090 (N_12090,N_11766,N_11841);
and U12091 (N_12091,N_11874,N_11853);
and U12092 (N_12092,N_11862,N_11855);
or U12093 (N_12093,N_11795,N_11771);
and U12094 (N_12094,N_11975,N_11778);
or U12095 (N_12095,N_11949,N_11905);
or U12096 (N_12096,N_11785,N_11792);
and U12097 (N_12097,N_11776,N_11999);
nand U12098 (N_12098,N_11920,N_11867);
xnor U12099 (N_12099,N_11985,N_11863);
xor U12100 (N_12100,N_11919,N_11953);
or U12101 (N_12101,N_11992,N_11843);
and U12102 (N_12102,N_11923,N_11873);
xor U12103 (N_12103,N_11827,N_11876);
nand U12104 (N_12104,N_11922,N_11759);
xor U12105 (N_12105,N_11818,N_11976);
xor U12106 (N_12106,N_11937,N_11840);
and U12107 (N_12107,N_11903,N_11809);
xor U12108 (N_12108,N_11906,N_11812);
xor U12109 (N_12109,N_11961,N_11824);
nor U12110 (N_12110,N_11765,N_11904);
xnor U12111 (N_12111,N_11907,N_11788);
or U12112 (N_12112,N_11851,N_11888);
and U12113 (N_12113,N_11800,N_11828);
xor U12114 (N_12114,N_11980,N_11816);
or U12115 (N_12115,N_11966,N_11988);
and U12116 (N_12116,N_11911,N_11895);
nor U12117 (N_12117,N_11801,N_11830);
or U12118 (N_12118,N_11916,N_11879);
and U12119 (N_12119,N_11918,N_11802);
or U12120 (N_12120,N_11957,N_11849);
or U12121 (N_12121,N_11783,N_11981);
xor U12122 (N_12122,N_11986,N_11990);
xnor U12123 (N_12123,N_11951,N_11815);
nand U12124 (N_12124,N_11967,N_11993);
and U12125 (N_12125,N_11878,N_11982);
nor U12126 (N_12126,N_11843,N_11994);
and U12127 (N_12127,N_11774,N_11970);
or U12128 (N_12128,N_11801,N_11888);
and U12129 (N_12129,N_11912,N_11873);
nor U12130 (N_12130,N_11967,N_11920);
nand U12131 (N_12131,N_11989,N_11982);
xor U12132 (N_12132,N_11896,N_11946);
or U12133 (N_12133,N_11983,N_11968);
nand U12134 (N_12134,N_11945,N_11943);
nand U12135 (N_12135,N_11846,N_11936);
xnor U12136 (N_12136,N_11895,N_11819);
nor U12137 (N_12137,N_11767,N_11970);
nand U12138 (N_12138,N_11901,N_11774);
nand U12139 (N_12139,N_11978,N_11996);
xor U12140 (N_12140,N_11792,N_11974);
nor U12141 (N_12141,N_11929,N_11977);
xor U12142 (N_12142,N_11919,N_11949);
nand U12143 (N_12143,N_11967,N_11927);
nand U12144 (N_12144,N_11911,N_11773);
nand U12145 (N_12145,N_11952,N_11907);
nand U12146 (N_12146,N_11861,N_11779);
nand U12147 (N_12147,N_11824,N_11987);
nand U12148 (N_12148,N_11755,N_11886);
and U12149 (N_12149,N_11794,N_11769);
nor U12150 (N_12150,N_11852,N_11870);
nand U12151 (N_12151,N_11788,N_11898);
xnor U12152 (N_12152,N_11793,N_11970);
nand U12153 (N_12153,N_11784,N_11998);
or U12154 (N_12154,N_11802,N_11850);
nand U12155 (N_12155,N_11970,N_11873);
xor U12156 (N_12156,N_11860,N_11825);
xnor U12157 (N_12157,N_11787,N_11912);
nand U12158 (N_12158,N_11851,N_11790);
xor U12159 (N_12159,N_11951,N_11905);
xor U12160 (N_12160,N_11854,N_11824);
nand U12161 (N_12161,N_11776,N_11784);
nand U12162 (N_12162,N_11823,N_11960);
nor U12163 (N_12163,N_11926,N_11889);
nor U12164 (N_12164,N_11897,N_11993);
or U12165 (N_12165,N_11828,N_11752);
and U12166 (N_12166,N_11840,N_11925);
or U12167 (N_12167,N_11914,N_11841);
or U12168 (N_12168,N_11995,N_11911);
nor U12169 (N_12169,N_11943,N_11983);
nor U12170 (N_12170,N_11764,N_11932);
xnor U12171 (N_12171,N_11961,N_11919);
and U12172 (N_12172,N_11785,N_11827);
nand U12173 (N_12173,N_11845,N_11885);
xnor U12174 (N_12174,N_11893,N_11899);
nor U12175 (N_12175,N_11936,N_11903);
or U12176 (N_12176,N_11945,N_11850);
and U12177 (N_12177,N_11791,N_11771);
xor U12178 (N_12178,N_11814,N_11912);
or U12179 (N_12179,N_11959,N_11889);
nor U12180 (N_12180,N_11883,N_11948);
nor U12181 (N_12181,N_11932,N_11996);
and U12182 (N_12182,N_11984,N_11922);
or U12183 (N_12183,N_11856,N_11835);
nor U12184 (N_12184,N_11837,N_11791);
and U12185 (N_12185,N_11836,N_11764);
nand U12186 (N_12186,N_11901,N_11988);
nand U12187 (N_12187,N_11782,N_11857);
xor U12188 (N_12188,N_11776,N_11992);
and U12189 (N_12189,N_11994,N_11954);
and U12190 (N_12190,N_11754,N_11825);
xnor U12191 (N_12191,N_11881,N_11835);
xor U12192 (N_12192,N_11862,N_11952);
and U12193 (N_12193,N_11928,N_11896);
and U12194 (N_12194,N_11907,N_11938);
or U12195 (N_12195,N_11885,N_11812);
xnor U12196 (N_12196,N_11833,N_11863);
nand U12197 (N_12197,N_11909,N_11981);
and U12198 (N_12198,N_11959,N_11769);
nor U12199 (N_12199,N_11917,N_11888);
nand U12200 (N_12200,N_11973,N_11805);
and U12201 (N_12201,N_11973,N_11955);
xnor U12202 (N_12202,N_11951,N_11853);
or U12203 (N_12203,N_11865,N_11812);
nor U12204 (N_12204,N_11977,N_11872);
or U12205 (N_12205,N_11823,N_11759);
and U12206 (N_12206,N_11958,N_11794);
and U12207 (N_12207,N_11953,N_11751);
xor U12208 (N_12208,N_11905,N_11918);
nor U12209 (N_12209,N_11786,N_11959);
xnor U12210 (N_12210,N_11805,N_11758);
nor U12211 (N_12211,N_11924,N_11906);
nor U12212 (N_12212,N_11903,N_11944);
xor U12213 (N_12213,N_11912,N_11939);
and U12214 (N_12214,N_11819,N_11801);
nand U12215 (N_12215,N_11810,N_11769);
xor U12216 (N_12216,N_11876,N_11959);
nand U12217 (N_12217,N_11901,N_11903);
or U12218 (N_12218,N_11838,N_11880);
xnor U12219 (N_12219,N_11807,N_11784);
nor U12220 (N_12220,N_11988,N_11938);
nand U12221 (N_12221,N_11761,N_11953);
and U12222 (N_12222,N_11937,N_11798);
nand U12223 (N_12223,N_11790,N_11823);
or U12224 (N_12224,N_11926,N_11873);
and U12225 (N_12225,N_11950,N_11880);
nor U12226 (N_12226,N_11975,N_11940);
nand U12227 (N_12227,N_11833,N_11775);
nor U12228 (N_12228,N_11757,N_11789);
and U12229 (N_12229,N_11925,N_11752);
or U12230 (N_12230,N_11916,N_11948);
or U12231 (N_12231,N_11761,N_11930);
xor U12232 (N_12232,N_11985,N_11917);
xnor U12233 (N_12233,N_11908,N_11793);
or U12234 (N_12234,N_11946,N_11801);
xor U12235 (N_12235,N_11826,N_11909);
and U12236 (N_12236,N_11852,N_11769);
or U12237 (N_12237,N_11867,N_11947);
or U12238 (N_12238,N_11902,N_11830);
or U12239 (N_12239,N_11820,N_11890);
nor U12240 (N_12240,N_11799,N_11796);
nand U12241 (N_12241,N_11790,N_11921);
nor U12242 (N_12242,N_11885,N_11957);
and U12243 (N_12243,N_11835,N_11791);
and U12244 (N_12244,N_11909,N_11975);
or U12245 (N_12245,N_11779,N_11873);
and U12246 (N_12246,N_11912,N_11997);
and U12247 (N_12247,N_11874,N_11847);
or U12248 (N_12248,N_11865,N_11894);
nand U12249 (N_12249,N_11765,N_11914);
nor U12250 (N_12250,N_12150,N_12054);
xnor U12251 (N_12251,N_12249,N_12130);
and U12252 (N_12252,N_12180,N_12203);
or U12253 (N_12253,N_12061,N_12233);
nand U12254 (N_12254,N_12078,N_12072);
nor U12255 (N_12255,N_12107,N_12163);
nand U12256 (N_12256,N_12147,N_12079);
nor U12257 (N_12257,N_12029,N_12143);
or U12258 (N_12258,N_12189,N_12223);
or U12259 (N_12259,N_12148,N_12243);
or U12260 (N_12260,N_12099,N_12036);
nor U12261 (N_12261,N_12020,N_12097);
nand U12262 (N_12262,N_12067,N_12214);
xor U12263 (N_12263,N_12226,N_12169);
and U12264 (N_12264,N_12083,N_12100);
nand U12265 (N_12265,N_12191,N_12154);
nor U12266 (N_12266,N_12155,N_12216);
xor U12267 (N_12267,N_12207,N_12140);
xnor U12268 (N_12268,N_12094,N_12239);
and U12269 (N_12269,N_12220,N_12158);
nor U12270 (N_12270,N_12034,N_12027);
nand U12271 (N_12271,N_12222,N_12016);
nor U12272 (N_12272,N_12175,N_12237);
and U12273 (N_12273,N_12227,N_12028);
or U12274 (N_12274,N_12219,N_12033);
xor U12275 (N_12275,N_12014,N_12129);
or U12276 (N_12276,N_12096,N_12005);
or U12277 (N_12277,N_12190,N_12132);
nand U12278 (N_12278,N_12045,N_12166);
nand U12279 (N_12279,N_12161,N_12185);
nand U12280 (N_12280,N_12095,N_12164);
or U12281 (N_12281,N_12184,N_12073);
and U12282 (N_12282,N_12170,N_12000);
and U12283 (N_12283,N_12023,N_12013);
and U12284 (N_12284,N_12011,N_12044);
nor U12285 (N_12285,N_12115,N_12225);
and U12286 (N_12286,N_12187,N_12048);
xor U12287 (N_12287,N_12002,N_12063);
or U12288 (N_12288,N_12046,N_12188);
and U12289 (N_12289,N_12176,N_12186);
and U12290 (N_12290,N_12121,N_12165);
xnor U12291 (N_12291,N_12127,N_12089);
or U12292 (N_12292,N_12229,N_12077);
nor U12293 (N_12293,N_12111,N_12181);
xor U12294 (N_12294,N_12232,N_12196);
xor U12295 (N_12295,N_12056,N_12245);
and U12296 (N_12296,N_12144,N_12137);
nor U12297 (N_12297,N_12106,N_12234);
and U12298 (N_12298,N_12134,N_12167);
or U12299 (N_12299,N_12200,N_12060);
nor U12300 (N_12300,N_12131,N_12218);
nand U12301 (N_12301,N_12209,N_12213);
and U12302 (N_12302,N_12123,N_12157);
and U12303 (N_12303,N_12066,N_12084);
nand U12304 (N_12304,N_12151,N_12179);
or U12305 (N_12305,N_12019,N_12092);
and U12306 (N_12306,N_12133,N_12086);
and U12307 (N_12307,N_12104,N_12153);
xnor U12308 (N_12308,N_12199,N_12247);
nor U12309 (N_12309,N_12030,N_12021);
or U12310 (N_12310,N_12244,N_12093);
xor U12311 (N_12311,N_12177,N_12145);
nand U12312 (N_12312,N_12112,N_12159);
or U12313 (N_12313,N_12202,N_12238);
nor U12314 (N_12314,N_12139,N_12241);
and U12315 (N_12315,N_12242,N_12003);
xor U12316 (N_12316,N_12022,N_12041);
xnor U12317 (N_12317,N_12110,N_12088);
and U12318 (N_12318,N_12136,N_12080);
and U12319 (N_12319,N_12015,N_12240);
or U12320 (N_12320,N_12235,N_12085);
xnor U12321 (N_12321,N_12074,N_12043);
nand U12322 (N_12322,N_12008,N_12038);
nor U12323 (N_12323,N_12040,N_12172);
nand U12324 (N_12324,N_12082,N_12171);
and U12325 (N_12325,N_12168,N_12206);
nor U12326 (N_12326,N_12217,N_12017);
and U12327 (N_12327,N_12201,N_12102);
nor U12328 (N_12328,N_12210,N_12012);
nand U12329 (N_12329,N_12215,N_12231);
or U12330 (N_12330,N_12055,N_12122);
nor U12331 (N_12331,N_12049,N_12156);
xor U12332 (N_12332,N_12010,N_12105);
nand U12333 (N_12333,N_12050,N_12059);
nor U12334 (N_12334,N_12146,N_12091);
nor U12335 (N_12335,N_12004,N_12071);
or U12336 (N_12336,N_12081,N_12009);
and U12337 (N_12337,N_12149,N_12087);
nand U12338 (N_12338,N_12192,N_12113);
or U12339 (N_12339,N_12114,N_12090);
nor U12340 (N_12340,N_12221,N_12135);
or U12341 (N_12341,N_12173,N_12212);
and U12342 (N_12342,N_12026,N_12018);
xor U12343 (N_12343,N_12236,N_12076);
or U12344 (N_12344,N_12119,N_12183);
or U12345 (N_12345,N_12024,N_12160);
xor U12346 (N_12346,N_12182,N_12195);
xnor U12347 (N_12347,N_12138,N_12198);
or U12348 (N_12348,N_12052,N_12053);
and U12349 (N_12349,N_12007,N_12051);
nand U12350 (N_12350,N_12116,N_12162);
nand U12351 (N_12351,N_12025,N_12037);
nand U12352 (N_12352,N_12062,N_12031);
xor U12353 (N_12353,N_12109,N_12047);
xor U12354 (N_12354,N_12211,N_12101);
nor U12355 (N_12355,N_12126,N_12058);
nand U12356 (N_12356,N_12125,N_12174);
nor U12357 (N_12357,N_12142,N_12124);
xor U12358 (N_12358,N_12178,N_12230);
and U12359 (N_12359,N_12197,N_12006);
or U12360 (N_12360,N_12039,N_12248);
xor U12361 (N_12361,N_12064,N_12208);
nor U12362 (N_12362,N_12065,N_12246);
nand U12363 (N_12363,N_12068,N_12042);
or U12364 (N_12364,N_12117,N_12204);
nor U12365 (N_12365,N_12032,N_12001);
xnor U12366 (N_12366,N_12194,N_12108);
or U12367 (N_12367,N_12069,N_12152);
and U12368 (N_12368,N_12120,N_12205);
nor U12369 (N_12369,N_12057,N_12118);
nand U12370 (N_12370,N_12103,N_12128);
and U12371 (N_12371,N_12141,N_12193);
and U12372 (N_12372,N_12098,N_12228);
nand U12373 (N_12373,N_12224,N_12070);
xnor U12374 (N_12374,N_12075,N_12035);
xnor U12375 (N_12375,N_12050,N_12240);
or U12376 (N_12376,N_12078,N_12241);
nand U12377 (N_12377,N_12012,N_12185);
nand U12378 (N_12378,N_12207,N_12085);
and U12379 (N_12379,N_12171,N_12189);
nand U12380 (N_12380,N_12127,N_12010);
xnor U12381 (N_12381,N_12200,N_12045);
nor U12382 (N_12382,N_12121,N_12181);
nand U12383 (N_12383,N_12151,N_12118);
xor U12384 (N_12384,N_12239,N_12204);
and U12385 (N_12385,N_12035,N_12155);
and U12386 (N_12386,N_12159,N_12062);
nand U12387 (N_12387,N_12135,N_12174);
xor U12388 (N_12388,N_12238,N_12224);
nor U12389 (N_12389,N_12156,N_12214);
and U12390 (N_12390,N_12127,N_12237);
nor U12391 (N_12391,N_12038,N_12129);
nand U12392 (N_12392,N_12158,N_12194);
nor U12393 (N_12393,N_12228,N_12221);
and U12394 (N_12394,N_12185,N_12039);
xnor U12395 (N_12395,N_12072,N_12090);
nand U12396 (N_12396,N_12169,N_12000);
and U12397 (N_12397,N_12208,N_12081);
nor U12398 (N_12398,N_12066,N_12187);
nand U12399 (N_12399,N_12220,N_12060);
xor U12400 (N_12400,N_12033,N_12029);
and U12401 (N_12401,N_12142,N_12216);
nor U12402 (N_12402,N_12129,N_12135);
xnor U12403 (N_12403,N_12157,N_12073);
or U12404 (N_12404,N_12169,N_12153);
xnor U12405 (N_12405,N_12207,N_12044);
nor U12406 (N_12406,N_12041,N_12122);
xor U12407 (N_12407,N_12060,N_12181);
nand U12408 (N_12408,N_12102,N_12209);
xor U12409 (N_12409,N_12011,N_12172);
or U12410 (N_12410,N_12156,N_12230);
and U12411 (N_12411,N_12166,N_12066);
and U12412 (N_12412,N_12187,N_12107);
xor U12413 (N_12413,N_12161,N_12219);
or U12414 (N_12414,N_12065,N_12226);
xnor U12415 (N_12415,N_12073,N_12171);
nor U12416 (N_12416,N_12103,N_12245);
and U12417 (N_12417,N_12236,N_12248);
or U12418 (N_12418,N_12215,N_12021);
nor U12419 (N_12419,N_12010,N_12245);
xor U12420 (N_12420,N_12064,N_12146);
nand U12421 (N_12421,N_12103,N_12239);
or U12422 (N_12422,N_12191,N_12004);
xor U12423 (N_12423,N_12241,N_12178);
nand U12424 (N_12424,N_12243,N_12225);
and U12425 (N_12425,N_12096,N_12185);
nand U12426 (N_12426,N_12230,N_12207);
or U12427 (N_12427,N_12080,N_12027);
nand U12428 (N_12428,N_12158,N_12233);
xor U12429 (N_12429,N_12099,N_12229);
nor U12430 (N_12430,N_12089,N_12117);
nor U12431 (N_12431,N_12249,N_12180);
xor U12432 (N_12432,N_12056,N_12217);
and U12433 (N_12433,N_12014,N_12211);
nor U12434 (N_12434,N_12133,N_12016);
and U12435 (N_12435,N_12017,N_12057);
xor U12436 (N_12436,N_12140,N_12081);
or U12437 (N_12437,N_12096,N_12176);
nor U12438 (N_12438,N_12029,N_12181);
xor U12439 (N_12439,N_12151,N_12099);
and U12440 (N_12440,N_12015,N_12025);
and U12441 (N_12441,N_12210,N_12236);
or U12442 (N_12442,N_12220,N_12193);
xnor U12443 (N_12443,N_12061,N_12123);
nor U12444 (N_12444,N_12061,N_12172);
xor U12445 (N_12445,N_12151,N_12002);
nor U12446 (N_12446,N_12007,N_12238);
or U12447 (N_12447,N_12237,N_12219);
xor U12448 (N_12448,N_12237,N_12113);
nor U12449 (N_12449,N_12176,N_12010);
xor U12450 (N_12450,N_12159,N_12247);
and U12451 (N_12451,N_12009,N_12055);
and U12452 (N_12452,N_12175,N_12033);
and U12453 (N_12453,N_12013,N_12140);
xor U12454 (N_12454,N_12164,N_12241);
xnor U12455 (N_12455,N_12214,N_12033);
nand U12456 (N_12456,N_12120,N_12059);
or U12457 (N_12457,N_12051,N_12231);
and U12458 (N_12458,N_12090,N_12134);
or U12459 (N_12459,N_12045,N_12014);
or U12460 (N_12460,N_12157,N_12011);
and U12461 (N_12461,N_12113,N_12015);
nor U12462 (N_12462,N_12161,N_12181);
and U12463 (N_12463,N_12214,N_12197);
xor U12464 (N_12464,N_12082,N_12087);
nor U12465 (N_12465,N_12244,N_12217);
nor U12466 (N_12466,N_12081,N_12109);
nor U12467 (N_12467,N_12218,N_12240);
nor U12468 (N_12468,N_12024,N_12169);
nor U12469 (N_12469,N_12117,N_12007);
nand U12470 (N_12470,N_12118,N_12115);
or U12471 (N_12471,N_12016,N_12228);
and U12472 (N_12472,N_12093,N_12206);
or U12473 (N_12473,N_12061,N_12057);
nand U12474 (N_12474,N_12072,N_12214);
xnor U12475 (N_12475,N_12035,N_12247);
xnor U12476 (N_12476,N_12148,N_12041);
or U12477 (N_12477,N_12048,N_12209);
nand U12478 (N_12478,N_12045,N_12120);
nand U12479 (N_12479,N_12241,N_12091);
and U12480 (N_12480,N_12132,N_12236);
nand U12481 (N_12481,N_12136,N_12091);
nand U12482 (N_12482,N_12226,N_12101);
nand U12483 (N_12483,N_12225,N_12130);
nand U12484 (N_12484,N_12024,N_12144);
nand U12485 (N_12485,N_12064,N_12131);
nor U12486 (N_12486,N_12104,N_12111);
or U12487 (N_12487,N_12135,N_12186);
nor U12488 (N_12488,N_12244,N_12119);
or U12489 (N_12489,N_12147,N_12083);
and U12490 (N_12490,N_12171,N_12035);
or U12491 (N_12491,N_12135,N_12131);
xor U12492 (N_12492,N_12171,N_12132);
and U12493 (N_12493,N_12082,N_12190);
nor U12494 (N_12494,N_12029,N_12239);
xor U12495 (N_12495,N_12107,N_12129);
nand U12496 (N_12496,N_12226,N_12084);
nor U12497 (N_12497,N_12134,N_12115);
nand U12498 (N_12498,N_12166,N_12033);
or U12499 (N_12499,N_12185,N_12124);
or U12500 (N_12500,N_12437,N_12379);
and U12501 (N_12501,N_12301,N_12396);
and U12502 (N_12502,N_12473,N_12337);
xor U12503 (N_12503,N_12429,N_12277);
and U12504 (N_12504,N_12276,N_12343);
nor U12505 (N_12505,N_12490,N_12481);
nand U12506 (N_12506,N_12392,N_12338);
and U12507 (N_12507,N_12326,N_12323);
nand U12508 (N_12508,N_12330,N_12311);
xnor U12509 (N_12509,N_12256,N_12305);
xor U12510 (N_12510,N_12350,N_12293);
nor U12511 (N_12511,N_12272,N_12358);
nor U12512 (N_12512,N_12278,N_12303);
and U12513 (N_12513,N_12496,N_12406);
or U12514 (N_12514,N_12365,N_12464);
nor U12515 (N_12515,N_12281,N_12373);
xnor U12516 (N_12516,N_12271,N_12442);
nor U12517 (N_12517,N_12485,N_12498);
nand U12518 (N_12518,N_12279,N_12466);
and U12519 (N_12519,N_12483,N_12454);
xnor U12520 (N_12520,N_12257,N_12424);
or U12521 (N_12521,N_12408,N_12459);
or U12522 (N_12522,N_12479,N_12477);
nand U12523 (N_12523,N_12369,N_12364);
xor U12524 (N_12524,N_12439,N_12474);
nor U12525 (N_12525,N_12268,N_12431);
and U12526 (N_12526,N_12266,N_12344);
nand U12527 (N_12527,N_12436,N_12486);
and U12528 (N_12528,N_12348,N_12352);
or U12529 (N_12529,N_12269,N_12388);
and U12530 (N_12530,N_12491,N_12289);
nand U12531 (N_12531,N_12488,N_12314);
nor U12532 (N_12532,N_12447,N_12254);
xnor U12533 (N_12533,N_12414,N_12399);
nor U12534 (N_12534,N_12467,N_12310);
nand U12535 (N_12535,N_12342,N_12291);
nand U12536 (N_12536,N_12374,N_12446);
xor U12537 (N_12537,N_12492,N_12312);
nor U12538 (N_12538,N_12449,N_12445);
and U12539 (N_12539,N_12426,N_12443);
nor U12540 (N_12540,N_12444,N_12400);
and U12541 (N_12541,N_12407,N_12340);
or U12542 (N_12542,N_12397,N_12335);
xor U12543 (N_12543,N_12355,N_12494);
nand U12544 (N_12544,N_12353,N_12255);
and U12545 (N_12545,N_12319,N_12371);
or U12546 (N_12546,N_12423,N_12292);
and U12547 (N_12547,N_12280,N_12497);
nand U12548 (N_12548,N_12458,N_12331);
or U12549 (N_12549,N_12290,N_12383);
or U12550 (N_12550,N_12283,N_12375);
nor U12551 (N_12551,N_12395,N_12327);
nor U12552 (N_12552,N_12463,N_12306);
nand U12553 (N_12553,N_12489,N_12302);
nand U12554 (N_12554,N_12333,N_12356);
or U12555 (N_12555,N_12387,N_12366);
nor U12556 (N_12556,N_12434,N_12336);
xor U12557 (N_12557,N_12461,N_12378);
or U12558 (N_12558,N_12260,N_12370);
and U12559 (N_12559,N_12413,N_12456);
nand U12560 (N_12560,N_12318,N_12297);
and U12561 (N_12561,N_12328,N_12422);
or U12562 (N_12562,N_12253,N_12274);
xnor U12563 (N_12563,N_12390,N_12261);
nand U12564 (N_12564,N_12465,N_12299);
or U12565 (N_12565,N_12264,N_12391);
or U12566 (N_12566,N_12307,N_12440);
nand U12567 (N_12567,N_12360,N_12401);
nand U12568 (N_12568,N_12361,N_12354);
xnor U12569 (N_12569,N_12287,N_12441);
nor U12570 (N_12570,N_12487,N_12359);
or U12571 (N_12571,N_12478,N_12480);
or U12572 (N_12572,N_12377,N_12329);
and U12573 (N_12573,N_12402,N_12252);
xor U12574 (N_12574,N_12304,N_12349);
and U12575 (N_12575,N_12398,N_12393);
or U12576 (N_12576,N_12448,N_12285);
or U12577 (N_12577,N_12316,N_12453);
or U12578 (N_12578,N_12286,N_12273);
and U12579 (N_12579,N_12457,N_12282);
or U12580 (N_12580,N_12409,N_12372);
xor U12581 (N_12581,N_12420,N_12263);
nor U12582 (N_12582,N_12321,N_12339);
and U12583 (N_12583,N_12403,N_12345);
nor U12584 (N_12584,N_12418,N_12362);
nand U12585 (N_12585,N_12433,N_12315);
and U12586 (N_12586,N_12427,N_12499);
nand U12587 (N_12587,N_12484,N_12300);
xor U12588 (N_12588,N_12432,N_12450);
nand U12589 (N_12589,N_12452,N_12482);
nand U12590 (N_12590,N_12324,N_12419);
and U12591 (N_12591,N_12363,N_12317);
nor U12592 (N_12592,N_12346,N_12411);
nand U12593 (N_12593,N_12389,N_12386);
xnor U12594 (N_12594,N_12295,N_12294);
nand U12595 (N_12595,N_12267,N_12430);
nor U12596 (N_12596,N_12435,N_12460);
xor U12597 (N_12597,N_12468,N_12475);
xor U12598 (N_12598,N_12258,N_12308);
and U12599 (N_12599,N_12428,N_12270);
or U12600 (N_12600,N_12404,N_12296);
and U12601 (N_12601,N_12438,N_12415);
xor U12602 (N_12602,N_12410,N_12288);
or U12603 (N_12603,N_12421,N_12376);
and U12604 (N_12604,N_12313,N_12262);
nor U12605 (N_12605,N_12381,N_12309);
nor U12606 (N_12606,N_12298,N_12469);
nor U12607 (N_12607,N_12259,N_12334);
or U12608 (N_12608,N_12380,N_12250);
nand U12609 (N_12609,N_12275,N_12251);
nor U12610 (N_12610,N_12382,N_12367);
nor U12611 (N_12611,N_12284,N_12385);
nor U12612 (N_12612,N_12416,N_12320);
and U12613 (N_12613,N_12394,N_12417);
nor U12614 (N_12614,N_12471,N_12405);
nor U12615 (N_12615,N_12322,N_12357);
nand U12616 (N_12616,N_12451,N_12265);
xor U12617 (N_12617,N_12325,N_12347);
or U12618 (N_12618,N_12495,N_12425);
nand U12619 (N_12619,N_12368,N_12351);
or U12620 (N_12620,N_12412,N_12384);
or U12621 (N_12621,N_12462,N_12455);
and U12622 (N_12622,N_12470,N_12472);
or U12623 (N_12623,N_12332,N_12493);
and U12624 (N_12624,N_12476,N_12341);
nand U12625 (N_12625,N_12258,N_12352);
or U12626 (N_12626,N_12412,N_12371);
xnor U12627 (N_12627,N_12350,N_12331);
nor U12628 (N_12628,N_12252,N_12466);
nor U12629 (N_12629,N_12261,N_12252);
nand U12630 (N_12630,N_12380,N_12347);
nor U12631 (N_12631,N_12337,N_12467);
xnor U12632 (N_12632,N_12482,N_12460);
or U12633 (N_12633,N_12264,N_12427);
and U12634 (N_12634,N_12312,N_12340);
nor U12635 (N_12635,N_12265,N_12477);
or U12636 (N_12636,N_12475,N_12268);
xnor U12637 (N_12637,N_12263,N_12481);
and U12638 (N_12638,N_12425,N_12263);
xor U12639 (N_12639,N_12469,N_12495);
nand U12640 (N_12640,N_12492,N_12472);
nand U12641 (N_12641,N_12438,N_12363);
or U12642 (N_12642,N_12438,N_12258);
and U12643 (N_12643,N_12453,N_12416);
and U12644 (N_12644,N_12361,N_12401);
nand U12645 (N_12645,N_12417,N_12459);
nor U12646 (N_12646,N_12476,N_12463);
and U12647 (N_12647,N_12287,N_12314);
nor U12648 (N_12648,N_12284,N_12260);
xnor U12649 (N_12649,N_12350,N_12482);
xnor U12650 (N_12650,N_12466,N_12344);
and U12651 (N_12651,N_12390,N_12288);
nor U12652 (N_12652,N_12436,N_12481);
nand U12653 (N_12653,N_12406,N_12296);
nor U12654 (N_12654,N_12329,N_12420);
or U12655 (N_12655,N_12364,N_12256);
nand U12656 (N_12656,N_12363,N_12268);
nor U12657 (N_12657,N_12257,N_12468);
nor U12658 (N_12658,N_12499,N_12368);
or U12659 (N_12659,N_12314,N_12281);
nor U12660 (N_12660,N_12434,N_12309);
and U12661 (N_12661,N_12289,N_12427);
nor U12662 (N_12662,N_12490,N_12370);
nand U12663 (N_12663,N_12358,N_12382);
nand U12664 (N_12664,N_12399,N_12260);
xnor U12665 (N_12665,N_12372,N_12341);
xnor U12666 (N_12666,N_12335,N_12401);
nor U12667 (N_12667,N_12353,N_12351);
xnor U12668 (N_12668,N_12436,N_12313);
nand U12669 (N_12669,N_12347,N_12312);
and U12670 (N_12670,N_12486,N_12281);
xor U12671 (N_12671,N_12277,N_12428);
nor U12672 (N_12672,N_12472,N_12428);
or U12673 (N_12673,N_12427,N_12376);
xnor U12674 (N_12674,N_12410,N_12427);
nand U12675 (N_12675,N_12473,N_12378);
or U12676 (N_12676,N_12269,N_12349);
or U12677 (N_12677,N_12401,N_12439);
or U12678 (N_12678,N_12468,N_12294);
nor U12679 (N_12679,N_12480,N_12342);
or U12680 (N_12680,N_12326,N_12389);
nor U12681 (N_12681,N_12283,N_12424);
nand U12682 (N_12682,N_12301,N_12318);
and U12683 (N_12683,N_12298,N_12309);
or U12684 (N_12684,N_12336,N_12264);
xnor U12685 (N_12685,N_12350,N_12282);
and U12686 (N_12686,N_12420,N_12337);
xor U12687 (N_12687,N_12303,N_12490);
or U12688 (N_12688,N_12380,N_12449);
or U12689 (N_12689,N_12441,N_12428);
nand U12690 (N_12690,N_12365,N_12411);
and U12691 (N_12691,N_12487,N_12464);
and U12692 (N_12692,N_12449,N_12453);
and U12693 (N_12693,N_12262,N_12450);
and U12694 (N_12694,N_12337,N_12391);
or U12695 (N_12695,N_12284,N_12352);
or U12696 (N_12696,N_12297,N_12272);
nand U12697 (N_12697,N_12432,N_12375);
xnor U12698 (N_12698,N_12482,N_12342);
nor U12699 (N_12699,N_12345,N_12357);
xor U12700 (N_12700,N_12478,N_12379);
or U12701 (N_12701,N_12250,N_12256);
nor U12702 (N_12702,N_12467,N_12456);
xnor U12703 (N_12703,N_12298,N_12352);
or U12704 (N_12704,N_12256,N_12347);
nor U12705 (N_12705,N_12473,N_12437);
nor U12706 (N_12706,N_12467,N_12322);
and U12707 (N_12707,N_12350,N_12312);
or U12708 (N_12708,N_12307,N_12487);
xnor U12709 (N_12709,N_12357,N_12400);
or U12710 (N_12710,N_12291,N_12323);
or U12711 (N_12711,N_12325,N_12339);
or U12712 (N_12712,N_12305,N_12311);
and U12713 (N_12713,N_12456,N_12411);
nand U12714 (N_12714,N_12472,N_12269);
or U12715 (N_12715,N_12484,N_12390);
xor U12716 (N_12716,N_12412,N_12264);
or U12717 (N_12717,N_12499,N_12332);
or U12718 (N_12718,N_12347,N_12342);
nand U12719 (N_12719,N_12360,N_12477);
and U12720 (N_12720,N_12369,N_12323);
nand U12721 (N_12721,N_12302,N_12383);
xnor U12722 (N_12722,N_12395,N_12447);
nor U12723 (N_12723,N_12320,N_12325);
nor U12724 (N_12724,N_12492,N_12283);
nor U12725 (N_12725,N_12496,N_12480);
and U12726 (N_12726,N_12395,N_12410);
and U12727 (N_12727,N_12292,N_12417);
and U12728 (N_12728,N_12332,N_12411);
xor U12729 (N_12729,N_12342,N_12382);
and U12730 (N_12730,N_12456,N_12352);
nand U12731 (N_12731,N_12310,N_12343);
nand U12732 (N_12732,N_12281,N_12491);
and U12733 (N_12733,N_12436,N_12318);
and U12734 (N_12734,N_12403,N_12250);
nand U12735 (N_12735,N_12288,N_12326);
nor U12736 (N_12736,N_12261,N_12431);
or U12737 (N_12737,N_12423,N_12419);
or U12738 (N_12738,N_12464,N_12449);
nor U12739 (N_12739,N_12412,N_12349);
xnor U12740 (N_12740,N_12381,N_12365);
and U12741 (N_12741,N_12367,N_12375);
or U12742 (N_12742,N_12291,N_12488);
nor U12743 (N_12743,N_12267,N_12297);
xnor U12744 (N_12744,N_12478,N_12407);
xnor U12745 (N_12745,N_12457,N_12438);
and U12746 (N_12746,N_12336,N_12417);
or U12747 (N_12747,N_12251,N_12450);
nor U12748 (N_12748,N_12466,N_12403);
nor U12749 (N_12749,N_12356,N_12408);
nand U12750 (N_12750,N_12734,N_12640);
xnor U12751 (N_12751,N_12604,N_12606);
nor U12752 (N_12752,N_12551,N_12601);
xor U12753 (N_12753,N_12558,N_12570);
and U12754 (N_12754,N_12523,N_12556);
xnor U12755 (N_12755,N_12643,N_12649);
or U12756 (N_12756,N_12704,N_12507);
and U12757 (N_12757,N_12662,N_12618);
nand U12758 (N_12758,N_12502,N_12557);
xor U12759 (N_12759,N_12532,N_12612);
and U12760 (N_12760,N_12732,N_12508);
nand U12761 (N_12761,N_12693,N_12729);
xor U12762 (N_12762,N_12644,N_12635);
nor U12763 (N_12763,N_12561,N_12653);
xor U12764 (N_12764,N_12578,N_12654);
xor U12765 (N_12765,N_12665,N_12672);
or U12766 (N_12766,N_12617,N_12607);
and U12767 (N_12767,N_12615,N_12509);
and U12768 (N_12768,N_12541,N_12554);
nor U12769 (N_12769,N_12681,N_12567);
and U12770 (N_12770,N_12642,N_12591);
and U12771 (N_12771,N_12608,N_12659);
or U12772 (N_12772,N_12718,N_12547);
xnor U12773 (N_12773,N_12631,N_12705);
xor U12774 (N_12774,N_12727,N_12589);
or U12775 (N_12775,N_12650,N_12548);
xnor U12776 (N_12776,N_12527,N_12731);
and U12777 (N_12777,N_12703,N_12549);
or U12778 (N_12778,N_12535,N_12524);
and U12779 (N_12779,N_12670,N_12588);
and U12780 (N_12780,N_12748,N_12710);
nor U12781 (N_12781,N_12577,N_12657);
xnor U12782 (N_12782,N_12689,N_12699);
or U12783 (N_12783,N_12593,N_12683);
nand U12784 (N_12784,N_12611,N_12628);
nand U12785 (N_12785,N_12540,N_12652);
nand U12786 (N_12786,N_12730,N_12582);
nand U12787 (N_12787,N_12583,N_12664);
and U12788 (N_12788,N_12696,N_12625);
and U12789 (N_12789,N_12723,N_12528);
nor U12790 (N_12790,N_12647,N_12544);
and U12791 (N_12791,N_12676,N_12537);
and U12792 (N_12792,N_12504,N_12715);
xor U12793 (N_12793,N_12517,N_12533);
nand U12794 (N_12794,N_12634,N_12741);
and U12795 (N_12795,N_12576,N_12663);
and U12796 (N_12796,N_12609,N_12566);
and U12797 (N_12797,N_12656,N_12673);
xor U12798 (N_12798,N_12678,N_12559);
xnor U12799 (N_12799,N_12706,N_12728);
nor U12800 (N_12800,N_12671,N_12580);
nand U12801 (N_12801,N_12695,N_12501);
nor U12802 (N_12802,N_12605,N_12568);
nand U12803 (N_12803,N_12655,N_12714);
nor U12804 (N_12804,N_12538,N_12667);
xor U12805 (N_12805,N_12546,N_12637);
and U12806 (N_12806,N_12692,N_12739);
or U12807 (N_12807,N_12686,N_12726);
or U12808 (N_12808,N_12563,N_12742);
nand U12809 (N_12809,N_12531,N_12529);
or U12810 (N_12810,N_12565,N_12702);
or U12811 (N_12811,N_12749,N_12674);
nor U12812 (N_12812,N_12719,N_12629);
xor U12813 (N_12813,N_12587,N_12519);
and U12814 (N_12814,N_12555,N_12594);
nand U12815 (N_12815,N_12627,N_12581);
nor U12816 (N_12816,N_12573,N_12722);
or U12817 (N_12817,N_12575,N_12511);
xor U12818 (N_12818,N_12720,N_12623);
and U12819 (N_12819,N_12688,N_12717);
nor U12820 (N_12820,N_12632,N_12633);
and U12821 (N_12821,N_12733,N_12569);
nand U12822 (N_12822,N_12709,N_12736);
nor U12823 (N_12823,N_12610,N_12698);
nand U12824 (N_12824,N_12694,N_12744);
nor U12825 (N_12825,N_12505,N_12539);
and U12826 (N_12826,N_12630,N_12701);
and U12827 (N_12827,N_12530,N_12595);
or U12828 (N_12828,N_12562,N_12592);
and U12829 (N_12829,N_12708,N_12735);
nand U12830 (N_12830,N_12666,N_12572);
xnor U12831 (N_12831,N_12645,N_12746);
and U12832 (N_12832,N_12603,N_12545);
and U12833 (N_12833,N_12685,N_12682);
nor U12834 (N_12834,N_12620,N_12747);
xor U12835 (N_12835,N_12571,N_12516);
or U12836 (N_12836,N_12542,N_12515);
or U12837 (N_12837,N_12668,N_12700);
or U12838 (N_12838,N_12721,N_12660);
nor U12839 (N_12839,N_12713,N_12584);
or U12840 (N_12840,N_12743,N_12574);
nand U12841 (N_12841,N_12712,N_12737);
nor U12842 (N_12842,N_12590,N_12684);
and U12843 (N_12843,N_12651,N_12602);
nor U12844 (N_12844,N_12513,N_12613);
or U12845 (N_12845,N_12680,N_12520);
nand U12846 (N_12846,N_12724,N_12596);
and U12847 (N_12847,N_12687,N_12536);
nand U12848 (N_12848,N_12707,N_12658);
or U12849 (N_12849,N_12740,N_12669);
nor U12850 (N_12850,N_12534,N_12697);
or U12851 (N_12851,N_12661,N_12512);
nor U12852 (N_12852,N_12677,N_12639);
and U12853 (N_12853,N_12543,N_12597);
and U12854 (N_12854,N_12518,N_12598);
xor U12855 (N_12855,N_12646,N_12599);
and U12856 (N_12856,N_12552,N_12622);
and U12857 (N_12857,N_12619,N_12525);
nor U12858 (N_12858,N_12564,N_12526);
nor U12859 (N_12859,N_12585,N_12616);
nand U12860 (N_12860,N_12621,N_12648);
nand U12861 (N_12861,N_12503,N_12738);
xnor U12862 (N_12862,N_12553,N_12716);
xor U12863 (N_12863,N_12600,N_12711);
and U12864 (N_12864,N_12638,N_12550);
or U12865 (N_12865,N_12636,N_12675);
nand U12866 (N_12866,N_12500,N_12614);
or U12867 (N_12867,N_12521,N_12691);
xnor U12868 (N_12868,N_12626,N_12679);
or U12869 (N_12869,N_12624,N_12579);
and U12870 (N_12870,N_12745,N_12690);
xor U12871 (N_12871,N_12725,N_12522);
xor U12872 (N_12872,N_12514,N_12560);
or U12873 (N_12873,N_12586,N_12510);
nand U12874 (N_12874,N_12506,N_12641);
xor U12875 (N_12875,N_12565,N_12597);
xnor U12876 (N_12876,N_12523,N_12578);
or U12877 (N_12877,N_12661,N_12526);
xor U12878 (N_12878,N_12612,N_12677);
nand U12879 (N_12879,N_12615,N_12667);
or U12880 (N_12880,N_12649,N_12725);
xor U12881 (N_12881,N_12554,N_12668);
or U12882 (N_12882,N_12643,N_12670);
nor U12883 (N_12883,N_12615,N_12624);
or U12884 (N_12884,N_12670,N_12606);
nand U12885 (N_12885,N_12552,N_12535);
nor U12886 (N_12886,N_12684,N_12708);
xnor U12887 (N_12887,N_12508,N_12501);
nand U12888 (N_12888,N_12712,N_12735);
and U12889 (N_12889,N_12615,N_12541);
and U12890 (N_12890,N_12533,N_12540);
nor U12891 (N_12891,N_12730,N_12743);
nor U12892 (N_12892,N_12681,N_12673);
or U12893 (N_12893,N_12646,N_12554);
nand U12894 (N_12894,N_12737,N_12635);
or U12895 (N_12895,N_12606,N_12531);
nand U12896 (N_12896,N_12594,N_12529);
or U12897 (N_12897,N_12651,N_12747);
nand U12898 (N_12898,N_12692,N_12597);
or U12899 (N_12899,N_12508,N_12676);
or U12900 (N_12900,N_12623,N_12531);
and U12901 (N_12901,N_12623,N_12713);
xnor U12902 (N_12902,N_12565,N_12669);
xnor U12903 (N_12903,N_12568,N_12632);
xor U12904 (N_12904,N_12587,N_12730);
nor U12905 (N_12905,N_12513,N_12610);
nor U12906 (N_12906,N_12610,N_12743);
nand U12907 (N_12907,N_12694,N_12548);
xnor U12908 (N_12908,N_12720,N_12746);
xnor U12909 (N_12909,N_12536,N_12501);
nand U12910 (N_12910,N_12522,N_12524);
and U12911 (N_12911,N_12586,N_12515);
xor U12912 (N_12912,N_12580,N_12565);
or U12913 (N_12913,N_12603,N_12675);
xnor U12914 (N_12914,N_12594,N_12558);
nand U12915 (N_12915,N_12552,N_12675);
nor U12916 (N_12916,N_12728,N_12541);
or U12917 (N_12917,N_12716,N_12524);
or U12918 (N_12918,N_12627,N_12662);
and U12919 (N_12919,N_12578,N_12690);
xor U12920 (N_12920,N_12725,N_12572);
xnor U12921 (N_12921,N_12686,N_12594);
nand U12922 (N_12922,N_12507,N_12601);
and U12923 (N_12923,N_12716,N_12640);
nor U12924 (N_12924,N_12726,N_12662);
and U12925 (N_12925,N_12517,N_12644);
and U12926 (N_12926,N_12547,N_12676);
xor U12927 (N_12927,N_12647,N_12567);
nand U12928 (N_12928,N_12511,N_12672);
nor U12929 (N_12929,N_12624,N_12645);
and U12930 (N_12930,N_12632,N_12585);
nand U12931 (N_12931,N_12605,N_12649);
and U12932 (N_12932,N_12528,N_12673);
or U12933 (N_12933,N_12746,N_12636);
xor U12934 (N_12934,N_12737,N_12604);
nand U12935 (N_12935,N_12522,N_12701);
or U12936 (N_12936,N_12697,N_12609);
and U12937 (N_12937,N_12729,N_12603);
and U12938 (N_12938,N_12557,N_12740);
nand U12939 (N_12939,N_12604,N_12725);
xnor U12940 (N_12940,N_12636,N_12582);
nor U12941 (N_12941,N_12709,N_12708);
nand U12942 (N_12942,N_12722,N_12685);
nand U12943 (N_12943,N_12708,N_12505);
nand U12944 (N_12944,N_12748,N_12729);
and U12945 (N_12945,N_12728,N_12536);
nor U12946 (N_12946,N_12660,N_12506);
or U12947 (N_12947,N_12618,N_12571);
and U12948 (N_12948,N_12556,N_12696);
or U12949 (N_12949,N_12610,N_12642);
nor U12950 (N_12950,N_12569,N_12711);
or U12951 (N_12951,N_12747,N_12672);
or U12952 (N_12952,N_12610,N_12572);
and U12953 (N_12953,N_12684,N_12553);
or U12954 (N_12954,N_12660,N_12556);
nor U12955 (N_12955,N_12706,N_12636);
xnor U12956 (N_12956,N_12517,N_12503);
nand U12957 (N_12957,N_12620,N_12502);
nor U12958 (N_12958,N_12666,N_12566);
nand U12959 (N_12959,N_12576,N_12574);
xnor U12960 (N_12960,N_12671,N_12672);
nor U12961 (N_12961,N_12645,N_12732);
nor U12962 (N_12962,N_12618,N_12749);
nand U12963 (N_12963,N_12621,N_12669);
and U12964 (N_12964,N_12623,N_12663);
xnor U12965 (N_12965,N_12632,N_12695);
and U12966 (N_12966,N_12670,N_12656);
and U12967 (N_12967,N_12717,N_12627);
and U12968 (N_12968,N_12550,N_12610);
nand U12969 (N_12969,N_12623,N_12708);
xor U12970 (N_12970,N_12643,N_12690);
or U12971 (N_12971,N_12589,N_12683);
nand U12972 (N_12972,N_12648,N_12723);
xnor U12973 (N_12973,N_12529,N_12694);
and U12974 (N_12974,N_12643,N_12503);
or U12975 (N_12975,N_12571,N_12581);
and U12976 (N_12976,N_12619,N_12669);
xor U12977 (N_12977,N_12732,N_12595);
and U12978 (N_12978,N_12539,N_12518);
nand U12979 (N_12979,N_12683,N_12746);
and U12980 (N_12980,N_12574,N_12626);
and U12981 (N_12981,N_12736,N_12584);
nor U12982 (N_12982,N_12694,N_12514);
and U12983 (N_12983,N_12604,N_12712);
xor U12984 (N_12984,N_12527,N_12708);
xor U12985 (N_12985,N_12551,N_12654);
nand U12986 (N_12986,N_12673,N_12603);
nor U12987 (N_12987,N_12683,N_12741);
and U12988 (N_12988,N_12688,N_12576);
nand U12989 (N_12989,N_12703,N_12733);
nand U12990 (N_12990,N_12589,N_12588);
nor U12991 (N_12991,N_12743,N_12644);
xor U12992 (N_12992,N_12663,N_12574);
xor U12993 (N_12993,N_12575,N_12539);
nor U12994 (N_12994,N_12565,N_12734);
and U12995 (N_12995,N_12629,N_12607);
or U12996 (N_12996,N_12584,N_12699);
nor U12997 (N_12997,N_12618,N_12730);
xnor U12998 (N_12998,N_12734,N_12511);
nor U12999 (N_12999,N_12608,N_12548);
nand U13000 (N_13000,N_12927,N_12991);
and U13001 (N_13001,N_12797,N_12849);
and U13002 (N_13002,N_12989,N_12924);
nand U13003 (N_13003,N_12948,N_12951);
or U13004 (N_13004,N_12888,N_12813);
nor U13005 (N_13005,N_12860,N_12981);
nand U13006 (N_13006,N_12852,N_12878);
xor U13007 (N_13007,N_12850,N_12937);
nand U13008 (N_13008,N_12844,N_12897);
nand U13009 (N_13009,N_12895,N_12758);
and U13010 (N_13010,N_12803,N_12912);
nand U13011 (N_13011,N_12785,N_12953);
xnor U13012 (N_13012,N_12770,N_12931);
or U13013 (N_13013,N_12908,N_12801);
xnor U13014 (N_13014,N_12827,N_12862);
and U13015 (N_13015,N_12756,N_12898);
nand U13016 (N_13016,N_12859,N_12822);
or U13017 (N_13017,N_12865,N_12752);
nand U13018 (N_13018,N_12846,N_12755);
or U13019 (N_13019,N_12762,N_12904);
nor U13020 (N_13020,N_12892,N_12766);
or U13021 (N_13021,N_12759,N_12979);
nor U13022 (N_13022,N_12962,N_12789);
and U13023 (N_13023,N_12876,N_12944);
and U13024 (N_13024,N_12969,N_12974);
nor U13025 (N_13025,N_12972,N_12788);
nor U13026 (N_13026,N_12796,N_12947);
or U13027 (N_13027,N_12916,N_12853);
nand U13028 (N_13028,N_12925,N_12955);
nor U13029 (N_13029,N_12999,N_12793);
and U13030 (N_13030,N_12926,N_12854);
and U13031 (N_13031,N_12775,N_12967);
nor U13032 (N_13032,N_12869,N_12896);
nor U13033 (N_13033,N_12891,N_12763);
nor U13034 (N_13034,N_12750,N_12984);
and U13035 (N_13035,N_12863,N_12890);
and U13036 (N_13036,N_12913,N_12781);
or U13037 (N_13037,N_12851,N_12780);
nand U13038 (N_13038,N_12817,N_12990);
or U13039 (N_13039,N_12855,N_12975);
nor U13040 (N_13040,N_12905,N_12870);
or U13041 (N_13041,N_12884,N_12773);
and U13042 (N_13042,N_12882,N_12834);
or U13043 (N_13043,N_12996,N_12887);
nor U13044 (N_13044,N_12977,N_12800);
nor U13045 (N_13045,N_12814,N_12815);
nor U13046 (N_13046,N_12848,N_12779);
or U13047 (N_13047,N_12958,N_12932);
xor U13048 (N_13048,N_12816,N_12899);
nor U13049 (N_13049,N_12982,N_12832);
nand U13050 (N_13050,N_12938,N_12807);
nand U13051 (N_13051,N_12945,N_12966);
xnor U13052 (N_13052,N_12943,N_12811);
nor U13053 (N_13053,N_12941,N_12872);
xnor U13054 (N_13054,N_12942,N_12946);
xnor U13055 (N_13055,N_12930,N_12983);
nor U13056 (N_13056,N_12771,N_12760);
nor U13057 (N_13057,N_12968,N_12956);
xnor U13058 (N_13058,N_12765,N_12768);
nor U13059 (N_13059,N_12821,N_12820);
and U13060 (N_13060,N_12954,N_12864);
and U13061 (N_13061,N_12911,N_12809);
xnor U13062 (N_13062,N_12929,N_12963);
or U13063 (N_13063,N_12802,N_12935);
nand U13064 (N_13064,N_12920,N_12901);
nand U13065 (N_13065,N_12808,N_12825);
and U13066 (N_13066,N_12933,N_12842);
and U13067 (N_13067,N_12810,N_12812);
xnor U13068 (N_13068,N_12783,N_12754);
and U13069 (N_13069,N_12995,N_12894);
nand U13070 (N_13070,N_12907,N_12799);
and U13071 (N_13071,N_12767,N_12866);
and U13072 (N_13072,N_12909,N_12880);
or U13073 (N_13073,N_12960,N_12764);
and U13074 (N_13074,N_12790,N_12871);
xor U13075 (N_13075,N_12965,N_12776);
xnor U13076 (N_13076,N_12804,N_12798);
or U13077 (N_13077,N_12993,N_12787);
nand U13078 (N_13078,N_12923,N_12873);
nor U13079 (N_13079,N_12961,N_12980);
and U13080 (N_13080,N_12847,N_12828);
nor U13081 (N_13081,N_12839,N_12903);
xnor U13082 (N_13082,N_12857,N_12753);
nor U13083 (N_13083,N_12777,N_12868);
or U13084 (N_13084,N_12893,N_12886);
or U13085 (N_13085,N_12879,N_12792);
nand U13086 (N_13086,N_12818,N_12794);
nand U13087 (N_13087,N_12885,N_12835);
xnor U13088 (N_13088,N_12978,N_12906);
nand U13089 (N_13089,N_12881,N_12914);
nor U13090 (N_13090,N_12970,N_12795);
or U13091 (N_13091,N_12964,N_12772);
or U13092 (N_13092,N_12921,N_12874);
xor U13093 (N_13093,N_12998,N_12806);
and U13094 (N_13094,N_12856,N_12900);
and U13095 (N_13095,N_12936,N_12845);
nand U13096 (N_13096,N_12952,N_12957);
xor U13097 (N_13097,N_12824,N_12784);
and U13098 (N_13098,N_12786,N_12830);
and U13099 (N_13099,N_12985,N_12823);
and U13100 (N_13100,N_12997,N_12987);
and U13101 (N_13101,N_12902,N_12992);
xnor U13102 (N_13102,N_12939,N_12994);
nor U13103 (N_13103,N_12858,N_12889);
nor U13104 (N_13104,N_12843,N_12829);
nand U13105 (N_13105,N_12837,N_12986);
xor U13106 (N_13106,N_12922,N_12976);
nor U13107 (N_13107,N_12836,N_12819);
xor U13108 (N_13108,N_12833,N_12831);
and U13109 (N_13109,N_12910,N_12861);
nand U13110 (N_13110,N_12917,N_12883);
xor U13111 (N_13111,N_12751,N_12950);
xnor U13112 (N_13112,N_12769,N_12774);
xor U13113 (N_13113,N_12867,N_12919);
and U13114 (N_13114,N_12791,N_12971);
nor U13115 (N_13115,N_12877,N_12973);
xor U13116 (N_13116,N_12949,N_12940);
or U13117 (N_13117,N_12934,N_12826);
nand U13118 (N_13118,N_12838,N_12875);
and U13119 (N_13119,N_12918,N_12915);
and U13120 (N_13120,N_12840,N_12959);
xnor U13121 (N_13121,N_12988,N_12805);
and U13122 (N_13122,N_12782,N_12757);
xnor U13123 (N_13123,N_12928,N_12778);
nand U13124 (N_13124,N_12841,N_12761);
nand U13125 (N_13125,N_12997,N_12906);
or U13126 (N_13126,N_12978,N_12907);
nor U13127 (N_13127,N_12750,N_12936);
or U13128 (N_13128,N_12859,N_12838);
xnor U13129 (N_13129,N_12806,N_12775);
nand U13130 (N_13130,N_12961,N_12933);
xor U13131 (N_13131,N_12930,N_12864);
and U13132 (N_13132,N_12990,N_12985);
nor U13133 (N_13133,N_12809,N_12826);
nor U13134 (N_13134,N_12811,N_12952);
and U13135 (N_13135,N_12818,N_12845);
xnor U13136 (N_13136,N_12782,N_12883);
or U13137 (N_13137,N_12821,N_12798);
xnor U13138 (N_13138,N_12975,N_12836);
nor U13139 (N_13139,N_12883,N_12876);
and U13140 (N_13140,N_12833,N_12923);
xnor U13141 (N_13141,N_12940,N_12799);
xnor U13142 (N_13142,N_12804,N_12777);
or U13143 (N_13143,N_12798,N_12832);
nor U13144 (N_13144,N_12852,N_12909);
nor U13145 (N_13145,N_12890,N_12956);
and U13146 (N_13146,N_12776,N_12876);
or U13147 (N_13147,N_12895,N_12909);
nand U13148 (N_13148,N_12942,N_12898);
nand U13149 (N_13149,N_12973,N_12959);
xor U13150 (N_13150,N_12780,N_12823);
nor U13151 (N_13151,N_12969,N_12929);
and U13152 (N_13152,N_12898,N_12964);
nand U13153 (N_13153,N_12811,N_12910);
or U13154 (N_13154,N_12873,N_12840);
nand U13155 (N_13155,N_12888,N_12938);
nand U13156 (N_13156,N_12854,N_12776);
nor U13157 (N_13157,N_12818,N_12831);
and U13158 (N_13158,N_12995,N_12974);
xor U13159 (N_13159,N_12757,N_12918);
or U13160 (N_13160,N_12859,N_12971);
xor U13161 (N_13161,N_12857,N_12927);
xor U13162 (N_13162,N_12875,N_12824);
or U13163 (N_13163,N_12974,N_12766);
nor U13164 (N_13164,N_12970,N_12856);
nor U13165 (N_13165,N_12999,N_12830);
and U13166 (N_13166,N_12956,N_12844);
or U13167 (N_13167,N_12990,N_12891);
nand U13168 (N_13168,N_12763,N_12931);
nor U13169 (N_13169,N_12981,N_12832);
and U13170 (N_13170,N_12949,N_12826);
nand U13171 (N_13171,N_12873,N_12850);
nor U13172 (N_13172,N_12819,N_12806);
xnor U13173 (N_13173,N_12792,N_12885);
xor U13174 (N_13174,N_12974,N_12949);
or U13175 (N_13175,N_12878,N_12790);
nor U13176 (N_13176,N_12987,N_12842);
xnor U13177 (N_13177,N_12892,N_12834);
nand U13178 (N_13178,N_12794,N_12995);
nor U13179 (N_13179,N_12904,N_12892);
xor U13180 (N_13180,N_12911,N_12959);
or U13181 (N_13181,N_12833,N_12860);
nor U13182 (N_13182,N_12751,N_12891);
nand U13183 (N_13183,N_12817,N_12920);
nor U13184 (N_13184,N_12931,N_12938);
or U13185 (N_13185,N_12909,N_12849);
or U13186 (N_13186,N_12810,N_12802);
nand U13187 (N_13187,N_12954,N_12892);
nand U13188 (N_13188,N_12855,N_12782);
and U13189 (N_13189,N_12918,N_12964);
nand U13190 (N_13190,N_12957,N_12825);
nand U13191 (N_13191,N_12905,N_12987);
and U13192 (N_13192,N_12948,N_12830);
nor U13193 (N_13193,N_12772,N_12963);
nor U13194 (N_13194,N_12790,N_12937);
and U13195 (N_13195,N_12897,N_12875);
and U13196 (N_13196,N_12877,N_12759);
or U13197 (N_13197,N_12862,N_12856);
or U13198 (N_13198,N_12817,N_12852);
and U13199 (N_13199,N_12856,N_12832);
nor U13200 (N_13200,N_12835,N_12950);
or U13201 (N_13201,N_12948,N_12959);
nand U13202 (N_13202,N_12968,N_12972);
xnor U13203 (N_13203,N_12780,N_12832);
nor U13204 (N_13204,N_12780,N_12991);
xnor U13205 (N_13205,N_12760,N_12935);
nand U13206 (N_13206,N_12994,N_12846);
and U13207 (N_13207,N_12887,N_12762);
or U13208 (N_13208,N_12802,N_12983);
xnor U13209 (N_13209,N_12890,N_12952);
xnor U13210 (N_13210,N_12863,N_12764);
xor U13211 (N_13211,N_12864,N_12852);
nor U13212 (N_13212,N_12991,N_12783);
and U13213 (N_13213,N_12842,N_12960);
nor U13214 (N_13214,N_12762,N_12924);
or U13215 (N_13215,N_12857,N_12804);
or U13216 (N_13216,N_12803,N_12870);
and U13217 (N_13217,N_12875,N_12887);
xor U13218 (N_13218,N_12785,N_12790);
nand U13219 (N_13219,N_12784,N_12945);
nor U13220 (N_13220,N_12926,N_12960);
nor U13221 (N_13221,N_12955,N_12792);
xor U13222 (N_13222,N_12809,N_12888);
nand U13223 (N_13223,N_12935,N_12977);
or U13224 (N_13224,N_12758,N_12874);
or U13225 (N_13225,N_12925,N_12976);
xnor U13226 (N_13226,N_12901,N_12795);
nand U13227 (N_13227,N_12979,N_12934);
nor U13228 (N_13228,N_12805,N_12758);
or U13229 (N_13229,N_12853,N_12950);
or U13230 (N_13230,N_12890,N_12942);
nor U13231 (N_13231,N_12993,N_12992);
xnor U13232 (N_13232,N_12854,N_12812);
and U13233 (N_13233,N_12774,N_12845);
or U13234 (N_13234,N_12852,N_12988);
or U13235 (N_13235,N_12795,N_12828);
or U13236 (N_13236,N_12910,N_12759);
xor U13237 (N_13237,N_12818,N_12888);
and U13238 (N_13238,N_12851,N_12951);
xor U13239 (N_13239,N_12761,N_12925);
nand U13240 (N_13240,N_12953,N_12994);
or U13241 (N_13241,N_12790,N_12772);
nor U13242 (N_13242,N_12933,N_12787);
xor U13243 (N_13243,N_12825,N_12897);
xnor U13244 (N_13244,N_12830,N_12915);
and U13245 (N_13245,N_12917,N_12919);
nand U13246 (N_13246,N_12796,N_12944);
nor U13247 (N_13247,N_12866,N_12800);
nor U13248 (N_13248,N_12764,N_12904);
and U13249 (N_13249,N_12944,N_12799);
or U13250 (N_13250,N_13118,N_13147);
nand U13251 (N_13251,N_13222,N_13246);
nor U13252 (N_13252,N_13052,N_13072);
or U13253 (N_13253,N_13114,N_13169);
nor U13254 (N_13254,N_13020,N_13190);
nor U13255 (N_13255,N_13101,N_13047);
nor U13256 (N_13256,N_13042,N_13127);
nor U13257 (N_13257,N_13007,N_13081);
or U13258 (N_13258,N_13093,N_13155);
nand U13259 (N_13259,N_13213,N_13128);
or U13260 (N_13260,N_13091,N_13158);
nor U13261 (N_13261,N_13117,N_13129);
or U13262 (N_13262,N_13006,N_13103);
xnor U13263 (N_13263,N_13034,N_13087);
or U13264 (N_13264,N_13249,N_13029);
nand U13265 (N_13265,N_13238,N_13184);
and U13266 (N_13266,N_13240,N_13046);
xnor U13267 (N_13267,N_13172,N_13242);
nor U13268 (N_13268,N_13108,N_13200);
xnor U13269 (N_13269,N_13236,N_13159);
or U13270 (N_13270,N_13002,N_13025);
nand U13271 (N_13271,N_13062,N_13116);
xor U13272 (N_13272,N_13031,N_13037);
nand U13273 (N_13273,N_13109,N_13056);
nor U13274 (N_13274,N_13148,N_13164);
xnor U13275 (N_13275,N_13067,N_13012);
nor U13276 (N_13276,N_13119,N_13088);
xor U13277 (N_13277,N_13106,N_13153);
nand U13278 (N_13278,N_13188,N_13104);
xor U13279 (N_13279,N_13059,N_13205);
xnor U13280 (N_13280,N_13035,N_13133);
nor U13281 (N_13281,N_13115,N_13137);
xor U13282 (N_13282,N_13241,N_13013);
or U13283 (N_13283,N_13234,N_13125);
nor U13284 (N_13284,N_13022,N_13175);
nand U13285 (N_13285,N_13124,N_13207);
and U13286 (N_13286,N_13112,N_13196);
or U13287 (N_13287,N_13017,N_13201);
and U13288 (N_13288,N_13045,N_13197);
nor U13289 (N_13289,N_13065,N_13185);
nor U13290 (N_13290,N_13076,N_13192);
nand U13291 (N_13291,N_13053,N_13083);
or U13292 (N_13292,N_13174,N_13086);
xor U13293 (N_13293,N_13211,N_13161);
nor U13294 (N_13294,N_13145,N_13066);
nand U13295 (N_13295,N_13064,N_13095);
xnor U13296 (N_13296,N_13220,N_13111);
and U13297 (N_13297,N_13039,N_13160);
nor U13298 (N_13298,N_13227,N_13226);
nor U13299 (N_13299,N_13179,N_13223);
xor U13300 (N_13300,N_13015,N_13237);
xnor U13301 (N_13301,N_13177,N_13085);
nor U13302 (N_13302,N_13215,N_13110);
xor U13303 (N_13303,N_13187,N_13193);
and U13304 (N_13304,N_13030,N_13043);
or U13305 (N_13305,N_13107,N_13026);
xnor U13306 (N_13306,N_13036,N_13166);
and U13307 (N_13307,N_13217,N_13136);
nor U13308 (N_13308,N_13231,N_13141);
xnor U13309 (N_13309,N_13142,N_13221);
nand U13310 (N_13310,N_13195,N_13028);
or U13311 (N_13311,N_13230,N_13044);
xnor U13312 (N_13312,N_13152,N_13040);
or U13313 (N_13313,N_13224,N_13154);
xor U13314 (N_13314,N_13009,N_13073);
nor U13315 (N_13315,N_13173,N_13167);
and U13316 (N_13316,N_13060,N_13132);
or U13317 (N_13317,N_13123,N_13178);
or U13318 (N_13318,N_13146,N_13171);
nor U13319 (N_13319,N_13079,N_13140);
xor U13320 (N_13320,N_13181,N_13113);
nor U13321 (N_13321,N_13170,N_13003);
and U13322 (N_13322,N_13027,N_13092);
nor U13323 (N_13323,N_13245,N_13105);
nor U13324 (N_13324,N_13089,N_13168);
xor U13325 (N_13325,N_13019,N_13248);
or U13326 (N_13326,N_13162,N_13038);
xnor U13327 (N_13327,N_13218,N_13074);
nand U13328 (N_13328,N_13219,N_13055);
nor U13329 (N_13329,N_13247,N_13202);
or U13330 (N_13330,N_13130,N_13057);
or U13331 (N_13331,N_13041,N_13008);
and U13332 (N_13332,N_13239,N_13024);
xnor U13333 (N_13333,N_13198,N_13143);
nor U13334 (N_13334,N_13122,N_13100);
or U13335 (N_13335,N_13082,N_13070);
and U13336 (N_13336,N_13176,N_13021);
and U13337 (N_13337,N_13084,N_13126);
or U13338 (N_13338,N_13183,N_13078);
nor U13339 (N_13339,N_13180,N_13016);
nand U13340 (N_13340,N_13229,N_13051);
or U13341 (N_13341,N_13120,N_13135);
nor U13342 (N_13342,N_13214,N_13058);
or U13343 (N_13343,N_13049,N_13182);
nand U13344 (N_13344,N_13165,N_13102);
and U13345 (N_13345,N_13208,N_13163);
and U13346 (N_13346,N_13134,N_13225);
xor U13347 (N_13347,N_13005,N_13150);
nand U13348 (N_13348,N_13097,N_13096);
or U13349 (N_13349,N_13075,N_13149);
nand U13350 (N_13350,N_13077,N_13191);
and U13351 (N_13351,N_13209,N_13189);
and U13352 (N_13352,N_13032,N_13071);
nand U13353 (N_13353,N_13048,N_13235);
or U13354 (N_13354,N_13228,N_13080);
nor U13355 (N_13355,N_13206,N_13018);
nand U13356 (N_13356,N_13069,N_13014);
or U13357 (N_13357,N_13151,N_13004);
xnor U13358 (N_13358,N_13068,N_13233);
and U13359 (N_13359,N_13194,N_13131);
nor U13360 (N_13360,N_13204,N_13098);
xor U13361 (N_13361,N_13232,N_13243);
nand U13362 (N_13362,N_13121,N_13186);
or U13363 (N_13363,N_13023,N_13244);
or U13364 (N_13364,N_13099,N_13033);
or U13365 (N_13365,N_13000,N_13138);
nand U13366 (N_13366,N_13063,N_13212);
nor U13367 (N_13367,N_13144,N_13001);
xor U13368 (N_13368,N_13094,N_13139);
nand U13369 (N_13369,N_13210,N_13216);
or U13370 (N_13370,N_13156,N_13061);
and U13371 (N_13371,N_13010,N_13090);
nor U13372 (N_13372,N_13157,N_13203);
nor U13373 (N_13373,N_13050,N_13011);
nand U13374 (N_13374,N_13199,N_13054);
xnor U13375 (N_13375,N_13085,N_13049);
nor U13376 (N_13376,N_13001,N_13183);
or U13377 (N_13377,N_13046,N_13122);
nor U13378 (N_13378,N_13188,N_13094);
or U13379 (N_13379,N_13164,N_13106);
nand U13380 (N_13380,N_13150,N_13108);
nor U13381 (N_13381,N_13049,N_13205);
or U13382 (N_13382,N_13199,N_13241);
xor U13383 (N_13383,N_13123,N_13173);
and U13384 (N_13384,N_13227,N_13043);
xor U13385 (N_13385,N_13168,N_13237);
and U13386 (N_13386,N_13243,N_13245);
xnor U13387 (N_13387,N_13007,N_13023);
and U13388 (N_13388,N_13055,N_13082);
nor U13389 (N_13389,N_13024,N_13060);
nor U13390 (N_13390,N_13104,N_13046);
and U13391 (N_13391,N_13150,N_13124);
or U13392 (N_13392,N_13009,N_13145);
nor U13393 (N_13393,N_13194,N_13159);
nand U13394 (N_13394,N_13104,N_13148);
or U13395 (N_13395,N_13009,N_13133);
nand U13396 (N_13396,N_13048,N_13117);
nor U13397 (N_13397,N_13163,N_13242);
and U13398 (N_13398,N_13061,N_13207);
nor U13399 (N_13399,N_13005,N_13123);
xor U13400 (N_13400,N_13102,N_13144);
or U13401 (N_13401,N_13019,N_13190);
nand U13402 (N_13402,N_13210,N_13088);
nand U13403 (N_13403,N_13199,N_13013);
nor U13404 (N_13404,N_13181,N_13143);
xor U13405 (N_13405,N_13197,N_13141);
nand U13406 (N_13406,N_13048,N_13184);
nand U13407 (N_13407,N_13027,N_13052);
nand U13408 (N_13408,N_13230,N_13112);
nand U13409 (N_13409,N_13206,N_13208);
and U13410 (N_13410,N_13193,N_13174);
nor U13411 (N_13411,N_13158,N_13096);
nand U13412 (N_13412,N_13073,N_13114);
xor U13413 (N_13413,N_13168,N_13035);
nand U13414 (N_13414,N_13062,N_13219);
nor U13415 (N_13415,N_13121,N_13107);
or U13416 (N_13416,N_13229,N_13172);
xnor U13417 (N_13417,N_13155,N_13207);
nor U13418 (N_13418,N_13118,N_13201);
nand U13419 (N_13419,N_13051,N_13057);
and U13420 (N_13420,N_13013,N_13137);
xnor U13421 (N_13421,N_13102,N_13023);
or U13422 (N_13422,N_13101,N_13207);
nand U13423 (N_13423,N_13051,N_13240);
or U13424 (N_13424,N_13150,N_13001);
or U13425 (N_13425,N_13170,N_13143);
or U13426 (N_13426,N_13008,N_13228);
nor U13427 (N_13427,N_13140,N_13036);
nor U13428 (N_13428,N_13020,N_13106);
nor U13429 (N_13429,N_13158,N_13174);
nand U13430 (N_13430,N_13195,N_13002);
and U13431 (N_13431,N_13210,N_13055);
xor U13432 (N_13432,N_13109,N_13046);
and U13433 (N_13433,N_13241,N_13131);
nand U13434 (N_13434,N_13129,N_13244);
and U13435 (N_13435,N_13057,N_13185);
and U13436 (N_13436,N_13149,N_13120);
nor U13437 (N_13437,N_13199,N_13153);
nor U13438 (N_13438,N_13158,N_13221);
or U13439 (N_13439,N_13003,N_13205);
xnor U13440 (N_13440,N_13172,N_13074);
nand U13441 (N_13441,N_13236,N_13050);
or U13442 (N_13442,N_13078,N_13202);
nor U13443 (N_13443,N_13014,N_13146);
nor U13444 (N_13444,N_13044,N_13175);
or U13445 (N_13445,N_13230,N_13224);
or U13446 (N_13446,N_13182,N_13003);
nor U13447 (N_13447,N_13019,N_13053);
xnor U13448 (N_13448,N_13024,N_13020);
nand U13449 (N_13449,N_13248,N_13229);
and U13450 (N_13450,N_13049,N_13005);
nor U13451 (N_13451,N_13075,N_13182);
nand U13452 (N_13452,N_13094,N_13117);
and U13453 (N_13453,N_13216,N_13130);
nand U13454 (N_13454,N_13138,N_13051);
nor U13455 (N_13455,N_13040,N_13108);
nand U13456 (N_13456,N_13094,N_13214);
xnor U13457 (N_13457,N_13042,N_13152);
and U13458 (N_13458,N_13146,N_13167);
nand U13459 (N_13459,N_13162,N_13129);
nand U13460 (N_13460,N_13146,N_13238);
and U13461 (N_13461,N_13062,N_13005);
xnor U13462 (N_13462,N_13140,N_13171);
and U13463 (N_13463,N_13020,N_13000);
and U13464 (N_13464,N_13211,N_13233);
nor U13465 (N_13465,N_13093,N_13120);
xor U13466 (N_13466,N_13245,N_13148);
and U13467 (N_13467,N_13043,N_13081);
xor U13468 (N_13468,N_13018,N_13040);
or U13469 (N_13469,N_13178,N_13220);
xor U13470 (N_13470,N_13200,N_13180);
nand U13471 (N_13471,N_13222,N_13153);
or U13472 (N_13472,N_13033,N_13210);
nor U13473 (N_13473,N_13146,N_13025);
and U13474 (N_13474,N_13216,N_13050);
nand U13475 (N_13475,N_13109,N_13007);
or U13476 (N_13476,N_13245,N_13130);
nand U13477 (N_13477,N_13105,N_13017);
nand U13478 (N_13478,N_13073,N_13069);
or U13479 (N_13479,N_13112,N_13177);
and U13480 (N_13480,N_13096,N_13202);
or U13481 (N_13481,N_13214,N_13171);
or U13482 (N_13482,N_13217,N_13187);
nor U13483 (N_13483,N_13077,N_13051);
and U13484 (N_13484,N_13212,N_13240);
nor U13485 (N_13485,N_13054,N_13055);
or U13486 (N_13486,N_13246,N_13242);
or U13487 (N_13487,N_13147,N_13096);
nand U13488 (N_13488,N_13211,N_13232);
or U13489 (N_13489,N_13091,N_13119);
xor U13490 (N_13490,N_13103,N_13119);
xnor U13491 (N_13491,N_13052,N_13064);
and U13492 (N_13492,N_13180,N_13030);
and U13493 (N_13493,N_13220,N_13237);
nand U13494 (N_13494,N_13171,N_13127);
nand U13495 (N_13495,N_13011,N_13082);
xor U13496 (N_13496,N_13085,N_13189);
nand U13497 (N_13497,N_13159,N_13117);
nor U13498 (N_13498,N_13000,N_13223);
nand U13499 (N_13499,N_13097,N_13177);
nand U13500 (N_13500,N_13451,N_13492);
nand U13501 (N_13501,N_13470,N_13438);
nor U13502 (N_13502,N_13432,N_13400);
or U13503 (N_13503,N_13414,N_13386);
nand U13504 (N_13504,N_13367,N_13435);
xor U13505 (N_13505,N_13411,N_13368);
or U13506 (N_13506,N_13258,N_13430);
xor U13507 (N_13507,N_13403,N_13315);
nor U13508 (N_13508,N_13316,N_13477);
nand U13509 (N_13509,N_13282,N_13397);
and U13510 (N_13510,N_13441,N_13482);
nor U13511 (N_13511,N_13318,N_13480);
xnor U13512 (N_13512,N_13495,N_13335);
xnor U13513 (N_13513,N_13278,N_13450);
and U13514 (N_13514,N_13377,N_13360);
nor U13515 (N_13515,N_13291,N_13322);
xor U13516 (N_13516,N_13486,N_13396);
and U13517 (N_13517,N_13341,N_13348);
xnor U13518 (N_13518,N_13271,N_13387);
xnor U13519 (N_13519,N_13463,N_13474);
nand U13520 (N_13520,N_13263,N_13268);
nor U13521 (N_13521,N_13385,N_13356);
xnor U13522 (N_13522,N_13459,N_13256);
and U13523 (N_13523,N_13293,N_13292);
or U13524 (N_13524,N_13375,N_13274);
and U13525 (N_13525,N_13443,N_13391);
or U13526 (N_13526,N_13415,N_13369);
nor U13527 (N_13527,N_13283,N_13267);
nand U13528 (N_13528,N_13326,N_13354);
or U13529 (N_13529,N_13493,N_13276);
and U13530 (N_13530,N_13461,N_13456);
nor U13531 (N_13531,N_13261,N_13376);
and U13532 (N_13532,N_13426,N_13295);
and U13533 (N_13533,N_13380,N_13296);
and U13534 (N_13534,N_13281,N_13306);
nand U13535 (N_13535,N_13405,N_13431);
nand U13536 (N_13536,N_13317,N_13457);
or U13537 (N_13537,N_13381,N_13420);
and U13538 (N_13538,N_13408,N_13313);
nand U13539 (N_13539,N_13422,N_13378);
xor U13540 (N_13540,N_13404,N_13494);
xnor U13541 (N_13541,N_13394,N_13273);
nand U13542 (N_13542,N_13328,N_13362);
nand U13543 (N_13543,N_13334,N_13301);
nand U13544 (N_13544,N_13323,N_13320);
nor U13545 (N_13545,N_13270,N_13458);
or U13546 (N_13546,N_13314,N_13330);
nand U13547 (N_13547,N_13433,N_13344);
xor U13548 (N_13548,N_13446,N_13416);
nand U13549 (N_13549,N_13303,N_13299);
xor U13550 (N_13550,N_13436,N_13260);
or U13551 (N_13551,N_13262,N_13253);
nand U13552 (N_13552,N_13285,N_13352);
nand U13553 (N_13553,N_13478,N_13442);
or U13554 (N_13554,N_13409,N_13349);
xnor U13555 (N_13555,N_13472,N_13250);
nand U13556 (N_13556,N_13329,N_13346);
or U13557 (N_13557,N_13465,N_13350);
or U13558 (N_13558,N_13275,N_13399);
nand U13559 (N_13559,N_13312,N_13427);
and U13560 (N_13560,N_13469,N_13255);
or U13561 (N_13561,N_13388,N_13277);
or U13562 (N_13562,N_13460,N_13357);
and U13563 (N_13563,N_13307,N_13491);
xor U13564 (N_13564,N_13257,N_13393);
xor U13565 (N_13565,N_13325,N_13345);
and U13566 (N_13566,N_13452,N_13382);
nor U13567 (N_13567,N_13288,N_13289);
nor U13568 (N_13568,N_13331,N_13252);
and U13569 (N_13569,N_13475,N_13424);
nor U13570 (N_13570,N_13290,N_13332);
and U13571 (N_13571,N_13497,N_13259);
xor U13572 (N_13572,N_13351,N_13410);
xor U13573 (N_13573,N_13342,N_13490);
xor U13574 (N_13574,N_13473,N_13333);
and U13575 (N_13575,N_13398,N_13266);
nand U13576 (N_13576,N_13496,N_13309);
and U13577 (N_13577,N_13355,N_13294);
xor U13578 (N_13578,N_13280,N_13302);
nor U13579 (N_13579,N_13379,N_13437);
xor U13580 (N_13580,N_13365,N_13372);
nor U13581 (N_13581,N_13374,N_13305);
nand U13582 (N_13582,N_13310,N_13358);
and U13583 (N_13583,N_13488,N_13265);
nand U13584 (N_13584,N_13324,N_13481);
or U13585 (N_13585,N_13370,N_13336);
or U13586 (N_13586,N_13449,N_13383);
nand U13587 (N_13587,N_13251,N_13384);
xor U13588 (N_13588,N_13466,N_13371);
xnor U13589 (N_13589,N_13254,N_13407);
nor U13590 (N_13590,N_13286,N_13347);
nor U13591 (N_13591,N_13343,N_13467);
nand U13592 (N_13592,N_13359,N_13439);
xor U13593 (N_13593,N_13339,N_13304);
nor U13594 (N_13594,N_13484,N_13468);
xor U13595 (N_13595,N_13327,N_13361);
nand U13596 (N_13596,N_13479,N_13401);
nor U13597 (N_13597,N_13498,N_13340);
nand U13598 (N_13598,N_13402,N_13406);
nand U13599 (N_13599,N_13298,N_13321);
or U13600 (N_13600,N_13499,N_13421);
and U13601 (N_13601,N_13363,N_13429);
or U13602 (N_13602,N_13269,N_13308);
or U13603 (N_13603,N_13366,N_13423);
nand U13604 (N_13604,N_13300,N_13489);
nand U13605 (N_13605,N_13434,N_13485);
nand U13606 (N_13606,N_13462,N_13425);
and U13607 (N_13607,N_13287,N_13373);
and U13608 (N_13608,N_13448,N_13476);
and U13609 (N_13609,N_13338,N_13428);
xor U13610 (N_13610,N_13364,N_13455);
xnor U13611 (N_13611,N_13413,N_13389);
nand U13612 (N_13612,N_13412,N_13353);
nor U13613 (N_13613,N_13337,N_13297);
and U13614 (N_13614,N_13447,N_13311);
xor U13615 (N_13615,N_13392,N_13464);
and U13616 (N_13616,N_13395,N_13264);
and U13617 (N_13617,N_13319,N_13390);
nor U13618 (N_13618,N_13419,N_13483);
xor U13619 (N_13619,N_13471,N_13440);
nand U13620 (N_13620,N_13444,N_13272);
or U13621 (N_13621,N_13454,N_13445);
and U13622 (N_13622,N_13284,N_13417);
and U13623 (N_13623,N_13279,N_13418);
nand U13624 (N_13624,N_13487,N_13453);
nor U13625 (N_13625,N_13263,N_13259);
or U13626 (N_13626,N_13385,N_13408);
and U13627 (N_13627,N_13412,N_13379);
nor U13628 (N_13628,N_13452,N_13348);
nand U13629 (N_13629,N_13470,N_13340);
nor U13630 (N_13630,N_13362,N_13301);
xnor U13631 (N_13631,N_13393,N_13365);
or U13632 (N_13632,N_13301,N_13458);
nor U13633 (N_13633,N_13264,N_13489);
or U13634 (N_13634,N_13293,N_13493);
or U13635 (N_13635,N_13496,N_13360);
and U13636 (N_13636,N_13309,N_13302);
nor U13637 (N_13637,N_13256,N_13423);
nor U13638 (N_13638,N_13370,N_13332);
xor U13639 (N_13639,N_13478,N_13406);
or U13640 (N_13640,N_13297,N_13447);
nor U13641 (N_13641,N_13408,N_13488);
and U13642 (N_13642,N_13327,N_13257);
nor U13643 (N_13643,N_13430,N_13471);
or U13644 (N_13644,N_13340,N_13376);
nor U13645 (N_13645,N_13362,N_13260);
or U13646 (N_13646,N_13303,N_13499);
or U13647 (N_13647,N_13448,N_13428);
or U13648 (N_13648,N_13476,N_13482);
nor U13649 (N_13649,N_13366,N_13335);
nor U13650 (N_13650,N_13432,N_13279);
xnor U13651 (N_13651,N_13479,N_13389);
xnor U13652 (N_13652,N_13418,N_13338);
xnor U13653 (N_13653,N_13303,N_13359);
or U13654 (N_13654,N_13434,N_13322);
nor U13655 (N_13655,N_13288,N_13330);
nor U13656 (N_13656,N_13475,N_13444);
and U13657 (N_13657,N_13355,N_13428);
xor U13658 (N_13658,N_13497,N_13365);
xor U13659 (N_13659,N_13388,N_13445);
and U13660 (N_13660,N_13302,N_13362);
or U13661 (N_13661,N_13391,N_13473);
nand U13662 (N_13662,N_13395,N_13300);
nand U13663 (N_13663,N_13277,N_13291);
nor U13664 (N_13664,N_13266,N_13390);
or U13665 (N_13665,N_13333,N_13374);
nor U13666 (N_13666,N_13452,N_13313);
xnor U13667 (N_13667,N_13328,N_13406);
nor U13668 (N_13668,N_13452,N_13356);
or U13669 (N_13669,N_13393,N_13292);
nand U13670 (N_13670,N_13309,N_13380);
nor U13671 (N_13671,N_13414,N_13464);
and U13672 (N_13672,N_13394,N_13417);
or U13673 (N_13673,N_13261,N_13419);
and U13674 (N_13674,N_13355,N_13482);
nand U13675 (N_13675,N_13476,N_13375);
nand U13676 (N_13676,N_13349,N_13289);
and U13677 (N_13677,N_13393,N_13294);
xor U13678 (N_13678,N_13489,N_13394);
or U13679 (N_13679,N_13485,N_13355);
nand U13680 (N_13680,N_13307,N_13321);
and U13681 (N_13681,N_13344,N_13318);
nor U13682 (N_13682,N_13453,N_13468);
nand U13683 (N_13683,N_13340,N_13275);
or U13684 (N_13684,N_13321,N_13258);
and U13685 (N_13685,N_13473,N_13417);
or U13686 (N_13686,N_13274,N_13397);
xor U13687 (N_13687,N_13494,N_13267);
nor U13688 (N_13688,N_13496,N_13482);
or U13689 (N_13689,N_13283,N_13297);
nor U13690 (N_13690,N_13451,N_13411);
nand U13691 (N_13691,N_13334,N_13290);
nand U13692 (N_13692,N_13355,N_13465);
and U13693 (N_13693,N_13313,N_13448);
xor U13694 (N_13694,N_13372,N_13432);
and U13695 (N_13695,N_13324,N_13451);
xnor U13696 (N_13696,N_13483,N_13257);
or U13697 (N_13697,N_13272,N_13459);
nor U13698 (N_13698,N_13481,N_13308);
and U13699 (N_13699,N_13310,N_13472);
nand U13700 (N_13700,N_13421,N_13495);
or U13701 (N_13701,N_13332,N_13397);
xnor U13702 (N_13702,N_13263,N_13333);
xnor U13703 (N_13703,N_13311,N_13491);
and U13704 (N_13704,N_13481,N_13389);
nor U13705 (N_13705,N_13387,N_13413);
and U13706 (N_13706,N_13391,N_13276);
nor U13707 (N_13707,N_13411,N_13371);
or U13708 (N_13708,N_13253,N_13263);
nor U13709 (N_13709,N_13460,N_13376);
xnor U13710 (N_13710,N_13405,N_13320);
and U13711 (N_13711,N_13474,N_13476);
xor U13712 (N_13712,N_13280,N_13311);
nand U13713 (N_13713,N_13315,N_13458);
or U13714 (N_13714,N_13267,N_13304);
nor U13715 (N_13715,N_13331,N_13354);
or U13716 (N_13716,N_13330,N_13358);
nand U13717 (N_13717,N_13336,N_13476);
or U13718 (N_13718,N_13475,N_13381);
and U13719 (N_13719,N_13350,N_13289);
xor U13720 (N_13720,N_13314,N_13387);
nand U13721 (N_13721,N_13273,N_13316);
and U13722 (N_13722,N_13475,N_13305);
or U13723 (N_13723,N_13367,N_13268);
and U13724 (N_13724,N_13367,N_13311);
nand U13725 (N_13725,N_13410,N_13412);
nor U13726 (N_13726,N_13341,N_13380);
nor U13727 (N_13727,N_13451,N_13465);
xnor U13728 (N_13728,N_13471,N_13487);
nor U13729 (N_13729,N_13361,N_13364);
and U13730 (N_13730,N_13398,N_13485);
nor U13731 (N_13731,N_13354,N_13364);
xor U13732 (N_13732,N_13382,N_13274);
nor U13733 (N_13733,N_13300,N_13415);
or U13734 (N_13734,N_13474,N_13413);
nor U13735 (N_13735,N_13276,N_13401);
nand U13736 (N_13736,N_13392,N_13307);
nor U13737 (N_13737,N_13285,N_13469);
or U13738 (N_13738,N_13347,N_13253);
xnor U13739 (N_13739,N_13384,N_13440);
and U13740 (N_13740,N_13251,N_13422);
xor U13741 (N_13741,N_13349,N_13373);
and U13742 (N_13742,N_13382,N_13476);
nor U13743 (N_13743,N_13343,N_13338);
nand U13744 (N_13744,N_13425,N_13413);
nor U13745 (N_13745,N_13322,N_13407);
xnor U13746 (N_13746,N_13285,N_13287);
nand U13747 (N_13747,N_13364,N_13277);
xor U13748 (N_13748,N_13318,N_13391);
or U13749 (N_13749,N_13447,N_13469);
or U13750 (N_13750,N_13608,N_13527);
and U13751 (N_13751,N_13578,N_13565);
nand U13752 (N_13752,N_13514,N_13714);
or U13753 (N_13753,N_13673,N_13625);
xor U13754 (N_13754,N_13723,N_13594);
and U13755 (N_13755,N_13664,N_13557);
nand U13756 (N_13756,N_13609,N_13611);
or U13757 (N_13757,N_13727,N_13501);
nand U13758 (N_13758,N_13571,N_13573);
or U13759 (N_13759,N_13600,N_13564);
nand U13760 (N_13760,N_13712,N_13599);
nand U13761 (N_13761,N_13643,N_13633);
xnor U13762 (N_13762,N_13551,N_13660);
nor U13763 (N_13763,N_13569,N_13702);
and U13764 (N_13764,N_13544,N_13529);
or U13765 (N_13765,N_13593,N_13606);
or U13766 (N_13766,N_13685,N_13553);
xnor U13767 (N_13767,N_13743,N_13699);
nor U13768 (N_13768,N_13696,N_13604);
nor U13769 (N_13769,N_13672,N_13724);
nor U13770 (N_13770,N_13646,N_13607);
or U13771 (N_13771,N_13510,N_13575);
or U13772 (N_13772,N_13733,N_13579);
nand U13773 (N_13773,N_13654,N_13563);
xor U13774 (N_13774,N_13560,N_13642);
xor U13775 (N_13775,N_13644,N_13509);
or U13776 (N_13776,N_13624,N_13531);
and U13777 (N_13777,N_13732,N_13570);
nand U13778 (N_13778,N_13647,N_13663);
and U13779 (N_13779,N_13650,N_13735);
and U13780 (N_13780,N_13523,N_13519);
xnor U13781 (N_13781,N_13535,N_13528);
xor U13782 (N_13782,N_13645,N_13541);
nand U13783 (N_13783,N_13503,N_13636);
and U13784 (N_13784,N_13628,N_13597);
nor U13785 (N_13785,N_13512,N_13617);
or U13786 (N_13786,N_13637,N_13681);
nand U13787 (N_13787,N_13708,N_13746);
xor U13788 (N_13788,N_13567,N_13547);
nor U13789 (N_13789,N_13588,N_13556);
nand U13790 (N_13790,N_13694,N_13677);
or U13791 (N_13791,N_13602,N_13716);
or U13792 (N_13792,N_13505,N_13533);
nand U13793 (N_13793,N_13518,N_13742);
and U13794 (N_13794,N_13630,N_13520);
nand U13795 (N_13795,N_13577,N_13639);
xnor U13796 (N_13796,N_13502,N_13500);
xor U13797 (N_13797,N_13591,N_13736);
nand U13798 (N_13798,N_13561,N_13581);
nand U13799 (N_13799,N_13725,N_13615);
and U13800 (N_13800,N_13666,N_13542);
or U13801 (N_13801,N_13709,N_13703);
nor U13802 (N_13802,N_13698,N_13707);
nand U13803 (N_13803,N_13513,N_13670);
or U13804 (N_13804,N_13536,N_13667);
xnor U13805 (N_13805,N_13676,N_13635);
or U13806 (N_13806,N_13697,N_13554);
and U13807 (N_13807,N_13525,N_13586);
nor U13808 (N_13808,N_13687,N_13747);
nor U13809 (N_13809,N_13534,N_13598);
nor U13810 (N_13810,N_13731,N_13506);
and U13811 (N_13811,N_13651,N_13576);
xor U13812 (N_13812,N_13640,N_13562);
and U13813 (N_13813,N_13610,N_13711);
and U13814 (N_13814,N_13558,N_13508);
nand U13815 (N_13815,N_13587,N_13661);
or U13816 (N_13816,N_13521,N_13526);
or U13817 (N_13817,N_13678,N_13620);
nand U13818 (N_13818,N_13739,N_13621);
nand U13819 (N_13819,N_13652,N_13713);
nor U13820 (N_13820,N_13705,N_13721);
or U13821 (N_13821,N_13734,N_13744);
xnor U13822 (N_13822,N_13717,N_13690);
nor U13823 (N_13823,N_13589,N_13616);
and U13824 (N_13824,N_13638,N_13552);
xor U13825 (N_13825,N_13719,N_13582);
nand U13826 (N_13826,N_13729,N_13504);
or U13827 (N_13827,N_13655,N_13710);
xnor U13828 (N_13828,N_13631,N_13566);
nor U13829 (N_13829,N_13726,N_13596);
xnor U13830 (N_13830,N_13511,N_13585);
and U13831 (N_13831,N_13543,N_13555);
nor U13832 (N_13832,N_13539,N_13691);
nor U13833 (N_13833,N_13656,N_13540);
nand U13834 (N_13834,N_13674,N_13613);
nand U13835 (N_13835,N_13641,N_13679);
nor U13836 (N_13836,N_13706,N_13745);
xnor U13837 (N_13837,N_13740,N_13595);
nor U13838 (N_13838,N_13590,N_13653);
and U13839 (N_13839,N_13675,N_13689);
xnor U13840 (N_13840,N_13626,N_13683);
or U13841 (N_13841,N_13737,N_13549);
xnor U13842 (N_13842,N_13738,N_13669);
or U13843 (N_13843,N_13583,N_13658);
nor U13844 (N_13844,N_13648,N_13668);
xnor U13845 (N_13845,N_13704,N_13548);
and U13846 (N_13846,N_13715,N_13627);
or U13847 (N_13847,N_13516,N_13601);
nor U13848 (N_13848,N_13572,N_13684);
and U13849 (N_13849,N_13688,N_13748);
nand U13850 (N_13850,N_13692,N_13718);
xnor U13851 (N_13851,N_13612,N_13722);
and U13852 (N_13852,N_13686,N_13659);
xnor U13853 (N_13853,N_13657,N_13532);
or U13854 (N_13854,N_13614,N_13507);
nor U13855 (N_13855,N_13671,N_13749);
xor U13856 (N_13856,N_13662,N_13649);
and U13857 (N_13857,N_13522,N_13700);
or U13858 (N_13858,N_13680,N_13568);
and U13859 (N_13859,N_13550,N_13623);
nor U13860 (N_13860,N_13665,N_13530);
or U13861 (N_13861,N_13693,N_13574);
nor U13862 (N_13862,N_13695,N_13728);
nor U13863 (N_13863,N_13741,N_13537);
nor U13864 (N_13864,N_13701,N_13629);
xnor U13865 (N_13865,N_13720,N_13517);
and U13866 (N_13866,N_13515,N_13622);
nand U13867 (N_13867,N_13592,N_13580);
xnor U13868 (N_13868,N_13584,N_13730);
nor U13869 (N_13869,N_13682,N_13538);
nor U13870 (N_13870,N_13634,N_13603);
nand U13871 (N_13871,N_13545,N_13559);
nor U13872 (N_13872,N_13618,N_13619);
and U13873 (N_13873,N_13605,N_13524);
or U13874 (N_13874,N_13632,N_13546);
or U13875 (N_13875,N_13645,N_13563);
or U13876 (N_13876,N_13578,N_13720);
nor U13877 (N_13877,N_13708,N_13677);
or U13878 (N_13878,N_13543,N_13564);
xor U13879 (N_13879,N_13658,N_13714);
nand U13880 (N_13880,N_13613,N_13721);
and U13881 (N_13881,N_13517,N_13682);
xnor U13882 (N_13882,N_13694,N_13558);
and U13883 (N_13883,N_13503,N_13635);
nand U13884 (N_13884,N_13587,N_13597);
and U13885 (N_13885,N_13511,N_13734);
and U13886 (N_13886,N_13710,N_13733);
or U13887 (N_13887,N_13544,N_13515);
nor U13888 (N_13888,N_13554,N_13616);
nor U13889 (N_13889,N_13615,N_13537);
xnor U13890 (N_13890,N_13747,N_13597);
xor U13891 (N_13891,N_13523,N_13500);
or U13892 (N_13892,N_13648,N_13537);
xnor U13893 (N_13893,N_13747,N_13531);
or U13894 (N_13894,N_13623,N_13706);
nor U13895 (N_13895,N_13709,N_13677);
nand U13896 (N_13896,N_13707,N_13642);
xnor U13897 (N_13897,N_13722,N_13621);
xnor U13898 (N_13898,N_13635,N_13610);
and U13899 (N_13899,N_13708,N_13580);
nor U13900 (N_13900,N_13598,N_13713);
or U13901 (N_13901,N_13704,N_13679);
nand U13902 (N_13902,N_13568,N_13638);
and U13903 (N_13903,N_13703,N_13748);
nand U13904 (N_13904,N_13746,N_13745);
nor U13905 (N_13905,N_13642,N_13610);
xor U13906 (N_13906,N_13624,N_13663);
nand U13907 (N_13907,N_13507,N_13679);
xor U13908 (N_13908,N_13684,N_13637);
or U13909 (N_13909,N_13596,N_13741);
nor U13910 (N_13910,N_13718,N_13647);
and U13911 (N_13911,N_13642,N_13584);
xnor U13912 (N_13912,N_13519,N_13589);
nand U13913 (N_13913,N_13569,N_13635);
or U13914 (N_13914,N_13542,N_13727);
nand U13915 (N_13915,N_13719,N_13518);
xnor U13916 (N_13916,N_13562,N_13514);
nand U13917 (N_13917,N_13545,N_13621);
nor U13918 (N_13918,N_13612,N_13648);
and U13919 (N_13919,N_13628,N_13743);
nor U13920 (N_13920,N_13571,N_13569);
or U13921 (N_13921,N_13739,N_13513);
nor U13922 (N_13922,N_13561,N_13653);
nand U13923 (N_13923,N_13708,N_13726);
and U13924 (N_13924,N_13698,N_13676);
nor U13925 (N_13925,N_13574,N_13715);
or U13926 (N_13926,N_13502,N_13570);
and U13927 (N_13927,N_13725,N_13602);
nand U13928 (N_13928,N_13720,N_13649);
xor U13929 (N_13929,N_13730,N_13511);
nor U13930 (N_13930,N_13549,N_13652);
nand U13931 (N_13931,N_13500,N_13506);
nand U13932 (N_13932,N_13641,N_13646);
and U13933 (N_13933,N_13631,N_13623);
and U13934 (N_13934,N_13648,N_13640);
nand U13935 (N_13935,N_13648,N_13658);
xnor U13936 (N_13936,N_13635,N_13708);
nand U13937 (N_13937,N_13602,N_13659);
xnor U13938 (N_13938,N_13539,N_13711);
xor U13939 (N_13939,N_13523,N_13621);
nand U13940 (N_13940,N_13592,N_13613);
and U13941 (N_13941,N_13612,N_13695);
xnor U13942 (N_13942,N_13726,N_13585);
nor U13943 (N_13943,N_13588,N_13699);
nand U13944 (N_13944,N_13736,N_13528);
or U13945 (N_13945,N_13640,N_13563);
and U13946 (N_13946,N_13584,N_13703);
or U13947 (N_13947,N_13605,N_13723);
nand U13948 (N_13948,N_13571,N_13708);
or U13949 (N_13949,N_13584,N_13530);
or U13950 (N_13950,N_13717,N_13618);
and U13951 (N_13951,N_13633,N_13651);
or U13952 (N_13952,N_13733,N_13522);
nand U13953 (N_13953,N_13683,N_13592);
xor U13954 (N_13954,N_13719,N_13531);
nand U13955 (N_13955,N_13728,N_13557);
xnor U13956 (N_13956,N_13699,N_13513);
and U13957 (N_13957,N_13645,N_13748);
xnor U13958 (N_13958,N_13522,N_13613);
xor U13959 (N_13959,N_13723,N_13679);
or U13960 (N_13960,N_13680,N_13728);
and U13961 (N_13961,N_13592,N_13626);
nor U13962 (N_13962,N_13612,N_13562);
and U13963 (N_13963,N_13621,N_13591);
xnor U13964 (N_13964,N_13591,N_13659);
nand U13965 (N_13965,N_13689,N_13717);
xor U13966 (N_13966,N_13535,N_13567);
nand U13967 (N_13967,N_13581,N_13628);
nand U13968 (N_13968,N_13595,N_13532);
xnor U13969 (N_13969,N_13578,N_13559);
and U13970 (N_13970,N_13572,N_13662);
xnor U13971 (N_13971,N_13561,N_13534);
or U13972 (N_13972,N_13582,N_13571);
nand U13973 (N_13973,N_13510,N_13628);
and U13974 (N_13974,N_13557,N_13733);
nor U13975 (N_13975,N_13511,N_13573);
xor U13976 (N_13976,N_13658,N_13594);
nand U13977 (N_13977,N_13620,N_13633);
and U13978 (N_13978,N_13600,N_13672);
nand U13979 (N_13979,N_13687,N_13691);
xnor U13980 (N_13980,N_13534,N_13662);
and U13981 (N_13981,N_13619,N_13652);
nand U13982 (N_13982,N_13587,N_13578);
and U13983 (N_13983,N_13737,N_13639);
nor U13984 (N_13984,N_13574,N_13556);
nand U13985 (N_13985,N_13567,N_13686);
nor U13986 (N_13986,N_13533,N_13717);
nor U13987 (N_13987,N_13717,N_13540);
and U13988 (N_13988,N_13508,N_13526);
nor U13989 (N_13989,N_13608,N_13687);
xor U13990 (N_13990,N_13514,N_13644);
nand U13991 (N_13991,N_13525,N_13721);
nor U13992 (N_13992,N_13653,N_13721);
xnor U13993 (N_13993,N_13675,N_13627);
nor U13994 (N_13994,N_13613,N_13600);
nand U13995 (N_13995,N_13709,N_13501);
xor U13996 (N_13996,N_13677,N_13522);
xnor U13997 (N_13997,N_13740,N_13553);
or U13998 (N_13998,N_13584,N_13735);
nor U13999 (N_13999,N_13558,N_13662);
nand U14000 (N_14000,N_13754,N_13946);
and U14001 (N_14001,N_13771,N_13949);
nor U14002 (N_14002,N_13940,N_13934);
and U14003 (N_14003,N_13799,N_13789);
and U14004 (N_14004,N_13860,N_13933);
nor U14005 (N_14005,N_13752,N_13883);
or U14006 (N_14006,N_13819,N_13865);
nand U14007 (N_14007,N_13906,N_13810);
nand U14008 (N_14008,N_13975,N_13976);
nor U14009 (N_14009,N_13972,N_13973);
and U14010 (N_14010,N_13825,N_13968);
xnor U14011 (N_14011,N_13838,N_13922);
nand U14012 (N_14012,N_13854,N_13872);
xor U14013 (N_14013,N_13790,N_13868);
or U14014 (N_14014,N_13891,N_13850);
or U14015 (N_14015,N_13966,N_13842);
or U14016 (N_14016,N_13924,N_13987);
nand U14017 (N_14017,N_13923,N_13928);
or U14018 (N_14018,N_13885,N_13858);
nor U14019 (N_14019,N_13775,N_13770);
or U14020 (N_14020,N_13892,N_13920);
nor U14021 (N_14021,N_13795,N_13958);
nor U14022 (N_14022,N_13916,N_13926);
or U14023 (N_14023,N_13828,N_13794);
or U14024 (N_14024,N_13846,N_13767);
nor U14025 (N_14025,N_13751,N_13985);
and U14026 (N_14026,N_13802,N_13970);
and U14027 (N_14027,N_13758,N_13899);
or U14028 (N_14028,N_13978,N_13941);
xnor U14029 (N_14029,N_13833,N_13932);
xnor U14030 (N_14030,N_13896,N_13874);
or U14031 (N_14031,N_13894,N_13855);
nand U14032 (N_14032,N_13929,N_13994);
nor U14033 (N_14033,N_13804,N_13768);
or U14034 (N_14034,N_13753,N_13847);
or U14035 (N_14035,N_13982,N_13818);
nor U14036 (N_14036,N_13829,N_13851);
nor U14037 (N_14037,N_13814,N_13957);
nor U14038 (N_14038,N_13859,N_13871);
nand U14039 (N_14039,N_13888,N_13852);
xor U14040 (N_14040,N_13988,N_13956);
nor U14041 (N_14041,N_13834,N_13950);
or U14042 (N_14042,N_13881,N_13911);
nor U14043 (N_14043,N_13884,N_13800);
and U14044 (N_14044,N_13953,N_13817);
nand U14045 (N_14045,N_13784,N_13843);
nor U14046 (N_14046,N_13866,N_13826);
xnor U14047 (N_14047,N_13918,N_13857);
xor U14048 (N_14048,N_13919,N_13897);
and U14049 (N_14049,N_13764,N_13787);
and U14050 (N_14050,N_13880,N_13965);
xnor U14051 (N_14051,N_13938,N_13772);
and U14052 (N_14052,N_13925,N_13796);
or U14053 (N_14053,N_13807,N_13763);
nor U14054 (N_14054,N_13889,N_13766);
xnor U14055 (N_14055,N_13990,N_13954);
xor U14056 (N_14056,N_13944,N_13902);
nand U14057 (N_14057,N_13979,N_13867);
xnor U14058 (N_14058,N_13806,N_13983);
nand U14059 (N_14059,N_13853,N_13831);
nor U14060 (N_14060,N_13797,N_13921);
or U14061 (N_14061,N_13769,N_13836);
nor U14062 (N_14062,N_13830,N_13820);
xnor U14063 (N_14063,N_13750,N_13844);
nand U14064 (N_14064,N_13912,N_13952);
xnor U14065 (N_14065,N_13783,N_13937);
xor U14066 (N_14066,N_13890,N_13822);
xor U14067 (N_14067,N_13986,N_13993);
xnor U14068 (N_14068,N_13913,N_13759);
xor U14069 (N_14069,N_13862,N_13960);
nand U14070 (N_14070,N_13882,N_13876);
nand U14071 (N_14071,N_13908,N_13887);
nand U14072 (N_14072,N_13879,N_13995);
or U14073 (N_14073,N_13963,N_13875);
nor U14074 (N_14074,N_13774,N_13832);
xnor U14075 (N_14075,N_13870,N_13984);
nand U14076 (N_14076,N_13809,N_13815);
nand U14077 (N_14077,N_13935,N_13861);
nand U14078 (N_14078,N_13808,N_13936);
and U14079 (N_14079,N_13792,N_13786);
nand U14080 (N_14080,N_13962,N_13878);
xor U14081 (N_14081,N_13930,N_13917);
nand U14082 (N_14082,N_13755,N_13863);
nor U14083 (N_14083,N_13910,N_13948);
nor U14084 (N_14084,N_13989,N_13848);
xor U14085 (N_14085,N_13779,N_13840);
nand U14086 (N_14086,N_13777,N_13942);
and U14087 (N_14087,N_13907,N_13856);
or U14088 (N_14088,N_13793,N_13904);
nand U14089 (N_14089,N_13886,N_13841);
nand U14090 (N_14090,N_13823,N_13757);
xnor U14091 (N_14091,N_13816,N_13901);
or U14092 (N_14092,N_13864,N_13959);
or U14093 (N_14093,N_13827,N_13801);
or U14094 (N_14094,N_13895,N_13805);
or U14095 (N_14095,N_13943,N_13931);
nand U14096 (N_14096,N_13893,N_13781);
and U14097 (N_14097,N_13803,N_13996);
nand U14098 (N_14098,N_13773,N_13900);
nor U14099 (N_14099,N_13997,N_13778);
xnor U14100 (N_14100,N_13811,N_13756);
xnor U14101 (N_14101,N_13877,N_13824);
nand U14102 (N_14102,N_13909,N_13969);
nand U14103 (N_14103,N_13782,N_13998);
or U14104 (N_14104,N_13914,N_13839);
or U14105 (N_14105,N_13798,N_13903);
and U14106 (N_14106,N_13905,N_13788);
nor U14107 (N_14107,N_13813,N_13999);
and U14108 (N_14108,N_13776,N_13967);
and U14109 (N_14109,N_13947,N_13873);
or U14110 (N_14110,N_13974,N_13761);
xor U14111 (N_14111,N_13837,N_13964);
or U14112 (N_14112,N_13981,N_13762);
xor U14113 (N_14113,N_13992,N_13760);
xnor U14114 (N_14114,N_13845,N_13821);
nand U14115 (N_14115,N_13785,N_13977);
and U14116 (N_14116,N_13765,N_13961);
and U14117 (N_14117,N_13971,N_13812);
and U14118 (N_14118,N_13849,N_13945);
nor U14119 (N_14119,N_13780,N_13955);
nor U14120 (N_14120,N_13915,N_13791);
nand U14121 (N_14121,N_13980,N_13835);
nor U14122 (N_14122,N_13927,N_13898);
nor U14123 (N_14123,N_13951,N_13869);
and U14124 (N_14124,N_13939,N_13991);
xnor U14125 (N_14125,N_13886,N_13775);
or U14126 (N_14126,N_13764,N_13869);
nand U14127 (N_14127,N_13876,N_13870);
and U14128 (N_14128,N_13990,N_13966);
xnor U14129 (N_14129,N_13819,N_13867);
or U14130 (N_14130,N_13904,N_13974);
and U14131 (N_14131,N_13819,N_13813);
or U14132 (N_14132,N_13847,N_13806);
nand U14133 (N_14133,N_13902,N_13817);
nand U14134 (N_14134,N_13838,N_13904);
xnor U14135 (N_14135,N_13914,N_13869);
xnor U14136 (N_14136,N_13885,N_13804);
and U14137 (N_14137,N_13884,N_13839);
nor U14138 (N_14138,N_13879,N_13898);
or U14139 (N_14139,N_13795,N_13893);
nand U14140 (N_14140,N_13842,N_13896);
and U14141 (N_14141,N_13794,N_13755);
and U14142 (N_14142,N_13859,N_13930);
nand U14143 (N_14143,N_13943,N_13754);
xnor U14144 (N_14144,N_13823,N_13879);
nor U14145 (N_14145,N_13976,N_13926);
nand U14146 (N_14146,N_13767,N_13872);
and U14147 (N_14147,N_13895,N_13817);
or U14148 (N_14148,N_13823,N_13934);
or U14149 (N_14149,N_13996,N_13773);
xor U14150 (N_14150,N_13903,N_13886);
or U14151 (N_14151,N_13967,N_13876);
nor U14152 (N_14152,N_13902,N_13900);
xor U14153 (N_14153,N_13956,N_13792);
xor U14154 (N_14154,N_13786,N_13866);
nand U14155 (N_14155,N_13793,N_13958);
or U14156 (N_14156,N_13793,N_13820);
xor U14157 (N_14157,N_13920,N_13845);
nand U14158 (N_14158,N_13957,N_13803);
and U14159 (N_14159,N_13939,N_13854);
xor U14160 (N_14160,N_13982,N_13979);
nor U14161 (N_14161,N_13755,N_13775);
nor U14162 (N_14162,N_13755,N_13820);
or U14163 (N_14163,N_13793,N_13932);
or U14164 (N_14164,N_13889,N_13767);
xnor U14165 (N_14165,N_13977,N_13837);
nand U14166 (N_14166,N_13951,N_13870);
xnor U14167 (N_14167,N_13764,N_13825);
and U14168 (N_14168,N_13893,N_13884);
nor U14169 (N_14169,N_13840,N_13941);
nand U14170 (N_14170,N_13984,N_13980);
and U14171 (N_14171,N_13988,N_13900);
nand U14172 (N_14172,N_13921,N_13972);
nand U14173 (N_14173,N_13908,N_13831);
nor U14174 (N_14174,N_13829,N_13803);
nand U14175 (N_14175,N_13918,N_13951);
nor U14176 (N_14176,N_13952,N_13999);
nor U14177 (N_14177,N_13988,N_13798);
nor U14178 (N_14178,N_13837,N_13840);
or U14179 (N_14179,N_13890,N_13762);
nand U14180 (N_14180,N_13952,N_13832);
nor U14181 (N_14181,N_13816,N_13825);
or U14182 (N_14182,N_13887,N_13758);
xor U14183 (N_14183,N_13813,N_13873);
xor U14184 (N_14184,N_13825,N_13902);
or U14185 (N_14185,N_13830,N_13751);
nor U14186 (N_14186,N_13999,N_13770);
xnor U14187 (N_14187,N_13758,N_13940);
or U14188 (N_14188,N_13890,N_13954);
nand U14189 (N_14189,N_13871,N_13907);
nor U14190 (N_14190,N_13965,N_13905);
or U14191 (N_14191,N_13996,N_13957);
nor U14192 (N_14192,N_13874,N_13997);
nand U14193 (N_14193,N_13829,N_13897);
xnor U14194 (N_14194,N_13873,N_13956);
nand U14195 (N_14195,N_13857,N_13915);
nor U14196 (N_14196,N_13752,N_13816);
xnor U14197 (N_14197,N_13798,N_13826);
nor U14198 (N_14198,N_13837,N_13901);
nand U14199 (N_14199,N_13811,N_13777);
and U14200 (N_14200,N_13956,N_13858);
or U14201 (N_14201,N_13956,N_13761);
or U14202 (N_14202,N_13999,N_13877);
or U14203 (N_14203,N_13975,N_13948);
nor U14204 (N_14204,N_13985,N_13895);
nor U14205 (N_14205,N_13845,N_13849);
nand U14206 (N_14206,N_13964,N_13906);
and U14207 (N_14207,N_13939,N_13834);
and U14208 (N_14208,N_13814,N_13969);
nand U14209 (N_14209,N_13932,N_13861);
nand U14210 (N_14210,N_13786,N_13916);
or U14211 (N_14211,N_13924,N_13978);
and U14212 (N_14212,N_13754,N_13952);
or U14213 (N_14213,N_13816,N_13947);
xnor U14214 (N_14214,N_13767,N_13989);
nor U14215 (N_14215,N_13923,N_13775);
or U14216 (N_14216,N_13857,N_13767);
xnor U14217 (N_14217,N_13932,N_13962);
xnor U14218 (N_14218,N_13986,N_13851);
and U14219 (N_14219,N_13878,N_13948);
nor U14220 (N_14220,N_13806,N_13814);
or U14221 (N_14221,N_13788,N_13867);
nand U14222 (N_14222,N_13805,N_13825);
xnor U14223 (N_14223,N_13752,N_13789);
xor U14224 (N_14224,N_13878,N_13762);
xor U14225 (N_14225,N_13888,N_13754);
xnor U14226 (N_14226,N_13918,N_13809);
and U14227 (N_14227,N_13840,N_13970);
or U14228 (N_14228,N_13979,N_13799);
xnor U14229 (N_14229,N_13763,N_13798);
or U14230 (N_14230,N_13815,N_13843);
nand U14231 (N_14231,N_13979,N_13904);
and U14232 (N_14232,N_13951,N_13963);
nor U14233 (N_14233,N_13925,N_13927);
nor U14234 (N_14234,N_13791,N_13998);
or U14235 (N_14235,N_13869,N_13754);
and U14236 (N_14236,N_13996,N_13944);
nor U14237 (N_14237,N_13936,N_13884);
or U14238 (N_14238,N_13983,N_13917);
xnor U14239 (N_14239,N_13882,N_13951);
nor U14240 (N_14240,N_13947,N_13829);
or U14241 (N_14241,N_13931,N_13865);
nand U14242 (N_14242,N_13945,N_13814);
xnor U14243 (N_14243,N_13914,N_13919);
nand U14244 (N_14244,N_13918,N_13835);
or U14245 (N_14245,N_13861,N_13781);
nor U14246 (N_14246,N_13777,N_13873);
nor U14247 (N_14247,N_13993,N_13908);
and U14248 (N_14248,N_13806,N_13928);
or U14249 (N_14249,N_13946,N_13781);
or U14250 (N_14250,N_14219,N_14163);
or U14251 (N_14251,N_14104,N_14034);
or U14252 (N_14252,N_14142,N_14127);
nand U14253 (N_14253,N_14113,N_14121);
or U14254 (N_14254,N_14095,N_14144);
and U14255 (N_14255,N_14009,N_14176);
or U14256 (N_14256,N_14040,N_14189);
nor U14257 (N_14257,N_14161,N_14173);
and U14258 (N_14258,N_14226,N_14096);
and U14259 (N_14259,N_14202,N_14013);
nand U14260 (N_14260,N_14086,N_14243);
nor U14261 (N_14261,N_14099,N_14087);
or U14262 (N_14262,N_14147,N_14111);
and U14263 (N_14263,N_14151,N_14048);
xnor U14264 (N_14264,N_14187,N_14084);
xnor U14265 (N_14265,N_14145,N_14108);
or U14266 (N_14266,N_14129,N_14184);
nand U14267 (N_14267,N_14124,N_14133);
nand U14268 (N_14268,N_14010,N_14165);
nand U14269 (N_14269,N_14126,N_14168);
and U14270 (N_14270,N_14230,N_14071);
and U14271 (N_14271,N_14088,N_14026);
nor U14272 (N_14272,N_14159,N_14122);
nor U14273 (N_14273,N_14069,N_14238);
or U14274 (N_14274,N_14244,N_14059);
nor U14275 (N_14275,N_14052,N_14123);
nor U14276 (N_14276,N_14208,N_14216);
nor U14277 (N_14277,N_14101,N_14190);
and U14278 (N_14278,N_14058,N_14228);
nor U14279 (N_14279,N_14150,N_14209);
nand U14280 (N_14280,N_14049,N_14178);
and U14281 (N_14281,N_14140,N_14054);
and U14282 (N_14282,N_14037,N_14091);
or U14283 (N_14283,N_14043,N_14152);
nor U14284 (N_14284,N_14195,N_14229);
or U14285 (N_14285,N_14005,N_14172);
xnor U14286 (N_14286,N_14130,N_14023);
or U14287 (N_14287,N_14249,N_14109);
nor U14288 (N_14288,N_14118,N_14128);
or U14289 (N_14289,N_14004,N_14085);
xor U14290 (N_14290,N_14039,N_14000);
nor U14291 (N_14291,N_14060,N_14138);
xor U14292 (N_14292,N_14207,N_14115);
nor U14293 (N_14293,N_14107,N_14021);
nand U14294 (N_14294,N_14082,N_14032);
xor U14295 (N_14295,N_14197,N_14092);
xnor U14296 (N_14296,N_14192,N_14193);
or U14297 (N_14297,N_14075,N_14210);
nand U14298 (N_14298,N_14100,N_14248);
and U14299 (N_14299,N_14204,N_14081);
or U14300 (N_14300,N_14031,N_14132);
or U14301 (N_14301,N_14076,N_14025);
nand U14302 (N_14302,N_14246,N_14239);
nand U14303 (N_14303,N_14055,N_14169);
or U14304 (N_14304,N_14149,N_14029);
and U14305 (N_14305,N_14131,N_14155);
or U14306 (N_14306,N_14218,N_14074);
or U14307 (N_14307,N_14064,N_14241);
nor U14308 (N_14308,N_14215,N_14030);
nand U14309 (N_14309,N_14094,N_14196);
nor U14310 (N_14310,N_14045,N_14233);
nand U14311 (N_14311,N_14047,N_14205);
xor U14312 (N_14312,N_14212,N_14186);
and U14313 (N_14313,N_14120,N_14027);
and U14314 (N_14314,N_14154,N_14102);
xor U14315 (N_14315,N_14072,N_14234);
xnor U14316 (N_14316,N_14182,N_14158);
and U14317 (N_14317,N_14139,N_14177);
and U14318 (N_14318,N_14106,N_14153);
xor U14319 (N_14319,N_14162,N_14056);
xor U14320 (N_14320,N_14028,N_14008);
nand U14321 (N_14321,N_14134,N_14146);
and U14322 (N_14322,N_14035,N_14175);
nand U14323 (N_14323,N_14116,N_14224);
nor U14324 (N_14324,N_14235,N_14174);
xnor U14325 (N_14325,N_14185,N_14214);
and U14326 (N_14326,N_14166,N_14232);
and U14327 (N_14327,N_14198,N_14194);
and U14328 (N_14328,N_14199,N_14170);
nor U14329 (N_14329,N_14135,N_14156);
or U14330 (N_14330,N_14062,N_14203);
and U14331 (N_14331,N_14223,N_14167);
or U14332 (N_14332,N_14070,N_14020);
nand U14333 (N_14333,N_14018,N_14042);
nor U14334 (N_14334,N_14024,N_14053);
and U14335 (N_14335,N_14022,N_14011);
xnor U14336 (N_14336,N_14077,N_14080);
and U14337 (N_14337,N_14119,N_14201);
and U14338 (N_14338,N_14157,N_14006);
or U14339 (N_14339,N_14007,N_14213);
xnor U14340 (N_14340,N_14180,N_14242);
xnor U14341 (N_14341,N_14017,N_14225);
and U14342 (N_14342,N_14044,N_14110);
or U14343 (N_14343,N_14211,N_14068);
and U14344 (N_14344,N_14061,N_14217);
nor U14345 (N_14345,N_14137,N_14220);
nand U14346 (N_14346,N_14093,N_14002);
and U14347 (N_14347,N_14014,N_14103);
nand U14348 (N_14348,N_14206,N_14083);
and U14349 (N_14349,N_14148,N_14143);
nand U14350 (N_14350,N_14036,N_14019);
nand U14351 (N_14351,N_14236,N_14181);
xor U14352 (N_14352,N_14038,N_14245);
xnor U14353 (N_14353,N_14171,N_14078);
nor U14354 (N_14354,N_14066,N_14046);
nor U14355 (N_14355,N_14136,N_14125);
and U14356 (N_14356,N_14117,N_14015);
nand U14357 (N_14357,N_14097,N_14237);
nor U14358 (N_14358,N_14067,N_14050);
xnor U14359 (N_14359,N_14098,N_14221);
or U14360 (N_14360,N_14231,N_14051);
nor U14361 (N_14361,N_14183,N_14063);
nand U14362 (N_14362,N_14112,N_14079);
nor U14363 (N_14363,N_14191,N_14041);
and U14364 (N_14364,N_14012,N_14200);
or U14365 (N_14365,N_14105,N_14089);
xnor U14366 (N_14366,N_14057,N_14033);
nor U14367 (N_14367,N_14065,N_14001);
nor U14368 (N_14368,N_14160,N_14247);
or U14369 (N_14369,N_14073,N_14227);
nand U14370 (N_14370,N_14188,N_14179);
nor U14371 (N_14371,N_14240,N_14164);
nand U14372 (N_14372,N_14090,N_14141);
or U14373 (N_14373,N_14222,N_14016);
or U14374 (N_14374,N_14114,N_14003);
xor U14375 (N_14375,N_14202,N_14167);
nor U14376 (N_14376,N_14113,N_14010);
nand U14377 (N_14377,N_14028,N_14082);
or U14378 (N_14378,N_14144,N_14186);
and U14379 (N_14379,N_14003,N_14240);
nor U14380 (N_14380,N_14112,N_14050);
nor U14381 (N_14381,N_14099,N_14196);
xnor U14382 (N_14382,N_14075,N_14135);
xor U14383 (N_14383,N_14153,N_14012);
xnor U14384 (N_14384,N_14182,N_14207);
xnor U14385 (N_14385,N_14022,N_14159);
nor U14386 (N_14386,N_14071,N_14154);
nor U14387 (N_14387,N_14086,N_14145);
nand U14388 (N_14388,N_14185,N_14032);
and U14389 (N_14389,N_14227,N_14174);
and U14390 (N_14390,N_14011,N_14084);
or U14391 (N_14391,N_14240,N_14104);
and U14392 (N_14392,N_14052,N_14174);
nor U14393 (N_14393,N_14249,N_14235);
xnor U14394 (N_14394,N_14034,N_14164);
xnor U14395 (N_14395,N_14089,N_14043);
nor U14396 (N_14396,N_14053,N_14080);
nand U14397 (N_14397,N_14160,N_14180);
nor U14398 (N_14398,N_14122,N_14047);
nand U14399 (N_14399,N_14112,N_14201);
nand U14400 (N_14400,N_14159,N_14114);
nor U14401 (N_14401,N_14151,N_14166);
nor U14402 (N_14402,N_14184,N_14133);
xnor U14403 (N_14403,N_14221,N_14047);
and U14404 (N_14404,N_14029,N_14126);
or U14405 (N_14405,N_14017,N_14135);
nor U14406 (N_14406,N_14009,N_14055);
nand U14407 (N_14407,N_14206,N_14178);
or U14408 (N_14408,N_14165,N_14038);
and U14409 (N_14409,N_14078,N_14112);
nor U14410 (N_14410,N_14111,N_14153);
nand U14411 (N_14411,N_14001,N_14043);
or U14412 (N_14412,N_14004,N_14083);
xor U14413 (N_14413,N_14170,N_14237);
nand U14414 (N_14414,N_14160,N_14050);
or U14415 (N_14415,N_14022,N_14077);
nor U14416 (N_14416,N_14032,N_14097);
xor U14417 (N_14417,N_14146,N_14136);
and U14418 (N_14418,N_14052,N_14067);
nand U14419 (N_14419,N_14236,N_14120);
or U14420 (N_14420,N_14166,N_14031);
xor U14421 (N_14421,N_14110,N_14035);
nor U14422 (N_14422,N_14055,N_14013);
nand U14423 (N_14423,N_14189,N_14044);
or U14424 (N_14424,N_14211,N_14239);
nand U14425 (N_14425,N_14001,N_14062);
nor U14426 (N_14426,N_14015,N_14237);
xnor U14427 (N_14427,N_14111,N_14101);
nand U14428 (N_14428,N_14165,N_14013);
xnor U14429 (N_14429,N_14048,N_14190);
xnor U14430 (N_14430,N_14203,N_14033);
or U14431 (N_14431,N_14002,N_14100);
nor U14432 (N_14432,N_14021,N_14056);
or U14433 (N_14433,N_14059,N_14052);
and U14434 (N_14434,N_14195,N_14185);
nor U14435 (N_14435,N_14150,N_14184);
or U14436 (N_14436,N_14192,N_14170);
xor U14437 (N_14437,N_14219,N_14214);
and U14438 (N_14438,N_14063,N_14210);
nand U14439 (N_14439,N_14198,N_14092);
or U14440 (N_14440,N_14059,N_14224);
xnor U14441 (N_14441,N_14188,N_14149);
xnor U14442 (N_14442,N_14061,N_14001);
or U14443 (N_14443,N_14182,N_14014);
nand U14444 (N_14444,N_14178,N_14023);
nor U14445 (N_14445,N_14242,N_14136);
nand U14446 (N_14446,N_14070,N_14149);
and U14447 (N_14447,N_14121,N_14031);
or U14448 (N_14448,N_14103,N_14195);
nand U14449 (N_14449,N_14249,N_14125);
nor U14450 (N_14450,N_14153,N_14183);
or U14451 (N_14451,N_14139,N_14099);
nand U14452 (N_14452,N_14213,N_14117);
nand U14453 (N_14453,N_14140,N_14188);
and U14454 (N_14454,N_14004,N_14180);
nand U14455 (N_14455,N_14207,N_14160);
or U14456 (N_14456,N_14176,N_14165);
nand U14457 (N_14457,N_14117,N_14127);
xnor U14458 (N_14458,N_14092,N_14094);
nor U14459 (N_14459,N_14102,N_14068);
or U14460 (N_14460,N_14069,N_14208);
and U14461 (N_14461,N_14070,N_14015);
and U14462 (N_14462,N_14135,N_14052);
or U14463 (N_14463,N_14051,N_14161);
nor U14464 (N_14464,N_14001,N_14033);
nor U14465 (N_14465,N_14055,N_14193);
and U14466 (N_14466,N_14133,N_14016);
and U14467 (N_14467,N_14234,N_14137);
and U14468 (N_14468,N_14168,N_14030);
and U14469 (N_14469,N_14199,N_14135);
and U14470 (N_14470,N_14153,N_14209);
or U14471 (N_14471,N_14238,N_14117);
or U14472 (N_14472,N_14200,N_14030);
nand U14473 (N_14473,N_14221,N_14051);
and U14474 (N_14474,N_14015,N_14227);
or U14475 (N_14475,N_14236,N_14145);
nor U14476 (N_14476,N_14021,N_14034);
xor U14477 (N_14477,N_14158,N_14238);
xor U14478 (N_14478,N_14131,N_14210);
and U14479 (N_14479,N_14047,N_14231);
xor U14480 (N_14480,N_14171,N_14087);
or U14481 (N_14481,N_14069,N_14175);
xnor U14482 (N_14482,N_14102,N_14176);
nor U14483 (N_14483,N_14105,N_14080);
nor U14484 (N_14484,N_14247,N_14035);
nand U14485 (N_14485,N_14206,N_14176);
or U14486 (N_14486,N_14120,N_14057);
or U14487 (N_14487,N_14122,N_14169);
nand U14488 (N_14488,N_14048,N_14174);
nand U14489 (N_14489,N_14142,N_14039);
nand U14490 (N_14490,N_14071,N_14166);
or U14491 (N_14491,N_14032,N_14020);
nor U14492 (N_14492,N_14123,N_14110);
nor U14493 (N_14493,N_14048,N_14185);
or U14494 (N_14494,N_14015,N_14132);
or U14495 (N_14495,N_14149,N_14047);
nand U14496 (N_14496,N_14025,N_14012);
or U14497 (N_14497,N_14142,N_14081);
nor U14498 (N_14498,N_14021,N_14128);
nor U14499 (N_14499,N_14179,N_14053);
xor U14500 (N_14500,N_14443,N_14489);
nor U14501 (N_14501,N_14376,N_14374);
and U14502 (N_14502,N_14430,N_14251);
nor U14503 (N_14503,N_14455,N_14316);
nand U14504 (N_14504,N_14420,N_14383);
or U14505 (N_14505,N_14260,N_14313);
and U14506 (N_14506,N_14451,N_14319);
nor U14507 (N_14507,N_14478,N_14291);
or U14508 (N_14508,N_14388,N_14437);
and U14509 (N_14509,N_14367,N_14457);
and U14510 (N_14510,N_14395,N_14447);
nor U14511 (N_14511,N_14336,N_14351);
nor U14512 (N_14512,N_14427,N_14378);
nor U14513 (N_14513,N_14481,N_14488);
nand U14514 (N_14514,N_14302,N_14497);
nand U14515 (N_14515,N_14352,N_14261);
or U14516 (N_14516,N_14359,N_14333);
or U14517 (N_14517,N_14450,N_14458);
nor U14518 (N_14518,N_14343,N_14360);
and U14519 (N_14519,N_14473,N_14477);
and U14520 (N_14520,N_14357,N_14328);
and U14521 (N_14521,N_14309,N_14256);
or U14522 (N_14522,N_14363,N_14446);
xor U14523 (N_14523,N_14331,N_14304);
nor U14524 (N_14524,N_14461,N_14305);
nor U14525 (N_14525,N_14252,N_14334);
and U14526 (N_14526,N_14298,N_14280);
xor U14527 (N_14527,N_14433,N_14371);
or U14528 (N_14528,N_14267,N_14327);
and U14529 (N_14529,N_14468,N_14475);
or U14530 (N_14530,N_14417,N_14425);
nor U14531 (N_14531,N_14315,N_14295);
xnor U14532 (N_14532,N_14423,N_14469);
nand U14533 (N_14533,N_14470,N_14426);
or U14534 (N_14534,N_14342,N_14472);
or U14535 (N_14535,N_14496,N_14255);
or U14536 (N_14536,N_14403,N_14467);
nand U14537 (N_14537,N_14414,N_14306);
or U14538 (N_14538,N_14284,N_14321);
or U14539 (N_14539,N_14325,N_14320);
nand U14540 (N_14540,N_14441,N_14381);
or U14541 (N_14541,N_14391,N_14289);
nand U14542 (N_14542,N_14275,N_14292);
xnor U14543 (N_14543,N_14375,N_14448);
nor U14544 (N_14544,N_14404,N_14462);
or U14545 (N_14545,N_14296,N_14397);
nor U14546 (N_14546,N_14384,N_14262);
or U14547 (N_14547,N_14372,N_14366);
and U14548 (N_14548,N_14364,N_14459);
nor U14549 (N_14549,N_14483,N_14377);
and U14550 (N_14550,N_14438,N_14283);
and U14551 (N_14551,N_14353,N_14393);
or U14552 (N_14552,N_14308,N_14281);
nand U14553 (N_14553,N_14449,N_14382);
nor U14554 (N_14554,N_14345,N_14491);
and U14555 (N_14555,N_14282,N_14408);
nor U14556 (N_14556,N_14499,N_14370);
or U14557 (N_14557,N_14286,N_14407);
nand U14558 (N_14558,N_14277,N_14299);
or U14559 (N_14559,N_14330,N_14390);
nand U14560 (N_14560,N_14338,N_14415);
or U14561 (N_14561,N_14350,N_14479);
nand U14562 (N_14562,N_14314,N_14294);
nand U14563 (N_14563,N_14268,N_14484);
nor U14564 (N_14564,N_14487,N_14263);
or U14565 (N_14565,N_14410,N_14394);
nand U14566 (N_14566,N_14402,N_14265);
and U14567 (N_14567,N_14419,N_14464);
nand U14568 (N_14568,N_14317,N_14411);
or U14569 (N_14569,N_14344,N_14264);
xnor U14570 (N_14570,N_14398,N_14482);
or U14571 (N_14571,N_14322,N_14271);
or U14572 (N_14572,N_14369,N_14358);
and U14573 (N_14573,N_14365,N_14361);
or U14574 (N_14574,N_14444,N_14399);
nor U14575 (N_14575,N_14498,N_14356);
and U14576 (N_14576,N_14288,N_14278);
nor U14577 (N_14577,N_14346,N_14290);
xnor U14578 (N_14578,N_14380,N_14412);
nor U14579 (N_14579,N_14465,N_14273);
or U14580 (N_14580,N_14386,N_14293);
xor U14581 (N_14581,N_14335,N_14416);
nor U14582 (N_14582,N_14349,N_14266);
or U14583 (N_14583,N_14396,N_14490);
nand U14584 (N_14584,N_14254,N_14259);
and U14585 (N_14585,N_14400,N_14494);
and U14586 (N_14586,N_14337,N_14318);
or U14587 (N_14587,N_14347,N_14418);
xnor U14588 (N_14588,N_14454,N_14435);
nand U14589 (N_14589,N_14354,N_14332);
or U14590 (N_14590,N_14387,N_14297);
xnor U14591 (N_14591,N_14274,N_14310);
or U14592 (N_14592,N_14401,N_14434);
or U14593 (N_14593,N_14431,N_14474);
xor U14594 (N_14594,N_14436,N_14406);
and U14595 (N_14595,N_14287,N_14452);
nand U14596 (N_14596,N_14456,N_14476);
nand U14597 (N_14597,N_14413,N_14439);
or U14598 (N_14598,N_14392,N_14300);
nor U14599 (N_14599,N_14348,N_14253);
or U14600 (N_14600,N_14373,N_14303);
xnor U14601 (N_14601,N_14269,N_14270);
nand U14602 (N_14602,N_14301,N_14453);
nand U14603 (N_14603,N_14341,N_14440);
and U14604 (N_14604,N_14424,N_14311);
xor U14605 (N_14605,N_14279,N_14492);
nor U14606 (N_14606,N_14485,N_14422);
or U14607 (N_14607,N_14257,N_14324);
and U14608 (N_14608,N_14285,N_14409);
and U14609 (N_14609,N_14272,N_14405);
xor U14610 (N_14610,N_14463,N_14429);
nor U14611 (N_14611,N_14486,N_14368);
nor U14612 (N_14612,N_14471,N_14493);
and U14613 (N_14613,N_14312,N_14307);
nand U14614 (N_14614,N_14340,N_14339);
and U14615 (N_14615,N_14276,N_14421);
nand U14616 (N_14616,N_14323,N_14460);
nand U14617 (N_14617,N_14355,N_14432);
xnor U14618 (N_14618,N_14329,N_14495);
nand U14619 (N_14619,N_14362,N_14385);
nor U14620 (N_14620,N_14326,N_14389);
or U14621 (N_14621,N_14442,N_14250);
or U14622 (N_14622,N_14258,N_14379);
nor U14623 (N_14623,N_14445,N_14480);
or U14624 (N_14624,N_14466,N_14428);
and U14625 (N_14625,N_14376,N_14342);
nor U14626 (N_14626,N_14461,N_14261);
or U14627 (N_14627,N_14406,N_14265);
nor U14628 (N_14628,N_14439,N_14395);
and U14629 (N_14629,N_14387,N_14467);
or U14630 (N_14630,N_14397,N_14269);
xnor U14631 (N_14631,N_14354,N_14414);
and U14632 (N_14632,N_14398,N_14349);
and U14633 (N_14633,N_14347,N_14404);
xor U14634 (N_14634,N_14393,N_14440);
nor U14635 (N_14635,N_14287,N_14473);
nand U14636 (N_14636,N_14252,N_14425);
nor U14637 (N_14637,N_14427,N_14496);
nand U14638 (N_14638,N_14468,N_14286);
and U14639 (N_14639,N_14267,N_14420);
xnor U14640 (N_14640,N_14401,N_14274);
xnor U14641 (N_14641,N_14335,N_14417);
nor U14642 (N_14642,N_14286,N_14483);
and U14643 (N_14643,N_14478,N_14343);
nor U14644 (N_14644,N_14434,N_14305);
xnor U14645 (N_14645,N_14324,N_14425);
xor U14646 (N_14646,N_14388,N_14330);
xor U14647 (N_14647,N_14256,N_14370);
nand U14648 (N_14648,N_14461,N_14301);
xnor U14649 (N_14649,N_14294,N_14359);
xor U14650 (N_14650,N_14319,N_14412);
nand U14651 (N_14651,N_14403,N_14297);
nand U14652 (N_14652,N_14498,N_14327);
or U14653 (N_14653,N_14430,N_14314);
xor U14654 (N_14654,N_14374,N_14280);
or U14655 (N_14655,N_14367,N_14270);
nand U14656 (N_14656,N_14452,N_14355);
nor U14657 (N_14657,N_14351,N_14307);
xor U14658 (N_14658,N_14284,N_14330);
nand U14659 (N_14659,N_14400,N_14292);
nand U14660 (N_14660,N_14359,N_14322);
or U14661 (N_14661,N_14402,N_14303);
nand U14662 (N_14662,N_14285,N_14440);
xnor U14663 (N_14663,N_14298,N_14412);
or U14664 (N_14664,N_14318,N_14388);
nor U14665 (N_14665,N_14494,N_14373);
nand U14666 (N_14666,N_14251,N_14273);
or U14667 (N_14667,N_14320,N_14360);
xor U14668 (N_14668,N_14475,N_14414);
nand U14669 (N_14669,N_14470,N_14273);
and U14670 (N_14670,N_14487,N_14333);
nor U14671 (N_14671,N_14367,N_14479);
and U14672 (N_14672,N_14285,N_14467);
nor U14673 (N_14673,N_14251,N_14474);
nand U14674 (N_14674,N_14331,N_14276);
and U14675 (N_14675,N_14258,N_14268);
nand U14676 (N_14676,N_14488,N_14435);
nand U14677 (N_14677,N_14430,N_14466);
nand U14678 (N_14678,N_14364,N_14485);
and U14679 (N_14679,N_14355,N_14275);
and U14680 (N_14680,N_14320,N_14464);
or U14681 (N_14681,N_14299,N_14465);
and U14682 (N_14682,N_14464,N_14452);
xnor U14683 (N_14683,N_14326,N_14361);
and U14684 (N_14684,N_14353,N_14433);
xor U14685 (N_14685,N_14406,N_14448);
nand U14686 (N_14686,N_14363,N_14380);
and U14687 (N_14687,N_14496,N_14482);
and U14688 (N_14688,N_14355,N_14374);
nand U14689 (N_14689,N_14389,N_14336);
and U14690 (N_14690,N_14421,N_14268);
or U14691 (N_14691,N_14488,N_14259);
or U14692 (N_14692,N_14278,N_14420);
xor U14693 (N_14693,N_14481,N_14348);
nor U14694 (N_14694,N_14413,N_14444);
and U14695 (N_14695,N_14358,N_14375);
nor U14696 (N_14696,N_14292,N_14495);
and U14697 (N_14697,N_14479,N_14377);
nand U14698 (N_14698,N_14269,N_14413);
and U14699 (N_14699,N_14482,N_14287);
nor U14700 (N_14700,N_14455,N_14445);
xor U14701 (N_14701,N_14324,N_14391);
nand U14702 (N_14702,N_14281,N_14254);
nand U14703 (N_14703,N_14401,N_14422);
xnor U14704 (N_14704,N_14434,N_14493);
xor U14705 (N_14705,N_14326,N_14273);
nor U14706 (N_14706,N_14399,N_14469);
nor U14707 (N_14707,N_14423,N_14470);
nor U14708 (N_14708,N_14467,N_14486);
nor U14709 (N_14709,N_14376,N_14395);
nand U14710 (N_14710,N_14367,N_14264);
or U14711 (N_14711,N_14263,N_14425);
xor U14712 (N_14712,N_14456,N_14443);
nor U14713 (N_14713,N_14381,N_14463);
nand U14714 (N_14714,N_14315,N_14356);
nor U14715 (N_14715,N_14495,N_14306);
or U14716 (N_14716,N_14259,N_14303);
xnor U14717 (N_14717,N_14417,N_14268);
or U14718 (N_14718,N_14373,N_14382);
or U14719 (N_14719,N_14497,N_14479);
nor U14720 (N_14720,N_14277,N_14418);
nor U14721 (N_14721,N_14416,N_14276);
xor U14722 (N_14722,N_14305,N_14445);
xor U14723 (N_14723,N_14427,N_14476);
and U14724 (N_14724,N_14315,N_14280);
xnor U14725 (N_14725,N_14408,N_14345);
xor U14726 (N_14726,N_14447,N_14456);
or U14727 (N_14727,N_14312,N_14459);
or U14728 (N_14728,N_14289,N_14429);
xnor U14729 (N_14729,N_14379,N_14422);
nand U14730 (N_14730,N_14337,N_14373);
xor U14731 (N_14731,N_14372,N_14377);
xnor U14732 (N_14732,N_14276,N_14303);
and U14733 (N_14733,N_14288,N_14465);
and U14734 (N_14734,N_14486,N_14340);
nand U14735 (N_14735,N_14251,N_14383);
nand U14736 (N_14736,N_14419,N_14395);
nand U14737 (N_14737,N_14388,N_14482);
and U14738 (N_14738,N_14492,N_14330);
and U14739 (N_14739,N_14409,N_14297);
or U14740 (N_14740,N_14405,N_14484);
nand U14741 (N_14741,N_14384,N_14276);
nand U14742 (N_14742,N_14416,N_14467);
nand U14743 (N_14743,N_14481,N_14400);
nor U14744 (N_14744,N_14362,N_14390);
nand U14745 (N_14745,N_14375,N_14409);
or U14746 (N_14746,N_14425,N_14407);
nand U14747 (N_14747,N_14314,N_14308);
or U14748 (N_14748,N_14443,N_14389);
or U14749 (N_14749,N_14373,N_14392);
xor U14750 (N_14750,N_14647,N_14694);
nor U14751 (N_14751,N_14617,N_14599);
nor U14752 (N_14752,N_14581,N_14635);
xor U14753 (N_14753,N_14667,N_14658);
nand U14754 (N_14754,N_14646,N_14552);
nor U14755 (N_14755,N_14651,N_14640);
nand U14756 (N_14756,N_14563,N_14678);
xnor U14757 (N_14757,N_14727,N_14573);
xor U14758 (N_14758,N_14601,N_14534);
xor U14759 (N_14759,N_14564,N_14560);
or U14760 (N_14760,N_14621,N_14548);
nor U14761 (N_14761,N_14590,N_14686);
xnor U14762 (N_14762,N_14521,N_14645);
nand U14763 (N_14763,N_14711,N_14541);
and U14764 (N_14764,N_14605,N_14712);
nor U14765 (N_14765,N_14510,N_14539);
or U14766 (N_14766,N_14574,N_14631);
and U14767 (N_14767,N_14503,N_14526);
xor U14768 (N_14768,N_14682,N_14629);
xnor U14769 (N_14769,N_14636,N_14662);
nor U14770 (N_14770,N_14738,N_14623);
and U14771 (N_14771,N_14668,N_14537);
and U14772 (N_14772,N_14693,N_14654);
xnor U14773 (N_14773,N_14559,N_14703);
nand U14774 (N_14774,N_14611,N_14737);
nand U14775 (N_14775,N_14557,N_14575);
nand U14776 (N_14776,N_14562,N_14749);
or U14777 (N_14777,N_14543,N_14642);
or U14778 (N_14778,N_14570,N_14596);
xor U14779 (N_14779,N_14698,N_14707);
nor U14780 (N_14780,N_14615,N_14660);
xor U14781 (N_14781,N_14530,N_14744);
nand U14782 (N_14782,N_14613,N_14592);
xor U14783 (N_14783,N_14593,N_14598);
or U14784 (N_14784,N_14536,N_14677);
and U14785 (N_14785,N_14718,N_14577);
and U14786 (N_14786,N_14696,N_14514);
or U14787 (N_14787,N_14533,N_14710);
nor U14788 (N_14788,N_14716,N_14715);
nor U14789 (N_14789,N_14544,N_14512);
nand U14790 (N_14790,N_14525,N_14729);
and U14791 (N_14791,N_14743,N_14723);
xnor U14792 (N_14792,N_14670,N_14506);
xnor U14793 (N_14793,N_14697,N_14622);
and U14794 (N_14794,N_14714,N_14532);
nand U14795 (N_14795,N_14553,N_14607);
xor U14796 (N_14796,N_14602,N_14620);
and U14797 (N_14797,N_14535,N_14556);
and U14798 (N_14798,N_14547,N_14673);
and U14799 (N_14799,N_14665,N_14614);
and U14800 (N_14800,N_14587,N_14604);
or U14801 (N_14801,N_14566,N_14666);
nor U14802 (N_14802,N_14683,N_14674);
or U14803 (N_14803,N_14511,N_14661);
nor U14804 (N_14804,N_14612,N_14679);
nand U14805 (N_14805,N_14721,N_14546);
xor U14806 (N_14806,N_14549,N_14681);
xor U14807 (N_14807,N_14583,N_14745);
or U14808 (N_14808,N_14644,N_14515);
nor U14809 (N_14809,N_14569,N_14639);
or U14810 (N_14810,N_14747,N_14641);
xnor U14811 (N_14811,N_14634,N_14695);
or U14812 (N_14812,N_14616,N_14702);
nor U14813 (N_14813,N_14627,N_14586);
xor U14814 (N_14814,N_14637,N_14701);
nor U14815 (N_14815,N_14656,N_14603);
or U14816 (N_14816,N_14568,N_14588);
and U14817 (N_14817,N_14584,N_14709);
xor U14818 (N_14818,N_14728,N_14507);
or U14819 (N_14819,N_14688,N_14519);
or U14820 (N_14820,N_14578,N_14731);
or U14821 (N_14821,N_14672,N_14531);
xnor U14822 (N_14822,N_14555,N_14746);
or U14823 (N_14823,N_14580,N_14739);
xnor U14824 (N_14824,N_14517,N_14748);
nor U14825 (N_14825,N_14504,N_14567);
nor U14826 (N_14826,N_14554,N_14505);
or U14827 (N_14827,N_14740,N_14609);
or U14828 (N_14828,N_14565,N_14619);
nand U14829 (N_14829,N_14725,N_14527);
nor U14830 (N_14830,N_14545,N_14671);
xor U14831 (N_14831,N_14523,N_14502);
or U14832 (N_14832,N_14520,N_14529);
xor U14833 (N_14833,N_14522,N_14579);
nand U14834 (N_14834,N_14628,N_14501);
and U14835 (N_14835,N_14676,N_14595);
and U14836 (N_14836,N_14691,N_14509);
and U14837 (N_14837,N_14659,N_14600);
and U14838 (N_14838,N_14708,N_14606);
or U14839 (N_14839,N_14730,N_14741);
nand U14840 (N_14840,N_14513,N_14690);
and U14841 (N_14841,N_14508,N_14540);
xor U14842 (N_14842,N_14551,N_14726);
xnor U14843 (N_14843,N_14518,N_14624);
nand U14844 (N_14844,N_14528,N_14632);
and U14845 (N_14845,N_14608,N_14524);
xnor U14846 (N_14846,N_14732,N_14582);
and U14847 (N_14847,N_14664,N_14663);
nand U14848 (N_14848,N_14638,N_14655);
nor U14849 (N_14849,N_14550,N_14652);
and U14850 (N_14850,N_14675,N_14643);
or U14851 (N_14851,N_14648,N_14500);
and U14852 (N_14852,N_14722,N_14653);
nor U14853 (N_14853,N_14657,N_14561);
and U14854 (N_14854,N_14717,N_14649);
and U14855 (N_14855,N_14633,N_14687);
and U14856 (N_14856,N_14571,N_14700);
and U14857 (N_14857,N_14735,N_14719);
xor U14858 (N_14858,N_14736,N_14576);
nor U14859 (N_14859,N_14585,N_14538);
nand U14860 (N_14860,N_14734,N_14594);
nand U14861 (N_14861,N_14572,N_14742);
nand U14862 (N_14862,N_14689,N_14692);
nor U14863 (N_14863,N_14610,N_14618);
and U14864 (N_14864,N_14699,N_14684);
nor U14865 (N_14865,N_14597,N_14589);
nand U14866 (N_14866,N_14558,N_14680);
or U14867 (N_14867,N_14591,N_14630);
or U14868 (N_14868,N_14685,N_14733);
nand U14869 (N_14869,N_14720,N_14705);
and U14870 (N_14870,N_14669,N_14706);
nand U14871 (N_14871,N_14724,N_14625);
xor U14872 (N_14872,N_14626,N_14713);
xor U14873 (N_14873,N_14650,N_14704);
and U14874 (N_14874,N_14516,N_14542);
nand U14875 (N_14875,N_14552,N_14538);
and U14876 (N_14876,N_14598,N_14670);
or U14877 (N_14877,N_14647,N_14640);
nand U14878 (N_14878,N_14593,N_14572);
nand U14879 (N_14879,N_14697,N_14510);
and U14880 (N_14880,N_14521,N_14571);
or U14881 (N_14881,N_14528,N_14737);
xnor U14882 (N_14882,N_14715,N_14592);
nor U14883 (N_14883,N_14621,N_14587);
nor U14884 (N_14884,N_14707,N_14582);
xnor U14885 (N_14885,N_14652,N_14634);
and U14886 (N_14886,N_14637,N_14746);
and U14887 (N_14887,N_14538,N_14714);
and U14888 (N_14888,N_14705,N_14545);
and U14889 (N_14889,N_14588,N_14574);
or U14890 (N_14890,N_14649,N_14675);
and U14891 (N_14891,N_14642,N_14617);
xnor U14892 (N_14892,N_14733,N_14686);
xor U14893 (N_14893,N_14681,N_14740);
or U14894 (N_14894,N_14546,N_14604);
and U14895 (N_14895,N_14636,N_14549);
and U14896 (N_14896,N_14604,N_14547);
nand U14897 (N_14897,N_14731,N_14726);
or U14898 (N_14898,N_14550,N_14531);
nand U14899 (N_14899,N_14640,N_14711);
or U14900 (N_14900,N_14576,N_14574);
and U14901 (N_14901,N_14653,N_14507);
nor U14902 (N_14902,N_14531,N_14742);
nor U14903 (N_14903,N_14749,N_14563);
or U14904 (N_14904,N_14555,N_14508);
and U14905 (N_14905,N_14605,N_14553);
and U14906 (N_14906,N_14673,N_14587);
nand U14907 (N_14907,N_14593,N_14587);
and U14908 (N_14908,N_14616,N_14598);
nor U14909 (N_14909,N_14607,N_14716);
xor U14910 (N_14910,N_14721,N_14748);
or U14911 (N_14911,N_14563,N_14618);
and U14912 (N_14912,N_14620,N_14647);
and U14913 (N_14913,N_14698,N_14690);
or U14914 (N_14914,N_14725,N_14732);
nor U14915 (N_14915,N_14716,N_14510);
or U14916 (N_14916,N_14590,N_14697);
xnor U14917 (N_14917,N_14679,N_14732);
nand U14918 (N_14918,N_14586,N_14673);
nand U14919 (N_14919,N_14634,N_14707);
nor U14920 (N_14920,N_14688,N_14638);
nor U14921 (N_14921,N_14687,N_14611);
xor U14922 (N_14922,N_14576,N_14510);
xnor U14923 (N_14923,N_14527,N_14693);
nor U14924 (N_14924,N_14631,N_14634);
nand U14925 (N_14925,N_14672,N_14642);
xnor U14926 (N_14926,N_14643,N_14687);
or U14927 (N_14927,N_14524,N_14641);
nor U14928 (N_14928,N_14715,N_14728);
xor U14929 (N_14929,N_14552,N_14648);
xor U14930 (N_14930,N_14540,N_14692);
and U14931 (N_14931,N_14642,N_14614);
nor U14932 (N_14932,N_14725,N_14666);
nand U14933 (N_14933,N_14646,N_14699);
or U14934 (N_14934,N_14512,N_14702);
xnor U14935 (N_14935,N_14556,N_14747);
and U14936 (N_14936,N_14592,N_14616);
nor U14937 (N_14937,N_14514,N_14703);
nor U14938 (N_14938,N_14639,N_14664);
xor U14939 (N_14939,N_14716,N_14519);
and U14940 (N_14940,N_14724,N_14682);
or U14941 (N_14941,N_14558,N_14713);
and U14942 (N_14942,N_14628,N_14544);
and U14943 (N_14943,N_14577,N_14532);
and U14944 (N_14944,N_14565,N_14748);
nand U14945 (N_14945,N_14599,N_14610);
nand U14946 (N_14946,N_14516,N_14630);
or U14947 (N_14947,N_14543,N_14548);
or U14948 (N_14948,N_14508,N_14704);
nor U14949 (N_14949,N_14583,N_14711);
nor U14950 (N_14950,N_14549,N_14525);
xor U14951 (N_14951,N_14513,N_14652);
xnor U14952 (N_14952,N_14560,N_14721);
or U14953 (N_14953,N_14502,N_14696);
or U14954 (N_14954,N_14529,N_14646);
nand U14955 (N_14955,N_14591,N_14730);
nor U14956 (N_14956,N_14543,N_14527);
and U14957 (N_14957,N_14733,N_14640);
xor U14958 (N_14958,N_14505,N_14515);
nand U14959 (N_14959,N_14636,N_14726);
xor U14960 (N_14960,N_14540,N_14728);
xnor U14961 (N_14961,N_14603,N_14744);
or U14962 (N_14962,N_14557,N_14508);
nor U14963 (N_14963,N_14510,N_14609);
or U14964 (N_14964,N_14692,N_14628);
and U14965 (N_14965,N_14506,N_14699);
xnor U14966 (N_14966,N_14603,N_14637);
xnor U14967 (N_14967,N_14581,N_14583);
or U14968 (N_14968,N_14529,N_14736);
and U14969 (N_14969,N_14502,N_14747);
and U14970 (N_14970,N_14745,N_14525);
or U14971 (N_14971,N_14530,N_14622);
xor U14972 (N_14972,N_14588,N_14603);
xnor U14973 (N_14973,N_14729,N_14658);
and U14974 (N_14974,N_14583,N_14692);
or U14975 (N_14975,N_14572,N_14708);
or U14976 (N_14976,N_14547,N_14602);
nand U14977 (N_14977,N_14675,N_14614);
and U14978 (N_14978,N_14505,N_14555);
or U14979 (N_14979,N_14588,N_14531);
xor U14980 (N_14980,N_14648,N_14728);
xor U14981 (N_14981,N_14640,N_14542);
nor U14982 (N_14982,N_14580,N_14606);
and U14983 (N_14983,N_14678,N_14580);
nor U14984 (N_14984,N_14569,N_14577);
and U14985 (N_14985,N_14710,N_14620);
xor U14986 (N_14986,N_14576,N_14673);
nand U14987 (N_14987,N_14541,N_14654);
or U14988 (N_14988,N_14633,N_14519);
nor U14989 (N_14989,N_14510,N_14578);
nand U14990 (N_14990,N_14650,N_14666);
nor U14991 (N_14991,N_14713,N_14593);
and U14992 (N_14992,N_14522,N_14696);
nor U14993 (N_14993,N_14627,N_14636);
nand U14994 (N_14994,N_14631,N_14526);
nor U14995 (N_14995,N_14662,N_14528);
nand U14996 (N_14996,N_14596,N_14675);
and U14997 (N_14997,N_14729,N_14565);
and U14998 (N_14998,N_14527,N_14523);
nand U14999 (N_14999,N_14729,N_14585);
or U15000 (N_15000,N_14853,N_14866);
nor U15001 (N_15001,N_14910,N_14871);
nand U15002 (N_15002,N_14868,N_14872);
or U15003 (N_15003,N_14880,N_14856);
nand U15004 (N_15004,N_14836,N_14979);
and U15005 (N_15005,N_14827,N_14977);
xnor U15006 (N_15006,N_14839,N_14790);
or U15007 (N_15007,N_14958,N_14787);
xor U15008 (N_15008,N_14819,N_14922);
nand U15009 (N_15009,N_14821,N_14881);
nor U15010 (N_15010,N_14884,N_14953);
or U15011 (N_15011,N_14993,N_14937);
or U15012 (N_15012,N_14899,N_14861);
xnor U15013 (N_15013,N_14998,N_14971);
and U15014 (N_15014,N_14931,N_14756);
nand U15015 (N_15015,N_14852,N_14994);
nand U15016 (N_15016,N_14810,N_14895);
and U15017 (N_15017,N_14923,N_14945);
nand U15018 (N_15018,N_14905,N_14833);
nand U15019 (N_15019,N_14893,N_14844);
nor U15020 (N_15020,N_14894,N_14890);
nand U15021 (N_15021,N_14802,N_14974);
xor U15022 (N_15022,N_14942,N_14939);
and U15023 (N_15023,N_14855,N_14764);
xnor U15024 (N_15024,N_14877,N_14999);
xor U15025 (N_15025,N_14938,N_14875);
nor U15026 (N_15026,N_14943,N_14759);
nand U15027 (N_15027,N_14948,N_14930);
and U15028 (N_15028,N_14978,N_14793);
and U15029 (N_15029,N_14825,N_14796);
and U15030 (N_15030,N_14799,N_14824);
nor U15031 (N_15031,N_14800,N_14924);
or U15032 (N_15032,N_14838,N_14865);
xnor U15033 (N_15033,N_14901,N_14753);
or U15034 (N_15034,N_14988,N_14961);
xnor U15035 (N_15035,N_14935,N_14878);
and U15036 (N_15036,N_14959,N_14830);
or U15037 (N_15037,N_14849,N_14752);
nor U15038 (N_15038,N_14768,N_14897);
nor U15039 (N_15039,N_14889,N_14826);
and U15040 (N_15040,N_14968,N_14774);
nor U15041 (N_15041,N_14987,N_14904);
or U15042 (N_15042,N_14927,N_14990);
and U15043 (N_15043,N_14820,N_14792);
or U15044 (N_15044,N_14760,N_14869);
nand U15045 (N_15045,N_14883,N_14912);
or U15046 (N_15046,N_14860,N_14777);
nor U15047 (N_15047,N_14850,N_14828);
or U15048 (N_15048,N_14786,N_14807);
and U15049 (N_15049,N_14892,N_14887);
xnor U15050 (N_15050,N_14929,N_14914);
and U15051 (N_15051,N_14863,N_14921);
or U15052 (N_15052,N_14908,N_14947);
nor U15053 (N_15053,N_14982,N_14829);
nor U15054 (N_15054,N_14925,N_14970);
nand U15055 (N_15055,N_14885,N_14870);
xor U15056 (N_15056,N_14915,N_14794);
and U15057 (N_15057,N_14791,N_14754);
xor U15058 (N_15058,N_14903,N_14812);
nor U15059 (N_15059,N_14803,N_14801);
xnor U15060 (N_15060,N_14842,N_14778);
nor U15061 (N_15061,N_14864,N_14769);
or U15062 (N_15062,N_14972,N_14751);
nand U15063 (N_15063,N_14804,N_14995);
or U15064 (N_15064,N_14831,N_14985);
nand U15065 (N_15065,N_14795,N_14837);
or U15066 (N_15066,N_14996,N_14811);
xnor U15067 (N_15067,N_14962,N_14976);
or U15068 (N_15068,N_14785,N_14991);
nor U15069 (N_15069,N_14960,N_14989);
xnor U15070 (N_15070,N_14859,N_14954);
or U15071 (N_15071,N_14967,N_14900);
nor U15072 (N_15072,N_14784,N_14834);
nor U15073 (N_15073,N_14808,N_14775);
nand U15074 (N_15074,N_14886,N_14771);
and U15075 (N_15075,N_14817,N_14873);
and U15076 (N_15076,N_14770,N_14944);
or U15077 (N_15077,N_14975,N_14815);
or U15078 (N_15078,N_14783,N_14832);
xnor U15079 (N_15079,N_14940,N_14858);
nor U15080 (N_15080,N_14762,N_14980);
nand U15081 (N_15081,N_14920,N_14766);
and U15082 (N_15082,N_14780,N_14907);
and U15083 (N_15083,N_14969,N_14896);
nor U15084 (N_15084,N_14765,N_14898);
nand U15085 (N_15085,N_14781,N_14957);
xnor U15086 (N_15086,N_14919,N_14917);
nand U15087 (N_15087,N_14755,N_14986);
nand U15088 (N_15088,N_14862,N_14902);
nand U15089 (N_15089,N_14973,N_14867);
nand U15090 (N_15090,N_14936,N_14916);
xor U15091 (N_15091,N_14984,N_14997);
or U15092 (N_15092,N_14963,N_14934);
or U15093 (N_15093,N_14965,N_14840);
xnor U15094 (N_15094,N_14846,N_14797);
or U15095 (N_15095,N_14798,N_14805);
or U15096 (N_15096,N_14882,N_14776);
or U15097 (N_15097,N_14822,N_14941);
nand U15098 (N_15098,N_14750,N_14763);
nand U15099 (N_15099,N_14757,N_14788);
nor U15100 (N_15100,N_14964,N_14951);
xnor U15101 (N_15101,N_14789,N_14818);
nand U15102 (N_15102,N_14933,N_14823);
nor U15103 (N_15103,N_14835,N_14857);
or U15104 (N_15104,N_14848,N_14932);
nand U15105 (N_15105,N_14949,N_14806);
or U15106 (N_15106,N_14876,N_14879);
nand U15107 (N_15107,N_14847,N_14955);
and U15108 (N_15108,N_14841,N_14913);
or U15109 (N_15109,N_14854,N_14845);
or U15110 (N_15110,N_14950,N_14843);
or U15111 (N_15111,N_14816,N_14891);
or U15112 (N_15112,N_14851,N_14814);
and U15113 (N_15113,N_14906,N_14779);
or U15114 (N_15114,N_14952,N_14773);
xor U15115 (N_15115,N_14992,N_14761);
or U15116 (N_15116,N_14926,N_14758);
and U15117 (N_15117,N_14928,N_14981);
or U15118 (N_15118,N_14782,N_14888);
and U15119 (N_15119,N_14772,N_14956);
nand U15120 (N_15120,N_14918,N_14813);
nand U15121 (N_15121,N_14966,N_14983);
or U15122 (N_15122,N_14767,N_14909);
nor U15123 (N_15123,N_14911,N_14946);
or U15124 (N_15124,N_14874,N_14809);
nand U15125 (N_15125,N_14755,N_14933);
xnor U15126 (N_15126,N_14840,N_14946);
xnor U15127 (N_15127,N_14959,N_14967);
nand U15128 (N_15128,N_14913,N_14858);
nand U15129 (N_15129,N_14911,N_14982);
and U15130 (N_15130,N_14874,N_14987);
xor U15131 (N_15131,N_14884,N_14979);
and U15132 (N_15132,N_14974,N_14965);
xnor U15133 (N_15133,N_14801,N_14802);
or U15134 (N_15134,N_14895,N_14772);
xnor U15135 (N_15135,N_14933,N_14882);
or U15136 (N_15136,N_14768,N_14942);
and U15137 (N_15137,N_14759,N_14824);
or U15138 (N_15138,N_14801,N_14794);
or U15139 (N_15139,N_14964,N_14888);
and U15140 (N_15140,N_14913,N_14987);
xnor U15141 (N_15141,N_14883,N_14847);
or U15142 (N_15142,N_14752,N_14957);
nand U15143 (N_15143,N_14802,N_14825);
xnor U15144 (N_15144,N_14954,N_14973);
nor U15145 (N_15145,N_14830,N_14885);
xor U15146 (N_15146,N_14837,N_14824);
xor U15147 (N_15147,N_14992,N_14760);
and U15148 (N_15148,N_14937,N_14944);
and U15149 (N_15149,N_14895,N_14947);
xnor U15150 (N_15150,N_14775,N_14960);
xor U15151 (N_15151,N_14780,N_14844);
nor U15152 (N_15152,N_14897,N_14959);
nand U15153 (N_15153,N_14778,N_14956);
or U15154 (N_15154,N_14981,N_14824);
xnor U15155 (N_15155,N_14760,N_14922);
or U15156 (N_15156,N_14763,N_14956);
xor U15157 (N_15157,N_14791,N_14772);
and U15158 (N_15158,N_14853,N_14932);
nor U15159 (N_15159,N_14815,N_14933);
or U15160 (N_15160,N_14798,N_14797);
nand U15161 (N_15161,N_14827,N_14825);
nor U15162 (N_15162,N_14927,N_14992);
xnor U15163 (N_15163,N_14931,N_14966);
xnor U15164 (N_15164,N_14918,N_14858);
xor U15165 (N_15165,N_14989,N_14866);
nor U15166 (N_15166,N_14762,N_14979);
nand U15167 (N_15167,N_14771,N_14777);
nand U15168 (N_15168,N_14838,N_14875);
and U15169 (N_15169,N_14855,N_14776);
nand U15170 (N_15170,N_14910,N_14750);
and U15171 (N_15171,N_14778,N_14915);
xor U15172 (N_15172,N_14864,N_14897);
nor U15173 (N_15173,N_14988,N_14908);
nor U15174 (N_15174,N_14834,N_14894);
or U15175 (N_15175,N_14960,N_14976);
and U15176 (N_15176,N_14998,N_14838);
and U15177 (N_15177,N_14911,N_14900);
or U15178 (N_15178,N_14875,N_14972);
or U15179 (N_15179,N_14785,N_14805);
nand U15180 (N_15180,N_14879,N_14788);
nor U15181 (N_15181,N_14773,N_14924);
xnor U15182 (N_15182,N_14869,N_14802);
nor U15183 (N_15183,N_14958,N_14932);
nor U15184 (N_15184,N_14769,N_14928);
and U15185 (N_15185,N_14848,N_14906);
and U15186 (N_15186,N_14756,N_14823);
and U15187 (N_15187,N_14915,N_14869);
or U15188 (N_15188,N_14802,N_14978);
xor U15189 (N_15189,N_14913,N_14992);
or U15190 (N_15190,N_14952,N_14986);
and U15191 (N_15191,N_14959,N_14969);
xor U15192 (N_15192,N_14756,N_14940);
and U15193 (N_15193,N_14781,N_14820);
or U15194 (N_15194,N_14754,N_14970);
or U15195 (N_15195,N_14838,N_14837);
nor U15196 (N_15196,N_14802,N_14848);
nor U15197 (N_15197,N_14841,N_14957);
nor U15198 (N_15198,N_14943,N_14917);
and U15199 (N_15199,N_14795,N_14927);
nand U15200 (N_15200,N_14795,N_14859);
nor U15201 (N_15201,N_14812,N_14860);
nand U15202 (N_15202,N_14862,N_14765);
and U15203 (N_15203,N_14989,N_14930);
or U15204 (N_15204,N_14905,N_14785);
nand U15205 (N_15205,N_14921,N_14966);
xnor U15206 (N_15206,N_14764,N_14829);
nor U15207 (N_15207,N_14771,N_14908);
xnor U15208 (N_15208,N_14761,N_14976);
nand U15209 (N_15209,N_14988,N_14968);
xnor U15210 (N_15210,N_14905,N_14808);
nor U15211 (N_15211,N_14806,N_14753);
and U15212 (N_15212,N_14931,N_14962);
xor U15213 (N_15213,N_14814,N_14890);
and U15214 (N_15214,N_14930,N_14789);
nand U15215 (N_15215,N_14905,N_14979);
and U15216 (N_15216,N_14925,N_14996);
nand U15217 (N_15217,N_14763,N_14819);
nand U15218 (N_15218,N_14874,N_14917);
nand U15219 (N_15219,N_14973,N_14935);
and U15220 (N_15220,N_14832,N_14936);
and U15221 (N_15221,N_14864,N_14869);
nor U15222 (N_15222,N_14833,N_14901);
or U15223 (N_15223,N_14814,N_14922);
or U15224 (N_15224,N_14919,N_14774);
or U15225 (N_15225,N_14798,N_14924);
xnor U15226 (N_15226,N_14759,N_14949);
and U15227 (N_15227,N_14990,N_14908);
nor U15228 (N_15228,N_14951,N_14773);
nand U15229 (N_15229,N_14778,N_14895);
nor U15230 (N_15230,N_14768,N_14814);
and U15231 (N_15231,N_14926,N_14798);
nor U15232 (N_15232,N_14917,N_14859);
or U15233 (N_15233,N_14937,N_14819);
nor U15234 (N_15234,N_14806,N_14870);
or U15235 (N_15235,N_14949,N_14882);
xnor U15236 (N_15236,N_14891,N_14750);
xor U15237 (N_15237,N_14974,N_14758);
or U15238 (N_15238,N_14794,N_14900);
xor U15239 (N_15239,N_14810,N_14871);
xor U15240 (N_15240,N_14755,N_14835);
or U15241 (N_15241,N_14825,N_14984);
nand U15242 (N_15242,N_14909,N_14872);
and U15243 (N_15243,N_14909,N_14822);
xor U15244 (N_15244,N_14797,N_14898);
nand U15245 (N_15245,N_14754,N_14935);
nor U15246 (N_15246,N_14924,N_14955);
xor U15247 (N_15247,N_14938,N_14832);
nand U15248 (N_15248,N_14994,N_14879);
and U15249 (N_15249,N_14879,N_14974);
xor U15250 (N_15250,N_15012,N_15249);
and U15251 (N_15251,N_15127,N_15182);
and U15252 (N_15252,N_15117,N_15145);
and U15253 (N_15253,N_15185,N_15139);
nand U15254 (N_15254,N_15025,N_15032);
and U15255 (N_15255,N_15248,N_15015);
or U15256 (N_15256,N_15237,N_15113);
or U15257 (N_15257,N_15246,N_15130);
or U15258 (N_15258,N_15043,N_15162);
nor U15259 (N_15259,N_15207,N_15171);
xor U15260 (N_15260,N_15047,N_15026);
nor U15261 (N_15261,N_15081,N_15222);
or U15262 (N_15262,N_15054,N_15191);
nor U15263 (N_15263,N_15247,N_15209);
and U15264 (N_15264,N_15101,N_15074);
nor U15265 (N_15265,N_15060,N_15124);
nand U15266 (N_15266,N_15045,N_15106);
nand U15267 (N_15267,N_15133,N_15046);
xor U15268 (N_15268,N_15038,N_15179);
nand U15269 (N_15269,N_15213,N_15175);
nand U15270 (N_15270,N_15143,N_15097);
and U15271 (N_15271,N_15192,N_15149);
nor U15272 (N_15272,N_15009,N_15227);
xnor U15273 (N_15273,N_15157,N_15165);
and U15274 (N_15274,N_15064,N_15123);
nor U15275 (N_15275,N_15159,N_15177);
and U15276 (N_15276,N_15108,N_15180);
or U15277 (N_15277,N_15083,N_15104);
nand U15278 (N_15278,N_15006,N_15041);
nand U15279 (N_15279,N_15232,N_15034);
and U15280 (N_15280,N_15228,N_15114);
xnor U15281 (N_15281,N_15073,N_15153);
nor U15282 (N_15282,N_15111,N_15118);
nor U15283 (N_15283,N_15071,N_15212);
and U15284 (N_15284,N_15161,N_15224);
and U15285 (N_15285,N_15067,N_15220);
and U15286 (N_15286,N_15103,N_15058);
nand U15287 (N_15287,N_15151,N_15094);
or U15288 (N_15288,N_15022,N_15203);
nand U15289 (N_15289,N_15154,N_15193);
nand U15290 (N_15290,N_15146,N_15137);
or U15291 (N_15291,N_15214,N_15100);
and U15292 (N_15292,N_15005,N_15126);
nand U15293 (N_15293,N_15017,N_15090);
nand U15294 (N_15294,N_15062,N_15226);
nor U15295 (N_15295,N_15234,N_15188);
or U15296 (N_15296,N_15070,N_15129);
nand U15297 (N_15297,N_15167,N_15229);
and U15298 (N_15298,N_15132,N_15093);
nand U15299 (N_15299,N_15077,N_15150);
nor U15300 (N_15300,N_15055,N_15076);
nor U15301 (N_15301,N_15197,N_15206);
xor U15302 (N_15302,N_15105,N_15186);
and U15303 (N_15303,N_15011,N_15138);
or U15304 (N_15304,N_15059,N_15181);
xnor U15305 (N_15305,N_15082,N_15172);
xnor U15306 (N_15306,N_15160,N_15163);
xor U15307 (N_15307,N_15152,N_15243);
nor U15308 (N_15308,N_15115,N_15035);
nand U15309 (N_15309,N_15078,N_15141);
and U15310 (N_15310,N_15190,N_15205);
and U15311 (N_15311,N_15166,N_15030);
nand U15312 (N_15312,N_15028,N_15116);
or U15313 (N_15313,N_15245,N_15242);
nand U15314 (N_15314,N_15052,N_15194);
and U15315 (N_15315,N_15027,N_15239);
or U15316 (N_15316,N_15004,N_15201);
nor U15317 (N_15317,N_15128,N_15072);
or U15318 (N_15318,N_15014,N_15217);
nor U15319 (N_15319,N_15087,N_15174);
xnor U15320 (N_15320,N_15208,N_15037);
xnor U15321 (N_15321,N_15241,N_15240);
or U15322 (N_15322,N_15048,N_15131);
nor U15323 (N_15323,N_15183,N_15235);
or U15324 (N_15324,N_15066,N_15039);
and U15325 (N_15325,N_15024,N_15075);
nor U15326 (N_15326,N_15135,N_15122);
and U15327 (N_15327,N_15091,N_15088);
xor U15328 (N_15328,N_15056,N_15063);
and U15329 (N_15329,N_15069,N_15156);
and U15330 (N_15330,N_15000,N_15218);
or U15331 (N_15331,N_15102,N_15168);
nand U15332 (N_15332,N_15142,N_15230);
and U15333 (N_15333,N_15008,N_15086);
or U15334 (N_15334,N_15215,N_15095);
and U15335 (N_15335,N_15136,N_15120);
and U15336 (N_15336,N_15158,N_15169);
nand U15337 (N_15337,N_15178,N_15110);
and U15338 (N_15338,N_15164,N_15018);
xnor U15339 (N_15339,N_15098,N_15170);
or U15340 (N_15340,N_15099,N_15199);
xnor U15341 (N_15341,N_15040,N_15001);
or U15342 (N_15342,N_15079,N_15148);
nand U15343 (N_15343,N_15019,N_15084);
nand U15344 (N_15344,N_15033,N_15121);
nand U15345 (N_15345,N_15211,N_15036);
or U15346 (N_15346,N_15031,N_15176);
nor U15347 (N_15347,N_15013,N_15210);
nor U15348 (N_15348,N_15080,N_15003);
and U15349 (N_15349,N_15042,N_15049);
and U15350 (N_15350,N_15196,N_15219);
nand U15351 (N_15351,N_15023,N_15198);
xnor U15352 (N_15352,N_15119,N_15200);
and U15353 (N_15353,N_15053,N_15134);
nand U15354 (N_15354,N_15225,N_15010);
xor U15355 (N_15355,N_15244,N_15184);
nor U15356 (N_15356,N_15107,N_15187);
nand U15357 (N_15357,N_15125,N_15021);
nor U15358 (N_15358,N_15089,N_15007);
nand U15359 (N_15359,N_15231,N_15050);
or U15360 (N_15360,N_15112,N_15155);
xor U15361 (N_15361,N_15109,N_15144);
or U15362 (N_15362,N_15236,N_15065);
and U15363 (N_15363,N_15140,N_15068);
or U15364 (N_15364,N_15233,N_15223);
and U15365 (N_15365,N_15195,N_15051);
xor U15366 (N_15366,N_15238,N_15204);
nor U15367 (N_15367,N_15189,N_15057);
and U15368 (N_15368,N_15173,N_15016);
or U15369 (N_15369,N_15061,N_15020);
and U15370 (N_15370,N_15096,N_15216);
and U15371 (N_15371,N_15044,N_15221);
nand U15372 (N_15372,N_15085,N_15147);
xnor U15373 (N_15373,N_15002,N_15092);
nand U15374 (N_15374,N_15029,N_15202);
and U15375 (N_15375,N_15135,N_15222);
or U15376 (N_15376,N_15019,N_15091);
nor U15377 (N_15377,N_15007,N_15155);
nor U15378 (N_15378,N_15050,N_15199);
xnor U15379 (N_15379,N_15035,N_15211);
nor U15380 (N_15380,N_15128,N_15190);
nand U15381 (N_15381,N_15060,N_15187);
nor U15382 (N_15382,N_15183,N_15238);
or U15383 (N_15383,N_15062,N_15134);
or U15384 (N_15384,N_15096,N_15211);
xor U15385 (N_15385,N_15061,N_15052);
xor U15386 (N_15386,N_15082,N_15171);
and U15387 (N_15387,N_15107,N_15164);
nor U15388 (N_15388,N_15229,N_15099);
or U15389 (N_15389,N_15023,N_15087);
nor U15390 (N_15390,N_15071,N_15222);
or U15391 (N_15391,N_15033,N_15097);
or U15392 (N_15392,N_15207,N_15133);
and U15393 (N_15393,N_15157,N_15131);
or U15394 (N_15394,N_15092,N_15247);
nand U15395 (N_15395,N_15157,N_15096);
or U15396 (N_15396,N_15049,N_15036);
xnor U15397 (N_15397,N_15240,N_15150);
or U15398 (N_15398,N_15158,N_15243);
xnor U15399 (N_15399,N_15182,N_15016);
nand U15400 (N_15400,N_15240,N_15077);
nand U15401 (N_15401,N_15227,N_15044);
and U15402 (N_15402,N_15122,N_15034);
and U15403 (N_15403,N_15104,N_15008);
nor U15404 (N_15404,N_15164,N_15083);
xor U15405 (N_15405,N_15220,N_15159);
xnor U15406 (N_15406,N_15170,N_15214);
nand U15407 (N_15407,N_15200,N_15197);
xor U15408 (N_15408,N_15094,N_15225);
nand U15409 (N_15409,N_15037,N_15153);
nand U15410 (N_15410,N_15022,N_15021);
nor U15411 (N_15411,N_15115,N_15217);
and U15412 (N_15412,N_15201,N_15168);
or U15413 (N_15413,N_15213,N_15177);
or U15414 (N_15414,N_15248,N_15247);
and U15415 (N_15415,N_15174,N_15129);
nor U15416 (N_15416,N_15106,N_15004);
nand U15417 (N_15417,N_15087,N_15086);
nor U15418 (N_15418,N_15186,N_15178);
nor U15419 (N_15419,N_15094,N_15121);
and U15420 (N_15420,N_15239,N_15124);
nand U15421 (N_15421,N_15142,N_15014);
xnor U15422 (N_15422,N_15136,N_15034);
or U15423 (N_15423,N_15076,N_15002);
xnor U15424 (N_15424,N_15098,N_15088);
and U15425 (N_15425,N_15031,N_15023);
nor U15426 (N_15426,N_15053,N_15086);
and U15427 (N_15427,N_15094,N_15192);
nor U15428 (N_15428,N_15042,N_15224);
nand U15429 (N_15429,N_15065,N_15240);
nor U15430 (N_15430,N_15169,N_15171);
nor U15431 (N_15431,N_15093,N_15224);
nor U15432 (N_15432,N_15046,N_15111);
or U15433 (N_15433,N_15182,N_15062);
xor U15434 (N_15434,N_15199,N_15159);
xor U15435 (N_15435,N_15174,N_15132);
nand U15436 (N_15436,N_15006,N_15126);
xnor U15437 (N_15437,N_15063,N_15211);
nor U15438 (N_15438,N_15096,N_15148);
xor U15439 (N_15439,N_15176,N_15018);
xor U15440 (N_15440,N_15198,N_15213);
xor U15441 (N_15441,N_15063,N_15246);
nor U15442 (N_15442,N_15190,N_15246);
nor U15443 (N_15443,N_15090,N_15114);
or U15444 (N_15444,N_15071,N_15192);
nand U15445 (N_15445,N_15052,N_15015);
nor U15446 (N_15446,N_15043,N_15178);
or U15447 (N_15447,N_15240,N_15101);
or U15448 (N_15448,N_15122,N_15143);
nor U15449 (N_15449,N_15067,N_15221);
nor U15450 (N_15450,N_15011,N_15071);
nand U15451 (N_15451,N_15015,N_15120);
nor U15452 (N_15452,N_15104,N_15043);
and U15453 (N_15453,N_15247,N_15005);
nand U15454 (N_15454,N_15086,N_15236);
xnor U15455 (N_15455,N_15033,N_15003);
nor U15456 (N_15456,N_15174,N_15007);
xnor U15457 (N_15457,N_15222,N_15066);
xnor U15458 (N_15458,N_15123,N_15096);
and U15459 (N_15459,N_15190,N_15009);
nand U15460 (N_15460,N_15242,N_15147);
nand U15461 (N_15461,N_15048,N_15036);
or U15462 (N_15462,N_15204,N_15031);
or U15463 (N_15463,N_15087,N_15191);
nand U15464 (N_15464,N_15054,N_15192);
nand U15465 (N_15465,N_15161,N_15112);
nand U15466 (N_15466,N_15074,N_15041);
and U15467 (N_15467,N_15118,N_15242);
nor U15468 (N_15468,N_15200,N_15232);
or U15469 (N_15469,N_15170,N_15103);
and U15470 (N_15470,N_15236,N_15100);
nor U15471 (N_15471,N_15074,N_15131);
and U15472 (N_15472,N_15021,N_15173);
and U15473 (N_15473,N_15191,N_15062);
or U15474 (N_15474,N_15066,N_15048);
nor U15475 (N_15475,N_15215,N_15146);
or U15476 (N_15476,N_15039,N_15172);
nor U15477 (N_15477,N_15109,N_15054);
nand U15478 (N_15478,N_15030,N_15242);
xor U15479 (N_15479,N_15074,N_15077);
xnor U15480 (N_15480,N_15155,N_15160);
or U15481 (N_15481,N_15234,N_15009);
nor U15482 (N_15482,N_15035,N_15159);
nand U15483 (N_15483,N_15080,N_15106);
nand U15484 (N_15484,N_15176,N_15024);
xnor U15485 (N_15485,N_15097,N_15166);
and U15486 (N_15486,N_15198,N_15197);
nor U15487 (N_15487,N_15129,N_15100);
nand U15488 (N_15488,N_15121,N_15084);
and U15489 (N_15489,N_15161,N_15071);
or U15490 (N_15490,N_15242,N_15125);
or U15491 (N_15491,N_15230,N_15059);
and U15492 (N_15492,N_15231,N_15214);
or U15493 (N_15493,N_15231,N_15194);
and U15494 (N_15494,N_15121,N_15038);
or U15495 (N_15495,N_15100,N_15037);
nand U15496 (N_15496,N_15045,N_15059);
nor U15497 (N_15497,N_15031,N_15051);
or U15498 (N_15498,N_15204,N_15077);
nor U15499 (N_15499,N_15052,N_15019);
or U15500 (N_15500,N_15359,N_15332);
or U15501 (N_15501,N_15350,N_15499);
or U15502 (N_15502,N_15284,N_15456);
xnor U15503 (N_15503,N_15321,N_15319);
xnor U15504 (N_15504,N_15264,N_15452);
and U15505 (N_15505,N_15370,N_15460);
nor U15506 (N_15506,N_15300,N_15334);
and U15507 (N_15507,N_15304,N_15291);
xnor U15508 (N_15508,N_15400,N_15262);
or U15509 (N_15509,N_15480,N_15384);
nor U15510 (N_15510,N_15437,N_15335);
and U15511 (N_15511,N_15316,N_15453);
nand U15512 (N_15512,N_15323,N_15357);
xor U15513 (N_15513,N_15446,N_15318);
or U15514 (N_15514,N_15467,N_15375);
or U15515 (N_15515,N_15411,N_15317);
xor U15516 (N_15516,N_15348,N_15362);
nor U15517 (N_15517,N_15256,N_15269);
nor U15518 (N_15518,N_15489,N_15346);
xnor U15519 (N_15519,N_15422,N_15325);
nor U15520 (N_15520,N_15443,N_15353);
or U15521 (N_15521,N_15483,N_15406);
xnor U15522 (N_15522,N_15268,N_15468);
xor U15523 (N_15523,N_15305,N_15409);
and U15524 (N_15524,N_15371,N_15293);
xor U15525 (N_15525,N_15486,N_15484);
nor U15526 (N_15526,N_15430,N_15276);
xnor U15527 (N_15527,N_15466,N_15498);
nor U15528 (N_15528,N_15395,N_15327);
or U15529 (N_15529,N_15296,N_15455);
nor U15530 (N_15530,N_15336,N_15420);
nor U15531 (N_15531,N_15394,N_15331);
or U15532 (N_15532,N_15355,N_15366);
and U15533 (N_15533,N_15282,N_15341);
or U15534 (N_15534,N_15476,N_15491);
xor U15535 (N_15535,N_15265,N_15495);
or U15536 (N_15536,N_15263,N_15429);
and U15537 (N_15537,N_15290,N_15352);
xor U15538 (N_15538,N_15413,N_15478);
nand U15539 (N_15539,N_15472,N_15497);
nor U15540 (N_15540,N_15396,N_15415);
or U15541 (N_15541,N_15294,N_15405);
or U15542 (N_15542,N_15458,N_15469);
or U15543 (N_15543,N_15340,N_15464);
or U15544 (N_15544,N_15278,N_15434);
and U15545 (N_15545,N_15351,N_15475);
nor U15546 (N_15546,N_15463,N_15380);
and U15547 (N_15547,N_15250,N_15283);
nor U15548 (N_15548,N_15465,N_15315);
xnor U15549 (N_15549,N_15295,N_15461);
nand U15550 (N_15550,N_15379,N_15492);
xnor U15551 (N_15551,N_15416,N_15337);
nand U15552 (N_15552,N_15436,N_15324);
xor U15553 (N_15553,N_15385,N_15426);
and U15554 (N_15554,N_15378,N_15273);
xnor U15555 (N_15555,N_15299,N_15462);
nor U15556 (N_15556,N_15428,N_15459);
nand U15557 (N_15557,N_15392,N_15349);
or U15558 (N_15558,N_15358,N_15306);
nand U15559 (N_15559,N_15354,N_15435);
nand U15560 (N_15560,N_15487,N_15389);
nand U15561 (N_15561,N_15281,N_15425);
and U15562 (N_15562,N_15345,N_15479);
nor U15563 (N_15563,N_15447,N_15441);
nand U15564 (N_15564,N_15387,N_15253);
nor U15565 (N_15565,N_15372,N_15407);
or U15566 (N_15566,N_15271,N_15450);
nand U15567 (N_15567,N_15454,N_15381);
nand U15568 (N_15568,N_15369,N_15342);
and U15569 (N_15569,N_15292,N_15403);
or U15570 (N_15570,N_15417,N_15485);
or U15571 (N_15571,N_15259,N_15251);
nand U15572 (N_15572,N_15307,N_15314);
nand U15573 (N_15573,N_15329,N_15393);
and U15574 (N_15574,N_15448,N_15373);
and U15575 (N_15575,N_15288,N_15286);
and U15576 (N_15576,N_15477,N_15418);
xnor U15577 (N_15577,N_15280,N_15449);
nand U15578 (N_15578,N_15360,N_15297);
or U15579 (N_15579,N_15279,N_15421);
and U15580 (N_15580,N_15488,N_15356);
xnor U15581 (N_15581,N_15258,N_15410);
or U15582 (N_15582,N_15438,N_15302);
nand U15583 (N_15583,N_15408,N_15433);
nor U15584 (N_15584,N_15289,N_15427);
xnor U15585 (N_15585,N_15255,N_15494);
and U15586 (N_15586,N_15338,N_15303);
xor U15587 (N_15587,N_15326,N_15308);
xnor U15588 (N_15588,N_15339,N_15386);
and U15589 (N_15589,N_15344,N_15301);
and U15590 (N_15590,N_15481,N_15287);
nor U15591 (N_15591,N_15388,N_15272);
nor U15592 (N_15592,N_15254,N_15270);
xnor U15593 (N_15593,N_15424,N_15374);
nor U15594 (N_15594,N_15414,N_15298);
nand U15595 (N_15595,N_15382,N_15363);
or U15596 (N_15596,N_15457,N_15343);
nor U15597 (N_15597,N_15367,N_15399);
xor U15598 (N_15598,N_15368,N_15361);
xnor U15599 (N_15599,N_15470,N_15440);
nand U15600 (N_15600,N_15451,N_15412);
xor U15601 (N_15601,N_15274,N_15390);
and U15602 (N_15602,N_15383,N_15333);
xor U15603 (N_15603,N_15322,N_15397);
or U15604 (N_15604,N_15496,N_15391);
nand U15605 (N_15605,N_15261,N_15252);
and U15606 (N_15606,N_15482,N_15398);
nand U15607 (N_15607,N_15419,N_15402);
and U15608 (N_15608,N_15257,N_15275);
nand U15609 (N_15609,N_15490,N_15328);
or U15610 (N_15610,N_15442,N_15310);
xor U15611 (N_15611,N_15260,N_15376);
xor U15612 (N_15612,N_15309,N_15266);
nand U15613 (N_15613,N_15404,N_15471);
or U15614 (N_15614,N_15444,N_15445);
or U15615 (N_15615,N_15365,N_15285);
nor U15616 (N_15616,N_15320,N_15377);
nor U15617 (N_15617,N_15423,N_15267);
nand U15618 (N_15618,N_15439,N_15401);
nand U15619 (N_15619,N_15311,N_15330);
xnor U15620 (N_15620,N_15493,N_15364);
or U15621 (N_15621,N_15473,N_15474);
and U15622 (N_15622,N_15347,N_15277);
nand U15623 (N_15623,N_15432,N_15431);
and U15624 (N_15624,N_15312,N_15313);
or U15625 (N_15625,N_15379,N_15468);
and U15626 (N_15626,N_15486,N_15448);
or U15627 (N_15627,N_15498,N_15484);
nor U15628 (N_15628,N_15387,N_15426);
nor U15629 (N_15629,N_15425,N_15263);
nor U15630 (N_15630,N_15445,N_15257);
xnor U15631 (N_15631,N_15295,N_15469);
and U15632 (N_15632,N_15325,N_15307);
nor U15633 (N_15633,N_15469,N_15318);
or U15634 (N_15634,N_15260,N_15492);
nand U15635 (N_15635,N_15331,N_15490);
or U15636 (N_15636,N_15322,N_15268);
and U15637 (N_15637,N_15415,N_15434);
nor U15638 (N_15638,N_15409,N_15321);
nor U15639 (N_15639,N_15342,N_15417);
nand U15640 (N_15640,N_15448,N_15463);
or U15641 (N_15641,N_15340,N_15419);
xor U15642 (N_15642,N_15412,N_15262);
xor U15643 (N_15643,N_15260,N_15384);
nor U15644 (N_15644,N_15472,N_15487);
xor U15645 (N_15645,N_15371,N_15325);
nand U15646 (N_15646,N_15259,N_15304);
nand U15647 (N_15647,N_15452,N_15323);
xor U15648 (N_15648,N_15272,N_15351);
and U15649 (N_15649,N_15369,N_15312);
and U15650 (N_15650,N_15496,N_15330);
nor U15651 (N_15651,N_15316,N_15262);
xor U15652 (N_15652,N_15319,N_15415);
and U15653 (N_15653,N_15343,N_15427);
nand U15654 (N_15654,N_15350,N_15496);
or U15655 (N_15655,N_15314,N_15408);
nor U15656 (N_15656,N_15395,N_15392);
nand U15657 (N_15657,N_15352,N_15423);
nand U15658 (N_15658,N_15325,N_15337);
nor U15659 (N_15659,N_15287,N_15445);
xnor U15660 (N_15660,N_15309,N_15375);
xnor U15661 (N_15661,N_15379,N_15334);
and U15662 (N_15662,N_15457,N_15297);
and U15663 (N_15663,N_15471,N_15427);
xnor U15664 (N_15664,N_15310,N_15264);
and U15665 (N_15665,N_15438,N_15259);
nand U15666 (N_15666,N_15432,N_15315);
or U15667 (N_15667,N_15485,N_15398);
and U15668 (N_15668,N_15384,N_15308);
or U15669 (N_15669,N_15371,N_15355);
xnor U15670 (N_15670,N_15370,N_15432);
xnor U15671 (N_15671,N_15254,N_15428);
nand U15672 (N_15672,N_15324,N_15355);
nor U15673 (N_15673,N_15382,N_15467);
and U15674 (N_15674,N_15496,N_15403);
and U15675 (N_15675,N_15449,N_15498);
and U15676 (N_15676,N_15411,N_15415);
or U15677 (N_15677,N_15478,N_15463);
xor U15678 (N_15678,N_15477,N_15254);
nor U15679 (N_15679,N_15290,N_15415);
or U15680 (N_15680,N_15379,N_15316);
nand U15681 (N_15681,N_15307,N_15359);
nor U15682 (N_15682,N_15391,N_15287);
nor U15683 (N_15683,N_15448,N_15262);
or U15684 (N_15684,N_15329,N_15352);
and U15685 (N_15685,N_15370,N_15409);
nand U15686 (N_15686,N_15295,N_15471);
xnor U15687 (N_15687,N_15332,N_15467);
nand U15688 (N_15688,N_15476,N_15432);
or U15689 (N_15689,N_15387,N_15341);
xnor U15690 (N_15690,N_15331,N_15368);
nor U15691 (N_15691,N_15340,N_15428);
or U15692 (N_15692,N_15379,N_15272);
nor U15693 (N_15693,N_15349,N_15324);
nand U15694 (N_15694,N_15282,N_15366);
or U15695 (N_15695,N_15252,N_15306);
or U15696 (N_15696,N_15382,N_15417);
or U15697 (N_15697,N_15369,N_15490);
and U15698 (N_15698,N_15336,N_15267);
nor U15699 (N_15699,N_15311,N_15272);
xnor U15700 (N_15700,N_15473,N_15385);
and U15701 (N_15701,N_15316,N_15410);
and U15702 (N_15702,N_15392,N_15413);
nand U15703 (N_15703,N_15283,N_15303);
xor U15704 (N_15704,N_15431,N_15273);
and U15705 (N_15705,N_15388,N_15315);
nor U15706 (N_15706,N_15453,N_15279);
nand U15707 (N_15707,N_15467,N_15298);
xor U15708 (N_15708,N_15448,N_15455);
nand U15709 (N_15709,N_15334,N_15358);
xor U15710 (N_15710,N_15381,N_15385);
nand U15711 (N_15711,N_15291,N_15418);
and U15712 (N_15712,N_15280,N_15408);
or U15713 (N_15713,N_15397,N_15263);
and U15714 (N_15714,N_15276,N_15322);
nand U15715 (N_15715,N_15453,N_15347);
nor U15716 (N_15716,N_15286,N_15454);
xor U15717 (N_15717,N_15436,N_15331);
xor U15718 (N_15718,N_15305,N_15387);
and U15719 (N_15719,N_15479,N_15409);
xor U15720 (N_15720,N_15377,N_15345);
and U15721 (N_15721,N_15400,N_15332);
nor U15722 (N_15722,N_15482,N_15495);
xnor U15723 (N_15723,N_15358,N_15381);
nor U15724 (N_15724,N_15258,N_15374);
nand U15725 (N_15725,N_15390,N_15462);
nor U15726 (N_15726,N_15292,N_15461);
or U15727 (N_15727,N_15268,N_15351);
nand U15728 (N_15728,N_15376,N_15332);
nand U15729 (N_15729,N_15299,N_15265);
and U15730 (N_15730,N_15368,N_15469);
and U15731 (N_15731,N_15296,N_15300);
and U15732 (N_15732,N_15347,N_15487);
xor U15733 (N_15733,N_15314,N_15351);
and U15734 (N_15734,N_15448,N_15457);
nand U15735 (N_15735,N_15374,N_15413);
xor U15736 (N_15736,N_15340,N_15321);
xor U15737 (N_15737,N_15443,N_15323);
nor U15738 (N_15738,N_15397,N_15405);
xnor U15739 (N_15739,N_15345,N_15411);
xnor U15740 (N_15740,N_15301,N_15273);
nor U15741 (N_15741,N_15268,N_15376);
xnor U15742 (N_15742,N_15341,N_15256);
xnor U15743 (N_15743,N_15318,N_15489);
nand U15744 (N_15744,N_15300,N_15454);
xnor U15745 (N_15745,N_15368,N_15453);
nor U15746 (N_15746,N_15263,N_15385);
or U15747 (N_15747,N_15446,N_15375);
nor U15748 (N_15748,N_15275,N_15461);
or U15749 (N_15749,N_15476,N_15453);
xnor U15750 (N_15750,N_15585,N_15655);
xnor U15751 (N_15751,N_15590,N_15625);
and U15752 (N_15752,N_15688,N_15607);
xor U15753 (N_15753,N_15701,N_15615);
nor U15754 (N_15754,N_15571,N_15593);
nand U15755 (N_15755,N_15641,N_15666);
nor U15756 (N_15756,N_15525,N_15669);
nor U15757 (N_15757,N_15578,N_15560);
nor U15758 (N_15758,N_15647,N_15668);
nor U15759 (N_15759,N_15680,N_15704);
or U15760 (N_15760,N_15714,N_15696);
nor U15761 (N_15761,N_15637,N_15504);
or U15762 (N_15762,N_15730,N_15558);
xor U15763 (N_15763,N_15532,N_15597);
nor U15764 (N_15764,N_15657,N_15576);
and U15765 (N_15765,N_15718,N_15731);
nor U15766 (N_15766,N_15501,N_15573);
and U15767 (N_15767,N_15632,N_15530);
xnor U15768 (N_15768,N_15724,N_15586);
nor U15769 (N_15769,N_15568,N_15639);
nand U15770 (N_15770,N_15687,N_15741);
and U15771 (N_15771,N_15613,N_15522);
nand U15772 (N_15772,N_15507,N_15596);
and U15773 (N_15773,N_15683,N_15664);
and U15774 (N_15774,N_15643,N_15513);
xnor U15775 (N_15775,N_15635,N_15689);
or U15776 (N_15776,N_15588,N_15660);
nand U15777 (N_15777,N_15654,N_15648);
nand U15778 (N_15778,N_15534,N_15744);
nand U15779 (N_15779,N_15739,N_15667);
and U15780 (N_15780,N_15567,N_15601);
or U15781 (N_15781,N_15652,N_15684);
or U15782 (N_15782,N_15545,N_15617);
nor U15783 (N_15783,N_15562,N_15519);
nor U15784 (N_15784,N_15506,N_15662);
or U15785 (N_15785,N_15604,N_15626);
or U15786 (N_15786,N_15670,N_15642);
and U15787 (N_15787,N_15727,N_15712);
xnor U15788 (N_15788,N_15638,N_15692);
xor U15789 (N_15789,N_15538,N_15653);
xnor U15790 (N_15790,N_15598,N_15691);
or U15791 (N_15791,N_15537,N_15551);
xor U15792 (N_15792,N_15546,N_15556);
xor U15793 (N_15793,N_15610,N_15690);
and U15794 (N_15794,N_15745,N_15516);
nor U15795 (N_15795,N_15528,N_15600);
and U15796 (N_15796,N_15678,N_15659);
nor U15797 (N_15797,N_15603,N_15665);
or U15798 (N_15798,N_15550,N_15624);
or U15799 (N_15799,N_15748,N_15552);
and U15800 (N_15800,N_15663,N_15723);
xnor U15801 (N_15801,N_15716,N_15502);
or U15802 (N_15802,N_15592,N_15735);
nor U15803 (N_15803,N_15612,N_15577);
nand U15804 (N_15804,N_15671,N_15557);
xnor U15805 (N_15805,N_15651,N_15728);
nand U15806 (N_15806,N_15589,N_15656);
or U15807 (N_15807,N_15531,N_15503);
nand U15808 (N_15808,N_15703,N_15646);
nor U15809 (N_15809,N_15661,N_15611);
or U15810 (N_15810,N_15594,N_15549);
xor U15811 (N_15811,N_15584,N_15742);
or U15812 (N_15812,N_15500,N_15720);
nand U15813 (N_15813,N_15693,N_15709);
and U15814 (N_15814,N_15582,N_15587);
and U15815 (N_15815,N_15633,N_15583);
nor U15816 (N_15816,N_15599,N_15512);
and U15817 (N_15817,N_15737,N_15614);
or U15818 (N_15818,N_15514,N_15574);
nor U15819 (N_15819,N_15677,N_15565);
nand U15820 (N_15820,N_15675,N_15685);
nand U15821 (N_15821,N_15559,N_15564);
nor U15822 (N_15822,N_15510,N_15616);
nand U15823 (N_15823,N_15535,N_15618);
nand U15824 (N_15824,N_15619,N_15605);
xnor U15825 (N_15825,N_15561,N_15520);
xnor U15826 (N_15826,N_15695,N_15711);
xnor U15827 (N_15827,N_15547,N_15729);
xor U15828 (N_15828,N_15623,N_15509);
or U15829 (N_15829,N_15524,N_15697);
or U15830 (N_15830,N_15553,N_15569);
or U15831 (N_15831,N_15521,N_15517);
and U15832 (N_15832,N_15621,N_15533);
xnor U15833 (N_15833,N_15539,N_15628);
and U15834 (N_15834,N_15640,N_15694);
and U15835 (N_15835,N_15726,N_15740);
nor U15836 (N_15836,N_15518,N_15725);
nand U15837 (N_15837,N_15644,N_15548);
xnor U15838 (N_15838,N_15555,N_15515);
or U15839 (N_15839,N_15679,N_15676);
xnor U15840 (N_15840,N_15710,N_15708);
nor U15841 (N_15841,N_15591,N_15734);
or U15842 (N_15842,N_15511,N_15747);
nor U15843 (N_15843,N_15722,N_15536);
or U15844 (N_15844,N_15681,N_15749);
xnor U15845 (N_15845,N_15658,N_15672);
nand U15846 (N_15846,N_15527,N_15575);
and U15847 (N_15847,N_15529,N_15715);
or U15848 (N_15848,N_15622,N_15700);
xnor U15849 (N_15849,N_15609,N_15543);
xor U15850 (N_15850,N_15627,N_15631);
and U15851 (N_15851,N_15645,N_15566);
nand U15852 (N_15852,N_15738,N_15698);
xnor U15853 (N_15853,N_15629,N_15706);
or U15854 (N_15854,N_15746,N_15733);
nand U15855 (N_15855,N_15581,N_15602);
or U15856 (N_15856,N_15713,N_15699);
nor U15857 (N_15857,N_15508,N_15736);
or U15858 (N_15858,N_15719,N_15702);
nor U15859 (N_15859,N_15717,N_15544);
nor U15860 (N_15860,N_15540,N_15542);
nor U15861 (N_15861,N_15572,N_15580);
xor U15862 (N_15862,N_15732,N_15743);
nand U15863 (N_15863,N_15630,N_15674);
xnor U15864 (N_15864,N_15686,N_15636);
nor U15865 (N_15865,N_15673,N_15505);
nand U15866 (N_15866,N_15595,N_15650);
or U15867 (N_15867,N_15634,N_15649);
nor U15868 (N_15868,N_15705,N_15707);
and U15869 (N_15869,N_15554,N_15526);
or U15870 (N_15870,N_15608,N_15721);
and U15871 (N_15871,N_15579,N_15606);
xor U15872 (N_15872,N_15570,N_15620);
nand U15873 (N_15873,N_15563,N_15682);
nand U15874 (N_15874,N_15541,N_15523);
nor U15875 (N_15875,N_15722,N_15551);
nor U15876 (N_15876,N_15568,N_15535);
nand U15877 (N_15877,N_15520,N_15610);
and U15878 (N_15878,N_15630,N_15724);
nand U15879 (N_15879,N_15555,N_15737);
or U15880 (N_15880,N_15591,N_15718);
nor U15881 (N_15881,N_15708,N_15561);
or U15882 (N_15882,N_15597,N_15748);
nand U15883 (N_15883,N_15651,N_15719);
xor U15884 (N_15884,N_15604,N_15605);
xor U15885 (N_15885,N_15562,N_15641);
nand U15886 (N_15886,N_15694,N_15592);
and U15887 (N_15887,N_15721,N_15577);
nor U15888 (N_15888,N_15709,N_15716);
nand U15889 (N_15889,N_15603,N_15563);
xor U15890 (N_15890,N_15649,N_15519);
nand U15891 (N_15891,N_15677,N_15557);
or U15892 (N_15892,N_15541,N_15568);
nor U15893 (N_15893,N_15706,N_15690);
or U15894 (N_15894,N_15524,N_15703);
nand U15895 (N_15895,N_15731,N_15738);
and U15896 (N_15896,N_15523,N_15560);
nand U15897 (N_15897,N_15647,N_15582);
or U15898 (N_15898,N_15530,N_15703);
or U15899 (N_15899,N_15615,N_15644);
or U15900 (N_15900,N_15616,N_15605);
and U15901 (N_15901,N_15673,N_15550);
or U15902 (N_15902,N_15657,N_15607);
xor U15903 (N_15903,N_15649,N_15619);
nand U15904 (N_15904,N_15657,N_15623);
nor U15905 (N_15905,N_15728,N_15593);
or U15906 (N_15906,N_15625,N_15637);
nor U15907 (N_15907,N_15650,N_15718);
xor U15908 (N_15908,N_15670,N_15640);
nor U15909 (N_15909,N_15580,N_15589);
and U15910 (N_15910,N_15748,N_15585);
or U15911 (N_15911,N_15555,N_15698);
nor U15912 (N_15912,N_15511,N_15714);
and U15913 (N_15913,N_15603,N_15693);
nor U15914 (N_15914,N_15702,N_15647);
or U15915 (N_15915,N_15548,N_15623);
nor U15916 (N_15916,N_15591,N_15535);
xor U15917 (N_15917,N_15654,N_15623);
or U15918 (N_15918,N_15711,N_15510);
nor U15919 (N_15919,N_15595,N_15503);
nor U15920 (N_15920,N_15717,N_15705);
nor U15921 (N_15921,N_15532,N_15736);
xnor U15922 (N_15922,N_15685,N_15578);
or U15923 (N_15923,N_15696,N_15515);
xor U15924 (N_15924,N_15500,N_15724);
nand U15925 (N_15925,N_15551,N_15546);
xnor U15926 (N_15926,N_15541,N_15688);
or U15927 (N_15927,N_15632,N_15625);
and U15928 (N_15928,N_15666,N_15728);
or U15929 (N_15929,N_15650,N_15712);
nor U15930 (N_15930,N_15502,N_15554);
nand U15931 (N_15931,N_15722,N_15544);
nor U15932 (N_15932,N_15610,N_15543);
nand U15933 (N_15933,N_15567,N_15697);
and U15934 (N_15934,N_15506,N_15502);
nor U15935 (N_15935,N_15509,N_15578);
nor U15936 (N_15936,N_15627,N_15730);
or U15937 (N_15937,N_15583,N_15520);
xor U15938 (N_15938,N_15562,N_15728);
nand U15939 (N_15939,N_15566,N_15576);
nor U15940 (N_15940,N_15715,N_15597);
nor U15941 (N_15941,N_15501,N_15643);
or U15942 (N_15942,N_15571,N_15738);
or U15943 (N_15943,N_15736,N_15693);
nor U15944 (N_15944,N_15519,N_15574);
nand U15945 (N_15945,N_15587,N_15557);
or U15946 (N_15946,N_15743,N_15684);
xnor U15947 (N_15947,N_15665,N_15667);
and U15948 (N_15948,N_15545,N_15745);
xnor U15949 (N_15949,N_15604,N_15738);
xor U15950 (N_15950,N_15522,N_15714);
nand U15951 (N_15951,N_15684,N_15666);
xnor U15952 (N_15952,N_15686,N_15646);
nor U15953 (N_15953,N_15568,N_15738);
nor U15954 (N_15954,N_15696,N_15697);
and U15955 (N_15955,N_15602,N_15564);
nand U15956 (N_15956,N_15732,N_15740);
nor U15957 (N_15957,N_15675,N_15542);
nand U15958 (N_15958,N_15503,N_15607);
and U15959 (N_15959,N_15579,N_15566);
nor U15960 (N_15960,N_15663,N_15659);
xnor U15961 (N_15961,N_15590,N_15723);
and U15962 (N_15962,N_15705,N_15578);
nand U15963 (N_15963,N_15542,N_15635);
nor U15964 (N_15964,N_15653,N_15655);
nor U15965 (N_15965,N_15675,N_15739);
and U15966 (N_15966,N_15581,N_15585);
xnor U15967 (N_15967,N_15531,N_15645);
nor U15968 (N_15968,N_15652,N_15534);
and U15969 (N_15969,N_15666,N_15716);
or U15970 (N_15970,N_15572,N_15681);
or U15971 (N_15971,N_15611,N_15662);
nand U15972 (N_15972,N_15629,N_15605);
nand U15973 (N_15973,N_15746,N_15688);
and U15974 (N_15974,N_15520,N_15700);
or U15975 (N_15975,N_15597,N_15679);
and U15976 (N_15976,N_15641,N_15576);
and U15977 (N_15977,N_15694,N_15722);
and U15978 (N_15978,N_15540,N_15579);
xnor U15979 (N_15979,N_15668,N_15693);
or U15980 (N_15980,N_15542,N_15692);
and U15981 (N_15981,N_15720,N_15542);
xor U15982 (N_15982,N_15542,N_15547);
xor U15983 (N_15983,N_15606,N_15520);
xor U15984 (N_15984,N_15510,N_15503);
or U15985 (N_15985,N_15676,N_15619);
nand U15986 (N_15986,N_15526,N_15601);
nand U15987 (N_15987,N_15559,N_15540);
and U15988 (N_15988,N_15654,N_15659);
or U15989 (N_15989,N_15500,N_15605);
and U15990 (N_15990,N_15553,N_15719);
xnor U15991 (N_15991,N_15529,N_15587);
xnor U15992 (N_15992,N_15594,N_15633);
or U15993 (N_15993,N_15688,N_15652);
xnor U15994 (N_15994,N_15670,N_15511);
nand U15995 (N_15995,N_15660,N_15713);
nor U15996 (N_15996,N_15508,N_15634);
nor U15997 (N_15997,N_15636,N_15556);
and U15998 (N_15998,N_15508,N_15681);
nand U15999 (N_15999,N_15546,N_15666);
xor U16000 (N_16000,N_15836,N_15769);
or U16001 (N_16001,N_15838,N_15925);
nand U16002 (N_16002,N_15803,N_15942);
and U16003 (N_16003,N_15891,N_15764);
and U16004 (N_16004,N_15859,N_15938);
or U16005 (N_16005,N_15845,N_15820);
or U16006 (N_16006,N_15789,N_15914);
xor U16007 (N_16007,N_15802,N_15856);
nor U16008 (N_16008,N_15844,N_15996);
nand U16009 (N_16009,N_15954,N_15953);
nor U16010 (N_16010,N_15916,N_15899);
nand U16011 (N_16011,N_15849,N_15784);
nand U16012 (N_16012,N_15816,N_15968);
nand U16013 (N_16013,N_15887,N_15755);
nor U16014 (N_16014,N_15994,N_15972);
nand U16015 (N_16015,N_15992,N_15834);
nand U16016 (N_16016,N_15810,N_15945);
xor U16017 (N_16017,N_15852,N_15943);
xnor U16018 (N_16018,N_15800,N_15877);
and U16019 (N_16019,N_15865,N_15772);
xnor U16020 (N_16020,N_15791,N_15867);
and U16021 (N_16021,N_15964,N_15828);
nor U16022 (N_16022,N_15957,N_15840);
or U16023 (N_16023,N_15804,N_15757);
or U16024 (N_16024,N_15777,N_15995);
xnor U16025 (N_16025,N_15897,N_15818);
nand U16026 (N_16026,N_15982,N_15811);
or U16027 (N_16027,N_15876,N_15926);
xor U16028 (N_16028,N_15770,N_15986);
or U16029 (N_16029,N_15944,N_15775);
xor U16030 (N_16030,N_15767,N_15919);
nand U16031 (N_16031,N_15907,N_15998);
nand U16032 (N_16032,N_15956,N_15947);
nand U16033 (N_16033,N_15962,N_15774);
nor U16034 (N_16034,N_15835,N_15955);
or U16035 (N_16035,N_15778,N_15888);
nor U16036 (N_16036,N_15868,N_15940);
or U16037 (N_16037,N_15922,N_15960);
and U16038 (N_16038,N_15894,N_15949);
nor U16039 (N_16039,N_15977,N_15915);
nor U16040 (N_16040,N_15824,N_15924);
and U16041 (N_16041,N_15843,N_15765);
nor U16042 (N_16042,N_15776,N_15930);
nor U16043 (N_16043,N_15861,N_15939);
and U16044 (N_16044,N_15928,N_15999);
and U16045 (N_16045,N_15902,N_15857);
nor U16046 (N_16046,N_15850,N_15978);
or U16047 (N_16047,N_15893,N_15950);
nor U16048 (N_16048,N_15961,N_15909);
nor U16049 (N_16049,N_15819,N_15799);
or U16050 (N_16050,N_15766,N_15837);
nor U16051 (N_16051,N_15906,N_15932);
nor U16052 (N_16052,N_15900,N_15948);
nand U16053 (N_16053,N_15763,N_15923);
or U16054 (N_16054,N_15771,N_15794);
nand U16055 (N_16055,N_15853,N_15882);
or U16056 (N_16056,N_15754,N_15815);
or U16057 (N_16057,N_15981,N_15935);
nor U16058 (N_16058,N_15991,N_15864);
nand U16059 (N_16059,N_15927,N_15896);
xor U16060 (N_16060,N_15933,N_15997);
xnor U16061 (N_16061,N_15831,N_15918);
xor U16062 (N_16062,N_15785,N_15797);
or U16063 (N_16063,N_15869,N_15990);
and U16064 (N_16064,N_15921,N_15751);
and U16065 (N_16065,N_15872,N_15885);
nand U16066 (N_16066,N_15946,N_15812);
xor U16067 (N_16067,N_15908,N_15993);
xor U16068 (N_16068,N_15912,N_15792);
or U16069 (N_16069,N_15971,N_15976);
nor U16070 (N_16070,N_15983,N_15790);
or U16071 (N_16071,N_15895,N_15760);
xor U16072 (N_16072,N_15905,N_15817);
or U16073 (N_16073,N_15959,N_15783);
or U16074 (N_16074,N_15762,N_15782);
or U16075 (N_16075,N_15805,N_15883);
nor U16076 (N_16076,N_15773,N_15854);
and U16077 (N_16077,N_15984,N_15833);
nand U16078 (N_16078,N_15911,N_15795);
xnor U16079 (N_16079,N_15750,N_15829);
or U16080 (N_16080,N_15788,N_15901);
or U16081 (N_16081,N_15987,N_15846);
nand U16082 (N_16082,N_15808,N_15858);
nor U16083 (N_16083,N_15860,N_15880);
xnor U16084 (N_16084,N_15855,N_15796);
or U16085 (N_16085,N_15752,N_15879);
xnor U16086 (N_16086,N_15871,N_15975);
and U16087 (N_16087,N_15958,N_15934);
or U16088 (N_16088,N_15969,N_15813);
nand U16089 (N_16089,N_15913,N_15874);
and U16090 (N_16090,N_15889,N_15866);
nor U16091 (N_16091,N_15941,N_15931);
nand U16092 (N_16092,N_15980,N_15839);
nor U16093 (N_16093,N_15830,N_15966);
or U16094 (N_16094,N_15758,N_15929);
nand U16095 (N_16095,N_15806,N_15862);
xor U16096 (N_16096,N_15965,N_15898);
nor U16097 (N_16097,N_15863,N_15979);
or U16098 (N_16098,N_15917,N_15779);
nor U16099 (N_16099,N_15825,N_15974);
and U16100 (N_16100,N_15793,N_15963);
or U16101 (N_16101,N_15952,N_15801);
nor U16102 (N_16102,N_15787,N_15756);
or U16103 (N_16103,N_15892,N_15851);
and U16104 (N_16104,N_15870,N_15985);
and U16105 (N_16105,N_15890,N_15951);
nor U16106 (N_16106,N_15827,N_15781);
nor U16107 (N_16107,N_15988,N_15878);
or U16108 (N_16108,N_15910,N_15920);
nand U16109 (N_16109,N_15904,N_15832);
nand U16110 (N_16110,N_15936,N_15759);
nand U16111 (N_16111,N_15847,N_15768);
nor U16112 (N_16112,N_15780,N_15886);
nor U16113 (N_16113,N_15798,N_15814);
xor U16114 (N_16114,N_15989,N_15875);
xnor U16115 (N_16115,N_15821,N_15761);
nor U16116 (N_16116,N_15967,N_15937);
xor U16117 (N_16117,N_15841,N_15823);
xnor U16118 (N_16118,N_15809,N_15753);
nor U16119 (N_16119,N_15848,N_15842);
and U16120 (N_16120,N_15970,N_15786);
nand U16121 (N_16121,N_15903,N_15973);
nand U16122 (N_16122,N_15873,N_15881);
or U16123 (N_16123,N_15826,N_15807);
or U16124 (N_16124,N_15822,N_15884);
or U16125 (N_16125,N_15805,N_15910);
nand U16126 (N_16126,N_15889,N_15781);
xnor U16127 (N_16127,N_15783,N_15875);
xnor U16128 (N_16128,N_15852,N_15901);
or U16129 (N_16129,N_15895,N_15881);
or U16130 (N_16130,N_15965,N_15766);
or U16131 (N_16131,N_15849,N_15923);
nand U16132 (N_16132,N_15928,N_15816);
nand U16133 (N_16133,N_15987,N_15924);
nor U16134 (N_16134,N_15946,N_15871);
nor U16135 (N_16135,N_15927,N_15873);
xor U16136 (N_16136,N_15958,N_15960);
and U16137 (N_16137,N_15847,N_15869);
nand U16138 (N_16138,N_15927,N_15941);
nand U16139 (N_16139,N_15838,N_15806);
and U16140 (N_16140,N_15875,N_15996);
and U16141 (N_16141,N_15948,N_15864);
xor U16142 (N_16142,N_15895,N_15775);
xor U16143 (N_16143,N_15925,N_15898);
nor U16144 (N_16144,N_15776,N_15969);
nor U16145 (N_16145,N_15811,N_15760);
or U16146 (N_16146,N_15835,N_15971);
and U16147 (N_16147,N_15991,N_15755);
or U16148 (N_16148,N_15820,N_15963);
or U16149 (N_16149,N_15756,N_15852);
nand U16150 (N_16150,N_15870,N_15843);
nand U16151 (N_16151,N_15866,N_15823);
xor U16152 (N_16152,N_15785,N_15782);
and U16153 (N_16153,N_15984,N_15780);
nand U16154 (N_16154,N_15829,N_15853);
or U16155 (N_16155,N_15980,N_15920);
xnor U16156 (N_16156,N_15866,N_15800);
nor U16157 (N_16157,N_15898,N_15918);
nor U16158 (N_16158,N_15983,N_15925);
nand U16159 (N_16159,N_15757,N_15882);
nand U16160 (N_16160,N_15793,N_15916);
nor U16161 (N_16161,N_15768,N_15842);
nand U16162 (N_16162,N_15939,N_15862);
nand U16163 (N_16163,N_15767,N_15879);
xnor U16164 (N_16164,N_15764,N_15848);
nand U16165 (N_16165,N_15786,N_15958);
or U16166 (N_16166,N_15976,N_15949);
nor U16167 (N_16167,N_15864,N_15930);
xnor U16168 (N_16168,N_15868,N_15820);
and U16169 (N_16169,N_15865,N_15992);
and U16170 (N_16170,N_15825,N_15976);
and U16171 (N_16171,N_15762,N_15792);
nand U16172 (N_16172,N_15777,N_15863);
nor U16173 (N_16173,N_15835,N_15808);
and U16174 (N_16174,N_15758,N_15975);
and U16175 (N_16175,N_15755,N_15981);
or U16176 (N_16176,N_15980,N_15998);
and U16177 (N_16177,N_15853,N_15865);
nor U16178 (N_16178,N_15889,N_15995);
xnor U16179 (N_16179,N_15896,N_15962);
and U16180 (N_16180,N_15859,N_15911);
or U16181 (N_16181,N_15815,N_15976);
or U16182 (N_16182,N_15943,N_15864);
and U16183 (N_16183,N_15957,N_15951);
xnor U16184 (N_16184,N_15839,N_15824);
and U16185 (N_16185,N_15809,N_15982);
nor U16186 (N_16186,N_15917,N_15924);
nor U16187 (N_16187,N_15958,N_15996);
nor U16188 (N_16188,N_15774,N_15879);
or U16189 (N_16189,N_15861,N_15845);
or U16190 (N_16190,N_15926,N_15936);
nand U16191 (N_16191,N_15910,N_15841);
nand U16192 (N_16192,N_15807,N_15987);
and U16193 (N_16193,N_15806,N_15849);
nand U16194 (N_16194,N_15962,N_15857);
and U16195 (N_16195,N_15920,N_15802);
nor U16196 (N_16196,N_15828,N_15877);
or U16197 (N_16197,N_15840,N_15811);
or U16198 (N_16198,N_15822,N_15942);
nor U16199 (N_16199,N_15815,N_15961);
and U16200 (N_16200,N_15792,N_15888);
or U16201 (N_16201,N_15753,N_15785);
nand U16202 (N_16202,N_15973,N_15986);
nor U16203 (N_16203,N_15926,N_15853);
xnor U16204 (N_16204,N_15937,N_15804);
or U16205 (N_16205,N_15840,N_15950);
nand U16206 (N_16206,N_15980,N_15897);
nor U16207 (N_16207,N_15942,N_15780);
or U16208 (N_16208,N_15966,N_15866);
and U16209 (N_16209,N_15941,N_15889);
xor U16210 (N_16210,N_15910,N_15821);
and U16211 (N_16211,N_15906,N_15885);
xnor U16212 (N_16212,N_15920,N_15799);
nand U16213 (N_16213,N_15873,N_15867);
and U16214 (N_16214,N_15800,N_15882);
xor U16215 (N_16215,N_15984,N_15811);
nor U16216 (N_16216,N_15804,N_15912);
nand U16217 (N_16217,N_15868,N_15983);
xnor U16218 (N_16218,N_15946,N_15844);
nand U16219 (N_16219,N_15779,N_15832);
xor U16220 (N_16220,N_15762,N_15825);
nor U16221 (N_16221,N_15910,N_15988);
and U16222 (N_16222,N_15992,N_15760);
and U16223 (N_16223,N_15962,N_15937);
xnor U16224 (N_16224,N_15933,N_15792);
and U16225 (N_16225,N_15983,N_15843);
nor U16226 (N_16226,N_15765,N_15943);
and U16227 (N_16227,N_15904,N_15789);
nor U16228 (N_16228,N_15840,N_15965);
nand U16229 (N_16229,N_15777,N_15812);
and U16230 (N_16230,N_15911,N_15907);
and U16231 (N_16231,N_15876,N_15961);
nor U16232 (N_16232,N_15893,N_15983);
nor U16233 (N_16233,N_15765,N_15857);
and U16234 (N_16234,N_15800,N_15902);
nand U16235 (N_16235,N_15753,N_15871);
xor U16236 (N_16236,N_15897,N_15899);
and U16237 (N_16237,N_15989,N_15786);
xor U16238 (N_16238,N_15785,N_15839);
nor U16239 (N_16239,N_15946,N_15802);
and U16240 (N_16240,N_15946,N_15872);
and U16241 (N_16241,N_15884,N_15892);
and U16242 (N_16242,N_15916,N_15999);
or U16243 (N_16243,N_15826,N_15871);
nand U16244 (N_16244,N_15990,N_15818);
and U16245 (N_16245,N_15969,N_15916);
and U16246 (N_16246,N_15897,N_15858);
or U16247 (N_16247,N_15928,N_15776);
nor U16248 (N_16248,N_15846,N_15790);
nand U16249 (N_16249,N_15953,N_15789);
or U16250 (N_16250,N_16242,N_16001);
xnor U16251 (N_16251,N_16206,N_16241);
or U16252 (N_16252,N_16198,N_16233);
nand U16253 (N_16253,N_16229,N_16162);
nor U16254 (N_16254,N_16091,N_16126);
or U16255 (N_16255,N_16076,N_16174);
or U16256 (N_16256,N_16215,N_16078);
and U16257 (N_16257,N_16041,N_16208);
nor U16258 (N_16258,N_16192,N_16043);
xor U16259 (N_16259,N_16203,N_16247);
xnor U16260 (N_16260,N_16142,N_16015);
or U16261 (N_16261,N_16140,N_16171);
nor U16262 (N_16262,N_16032,N_16115);
nor U16263 (N_16263,N_16202,N_16021);
xor U16264 (N_16264,N_16074,N_16098);
or U16265 (N_16265,N_16124,N_16178);
and U16266 (N_16266,N_16217,N_16114);
nor U16267 (N_16267,N_16009,N_16244);
nor U16268 (N_16268,N_16022,N_16096);
nor U16269 (N_16269,N_16038,N_16218);
and U16270 (N_16270,N_16050,N_16085);
nand U16271 (N_16271,N_16045,N_16219);
and U16272 (N_16272,N_16137,N_16092);
nor U16273 (N_16273,N_16030,N_16118);
xnor U16274 (N_16274,N_16157,N_16191);
and U16275 (N_16275,N_16061,N_16230);
or U16276 (N_16276,N_16190,N_16058);
or U16277 (N_16277,N_16000,N_16214);
and U16278 (N_16278,N_16213,N_16161);
or U16279 (N_16279,N_16158,N_16103);
nand U16280 (N_16280,N_16194,N_16236);
nor U16281 (N_16281,N_16051,N_16232);
nand U16282 (N_16282,N_16201,N_16006);
nor U16283 (N_16283,N_16133,N_16231);
nand U16284 (N_16284,N_16054,N_16227);
or U16285 (N_16285,N_16052,N_16117);
and U16286 (N_16286,N_16120,N_16189);
nor U16287 (N_16287,N_16169,N_16246);
or U16288 (N_16288,N_16093,N_16175);
nor U16289 (N_16289,N_16018,N_16135);
or U16290 (N_16290,N_16221,N_16176);
nand U16291 (N_16291,N_16020,N_16111);
xor U16292 (N_16292,N_16210,N_16173);
nor U16293 (N_16293,N_16240,N_16187);
and U16294 (N_16294,N_16183,N_16235);
xnor U16295 (N_16295,N_16237,N_16195);
xor U16296 (N_16296,N_16160,N_16087);
xor U16297 (N_16297,N_16079,N_16121);
nand U16298 (N_16298,N_16146,N_16168);
or U16299 (N_16299,N_16172,N_16025);
and U16300 (N_16300,N_16044,N_16166);
nor U16301 (N_16301,N_16127,N_16012);
xnor U16302 (N_16302,N_16077,N_16159);
xnor U16303 (N_16303,N_16019,N_16035);
nand U16304 (N_16304,N_16123,N_16097);
and U16305 (N_16305,N_16182,N_16239);
or U16306 (N_16306,N_16040,N_16071);
or U16307 (N_16307,N_16101,N_16105);
or U16308 (N_16308,N_16086,N_16132);
and U16309 (N_16309,N_16037,N_16148);
xor U16310 (N_16310,N_16197,N_16099);
nand U16311 (N_16311,N_16004,N_16023);
or U16312 (N_16312,N_16204,N_16067);
nand U16313 (N_16313,N_16149,N_16185);
nor U16314 (N_16314,N_16147,N_16131);
and U16315 (N_16315,N_16144,N_16116);
or U16316 (N_16316,N_16072,N_16179);
and U16317 (N_16317,N_16139,N_16082);
xnor U16318 (N_16318,N_16109,N_16193);
or U16319 (N_16319,N_16106,N_16164);
xnor U16320 (N_16320,N_16141,N_16170);
xnor U16321 (N_16321,N_16005,N_16152);
and U16322 (N_16322,N_16167,N_16112);
or U16323 (N_16323,N_16177,N_16129);
nand U16324 (N_16324,N_16226,N_16228);
xnor U16325 (N_16325,N_16069,N_16029);
nand U16326 (N_16326,N_16095,N_16138);
xor U16327 (N_16327,N_16184,N_16134);
and U16328 (N_16328,N_16122,N_16163);
nor U16329 (N_16329,N_16108,N_16066);
xor U16330 (N_16330,N_16199,N_16243);
nor U16331 (N_16331,N_16034,N_16211);
xnor U16332 (N_16332,N_16008,N_16102);
xnor U16333 (N_16333,N_16154,N_16107);
and U16334 (N_16334,N_16212,N_16225);
or U16335 (N_16335,N_16026,N_16049);
nand U16336 (N_16336,N_16186,N_16180);
nand U16337 (N_16337,N_16081,N_16057);
nand U16338 (N_16338,N_16031,N_16059);
and U16339 (N_16339,N_16073,N_16010);
xnor U16340 (N_16340,N_16223,N_16188);
nor U16341 (N_16341,N_16064,N_16165);
or U16342 (N_16342,N_16100,N_16039);
nor U16343 (N_16343,N_16088,N_16065);
xor U16344 (N_16344,N_16205,N_16216);
nor U16345 (N_16345,N_16011,N_16024);
nor U16346 (N_16346,N_16094,N_16153);
nand U16347 (N_16347,N_16207,N_16036);
xor U16348 (N_16348,N_16003,N_16053);
and U16349 (N_16349,N_16104,N_16042);
nand U16350 (N_16350,N_16248,N_16062);
xnor U16351 (N_16351,N_16028,N_16027);
nand U16352 (N_16352,N_16068,N_16234);
xor U16353 (N_16353,N_16016,N_16151);
or U16354 (N_16354,N_16013,N_16083);
nand U16355 (N_16355,N_16002,N_16048);
nand U16356 (N_16356,N_16063,N_16014);
or U16357 (N_16357,N_16113,N_16033);
or U16358 (N_16358,N_16130,N_16181);
nor U16359 (N_16359,N_16007,N_16220);
nor U16360 (N_16360,N_16110,N_16119);
nand U16361 (N_16361,N_16155,N_16245);
and U16362 (N_16362,N_16196,N_16143);
nor U16363 (N_16363,N_16238,N_16047);
and U16364 (N_16364,N_16055,N_16125);
and U16365 (N_16365,N_16200,N_16084);
nor U16366 (N_16366,N_16075,N_16080);
xor U16367 (N_16367,N_16089,N_16150);
or U16368 (N_16368,N_16070,N_16090);
and U16369 (N_16369,N_16249,N_16209);
nand U16370 (N_16370,N_16046,N_16224);
and U16371 (N_16371,N_16145,N_16222);
and U16372 (N_16372,N_16060,N_16056);
nand U16373 (N_16373,N_16128,N_16017);
nand U16374 (N_16374,N_16156,N_16136);
and U16375 (N_16375,N_16068,N_16056);
and U16376 (N_16376,N_16017,N_16010);
xor U16377 (N_16377,N_16116,N_16234);
or U16378 (N_16378,N_16134,N_16040);
nand U16379 (N_16379,N_16151,N_16202);
and U16380 (N_16380,N_16161,N_16193);
and U16381 (N_16381,N_16145,N_16249);
nor U16382 (N_16382,N_16210,N_16229);
xnor U16383 (N_16383,N_16074,N_16081);
nor U16384 (N_16384,N_16020,N_16162);
and U16385 (N_16385,N_16051,N_16002);
xnor U16386 (N_16386,N_16035,N_16201);
or U16387 (N_16387,N_16219,N_16050);
nor U16388 (N_16388,N_16037,N_16028);
nand U16389 (N_16389,N_16236,N_16138);
or U16390 (N_16390,N_16061,N_16004);
nand U16391 (N_16391,N_16094,N_16095);
and U16392 (N_16392,N_16229,N_16190);
or U16393 (N_16393,N_16149,N_16192);
xnor U16394 (N_16394,N_16191,N_16237);
and U16395 (N_16395,N_16173,N_16240);
nor U16396 (N_16396,N_16228,N_16121);
or U16397 (N_16397,N_16054,N_16166);
or U16398 (N_16398,N_16230,N_16034);
nand U16399 (N_16399,N_16172,N_16132);
or U16400 (N_16400,N_16086,N_16091);
xor U16401 (N_16401,N_16151,N_16225);
nor U16402 (N_16402,N_16065,N_16201);
and U16403 (N_16403,N_16234,N_16205);
nand U16404 (N_16404,N_16144,N_16041);
nand U16405 (N_16405,N_16000,N_16243);
nor U16406 (N_16406,N_16091,N_16214);
xor U16407 (N_16407,N_16214,N_16085);
and U16408 (N_16408,N_16065,N_16155);
nor U16409 (N_16409,N_16193,N_16085);
nand U16410 (N_16410,N_16077,N_16243);
nor U16411 (N_16411,N_16012,N_16052);
xnor U16412 (N_16412,N_16127,N_16154);
nand U16413 (N_16413,N_16239,N_16100);
nand U16414 (N_16414,N_16247,N_16085);
nand U16415 (N_16415,N_16205,N_16105);
or U16416 (N_16416,N_16196,N_16126);
nor U16417 (N_16417,N_16140,N_16144);
xnor U16418 (N_16418,N_16228,N_16023);
or U16419 (N_16419,N_16241,N_16091);
nand U16420 (N_16420,N_16110,N_16044);
xor U16421 (N_16421,N_16236,N_16119);
or U16422 (N_16422,N_16025,N_16088);
and U16423 (N_16423,N_16109,N_16008);
or U16424 (N_16424,N_16118,N_16188);
or U16425 (N_16425,N_16054,N_16080);
or U16426 (N_16426,N_16023,N_16093);
and U16427 (N_16427,N_16215,N_16223);
xor U16428 (N_16428,N_16032,N_16022);
or U16429 (N_16429,N_16228,N_16119);
nand U16430 (N_16430,N_16048,N_16177);
nand U16431 (N_16431,N_16162,N_16156);
and U16432 (N_16432,N_16067,N_16051);
and U16433 (N_16433,N_16013,N_16131);
nand U16434 (N_16434,N_16120,N_16069);
and U16435 (N_16435,N_16137,N_16127);
nand U16436 (N_16436,N_16164,N_16096);
or U16437 (N_16437,N_16164,N_16117);
nand U16438 (N_16438,N_16173,N_16207);
and U16439 (N_16439,N_16124,N_16007);
nand U16440 (N_16440,N_16188,N_16065);
nand U16441 (N_16441,N_16039,N_16237);
and U16442 (N_16442,N_16000,N_16015);
nand U16443 (N_16443,N_16039,N_16230);
nand U16444 (N_16444,N_16218,N_16019);
and U16445 (N_16445,N_16246,N_16206);
nand U16446 (N_16446,N_16230,N_16237);
nor U16447 (N_16447,N_16051,N_16173);
and U16448 (N_16448,N_16030,N_16076);
or U16449 (N_16449,N_16042,N_16003);
or U16450 (N_16450,N_16058,N_16096);
or U16451 (N_16451,N_16147,N_16135);
or U16452 (N_16452,N_16112,N_16063);
nand U16453 (N_16453,N_16120,N_16191);
and U16454 (N_16454,N_16068,N_16055);
nand U16455 (N_16455,N_16161,N_16040);
nor U16456 (N_16456,N_16106,N_16199);
nand U16457 (N_16457,N_16076,N_16227);
xor U16458 (N_16458,N_16049,N_16020);
nand U16459 (N_16459,N_16078,N_16101);
xor U16460 (N_16460,N_16021,N_16157);
and U16461 (N_16461,N_16059,N_16249);
nor U16462 (N_16462,N_16032,N_16090);
nor U16463 (N_16463,N_16210,N_16224);
nand U16464 (N_16464,N_16055,N_16168);
xnor U16465 (N_16465,N_16149,N_16055);
xnor U16466 (N_16466,N_16097,N_16106);
xor U16467 (N_16467,N_16045,N_16147);
nor U16468 (N_16468,N_16106,N_16151);
xnor U16469 (N_16469,N_16087,N_16086);
nor U16470 (N_16470,N_16224,N_16162);
and U16471 (N_16471,N_16084,N_16207);
xor U16472 (N_16472,N_16075,N_16172);
and U16473 (N_16473,N_16019,N_16108);
xnor U16474 (N_16474,N_16225,N_16002);
nor U16475 (N_16475,N_16065,N_16176);
and U16476 (N_16476,N_16102,N_16050);
xnor U16477 (N_16477,N_16093,N_16134);
and U16478 (N_16478,N_16128,N_16041);
and U16479 (N_16479,N_16185,N_16084);
nand U16480 (N_16480,N_16122,N_16162);
nor U16481 (N_16481,N_16092,N_16206);
and U16482 (N_16482,N_16199,N_16080);
and U16483 (N_16483,N_16240,N_16178);
or U16484 (N_16484,N_16092,N_16155);
and U16485 (N_16485,N_16103,N_16105);
and U16486 (N_16486,N_16015,N_16143);
or U16487 (N_16487,N_16026,N_16159);
or U16488 (N_16488,N_16090,N_16012);
and U16489 (N_16489,N_16151,N_16023);
nand U16490 (N_16490,N_16249,N_16056);
nor U16491 (N_16491,N_16186,N_16223);
nor U16492 (N_16492,N_16102,N_16066);
nor U16493 (N_16493,N_16208,N_16022);
and U16494 (N_16494,N_16093,N_16143);
nor U16495 (N_16495,N_16149,N_16230);
xnor U16496 (N_16496,N_16088,N_16102);
or U16497 (N_16497,N_16127,N_16074);
xor U16498 (N_16498,N_16031,N_16202);
nor U16499 (N_16499,N_16215,N_16178);
xnor U16500 (N_16500,N_16298,N_16266);
nor U16501 (N_16501,N_16405,N_16457);
and U16502 (N_16502,N_16263,N_16288);
and U16503 (N_16503,N_16350,N_16324);
and U16504 (N_16504,N_16334,N_16312);
xnor U16505 (N_16505,N_16465,N_16274);
nor U16506 (N_16506,N_16372,N_16325);
or U16507 (N_16507,N_16432,N_16481);
nor U16508 (N_16508,N_16291,N_16292);
nor U16509 (N_16509,N_16401,N_16307);
nand U16510 (N_16510,N_16458,N_16430);
or U16511 (N_16511,N_16271,N_16279);
nand U16512 (N_16512,N_16293,N_16282);
xnor U16513 (N_16513,N_16367,N_16394);
xnor U16514 (N_16514,N_16355,N_16252);
nor U16515 (N_16515,N_16370,N_16384);
nor U16516 (N_16516,N_16494,N_16303);
or U16517 (N_16517,N_16328,N_16378);
xnor U16518 (N_16518,N_16289,N_16301);
or U16519 (N_16519,N_16447,N_16297);
and U16520 (N_16520,N_16414,N_16424);
nor U16521 (N_16521,N_16330,N_16471);
nor U16522 (N_16522,N_16389,N_16374);
nand U16523 (N_16523,N_16285,N_16295);
xnor U16524 (N_16524,N_16349,N_16393);
or U16525 (N_16525,N_16273,N_16290);
and U16526 (N_16526,N_16264,N_16478);
or U16527 (N_16527,N_16397,N_16251);
and U16528 (N_16528,N_16383,N_16278);
xnor U16529 (N_16529,N_16352,N_16491);
and U16530 (N_16530,N_16333,N_16423);
and U16531 (N_16531,N_16420,N_16421);
and U16532 (N_16532,N_16365,N_16310);
and U16533 (N_16533,N_16443,N_16396);
or U16534 (N_16534,N_16489,N_16428);
xor U16535 (N_16535,N_16351,N_16323);
nor U16536 (N_16536,N_16467,N_16390);
nor U16537 (N_16537,N_16487,N_16322);
xor U16538 (N_16538,N_16498,N_16475);
xor U16539 (N_16539,N_16431,N_16371);
and U16540 (N_16540,N_16402,N_16495);
and U16541 (N_16541,N_16422,N_16344);
and U16542 (N_16542,N_16456,N_16366);
and U16543 (N_16543,N_16412,N_16373);
and U16544 (N_16544,N_16296,N_16376);
nand U16545 (N_16545,N_16382,N_16259);
xor U16546 (N_16546,N_16362,N_16433);
xnor U16547 (N_16547,N_16477,N_16476);
xnor U16548 (N_16548,N_16315,N_16353);
or U16549 (N_16549,N_16473,N_16463);
and U16550 (N_16550,N_16284,N_16419);
nor U16551 (N_16551,N_16321,N_16357);
nor U16552 (N_16552,N_16260,N_16346);
and U16553 (N_16553,N_16415,N_16338);
xnor U16554 (N_16554,N_16388,N_16269);
nand U16555 (N_16555,N_16462,N_16455);
xor U16556 (N_16556,N_16257,N_16381);
or U16557 (N_16557,N_16482,N_16261);
or U16558 (N_16558,N_16272,N_16361);
nor U16559 (N_16559,N_16270,N_16375);
xnor U16560 (N_16560,N_16446,N_16453);
nor U16561 (N_16561,N_16468,N_16434);
and U16562 (N_16562,N_16395,N_16400);
nand U16563 (N_16563,N_16363,N_16277);
nor U16564 (N_16564,N_16320,N_16354);
nand U16565 (N_16565,N_16440,N_16464);
xor U16566 (N_16566,N_16398,N_16470);
nor U16567 (N_16567,N_16299,N_16496);
or U16568 (N_16568,N_16450,N_16441);
and U16569 (N_16569,N_16488,N_16302);
nand U16570 (N_16570,N_16347,N_16331);
xor U16571 (N_16571,N_16369,N_16332);
xor U16572 (N_16572,N_16360,N_16368);
and U16573 (N_16573,N_16265,N_16474);
nor U16574 (N_16574,N_16427,N_16311);
or U16575 (N_16575,N_16403,N_16317);
and U16576 (N_16576,N_16339,N_16444);
nand U16577 (N_16577,N_16436,N_16255);
and U16578 (N_16578,N_16280,N_16460);
and U16579 (N_16579,N_16267,N_16439);
nor U16580 (N_16580,N_16268,N_16314);
and U16581 (N_16581,N_16313,N_16413);
xor U16582 (N_16582,N_16254,N_16319);
or U16583 (N_16583,N_16306,N_16429);
and U16584 (N_16584,N_16286,N_16304);
xnor U16585 (N_16585,N_16341,N_16416);
and U16586 (N_16586,N_16392,N_16484);
nand U16587 (N_16587,N_16483,N_16345);
nand U16588 (N_16588,N_16276,N_16262);
nor U16589 (N_16589,N_16318,N_16448);
and U16590 (N_16590,N_16283,N_16256);
xor U16591 (N_16591,N_16380,N_16442);
nor U16592 (N_16592,N_16329,N_16445);
or U16593 (N_16593,N_16454,N_16348);
xor U16594 (N_16594,N_16472,N_16438);
xnor U16595 (N_16595,N_16449,N_16308);
xor U16596 (N_16596,N_16343,N_16406);
nand U16597 (N_16597,N_16281,N_16451);
and U16598 (N_16598,N_16409,N_16326);
xnor U16599 (N_16599,N_16335,N_16287);
nor U16600 (N_16600,N_16337,N_16387);
nor U16601 (N_16601,N_16469,N_16407);
nand U16602 (N_16602,N_16385,N_16466);
xor U16603 (N_16603,N_16316,N_16356);
and U16604 (N_16604,N_16417,N_16309);
nand U16605 (N_16605,N_16499,N_16461);
xor U16606 (N_16606,N_16391,N_16459);
and U16607 (N_16607,N_16490,N_16253);
xnor U16608 (N_16608,N_16300,N_16258);
nand U16609 (N_16609,N_16399,N_16408);
nor U16610 (N_16610,N_16437,N_16250);
nand U16611 (N_16611,N_16435,N_16294);
nor U16612 (N_16612,N_16359,N_16418);
and U16613 (N_16613,N_16275,N_16410);
nor U16614 (N_16614,N_16486,N_16305);
xnor U16615 (N_16615,N_16411,N_16492);
xor U16616 (N_16616,N_16386,N_16404);
or U16617 (N_16617,N_16425,N_16426);
xor U16618 (N_16618,N_16379,N_16377);
and U16619 (N_16619,N_16340,N_16358);
xnor U16620 (N_16620,N_16327,N_16497);
or U16621 (N_16621,N_16493,N_16342);
nand U16622 (N_16622,N_16480,N_16485);
nor U16623 (N_16623,N_16452,N_16364);
nand U16624 (N_16624,N_16336,N_16479);
nand U16625 (N_16625,N_16457,N_16280);
nor U16626 (N_16626,N_16369,N_16251);
or U16627 (N_16627,N_16490,N_16365);
and U16628 (N_16628,N_16256,N_16438);
and U16629 (N_16629,N_16330,N_16482);
nor U16630 (N_16630,N_16324,N_16412);
nor U16631 (N_16631,N_16339,N_16273);
nand U16632 (N_16632,N_16423,N_16297);
nand U16633 (N_16633,N_16251,N_16424);
nand U16634 (N_16634,N_16369,N_16383);
or U16635 (N_16635,N_16489,N_16321);
xor U16636 (N_16636,N_16422,N_16283);
and U16637 (N_16637,N_16308,N_16258);
nor U16638 (N_16638,N_16356,N_16265);
or U16639 (N_16639,N_16495,N_16420);
or U16640 (N_16640,N_16392,N_16265);
and U16641 (N_16641,N_16430,N_16361);
nand U16642 (N_16642,N_16257,N_16253);
or U16643 (N_16643,N_16345,N_16289);
or U16644 (N_16644,N_16252,N_16330);
nor U16645 (N_16645,N_16331,N_16475);
nand U16646 (N_16646,N_16463,N_16271);
and U16647 (N_16647,N_16255,N_16299);
xnor U16648 (N_16648,N_16470,N_16267);
and U16649 (N_16649,N_16315,N_16478);
nand U16650 (N_16650,N_16457,N_16364);
nor U16651 (N_16651,N_16401,N_16377);
nand U16652 (N_16652,N_16385,N_16263);
xnor U16653 (N_16653,N_16421,N_16337);
and U16654 (N_16654,N_16406,N_16309);
xor U16655 (N_16655,N_16338,N_16263);
nor U16656 (N_16656,N_16325,N_16337);
and U16657 (N_16657,N_16476,N_16399);
xor U16658 (N_16658,N_16343,N_16394);
or U16659 (N_16659,N_16479,N_16397);
or U16660 (N_16660,N_16341,N_16397);
nor U16661 (N_16661,N_16370,N_16265);
xnor U16662 (N_16662,N_16452,N_16422);
nand U16663 (N_16663,N_16304,N_16300);
or U16664 (N_16664,N_16360,N_16398);
nand U16665 (N_16665,N_16388,N_16275);
or U16666 (N_16666,N_16397,N_16286);
or U16667 (N_16667,N_16261,N_16445);
nor U16668 (N_16668,N_16329,N_16308);
and U16669 (N_16669,N_16447,N_16299);
nor U16670 (N_16670,N_16348,N_16493);
or U16671 (N_16671,N_16392,N_16301);
nand U16672 (N_16672,N_16369,N_16365);
and U16673 (N_16673,N_16286,N_16270);
nand U16674 (N_16674,N_16442,N_16381);
or U16675 (N_16675,N_16466,N_16317);
nor U16676 (N_16676,N_16426,N_16469);
and U16677 (N_16677,N_16374,N_16410);
or U16678 (N_16678,N_16384,N_16471);
and U16679 (N_16679,N_16307,N_16433);
nor U16680 (N_16680,N_16261,N_16497);
nor U16681 (N_16681,N_16391,N_16332);
and U16682 (N_16682,N_16442,N_16397);
nor U16683 (N_16683,N_16290,N_16445);
and U16684 (N_16684,N_16268,N_16337);
or U16685 (N_16685,N_16372,N_16366);
nand U16686 (N_16686,N_16367,N_16488);
nand U16687 (N_16687,N_16269,N_16306);
xnor U16688 (N_16688,N_16321,N_16434);
and U16689 (N_16689,N_16301,N_16464);
and U16690 (N_16690,N_16347,N_16438);
xnor U16691 (N_16691,N_16264,N_16498);
or U16692 (N_16692,N_16388,N_16310);
nor U16693 (N_16693,N_16300,N_16358);
nand U16694 (N_16694,N_16387,N_16312);
nand U16695 (N_16695,N_16278,N_16326);
or U16696 (N_16696,N_16451,N_16356);
nor U16697 (N_16697,N_16296,N_16256);
nor U16698 (N_16698,N_16396,N_16366);
nand U16699 (N_16699,N_16261,N_16414);
nor U16700 (N_16700,N_16382,N_16407);
nand U16701 (N_16701,N_16326,N_16286);
xor U16702 (N_16702,N_16440,N_16394);
and U16703 (N_16703,N_16360,N_16316);
nand U16704 (N_16704,N_16421,N_16378);
nor U16705 (N_16705,N_16345,N_16260);
nor U16706 (N_16706,N_16306,N_16484);
xor U16707 (N_16707,N_16435,N_16331);
and U16708 (N_16708,N_16487,N_16352);
and U16709 (N_16709,N_16498,N_16357);
and U16710 (N_16710,N_16404,N_16251);
xor U16711 (N_16711,N_16410,N_16468);
or U16712 (N_16712,N_16469,N_16453);
xor U16713 (N_16713,N_16476,N_16376);
and U16714 (N_16714,N_16355,N_16425);
or U16715 (N_16715,N_16299,N_16335);
and U16716 (N_16716,N_16321,N_16272);
and U16717 (N_16717,N_16430,N_16465);
xnor U16718 (N_16718,N_16444,N_16356);
nand U16719 (N_16719,N_16379,N_16401);
nor U16720 (N_16720,N_16473,N_16389);
and U16721 (N_16721,N_16295,N_16447);
nor U16722 (N_16722,N_16355,N_16465);
nand U16723 (N_16723,N_16252,N_16415);
and U16724 (N_16724,N_16493,N_16401);
xnor U16725 (N_16725,N_16333,N_16336);
xnor U16726 (N_16726,N_16252,N_16387);
and U16727 (N_16727,N_16430,N_16275);
and U16728 (N_16728,N_16284,N_16278);
and U16729 (N_16729,N_16481,N_16261);
nor U16730 (N_16730,N_16394,N_16330);
nand U16731 (N_16731,N_16272,N_16426);
xnor U16732 (N_16732,N_16419,N_16359);
and U16733 (N_16733,N_16344,N_16272);
or U16734 (N_16734,N_16454,N_16272);
or U16735 (N_16735,N_16477,N_16311);
nand U16736 (N_16736,N_16469,N_16292);
nand U16737 (N_16737,N_16360,N_16362);
xnor U16738 (N_16738,N_16455,N_16400);
xor U16739 (N_16739,N_16433,N_16280);
nor U16740 (N_16740,N_16340,N_16412);
or U16741 (N_16741,N_16386,N_16356);
or U16742 (N_16742,N_16307,N_16273);
nand U16743 (N_16743,N_16470,N_16477);
nand U16744 (N_16744,N_16324,N_16428);
xnor U16745 (N_16745,N_16425,N_16266);
or U16746 (N_16746,N_16488,N_16351);
xor U16747 (N_16747,N_16297,N_16359);
and U16748 (N_16748,N_16479,N_16476);
nand U16749 (N_16749,N_16328,N_16394);
xor U16750 (N_16750,N_16577,N_16673);
and U16751 (N_16751,N_16724,N_16740);
and U16752 (N_16752,N_16638,N_16685);
nand U16753 (N_16753,N_16611,N_16737);
nor U16754 (N_16754,N_16690,N_16525);
or U16755 (N_16755,N_16701,N_16502);
or U16756 (N_16756,N_16559,N_16610);
nand U16757 (N_16757,N_16530,N_16595);
nand U16758 (N_16758,N_16676,N_16663);
and U16759 (N_16759,N_16527,N_16608);
nor U16760 (N_16760,N_16579,N_16572);
or U16761 (N_16761,N_16655,N_16639);
and U16762 (N_16762,N_16548,N_16513);
nor U16763 (N_16763,N_16561,N_16686);
or U16764 (N_16764,N_16576,N_16588);
xor U16765 (N_16765,N_16546,N_16531);
nand U16766 (N_16766,N_16568,N_16712);
nand U16767 (N_16767,N_16693,N_16619);
nor U16768 (N_16768,N_16698,N_16651);
xor U16769 (N_16769,N_16631,N_16599);
xor U16770 (N_16770,N_16671,N_16634);
nor U16771 (N_16771,N_16700,N_16627);
nand U16772 (N_16772,N_16594,N_16543);
nor U16773 (N_16773,N_16541,N_16677);
nand U16774 (N_16774,N_16665,N_16532);
nor U16775 (N_16775,N_16522,N_16739);
or U16776 (N_16776,N_16534,N_16567);
and U16777 (N_16777,N_16715,N_16720);
or U16778 (N_16778,N_16591,N_16643);
xor U16779 (N_16779,N_16584,N_16741);
and U16780 (N_16780,N_16649,N_16695);
nor U16781 (N_16781,N_16733,N_16672);
nand U16782 (N_16782,N_16536,N_16708);
xnor U16783 (N_16783,N_16633,N_16512);
nand U16784 (N_16784,N_16683,N_16607);
nor U16785 (N_16785,N_16544,N_16694);
nor U16786 (N_16786,N_16731,N_16551);
xnor U16787 (N_16787,N_16510,N_16601);
nor U16788 (N_16788,N_16636,N_16552);
and U16789 (N_16789,N_16635,N_16521);
nand U16790 (N_16790,N_16706,N_16705);
nand U16791 (N_16791,N_16605,N_16614);
nand U16792 (N_16792,N_16666,N_16507);
or U16793 (N_16793,N_16656,N_16501);
nor U16794 (N_16794,N_16660,N_16503);
nand U16795 (N_16795,N_16674,N_16585);
xnor U16796 (N_16796,N_16620,N_16689);
and U16797 (N_16797,N_16563,N_16542);
xnor U16798 (N_16798,N_16748,N_16680);
nor U16799 (N_16799,N_16696,N_16621);
and U16800 (N_16800,N_16511,N_16730);
and U16801 (N_16801,N_16648,N_16574);
nand U16802 (N_16802,N_16570,N_16734);
xor U16803 (N_16803,N_16713,N_16725);
nand U16804 (N_16804,N_16704,N_16622);
or U16805 (N_16805,N_16628,N_16571);
nor U16806 (N_16806,N_16520,N_16573);
or U16807 (N_16807,N_16617,N_16729);
xnor U16808 (N_16808,N_16644,N_16533);
and U16809 (N_16809,N_16587,N_16659);
nand U16810 (N_16810,N_16661,N_16602);
xnor U16811 (N_16811,N_16745,N_16684);
nor U16812 (N_16812,N_16717,N_16664);
or U16813 (N_16813,N_16647,N_16538);
and U16814 (N_16814,N_16514,N_16557);
xnor U16815 (N_16815,N_16699,N_16509);
nand U16816 (N_16816,N_16586,N_16735);
and U16817 (N_16817,N_16670,N_16679);
xnor U16818 (N_16818,N_16682,N_16711);
nor U16819 (N_16819,N_16598,N_16692);
nor U16820 (N_16820,N_16609,N_16709);
or U16821 (N_16821,N_16569,N_16593);
nand U16822 (N_16822,N_16504,N_16596);
xor U16823 (N_16823,N_16558,N_16668);
xnor U16824 (N_16824,N_16640,N_16600);
or U16825 (N_16825,N_16565,N_16518);
xnor U16826 (N_16826,N_16629,N_16669);
nor U16827 (N_16827,N_16560,N_16681);
xor U16828 (N_16828,N_16732,N_16582);
or U16829 (N_16829,N_16604,N_16714);
xnor U16830 (N_16830,N_16603,N_16539);
and U16831 (N_16831,N_16589,N_16500);
xnor U16832 (N_16832,N_16718,N_16526);
nor U16833 (N_16833,N_16616,N_16710);
or U16834 (N_16834,N_16675,N_16632);
nand U16835 (N_16835,N_16667,N_16624);
or U16836 (N_16836,N_16612,N_16678);
nor U16837 (N_16837,N_16652,N_16637);
nor U16838 (N_16838,N_16555,N_16550);
or U16839 (N_16839,N_16646,N_16657);
or U16840 (N_16840,N_16515,N_16688);
xor U16841 (N_16841,N_16540,N_16581);
xor U16842 (N_16842,N_16554,N_16736);
xnor U16843 (N_16843,N_16746,N_16556);
nand U16844 (N_16844,N_16642,N_16726);
and U16845 (N_16845,N_16723,N_16691);
or U16846 (N_16846,N_16564,N_16528);
and U16847 (N_16847,N_16583,N_16506);
or U16848 (N_16848,N_16562,N_16590);
or U16849 (N_16849,N_16722,N_16580);
xnor U16850 (N_16850,N_16529,N_16623);
xnor U16851 (N_16851,N_16549,N_16626);
and U16852 (N_16852,N_16728,N_16742);
nor U16853 (N_16853,N_16650,N_16592);
nor U16854 (N_16854,N_16641,N_16575);
nand U16855 (N_16855,N_16703,N_16645);
and U16856 (N_16856,N_16719,N_16505);
and U16857 (N_16857,N_16716,N_16744);
xor U16858 (N_16858,N_16508,N_16545);
nand U16859 (N_16859,N_16566,N_16630);
or U16860 (N_16860,N_16615,N_16727);
nor U16861 (N_16861,N_16658,N_16517);
nand U16862 (N_16862,N_16535,N_16707);
or U16863 (N_16863,N_16537,N_16721);
xor U16864 (N_16864,N_16653,N_16743);
xnor U16865 (N_16865,N_16702,N_16738);
or U16866 (N_16866,N_16519,N_16524);
and U16867 (N_16867,N_16597,N_16578);
nor U16868 (N_16868,N_16687,N_16516);
and U16869 (N_16869,N_16654,N_16523);
or U16870 (N_16870,N_16618,N_16613);
xor U16871 (N_16871,N_16749,N_16747);
nand U16872 (N_16872,N_16662,N_16625);
nor U16873 (N_16873,N_16606,N_16553);
nor U16874 (N_16874,N_16547,N_16697);
nor U16875 (N_16875,N_16519,N_16686);
xor U16876 (N_16876,N_16651,N_16659);
and U16877 (N_16877,N_16531,N_16704);
and U16878 (N_16878,N_16520,N_16588);
nor U16879 (N_16879,N_16619,N_16584);
nor U16880 (N_16880,N_16604,N_16517);
and U16881 (N_16881,N_16629,N_16562);
nand U16882 (N_16882,N_16563,N_16721);
or U16883 (N_16883,N_16567,N_16663);
nor U16884 (N_16884,N_16607,N_16615);
xnor U16885 (N_16885,N_16570,N_16510);
and U16886 (N_16886,N_16603,N_16740);
or U16887 (N_16887,N_16500,N_16614);
or U16888 (N_16888,N_16612,N_16692);
or U16889 (N_16889,N_16700,N_16622);
nand U16890 (N_16890,N_16582,N_16735);
nor U16891 (N_16891,N_16727,N_16656);
or U16892 (N_16892,N_16547,N_16539);
nand U16893 (N_16893,N_16640,N_16540);
and U16894 (N_16894,N_16631,N_16726);
nor U16895 (N_16895,N_16653,N_16501);
and U16896 (N_16896,N_16546,N_16532);
or U16897 (N_16897,N_16644,N_16697);
xor U16898 (N_16898,N_16726,N_16732);
or U16899 (N_16899,N_16711,N_16603);
or U16900 (N_16900,N_16647,N_16744);
or U16901 (N_16901,N_16546,N_16672);
and U16902 (N_16902,N_16552,N_16731);
and U16903 (N_16903,N_16722,N_16648);
xnor U16904 (N_16904,N_16613,N_16632);
xnor U16905 (N_16905,N_16553,N_16528);
nor U16906 (N_16906,N_16726,N_16568);
and U16907 (N_16907,N_16582,N_16686);
and U16908 (N_16908,N_16610,N_16659);
nand U16909 (N_16909,N_16644,N_16548);
and U16910 (N_16910,N_16518,N_16563);
nand U16911 (N_16911,N_16711,N_16702);
xnor U16912 (N_16912,N_16615,N_16651);
nand U16913 (N_16913,N_16545,N_16580);
and U16914 (N_16914,N_16596,N_16748);
or U16915 (N_16915,N_16681,N_16618);
and U16916 (N_16916,N_16719,N_16500);
or U16917 (N_16917,N_16654,N_16698);
nand U16918 (N_16918,N_16567,N_16560);
or U16919 (N_16919,N_16730,N_16682);
xnor U16920 (N_16920,N_16735,N_16550);
nand U16921 (N_16921,N_16701,N_16635);
nand U16922 (N_16922,N_16648,N_16678);
or U16923 (N_16923,N_16503,N_16523);
nand U16924 (N_16924,N_16701,N_16652);
and U16925 (N_16925,N_16689,N_16539);
nand U16926 (N_16926,N_16660,N_16714);
xnor U16927 (N_16927,N_16728,N_16627);
nand U16928 (N_16928,N_16667,N_16642);
nand U16929 (N_16929,N_16648,N_16716);
and U16930 (N_16930,N_16586,N_16733);
nand U16931 (N_16931,N_16547,N_16712);
xor U16932 (N_16932,N_16548,N_16545);
nor U16933 (N_16933,N_16529,N_16507);
xnor U16934 (N_16934,N_16701,N_16556);
xnor U16935 (N_16935,N_16682,N_16639);
nand U16936 (N_16936,N_16543,N_16585);
and U16937 (N_16937,N_16510,N_16524);
nor U16938 (N_16938,N_16701,N_16739);
or U16939 (N_16939,N_16695,N_16578);
xor U16940 (N_16940,N_16745,N_16748);
or U16941 (N_16941,N_16688,N_16652);
and U16942 (N_16942,N_16604,N_16702);
nor U16943 (N_16943,N_16701,N_16526);
or U16944 (N_16944,N_16553,N_16608);
nand U16945 (N_16945,N_16653,N_16537);
nand U16946 (N_16946,N_16743,N_16511);
nor U16947 (N_16947,N_16708,N_16562);
and U16948 (N_16948,N_16694,N_16645);
xor U16949 (N_16949,N_16503,N_16561);
xor U16950 (N_16950,N_16571,N_16593);
and U16951 (N_16951,N_16634,N_16642);
and U16952 (N_16952,N_16668,N_16563);
nor U16953 (N_16953,N_16676,N_16629);
or U16954 (N_16954,N_16708,N_16540);
nand U16955 (N_16955,N_16694,N_16517);
nand U16956 (N_16956,N_16748,N_16605);
nor U16957 (N_16957,N_16712,N_16535);
xor U16958 (N_16958,N_16553,N_16678);
nor U16959 (N_16959,N_16639,N_16728);
nand U16960 (N_16960,N_16656,N_16674);
nand U16961 (N_16961,N_16693,N_16616);
xor U16962 (N_16962,N_16501,N_16669);
and U16963 (N_16963,N_16689,N_16512);
and U16964 (N_16964,N_16505,N_16606);
and U16965 (N_16965,N_16575,N_16599);
or U16966 (N_16966,N_16657,N_16628);
and U16967 (N_16967,N_16736,N_16609);
xor U16968 (N_16968,N_16699,N_16701);
nand U16969 (N_16969,N_16697,N_16722);
and U16970 (N_16970,N_16534,N_16718);
nand U16971 (N_16971,N_16639,N_16717);
nor U16972 (N_16972,N_16662,N_16523);
xnor U16973 (N_16973,N_16561,N_16575);
nand U16974 (N_16974,N_16501,N_16606);
xnor U16975 (N_16975,N_16738,N_16643);
nor U16976 (N_16976,N_16601,N_16635);
nand U16977 (N_16977,N_16741,N_16567);
xnor U16978 (N_16978,N_16627,N_16726);
nand U16979 (N_16979,N_16728,N_16516);
and U16980 (N_16980,N_16569,N_16567);
nor U16981 (N_16981,N_16625,N_16530);
or U16982 (N_16982,N_16500,N_16647);
or U16983 (N_16983,N_16500,N_16554);
and U16984 (N_16984,N_16558,N_16589);
nor U16985 (N_16985,N_16630,N_16527);
or U16986 (N_16986,N_16658,N_16503);
nand U16987 (N_16987,N_16596,N_16582);
nand U16988 (N_16988,N_16708,N_16692);
xor U16989 (N_16989,N_16655,N_16702);
or U16990 (N_16990,N_16602,N_16643);
and U16991 (N_16991,N_16654,N_16623);
nor U16992 (N_16992,N_16554,N_16647);
nand U16993 (N_16993,N_16688,N_16583);
or U16994 (N_16994,N_16595,N_16560);
nor U16995 (N_16995,N_16625,N_16510);
nand U16996 (N_16996,N_16644,N_16518);
or U16997 (N_16997,N_16666,N_16709);
and U16998 (N_16998,N_16638,N_16609);
nor U16999 (N_16999,N_16727,N_16558);
or U17000 (N_17000,N_16844,N_16832);
nor U17001 (N_17001,N_16939,N_16879);
or U17002 (N_17002,N_16881,N_16859);
and U17003 (N_17003,N_16958,N_16760);
and U17004 (N_17004,N_16945,N_16792);
nand U17005 (N_17005,N_16996,N_16767);
nand U17006 (N_17006,N_16892,N_16826);
nor U17007 (N_17007,N_16759,N_16842);
nand U17008 (N_17008,N_16751,N_16815);
xor U17009 (N_17009,N_16960,N_16835);
xor U17010 (N_17010,N_16761,N_16757);
nand U17011 (N_17011,N_16912,N_16846);
nand U17012 (N_17012,N_16908,N_16750);
or U17013 (N_17013,N_16920,N_16957);
xor U17014 (N_17014,N_16976,N_16982);
xnor U17015 (N_17015,N_16768,N_16771);
and U17016 (N_17016,N_16901,N_16813);
nand U17017 (N_17017,N_16949,N_16882);
and U17018 (N_17018,N_16947,N_16865);
xnor U17019 (N_17019,N_16875,N_16852);
and U17020 (N_17020,N_16829,N_16822);
nand U17021 (N_17021,N_16955,N_16825);
nor U17022 (N_17022,N_16812,N_16790);
xor U17023 (N_17023,N_16791,N_16854);
nor U17024 (N_17024,N_16911,N_16827);
nor U17025 (N_17025,N_16872,N_16793);
nand U17026 (N_17026,N_16988,N_16797);
nor U17027 (N_17027,N_16994,N_16828);
xor U17028 (N_17028,N_16824,N_16874);
and U17029 (N_17029,N_16878,N_16926);
and U17030 (N_17030,N_16948,N_16765);
and U17031 (N_17031,N_16845,N_16801);
or U17032 (N_17032,N_16834,N_16820);
and U17033 (N_17033,N_16968,N_16795);
xor U17034 (N_17034,N_16823,N_16889);
xor U17035 (N_17035,N_16869,N_16989);
xor U17036 (N_17036,N_16794,N_16995);
xnor U17037 (N_17037,N_16928,N_16941);
or U17038 (N_17038,N_16921,N_16758);
nand U17039 (N_17039,N_16856,N_16787);
or U17040 (N_17040,N_16756,N_16800);
or U17041 (N_17041,N_16980,N_16780);
and U17042 (N_17042,N_16783,N_16764);
or U17043 (N_17043,N_16979,N_16905);
and U17044 (N_17044,N_16898,N_16867);
xor U17045 (N_17045,N_16893,N_16753);
nand U17046 (N_17046,N_16931,N_16873);
nor U17047 (N_17047,N_16883,N_16833);
nand U17048 (N_17048,N_16839,N_16909);
and U17049 (N_17049,N_16933,N_16885);
or U17050 (N_17050,N_16805,N_16809);
and U17051 (N_17051,N_16857,N_16913);
xnor U17052 (N_17052,N_16891,N_16789);
nand U17053 (N_17053,N_16977,N_16918);
xnor U17054 (N_17054,N_16944,N_16992);
or U17055 (N_17055,N_16965,N_16887);
and U17056 (N_17056,N_16915,N_16990);
and U17057 (N_17057,N_16776,N_16927);
and U17058 (N_17058,N_16935,N_16774);
or U17059 (N_17059,N_16769,N_16802);
nand U17060 (N_17060,N_16837,N_16840);
xor U17061 (N_17061,N_16855,N_16876);
and U17062 (N_17062,N_16858,N_16984);
xnor U17063 (N_17063,N_16903,N_16849);
and U17064 (N_17064,N_16808,N_16773);
and U17065 (N_17065,N_16967,N_16972);
and U17066 (N_17066,N_16902,N_16974);
or U17067 (N_17067,N_16798,N_16969);
or U17068 (N_17068,N_16810,N_16763);
nand U17069 (N_17069,N_16914,N_16803);
nor U17070 (N_17070,N_16953,N_16987);
xor U17071 (N_17071,N_16752,N_16843);
xor U17072 (N_17072,N_16954,N_16923);
nor U17073 (N_17073,N_16811,N_16777);
xnor U17074 (N_17074,N_16904,N_16806);
nor U17075 (N_17075,N_16938,N_16755);
xor U17076 (N_17076,N_16880,N_16853);
or U17077 (N_17077,N_16831,N_16838);
or U17078 (N_17078,N_16860,N_16924);
xnor U17079 (N_17079,N_16899,N_16807);
xor U17080 (N_17080,N_16985,N_16925);
nand U17081 (N_17081,N_16804,N_16999);
nor U17082 (N_17082,N_16951,N_16970);
nand U17083 (N_17083,N_16934,N_16907);
nor U17084 (N_17084,N_16784,N_16981);
or U17085 (N_17085,N_16896,N_16781);
and U17086 (N_17086,N_16952,N_16870);
and U17087 (N_17087,N_16866,N_16788);
nand U17088 (N_17088,N_16862,N_16962);
nor U17089 (N_17089,N_16785,N_16978);
and U17090 (N_17090,N_16848,N_16894);
xor U17091 (N_17091,N_16766,N_16775);
or U17092 (N_17092,N_16779,N_16910);
and U17093 (N_17093,N_16847,N_16991);
or U17094 (N_17094,N_16937,N_16917);
nor U17095 (N_17095,N_16993,N_16932);
and U17096 (N_17096,N_16818,N_16886);
nand U17097 (N_17097,N_16983,N_16772);
nor U17098 (N_17098,N_16836,N_16861);
nor U17099 (N_17099,N_16963,N_16830);
nand U17100 (N_17100,N_16816,N_16959);
xnor U17101 (N_17101,N_16762,N_16850);
or U17102 (N_17102,N_16821,N_16930);
nor U17103 (N_17103,N_16922,N_16900);
and U17104 (N_17104,N_16864,N_16956);
xnor U17105 (N_17105,N_16998,N_16778);
nor U17106 (N_17106,N_16919,N_16895);
or U17107 (N_17107,N_16966,N_16916);
and U17108 (N_17108,N_16817,N_16929);
nand U17109 (N_17109,N_16786,N_16863);
nor U17110 (N_17110,N_16971,N_16796);
xor U17111 (N_17111,N_16943,N_16782);
xnor U17112 (N_17112,N_16890,N_16819);
or U17113 (N_17113,N_16950,N_16973);
and U17114 (N_17114,N_16964,N_16814);
nand U17115 (N_17115,N_16841,N_16946);
nor U17116 (N_17116,N_16770,N_16877);
nor U17117 (N_17117,N_16986,N_16997);
nor U17118 (N_17118,N_16851,N_16897);
nand U17119 (N_17119,N_16975,N_16884);
xnor U17120 (N_17120,N_16871,N_16942);
or U17121 (N_17121,N_16906,N_16868);
or U17122 (N_17122,N_16799,N_16888);
nand U17123 (N_17123,N_16961,N_16936);
xnor U17124 (N_17124,N_16754,N_16940);
or U17125 (N_17125,N_16949,N_16865);
and U17126 (N_17126,N_16890,N_16844);
nand U17127 (N_17127,N_16986,N_16840);
or U17128 (N_17128,N_16967,N_16801);
nor U17129 (N_17129,N_16902,N_16895);
nand U17130 (N_17130,N_16913,N_16785);
xnor U17131 (N_17131,N_16808,N_16870);
or U17132 (N_17132,N_16926,N_16914);
nor U17133 (N_17133,N_16867,N_16973);
or U17134 (N_17134,N_16762,N_16933);
nor U17135 (N_17135,N_16793,N_16926);
nor U17136 (N_17136,N_16846,N_16903);
xor U17137 (N_17137,N_16952,N_16891);
or U17138 (N_17138,N_16985,N_16921);
xnor U17139 (N_17139,N_16945,N_16949);
nor U17140 (N_17140,N_16971,N_16775);
and U17141 (N_17141,N_16997,N_16926);
nand U17142 (N_17142,N_16752,N_16763);
or U17143 (N_17143,N_16845,N_16817);
or U17144 (N_17144,N_16952,N_16959);
and U17145 (N_17145,N_16757,N_16854);
xnor U17146 (N_17146,N_16933,N_16807);
and U17147 (N_17147,N_16757,N_16916);
nor U17148 (N_17148,N_16784,N_16974);
or U17149 (N_17149,N_16819,N_16939);
nor U17150 (N_17150,N_16902,N_16790);
xnor U17151 (N_17151,N_16997,N_16858);
and U17152 (N_17152,N_16848,N_16890);
xnor U17153 (N_17153,N_16926,N_16916);
nand U17154 (N_17154,N_16960,N_16924);
xnor U17155 (N_17155,N_16808,N_16816);
xor U17156 (N_17156,N_16776,N_16938);
or U17157 (N_17157,N_16930,N_16825);
nor U17158 (N_17158,N_16814,N_16855);
xor U17159 (N_17159,N_16878,N_16997);
and U17160 (N_17160,N_16805,N_16800);
or U17161 (N_17161,N_16991,N_16998);
xor U17162 (N_17162,N_16836,N_16885);
nand U17163 (N_17163,N_16972,N_16776);
and U17164 (N_17164,N_16891,N_16762);
or U17165 (N_17165,N_16947,N_16929);
nor U17166 (N_17166,N_16877,N_16935);
and U17167 (N_17167,N_16889,N_16912);
xnor U17168 (N_17168,N_16852,N_16992);
nand U17169 (N_17169,N_16972,N_16876);
nand U17170 (N_17170,N_16881,N_16929);
or U17171 (N_17171,N_16756,N_16782);
xnor U17172 (N_17172,N_16922,N_16773);
and U17173 (N_17173,N_16989,N_16752);
and U17174 (N_17174,N_16842,N_16982);
xor U17175 (N_17175,N_16848,N_16956);
or U17176 (N_17176,N_16921,N_16780);
or U17177 (N_17177,N_16794,N_16942);
or U17178 (N_17178,N_16753,N_16853);
nand U17179 (N_17179,N_16991,N_16964);
nor U17180 (N_17180,N_16887,N_16821);
nor U17181 (N_17181,N_16949,N_16775);
nand U17182 (N_17182,N_16809,N_16848);
nand U17183 (N_17183,N_16971,N_16828);
or U17184 (N_17184,N_16916,N_16953);
xnor U17185 (N_17185,N_16863,N_16774);
nand U17186 (N_17186,N_16803,N_16776);
and U17187 (N_17187,N_16997,N_16914);
or U17188 (N_17188,N_16834,N_16844);
nor U17189 (N_17189,N_16977,N_16910);
or U17190 (N_17190,N_16975,N_16890);
and U17191 (N_17191,N_16834,N_16978);
nand U17192 (N_17192,N_16942,N_16977);
xnor U17193 (N_17193,N_16839,N_16874);
or U17194 (N_17194,N_16888,N_16971);
nand U17195 (N_17195,N_16915,N_16757);
nand U17196 (N_17196,N_16854,N_16805);
or U17197 (N_17197,N_16865,N_16955);
and U17198 (N_17198,N_16968,N_16915);
nor U17199 (N_17199,N_16807,N_16843);
and U17200 (N_17200,N_16901,N_16924);
and U17201 (N_17201,N_16763,N_16889);
nor U17202 (N_17202,N_16940,N_16821);
xor U17203 (N_17203,N_16936,N_16980);
and U17204 (N_17204,N_16979,N_16958);
xnor U17205 (N_17205,N_16939,N_16993);
or U17206 (N_17206,N_16801,N_16930);
and U17207 (N_17207,N_16918,N_16808);
xnor U17208 (N_17208,N_16825,N_16821);
nor U17209 (N_17209,N_16830,N_16759);
or U17210 (N_17210,N_16970,N_16754);
nor U17211 (N_17211,N_16875,N_16925);
nor U17212 (N_17212,N_16957,N_16938);
and U17213 (N_17213,N_16817,N_16755);
or U17214 (N_17214,N_16868,N_16867);
or U17215 (N_17215,N_16884,N_16806);
nand U17216 (N_17216,N_16904,N_16977);
or U17217 (N_17217,N_16802,N_16807);
nor U17218 (N_17218,N_16910,N_16891);
and U17219 (N_17219,N_16889,N_16770);
and U17220 (N_17220,N_16764,N_16792);
xnor U17221 (N_17221,N_16909,N_16804);
and U17222 (N_17222,N_16758,N_16855);
and U17223 (N_17223,N_16847,N_16935);
nor U17224 (N_17224,N_16855,N_16928);
xnor U17225 (N_17225,N_16971,N_16890);
nor U17226 (N_17226,N_16944,N_16918);
nor U17227 (N_17227,N_16831,N_16809);
nand U17228 (N_17228,N_16879,N_16831);
nor U17229 (N_17229,N_16919,N_16929);
nand U17230 (N_17230,N_16819,N_16928);
and U17231 (N_17231,N_16825,N_16997);
nor U17232 (N_17232,N_16838,N_16808);
xnor U17233 (N_17233,N_16811,N_16913);
and U17234 (N_17234,N_16822,N_16890);
nor U17235 (N_17235,N_16908,N_16832);
nor U17236 (N_17236,N_16952,N_16936);
nor U17237 (N_17237,N_16993,N_16982);
xnor U17238 (N_17238,N_16872,N_16955);
nor U17239 (N_17239,N_16851,N_16788);
nand U17240 (N_17240,N_16786,N_16933);
xnor U17241 (N_17241,N_16752,N_16818);
xnor U17242 (N_17242,N_16904,N_16758);
nor U17243 (N_17243,N_16972,N_16808);
xor U17244 (N_17244,N_16883,N_16954);
xnor U17245 (N_17245,N_16902,N_16935);
or U17246 (N_17246,N_16763,N_16967);
and U17247 (N_17247,N_16902,N_16761);
and U17248 (N_17248,N_16982,N_16929);
nor U17249 (N_17249,N_16957,N_16780);
nor U17250 (N_17250,N_17081,N_17025);
nand U17251 (N_17251,N_17184,N_17163);
nor U17252 (N_17252,N_17073,N_17030);
nor U17253 (N_17253,N_17202,N_17118);
nor U17254 (N_17254,N_17049,N_17095);
or U17255 (N_17255,N_17080,N_17132);
and U17256 (N_17256,N_17137,N_17078);
nor U17257 (N_17257,N_17089,N_17044);
and U17258 (N_17258,N_17246,N_17210);
and U17259 (N_17259,N_17070,N_17139);
xor U17260 (N_17260,N_17020,N_17186);
and U17261 (N_17261,N_17160,N_17148);
nand U17262 (N_17262,N_17023,N_17229);
or U17263 (N_17263,N_17034,N_17093);
nand U17264 (N_17264,N_17112,N_17119);
xnor U17265 (N_17265,N_17230,N_17052);
and U17266 (N_17266,N_17159,N_17192);
and U17267 (N_17267,N_17241,N_17190);
nor U17268 (N_17268,N_17145,N_17104);
xnor U17269 (N_17269,N_17225,N_17054);
and U17270 (N_17270,N_17167,N_17214);
xor U17271 (N_17271,N_17059,N_17183);
nand U17272 (N_17272,N_17133,N_17075);
and U17273 (N_17273,N_17152,N_17015);
xnor U17274 (N_17274,N_17124,N_17117);
and U17275 (N_17275,N_17008,N_17142);
or U17276 (N_17276,N_17084,N_17082);
or U17277 (N_17277,N_17013,N_17146);
nor U17278 (N_17278,N_17106,N_17243);
xor U17279 (N_17279,N_17002,N_17024);
nand U17280 (N_17280,N_17021,N_17177);
and U17281 (N_17281,N_17079,N_17200);
nor U17282 (N_17282,N_17108,N_17061);
nor U17283 (N_17283,N_17219,N_17074);
or U17284 (N_17284,N_17140,N_17220);
xnor U17285 (N_17285,N_17068,N_17016);
xnor U17286 (N_17286,N_17009,N_17028);
nand U17287 (N_17287,N_17092,N_17236);
xnor U17288 (N_17288,N_17218,N_17062);
nand U17289 (N_17289,N_17111,N_17182);
nor U17290 (N_17290,N_17102,N_17050);
nand U17291 (N_17291,N_17097,N_17179);
and U17292 (N_17292,N_17029,N_17155);
xor U17293 (N_17293,N_17063,N_17101);
xor U17294 (N_17294,N_17131,N_17001);
and U17295 (N_17295,N_17171,N_17127);
xor U17296 (N_17296,N_17223,N_17027);
and U17297 (N_17297,N_17178,N_17085);
or U17298 (N_17298,N_17043,N_17245);
xor U17299 (N_17299,N_17208,N_17161);
nor U17300 (N_17300,N_17187,N_17135);
or U17301 (N_17301,N_17116,N_17240);
nand U17302 (N_17302,N_17077,N_17031);
nand U17303 (N_17303,N_17128,N_17017);
and U17304 (N_17304,N_17136,N_17056);
and U17305 (N_17305,N_17006,N_17189);
or U17306 (N_17306,N_17231,N_17134);
nand U17307 (N_17307,N_17126,N_17150);
xnor U17308 (N_17308,N_17238,N_17222);
nand U17309 (N_17309,N_17237,N_17055);
and U17310 (N_17310,N_17157,N_17072);
nor U17311 (N_17311,N_17109,N_17249);
and U17312 (N_17312,N_17114,N_17064);
or U17313 (N_17313,N_17065,N_17239);
or U17314 (N_17314,N_17162,N_17242);
and U17315 (N_17315,N_17156,N_17228);
and U17316 (N_17316,N_17120,N_17198);
xnor U17317 (N_17317,N_17197,N_17069);
xor U17318 (N_17318,N_17195,N_17019);
xnor U17319 (N_17319,N_17244,N_17010);
or U17320 (N_17320,N_17033,N_17129);
xor U17321 (N_17321,N_17181,N_17088);
xor U17322 (N_17322,N_17103,N_17206);
and U17323 (N_17323,N_17221,N_17005);
or U17324 (N_17324,N_17076,N_17046);
or U17325 (N_17325,N_17170,N_17234);
nor U17326 (N_17326,N_17026,N_17121);
or U17327 (N_17327,N_17012,N_17110);
nand U17328 (N_17328,N_17226,N_17174);
nor U17329 (N_17329,N_17122,N_17185);
xor U17330 (N_17330,N_17047,N_17051);
xor U17331 (N_17331,N_17175,N_17071);
nand U17332 (N_17332,N_17138,N_17213);
or U17333 (N_17333,N_17196,N_17048);
nand U17334 (N_17334,N_17060,N_17215);
xor U17335 (N_17335,N_17057,N_17173);
or U17336 (N_17336,N_17039,N_17194);
or U17337 (N_17337,N_17053,N_17172);
nor U17338 (N_17338,N_17217,N_17004);
xnor U17339 (N_17339,N_17169,N_17003);
or U17340 (N_17340,N_17168,N_17058);
or U17341 (N_17341,N_17153,N_17212);
or U17342 (N_17342,N_17066,N_17115);
nand U17343 (N_17343,N_17188,N_17227);
nand U17344 (N_17344,N_17098,N_17038);
nor U17345 (N_17345,N_17147,N_17099);
nor U17346 (N_17346,N_17040,N_17141);
and U17347 (N_17347,N_17224,N_17232);
and U17348 (N_17348,N_17000,N_17233);
or U17349 (N_17349,N_17094,N_17216);
or U17350 (N_17350,N_17247,N_17204);
nor U17351 (N_17351,N_17087,N_17107);
xor U17352 (N_17352,N_17180,N_17113);
nand U17353 (N_17353,N_17191,N_17165);
or U17354 (N_17354,N_17201,N_17164);
xnor U17355 (N_17355,N_17176,N_17144);
xor U17356 (N_17356,N_17149,N_17154);
nor U17357 (N_17357,N_17248,N_17130);
and U17358 (N_17358,N_17158,N_17090);
nand U17359 (N_17359,N_17011,N_17032);
and U17360 (N_17360,N_17203,N_17014);
nand U17361 (N_17361,N_17007,N_17091);
nor U17362 (N_17362,N_17018,N_17199);
xnor U17363 (N_17363,N_17096,N_17125);
nor U17364 (N_17364,N_17151,N_17205);
xor U17365 (N_17365,N_17209,N_17105);
or U17366 (N_17366,N_17143,N_17036);
and U17367 (N_17367,N_17235,N_17166);
xnor U17368 (N_17368,N_17211,N_17100);
nor U17369 (N_17369,N_17045,N_17193);
or U17370 (N_17370,N_17041,N_17035);
xnor U17371 (N_17371,N_17083,N_17086);
or U17372 (N_17372,N_17207,N_17022);
nand U17373 (N_17373,N_17067,N_17042);
nor U17374 (N_17374,N_17037,N_17123);
or U17375 (N_17375,N_17114,N_17003);
or U17376 (N_17376,N_17157,N_17066);
or U17377 (N_17377,N_17194,N_17245);
nand U17378 (N_17378,N_17179,N_17076);
nand U17379 (N_17379,N_17019,N_17105);
nand U17380 (N_17380,N_17108,N_17041);
or U17381 (N_17381,N_17058,N_17247);
xnor U17382 (N_17382,N_17059,N_17025);
or U17383 (N_17383,N_17244,N_17115);
nor U17384 (N_17384,N_17000,N_17139);
or U17385 (N_17385,N_17177,N_17169);
nor U17386 (N_17386,N_17078,N_17190);
xor U17387 (N_17387,N_17087,N_17098);
or U17388 (N_17388,N_17061,N_17014);
or U17389 (N_17389,N_17214,N_17194);
nor U17390 (N_17390,N_17176,N_17159);
and U17391 (N_17391,N_17002,N_17226);
or U17392 (N_17392,N_17166,N_17011);
or U17393 (N_17393,N_17157,N_17247);
nand U17394 (N_17394,N_17021,N_17061);
nor U17395 (N_17395,N_17129,N_17025);
nor U17396 (N_17396,N_17067,N_17095);
or U17397 (N_17397,N_17064,N_17000);
or U17398 (N_17398,N_17045,N_17107);
nand U17399 (N_17399,N_17174,N_17236);
nor U17400 (N_17400,N_17052,N_17098);
and U17401 (N_17401,N_17008,N_17115);
nand U17402 (N_17402,N_17129,N_17215);
xor U17403 (N_17403,N_17135,N_17224);
xnor U17404 (N_17404,N_17062,N_17089);
or U17405 (N_17405,N_17069,N_17180);
nand U17406 (N_17406,N_17121,N_17040);
or U17407 (N_17407,N_17046,N_17167);
and U17408 (N_17408,N_17113,N_17009);
and U17409 (N_17409,N_17042,N_17134);
nand U17410 (N_17410,N_17117,N_17102);
or U17411 (N_17411,N_17140,N_17006);
or U17412 (N_17412,N_17246,N_17173);
xnor U17413 (N_17413,N_17214,N_17048);
and U17414 (N_17414,N_17001,N_17017);
nand U17415 (N_17415,N_17226,N_17009);
and U17416 (N_17416,N_17054,N_17184);
or U17417 (N_17417,N_17207,N_17172);
nor U17418 (N_17418,N_17174,N_17137);
and U17419 (N_17419,N_17241,N_17214);
and U17420 (N_17420,N_17144,N_17094);
or U17421 (N_17421,N_17069,N_17220);
nand U17422 (N_17422,N_17198,N_17196);
and U17423 (N_17423,N_17175,N_17051);
xnor U17424 (N_17424,N_17070,N_17159);
nand U17425 (N_17425,N_17054,N_17062);
or U17426 (N_17426,N_17124,N_17245);
and U17427 (N_17427,N_17052,N_17082);
xnor U17428 (N_17428,N_17132,N_17185);
nor U17429 (N_17429,N_17043,N_17200);
xor U17430 (N_17430,N_17033,N_17149);
nand U17431 (N_17431,N_17098,N_17058);
xor U17432 (N_17432,N_17231,N_17114);
nand U17433 (N_17433,N_17071,N_17092);
nor U17434 (N_17434,N_17081,N_17049);
and U17435 (N_17435,N_17187,N_17023);
or U17436 (N_17436,N_17235,N_17066);
and U17437 (N_17437,N_17017,N_17036);
or U17438 (N_17438,N_17147,N_17038);
xor U17439 (N_17439,N_17193,N_17128);
or U17440 (N_17440,N_17023,N_17069);
xor U17441 (N_17441,N_17149,N_17234);
nand U17442 (N_17442,N_17110,N_17155);
nand U17443 (N_17443,N_17147,N_17049);
xor U17444 (N_17444,N_17202,N_17140);
nor U17445 (N_17445,N_17087,N_17136);
nor U17446 (N_17446,N_17049,N_17058);
xor U17447 (N_17447,N_17243,N_17103);
nand U17448 (N_17448,N_17151,N_17021);
xnor U17449 (N_17449,N_17158,N_17172);
nor U17450 (N_17450,N_17213,N_17172);
nor U17451 (N_17451,N_17225,N_17187);
or U17452 (N_17452,N_17056,N_17071);
or U17453 (N_17453,N_17212,N_17216);
xor U17454 (N_17454,N_17227,N_17070);
nand U17455 (N_17455,N_17029,N_17130);
and U17456 (N_17456,N_17123,N_17073);
and U17457 (N_17457,N_17024,N_17230);
xor U17458 (N_17458,N_17166,N_17120);
nor U17459 (N_17459,N_17094,N_17117);
nand U17460 (N_17460,N_17185,N_17079);
nand U17461 (N_17461,N_17157,N_17103);
xor U17462 (N_17462,N_17132,N_17064);
nor U17463 (N_17463,N_17231,N_17218);
nand U17464 (N_17464,N_17095,N_17174);
and U17465 (N_17465,N_17009,N_17220);
or U17466 (N_17466,N_17212,N_17237);
or U17467 (N_17467,N_17158,N_17080);
and U17468 (N_17468,N_17064,N_17204);
and U17469 (N_17469,N_17076,N_17056);
xnor U17470 (N_17470,N_17224,N_17156);
or U17471 (N_17471,N_17088,N_17075);
xor U17472 (N_17472,N_17212,N_17045);
or U17473 (N_17473,N_17008,N_17176);
xor U17474 (N_17474,N_17049,N_17007);
or U17475 (N_17475,N_17221,N_17156);
nor U17476 (N_17476,N_17082,N_17089);
nand U17477 (N_17477,N_17043,N_17164);
and U17478 (N_17478,N_17130,N_17181);
nand U17479 (N_17479,N_17158,N_17180);
xor U17480 (N_17480,N_17235,N_17104);
nor U17481 (N_17481,N_17223,N_17111);
nand U17482 (N_17482,N_17012,N_17217);
xnor U17483 (N_17483,N_17080,N_17138);
and U17484 (N_17484,N_17050,N_17120);
nor U17485 (N_17485,N_17181,N_17115);
xor U17486 (N_17486,N_17154,N_17106);
and U17487 (N_17487,N_17218,N_17038);
nor U17488 (N_17488,N_17215,N_17003);
or U17489 (N_17489,N_17139,N_17154);
and U17490 (N_17490,N_17091,N_17088);
and U17491 (N_17491,N_17227,N_17023);
and U17492 (N_17492,N_17081,N_17178);
nand U17493 (N_17493,N_17245,N_17200);
xnor U17494 (N_17494,N_17165,N_17173);
xor U17495 (N_17495,N_17030,N_17144);
nand U17496 (N_17496,N_17043,N_17068);
nor U17497 (N_17497,N_17182,N_17174);
and U17498 (N_17498,N_17024,N_17164);
and U17499 (N_17499,N_17082,N_17218);
nand U17500 (N_17500,N_17339,N_17253);
xor U17501 (N_17501,N_17336,N_17313);
nand U17502 (N_17502,N_17435,N_17482);
xor U17503 (N_17503,N_17346,N_17382);
xor U17504 (N_17504,N_17439,N_17412);
or U17505 (N_17505,N_17283,N_17415);
and U17506 (N_17506,N_17259,N_17368);
xnor U17507 (N_17507,N_17442,N_17457);
xnor U17508 (N_17508,N_17342,N_17320);
nor U17509 (N_17509,N_17443,N_17341);
or U17510 (N_17510,N_17327,N_17483);
nor U17511 (N_17511,N_17325,N_17498);
and U17512 (N_17512,N_17445,N_17438);
xnor U17513 (N_17513,N_17413,N_17315);
nor U17514 (N_17514,N_17321,N_17486);
nand U17515 (N_17515,N_17296,N_17366);
nor U17516 (N_17516,N_17251,N_17453);
nand U17517 (N_17517,N_17417,N_17372);
or U17518 (N_17518,N_17426,N_17396);
nor U17519 (N_17519,N_17495,N_17287);
and U17520 (N_17520,N_17356,N_17392);
or U17521 (N_17521,N_17385,N_17422);
nand U17522 (N_17522,N_17295,N_17257);
and U17523 (N_17523,N_17252,N_17390);
xnor U17524 (N_17524,N_17414,N_17352);
nor U17525 (N_17525,N_17303,N_17317);
nand U17526 (N_17526,N_17284,N_17319);
nand U17527 (N_17527,N_17416,N_17281);
nand U17528 (N_17528,N_17371,N_17465);
nand U17529 (N_17529,N_17496,N_17309);
xor U17530 (N_17530,N_17293,N_17467);
nand U17531 (N_17531,N_17298,N_17472);
and U17532 (N_17532,N_17263,N_17369);
xnor U17533 (N_17533,N_17481,N_17407);
nand U17534 (N_17534,N_17334,N_17494);
nand U17535 (N_17535,N_17423,N_17469);
or U17536 (N_17536,N_17456,N_17376);
nand U17537 (N_17537,N_17421,N_17305);
xnor U17538 (N_17538,N_17289,N_17280);
nand U17539 (N_17539,N_17454,N_17434);
nand U17540 (N_17540,N_17420,N_17492);
nand U17541 (N_17541,N_17398,N_17260);
or U17542 (N_17542,N_17402,N_17357);
xnor U17543 (N_17543,N_17447,N_17410);
xnor U17544 (N_17544,N_17405,N_17328);
nor U17545 (N_17545,N_17459,N_17288);
nor U17546 (N_17546,N_17449,N_17479);
or U17547 (N_17547,N_17347,N_17265);
xor U17548 (N_17548,N_17354,N_17406);
xnor U17549 (N_17549,N_17306,N_17437);
or U17550 (N_17550,N_17485,N_17345);
nand U17551 (N_17551,N_17411,N_17468);
xnor U17552 (N_17552,N_17489,N_17432);
nand U17553 (N_17553,N_17478,N_17463);
nand U17554 (N_17554,N_17264,N_17391);
or U17555 (N_17555,N_17379,N_17292);
nand U17556 (N_17556,N_17256,N_17466);
xnor U17557 (N_17557,N_17428,N_17349);
nand U17558 (N_17558,N_17361,N_17300);
nor U17559 (N_17559,N_17254,N_17312);
nand U17560 (N_17560,N_17408,N_17272);
or U17561 (N_17561,N_17353,N_17424);
xor U17562 (N_17562,N_17344,N_17395);
nand U17563 (N_17563,N_17316,N_17487);
and U17564 (N_17564,N_17324,N_17304);
nand U17565 (N_17565,N_17355,N_17318);
nand U17566 (N_17566,N_17294,N_17340);
and U17567 (N_17567,N_17343,N_17470);
or U17568 (N_17568,N_17399,N_17360);
or U17569 (N_17569,N_17330,N_17290);
or U17570 (N_17570,N_17490,N_17326);
nor U17571 (N_17571,N_17493,N_17475);
nand U17572 (N_17572,N_17394,N_17427);
nor U17573 (N_17573,N_17268,N_17279);
and U17574 (N_17574,N_17365,N_17451);
nor U17575 (N_17575,N_17429,N_17380);
or U17576 (N_17576,N_17364,N_17389);
or U17577 (N_17577,N_17266,N_17461);
nor U17578 (N_17578,N_17448,N_17378);
nor U17579 (N_17579,N_17446,N_17358);
xor U17580 (N_17580,N_17491,N_17350);
nor U17581 (N_17581,N_17262,N_17297);
and U17582 (N_17582,N_17261,N_17323);
nor U17583 (N_17583,N_17436,N_17258);
nor U17584 (N_17584,N_17308,N_17477);
xnor U17585 (N_17585,N_17488,N_17274);
and U17586 (N_17586,N_17278,N_17450);
or U17587 (N_17587,N_17383,N_17425);
nand U17588 (N_17588,N_17433,N_17374);
nand U17589 (N_17589,N_17286,N_17419);
nand U17590 (N_17590,N_17277,N_17291);
or U17591 (N_17591,N_17388,N_17359);
or U17592 (N_17592,N_17431,N_17386);
nor U17593 (N_17593,N_17418,N_17307);
or U17594 (N_17594,N_17273,N_17282);
nor U17595 (N_17595,N_17458,N_17362);
and U17596 (N_17596,N_17460,N_17370);
xnor U17597 (N_17597,N_17335,N_17276);
or U17598 (N_17598,N_17484,N_17471);
xnor U17599 (N_17599,N_17387,N_17267);
or U17600 (N_17600,N_17299,N_17462);
or U17601 (N_17601,N_17269,N_17499);
and U17602 (N_17602,N_17363,N_17440);
xor U17603 (N_17603,N_17275,N_17444);
xor U17604 (N_17604,N_17301,N_17285);
xor U17605 (N_17605,N_17452,N_17480);
nand U17606 (N_17606,N_17322,N_17497);
nand U17607 (N_17607,N_17375,N_17250);
xnor U17608 (N_17608,N_17271,N_17377);
and U17609 (N_17609,N_17310,N_17255);
nor U17610 (N_17610,N_17314,N_17384);
and U17611 (N_17611,N_17474,N_17403);
xnor U17612 (N_17612,N_17270,N_17409);
nand U17613 (N_17613,N_17332,N_17393);
and U17614 (N_17614,N_17367,N_17455);
or U17615 (N_17615,N_17333,N_17311);
nand U17616 (N_17616,N_17302,N_17351);
or U17617 (N_17617,N_17400,N_17430);
or U17618 (N_17618,N_17464,N_17337);
and U17619 (N_17619,N_17373,N_17397);
xnor U17620 (N_17620,N_17404,N_17348);
or U17621 (N_17621,N_17473,N_17441);
nand U17622 (N_17622,N_17338,N_17331);
nand U17623 (N_17623,N_17381,N_17329);
and U17624 (N_17624,N_17401,N_17476);
xnor U17625 (N_17625,N_17434,N_17426);
xor U17626 (N_17626,N_17388,N_17273);
xnor U17627 (N_17627,N_17428,N_17392);
and U17628 (N_17628,N_17417,N_17435);
or U17629 (N_17629,N_17385,N_17372);
nor U17630 (N_17630,N_17365,N_17370);
xnor U17631 (N_17631,N_17274,N_17310);
and U17632 (N_17632,N_17270,N_17337);
nand U17633 (N_17633,N_17305,N_17392);
nor U17634 (N_17634,N_17391,N_17418);
nor U17635 (N_17635,N_17437,N_17393);
nor U17636 (N_17636,N_17324,N_17499);
xnor U17637 (N_17637,N_17350,N_17278);
nand U17638 (N_17638,N_17364,N_17496);
xor U17639 (N_17639,N_17465,N_17383);
nor U17640 (N_17640,N_17297,N_17411);
or U17641 (N_17641,N_17325,N_17496);
xnor U17642 (N_17642,N_17444,N_17442);
xor U17643 (N_17643,N_17473,N_17498);
or U17644 (N_17644,N_17492,N_17483);
and U17645 (N_17645,N_17480,N_17256);
nand U17646 (N_17646,N_17370,N_17498);
and U17647 (N_17647,N_17357,N_17320);
nor U17648 (N_17648,N_17479,N_17444);
nand U17649 (N_17649,N_17467,N_17469);
and U17650 (N_17650,N_17384,N_17400);
nand U17651 (N_17651,N_17367,N_17282);
nor U17652 (N_17652,N_17418,N_17367);
and U17653 (N_17653,N_17313,N_17456);
xnor U17654 (N_17654,N_17279,N_17265);
or U17655 (N_17655,N_17495,N_17405);
or U17656 (N_17656,N_17320,N_17258);
nand U17657 (N_17657,N_17334,N_17490);
nand U17658 (N_17658,N_17345,N_17304);
nand U17659 (N_17659,N_17400,N_17276);
nor U17660 (N_17660,N_17354,N_17457);
or U17661 (N_17661,N_17487,N_17489);
or U17662 (N_17662,N_17310,N_17449);
nor U17663 (N_17663,N_17303,N_17452);
and U17664 (N_17664,N_17467,N_17364);
nor U17665 (N_17665,N_17404,N_17365);
or U17666 (N_17666,N_17418,N_17497);
or U17667 (N_17667,N_17254,N_17309);
xnor U17668 (N_17668,N_17343,N_17299);
or U17669 (N_17669,N_17402,N_17450);
or U17670 (N_17670,N_17366,N_17330);
nand U17671 (N_17671,N_17420,N_17298);
and U17672 (N_17672,N_17349,N_17405);
xnor U17673 (N_17673,N_17463,N_17400);
nand U17674 (N_17674,N_17356,N_17307);
nand U17675 (N_17675,N_17353,N_17420);
nand U17676 (N_17676,N_17400,N_17407);
nor U17677 (N_17677,N_17460,N_17258);
or U17678 (N_17678,N_17293,N_17296);
or U17679 (N_17679,N_17264,N_17284);
or U17680 (N_17680,N_17296,N_17260);
xnor U17681 (N_17681,N_17316,N_17358);
or U17682 (N_17682,N_17346,N_17385);
and U17683 (N_17683,N_17373,N_17339);
xor U17684 (N_17684,N_17252,N_17490);
xnor U17685 (N_17685,N_17420,N_17495);
nor U17686 (N_17686,N_17371,N_17404);
nand U17687 (N_17687,N_17347,N_17274);
xor U17688 (N_17688,N_17475,N_17271);
nor U17689 (N_17689,N_17489,N_17339);
xor U17690 (N_17690,N_17379,N_17261);
xnor U17691 (N_17691,N_17263,N_17381);
nor U17692 (N_17692,N_17279,N_17429);
and U17693 (N_17693,N_17452,N_17486);
nor U17694 (N_17694,N_17436,N_17420);
xnor U17695 (N_17695,N_17273,N_17442);
nand U17696 (N_17696,N_17380,N_17317);
xnor U17697 (N_17697,N_17479,N_17493);
and U17698 (N_17698,N_17488,N_17334);
nor U17699 (N_17699,N_17364,N_17447);
and U17700 (N_17700,N_17326,N_17361);
and U17701 (N_17701,N_17364,N_17490);
nand U17702 (N_17702,N_17381,N_17471);
nor U17703 (N_17703,N_17373,N_17287);
or U17704 (N_17704,N_17497,N_17358);
xor U17705 (N_17705,N_17303,N_17326);
nor U17706 (N_17706,N_17270,N_17358);
xnor U17707 (N_17707,N_17482,N_17438);
xnor U17708 (N_17708,N_17380,N_17403);
or U17709 (N_17709,N_17260,N_17400);
or U17710 (N_17710,N_17297,N_17359);
nor U17711 (N_17711,N_17423,N_17485);
nand U17712 (N_17712,N_17432,N_17358);
or U17713 (N_17713,N_17472,N_17325);
or U17714 (N_17714,N_17447,N_17459);
nor U17715 (N_17715,N_17423,N_17305);
and U17716 (N_17716,N_17437,N_17270);
nand U17717 (N_17717,N_17469,N_17363);
nand U17718 (N_17718,N_17290,N_17405);
nand U17719 (N_17719,N_17469,N_17361);
or U17720 (N_17720,N_17435,N_17284);
nand U17721 (N_17721,N_17390,N_17370);
and U17722 (N_17722,N_17358,N_17402);
and U17723 (N_17723,N_17305,N_17297);
and U17724 (N_17724,N_17382,N_17442);
nor U17725 (N_17725,N_17416,N_17277);
nand U17726 (N_17726,N_17330,N_17315);
or U17727 (N_17727,N_17322,N_17297);
nor U17728 (N_17728,N_17347,N_17283);
nand U17729 (N_17729,N_17386,N_17322);
and U17730 (N_17730,N_17268,N_17254);
or U17731 (N_17731,N_17463,N_17355);
or U17732 (N_17732,N_17412,N_17489);
nor U17733 (N_17733,N_17255,N_17378);
nand U17734 (N_17734,N_17373,N_17443);
or U17735 (N_17735,N_17348,N_17265);
nand U17736 (N_17736,N_17261,N_17431);
and U17737 (N_17737,N_17484,N_17385);
and U17738 (N_17738,N_17392,N_17362);
or U17739 (N_17739,N_17391,N_17334);
xor U17740 (N_17740,N_17378,N_17282);
xnor U17741 (N_17741,N_17259,N_17489);
xor U17742 (N_17742,N_17373,N_17453);
and U17743 (N_17743,N_17442,N_17378);
nor U17744 (N_17744,N_17429,N_17414);
nand U17745 (N_17745,N_17486,N_17372);
or U17746 (N_17746,N_17417,N_17461);
xnor U17747 (N_17747,N_17328,N_17396);
and U17748 (N_17748,N_17276,N_17310);
xor U17749 (N_17749,N_17359,N_17378);
nor U17750 (N_17750,N_17582,N_17574);
nand U17751 (N_17751,N_17736,N_17650);
nor U17752 (N_17752,N_17543,N_17592);
nor U17753 (N_17753,N_17531,N_17730);
and U17754 (N_17754,N_17746,N_17708);
nor U17755 (N_17755,N_17699,N_17537);
or U17756 (N_17756,N_17559,N_17720);
or U17757 (N_17757,N_17682,N_17677);
nand U17758 (N_17758,N_17716,N_17539);
nor U17759 (N_17759,N_17642,N_17684);
xor U17760 (N_17760,N_17554,N_17738);
nor U17761 (N_17761,N_17610,N_17611);
or U17762 (N_17762,N_17533,N_17643);
xnor U17763 (N_17763,N_17671,N_17581);
nand U17764 (N_17764,N_17673,N_17651);
nor U17765 (N_17765,N_17664,N_17548);
nand U17766 (N_17766,N_17656,N_17696);
or U17767 (N_17767,N_17733,N_17641);
xor U17768 (N_17768,N_17702,N_17535);
nand U17769 (N_17769,N_17549,N_17508);
or U17770 (N_17770,N_17542,N_17686);
or U17771 (N_17771,N_17711,N_17676);
nor U17772 (N_17772,N_17705,N_17749);
nor U17773 (N_17773,N_17516,N_17534);
nor U17774 (N_17774,N_17694,N_17727);
or U17775 (N_17775,N_17707,N_17504);
xnor U17776 (N_17776,N_17675,N_17713);
and U17777 (N_17777,N_17566,N_17739);
nor U17778 (N_17778,N_17547,N_17612);
xor U17779 (N_17779,N_17595,N_17583);
or U17780 (N_17780,N_17678,N_17502);
and U17781 (N_17781,N_17538,N_17695);
nor U17782 (N_17782,N_17556,N_17584);
or U17783 (N_17783,N_17687,N_17629);
xor U17784 (N_17784,N_17741,N_17725);
nand U17785 (N_17785,N_17514,N_17567);
and U17786 (N_17786,N_17679,N_17526);
and U17787 (N_17787,N_17580,N_17748);
and U17788 (N_17788,N_17555,N_17619);
xnor U17789 (N_17789,N_17659,N_17557);
nor U17790 (N_17790,N_17530,N_17623);
nor U17791 (N_17791,N_17621,N_17525);
and U17792 (N_17792,N_17731,N_17562);
nand U17793 (N_17793,N_17532,N_17624);
or U17794 (N_17794,N_17510,N_17578);
or U17795 (N_17795,N_17710,N_17545);
nand U17796 (N_17796,N_17600,N_17615);
nor U17797 (N_17797,N_17597,N_17568);
or U17798 (N_17798,N_17631,N_17518);
or U17799 (N_17799,N_17717,N_17552);
and U17800 (N_17800,N_17709,N_17575);
xnor U17801 (N_17801,N_17569,N_17617);
or U17802 (N_17802,N_17669,N_17590);
nand U17803 (N_17803,N_17561,N_17647);
xnor U17804 (N_17804,N_17640,N_17521);
nor U17805 (N_17805,N_17718,N_17744);
nand U17806 (N_17806,N_17564,N_17594);
and U17807 (N_17807,N_17740,N_17745);
or U17808 (N_17808,N_17704,N_17614);
nand U17809 (N_17809,N_17726,N_17637);
nor U17810 (N_17810,N_17625,N_17729);
nor U17811 (N_17811,N_17692,N_17700);
and U17812 (N_17812,N_17654,N_17529);
and U17813 (N_17813,N_17691,N_17620);
xnor U17814 (N_17814,N_17528,N_17724);
or U17815 (N_17815,N_17616,N_17734);
or U17816 (N_17816,N_17645,N_17500);
xnor U17817 (N_17817,N_17509,N_17553);
or U17818 (N_17818,N_17608,N_17573);
nor U17819 (N_17819,N_17506,N_17701);
nor U17820 (N_17820,N_17536,N_17630);
nand U17821 (N_17821,N_17618,N_17681);
and U17822 (N_17822,N_17572,N_17546);
nor U17823 (N_17823,N_17660,N_17698);
or U17824 (N_17824,N_17663,N_17587);
nand U17825 (N_17825,N_17633,N_17639);
xor U17826 (N_17826,N_17605,N_17517);
nor U17827 (N_17827,N_17541,N_17742);
nor U17828 (N_17828,N_17551,N_17712);
and U17829 (N_17829,N_17644,N_17527);
or U17830 (N_17830,N_17680,N_17719);
nor U17831 (N_17831,N_17604,N_17683);
nand U17832 (N_17832,N_17693,N_17560);
nor U17833 (N_17833,N_17593,N_17653);
nor U17834 (N_17834,N_17628,N_17588);
nor U17835 (N_17835,N_17522,N_17632);
and U17836 (N_17836,N_17685,N_17607);
nor U17837 (N_17837,N_17737,N_17576);
nand U17838 (N_17838,N_17638,N_17703);
nor U17839 (N_17839,N_17507,N_17571);
and U17840 (N_17840,N_17688,N_17511);
or U17841 (N_17841,N_17723,N_17697);
xnor U17842 (N_17842,N_17667,N_17646);
nand U17843 (N_17843,N_17732,N_17657);
nor U17844 (N_17844,N_17666,N_17513);
and U17845 (N_17845,N_17635,N_17558);
and U17846 (N_17846,N_17603,N_17722);
nand U17847 (N_17847,N_17550,N_17598);
and U17848 (N_17848,N_17599,N_17577);
nand U17849 (N_17849,N_17512,N_17540);
xnor U17850 (N_17850,N_17520,N_17613);
and U17851 (N_17851,N_17626,N_17747);
or U17852 (N_17852,N_17672,N_17501);
nand U17853 (N_17853,N_17655,N_17658);
or U17854 (N_17854,N_17649,N_17579);
nor U17855 (N_17855,N_17689,N_17503);
nand U17856 (N_17856,N_17565,N_17743);
xnor U17857 (N_17857,N_17586,N_17570);
and U17858 (N_17858,N_17606,N_17721);
nor U17859 (N_17859,N_17648,N_17622);
and U17860 (N_17860,N_17636,N_17665);
xnor U17861 (N_17861,N_17662,N_17505);
nor U17862 (N_17862,N_17668,N_17735);
nand U17863 (N_17863,N_17670,N_17523);
or U17864 (N_17864,N_17515,N_17661);
xor U17865 (N_17865,N_17715,N_17602);
nor U17866 (N_17866,N_17652,N_17601);
and U17867 (N_17867,N_17728,N_17714);
and U17868 (N_17868,N_17589,N_17524);
or U17869 (N_17869,N_17563,N_17596);
or U17870 (N_17870,N_17519,N_17706);
nand U17871 (N_17871,N_17627,N_17585);
nor U17872 (N_17872,N_17544,N_17634);
and U17873 (N_17873,N_17591,N_17690);
xor U17874 (N_17874,N_17674,N_17609);
or U17875 (N_17875,N_17701,N_17747);
or U17876 (N_17876,N_17570,N_17717);
nor U17877 (N_17877,N_17622,N_17552);
and U17878 (N_17878,N_17538,N_17702);
and U17879 (N_17879,N_17616,N_17593);
and U17880 (N_17880,N_17500,N_17650);
or U17881 (N_17881,N_17613,N_17712);
xor U17882 (N_17882,N_17558,N_17608);
and U17883 (N_17883,N_17629,N_17575);
and U17884 (N_17884,N_17555,N_17559);
and U17885 (N_17885,N_17636,N_17667);
nand U17886 (N_17886,N_17523,N_17689);
xnor U17887 (N_17887,N_17658,N_17572);
or U17888 (N_17888,N_17515,N_17624);
nor U17889 (N_17889,N_17625,N_17635);
nor U17890 (N_17890,N_17611,N_17627);
or U17891 (N_17891,N_17738,N_17649);
nor U17892 (N_17892,N_17529,N_17638);
xnor U17893 (N_17893,N_17643,N_17615);
and U17894 (N_17894,N_17537,N_17719);
or U17895 (N_17895,N_17543,N_17549);
nand U17896 (N_17896,N_17727,N_17673);
or U17897 (N_17897,N_17747,N_17567);
or U17898 (N_17898,N_17525,N_17591);
nor U17899 (N_17899,N_17696,N_17567);
nand U17900 (N_17900,N_17719,N_17541);
xor U17901 (N_17901,N_17560,N_17543);
nor U17902 (N_17902,N_17744,N_17558);
xor U17903 (N_17903,N_17529,N_17554);
xnor U17904 (N_17904,N_17545,N_17604);
and U17905 (N_17905,N_17742,N_17663);
or U17906 (N_17906,N_17672,N_17727);
nand U17907 (N_17907,N_17738,N_17645);
or U17908 (N_17908,N_17633,N_17657);
xor U17909 (N_17909,N_17746,N_17531);
and U17910 (N_17910,N_17694,N_17726);
and U17911 (N_17911,N_17539,N_17745);
or U17912 (N_17912,N_17699,N_17568);
nand U17913 (N_17913,N_17605,N_17731);
and U17914 (N_17914,N_17668,N_17744);
nand U17915 (N_17915,N_17600,N_17537);
xor U17916 (N_17916,N_17573,N_17748);
xnor U17917 (N_17917,N_17628,N_17506);
nor U17918 (N_17918,N_17655,N_17614);
nor U17919 (N_17919,N_17712,N_17558);
nand U17920 (N_17920,N_17703,N_17578);
and U17921 (N_17921,N_17668,N_17663);
or U17922 (N_17922,N_17543,N_17701);
nor U17923 (N_17923,N_17728,N_17705);
or U17924 (N_17924,N_17742,N_17617);
and U17925 (N_17925,N_17679,N_17629);
or U17926 (N_17926,N_17643,N_17504);
and U17927 (N_17927,N_17681,N_17742);
or U17928 (N_17928,N_17578,N_17528);
nand U17929 (N_17929,N_17669,N_17637);
or U17930 (N_17930,N_17559,N_17602);
xor U17931 (N_17931,N_17686,N_17522);
nand U17932 (N_17932,N_17706,N_17646);
xnor U17933 (N_17933,N_17576,N_17604);
or U17934 (N_17934,N_17730,N_17561);
nor U17935 (N_17935,N_17709,N_17536);
nand U17936 (N_17936,N_17707,N_17516);
xnor U17937 (N_17937,N_17723,N_17572);
xnor U17938 (N_17938,N_17703,N_17732);
or U17939 (N_17939,N_17737,N_17539);
and U17940 (N_17940,N_17563,N_17588);
or U17941 (N_17941,N_17553,N_17628);
and U17942 (N_17942,N_17635,N_17725);
or U17943 (N_17943,N_17581,N_17723);
and U17944 (N_17944,N_17582,N_17674);
nand U17945 (N_17945,N_17688,N_17549);
nor U17946 (N_17946,N_17721,N_17603);
nor U17947 (N_17947,N_17642,N_17578);
xnor U17948 (N_17948,N_17625,N_17712);
nand U17949 (N_17949,N_17651,N_17621);
xor U17950 (N_17950,N_17587,N_17690);
nor U17951 (N_17951,N_17573,N_17649);
and U17952 (N_17952,N_17699,N_17528);
nand U17953 (N_17953,N_17674,N_17547);
nor U17954 (N_17954,N_17640,N_17572);
nand U17955 (N_17955,N_17683,N_17620);
or U17956 (N_17956,N_17614,N_17563);
or U17957 (N_17957,N_17620,N_17505);
nand U17958 (N_17958,N_17715,N_17740);
xor U17959 (N_17959,N_17654,N_17728);
nor U17960 (N_17960,N_17664,N_17660);
xor U17961 (N_17961,N_17617,N_17736);
nor U17962 (N_17962,N_17521,N_17652);
or U17963 (N_17963,N_17608,N_17504);
nor U17964 (N_17964,N_17617,N_17740);
and U17965 (N_17965,N_17583,N_17644);
nand U17966 (N_17966,N_17743,N_17739);
nor U17967 (N_17967,N_17702,N_17701);
xor U17968 (N_17968,N_17525,N_17661);
nand U17969 (N_17969,N_17640,N_17654);
or U17970 (N_17970,N_17556,N_17573);
nand U17971 (N_17971,N_17711,N_17728);
nand U17972 (N_17972,N_17554,N_17617);
xnor U17973 (N_17973,N_17706,N_17730);
and U17974 (N_17974,N_17661,N_17706);
or U17975 (N_17975,N_17656,N_17534);
xnor U17976 (N_17976,N_17729,N_17696);
xor U17977 (N_17977,N_17696,N_17734);
nor U17978 (N_17978,N_17659,N_17738);
or U17979 (N_17979,N_17546,N_17511);
nor U17980 (N_17980,N_17568,N_17552);
nor U17981 (N_17981,N_17704,N_17707);
nand U17982 (N_17982,N_17727,N_17652);
nor U17983 (N_17983,N_17638,N_17708);
nand U17984 (N_17984,N_17738,N_17721);
or U17985 (N_17985,N_17714,N_17500);
xor U17986 (N_17986,N_17544,N_17659);
and U17987 (N_17987,N_17558,N_17535);
or U17988 (N_17988,N_17652,N_17714);
xnor U17989 (N_17989,N_17625,N_17545);
or U17990 (N_17990,N_17510,N_17733);
or U17991 (N_17991,N_17655,N_17596);
xor U17992 (N_17992,N_17717,N_17636);
nand U17993 (N_17993,N_17578,N_17686);
nor U17994 (N_17994,N_17578,N_17591);
nor U17995 (N_17995,N_17567,N_17634);
or U17996 (N_17996,N_17520,N_17573);
nor U17997 (N_17997,N_17738,N_17677);
and U17998 (N_17998,N_17559,N_17608);
or U17999 (N_17999,N_17510,N_17586);
or U18000 (N_18000,N_17994,N_17951);
and U18001 (N_18001,N_17807,N_17812);
nor U18002 (N_18002,N_17753,N_17840);
xnor U18003 (N_18003,N_17973,N_17824);
nand U18004 (N_18004,N_17910,N_17974);
or U18005 (N_18005,N_17943,N_17938);
nor U18006 (N_18006,N_17887,N_17911);
nand U18007 (N_18007,N_17995,N_17772);
and U18008 (N_18008,N_17971,N_17789);
nand U18009 (N_18009,N_17884,N_17852);
and U18010 (N_18010,N_17932,N_17888);
and U18011 (N_18011,N_17841,N_17865);
nand U18012 (N_18012,N_17766,N_17831);
xnor U18013 (N_18013,N_17979,N_17886);
or U18014 (N_18014,N_17760,N_17958);
and U18015 (N_18015,N_17845,N_17809);
and U18016 (N_18016,N_17872,N_17790);
nor U18017 (N_18017,N_17913,N_17944);
or U18018 (N_18018,N_17774,N_17785);
and U18019 (N_18019,N_17817,N_17851);
nand U18020 (N_18020,N_17870,N_17961);
xor U18021 (N_18021,N_17839,N_17819);
and U18022 (N_18022,N_17952,N_17877);
nand U18023 (N_18023,N_17863,N_17968);
nor U18024 (N_18024,N_17988,N_17883);
nor U18025 (N_18025,N_17837,N_17823);
nand U18026 (N_18026,N_17779,N_17975);
nand U18027 (N_18027,N_17929,N_17927);
nand U18028 (N_18028,N_17868,N_17876);
and U18029 (N_18029,N_17818,N_17964);
and U18030 (N_18030,N_17891,N_17900);
nand U18031 (N_18031,N_17759,N_17866);
nand U18032 (N_18032,N_17786,N_17916);
or U18033 (N_18033,N_17889,N_17764);
and U18034 (N_18034,N_17821,N_17776);
nand U18035 (N_18035,N_17836,N_17761);
and U18036 (N_18036,N_17792,N_17834);
xnor U18037 (N_18037,N_17903,N_17780);
and U18038 (N_18038,N_17783,N_17893);
and U18039 (N_18039,N_17775,N_17918);
xor U18040 (N_18040,N_17989,N_17970);
nand U18041 (N_18041,N_17940,N_17885);
or U18042 (N_18042,N_17922,N_17985);
nand U18043 (N_18043,N_17859,N_17782);
nand U18044 (N_18044,N_17934,N_17805);
nand U18045 (N_18045,N_17757,N_17867);
or U18046 (N_18046,N_17925,N_17962);
nor U18047 (N_18047,N_17983,N_17978);
xnor U18048 (N_18048,N_17763,N_17976);
nand U18049 (N_18049,N_17890,N_17827);
nor U18050 (N_18050,N_17750,N_17882);
and U18051 (N_18051,N_17857,N_17806);
and U18052 (N_18052,N_17767,N_17858);
nand U18053 (N_18053,N_17998,N_17802);
or U18054 (N_18054,N_17898,N_17803);
nor U18055 (N_18055,N_17933,N_17904);
nand U18056 (N_18056,N_17822,N_17751);
nor U18057 (N_18057,N_17773,N_17919);
or U18058 (N_18058,N_17873,N_17784);
nand U18059 (N_18059,N_17941,N_17928);
and U18060 (N_18060,N_17993,N_17980);
or U18061 (N_18061,N_17999,N_17871);
xnor U18062 (N_18062,N_17847,N_17788);
nand U18063 (N_18063,N_17829,N_17917);
or U18064 (N_18064,N_17752,N_17849);
nor U18065 (N_18065,N_17756,N_17797);
and U18066 (N_18066,N_17956,N_17768);
nand U18067 (N_18067,N_17820,N_17825);
or U18068 (N_18068,N_17930,N_17869);
xnor U18069 (N_18069,N_17905,N_17948);
nand U18070 (N_18070,N_17897,N_17770);
nor U18071 (N_18071,N_17828,N_17984);
nand U18072 (N_18072,N_17915,N_17950);
xor U18073 (N_18073,N_17754,N_17798);
or U18074 (N_18074,N_17926,N_17935);
nor U18075 (N_18075,N_17896,N_17864);
and U18076 (N_18076,N_17875,N_17791);
nand U18077 (N_18077,N_17856,N_17957);
nand U18078 (N_18078,N_17843,N_17992);
nand U18079 (N_18079,N_17846,N_17967);
or U18080 (N_18080,N_17954,N_17924);
xor U18081 (N_18081,N_17781,N_17842);
and U18082 (N_18082,N_17982,N_17920);
nor U18083 (N_18083,N_17879,N_17912);
nor U18084 (N_18084,N_17909,N_17794);
nand U18085 (N_18085,N_17937,N_17808);
xor U18086 (N_18086,N_17850,N_17947);
nor U18087 (N_18087,N_17907,N_17874);
nand U18088 (N_18088,N_17804,N_17965);
nor U18089 (N_18089,N_17906,N_17953);
nor U18090 (N_18090,N_17908,N_17801);
nand U18091 (N_18091,N_17799,N_17796);
or U18092 (N_18092,N_17977,N_17878);
xor U18093 (N_18093,N_17966,N_17931);
and U18094 (N_18094,N_17832,N_17771);
xnor U18095 (N_18095,N_17815,N_17861);
nor U18096 (N_18096,N_17899,N_17945);
nor U18097 (N_18097,N_17830,N_17810);
and U18098 (N_18098,N_17787,N_17811);
nand U18099 (N_18099,N_17959,N_17939);
and U18100 (N_18100,N_17987,N_17769);
and U18101 (N_18101,N_17755,N_17960);
and U18102 (N_18102,N_17986,N_17969);
nand U18103 (N_18103,N_17990,N_17895);
and U18104 (N_18104,N_17914,N_17894);
and U18105 (N_18105,N_17854,N_17991);
or U18106 (N_18106,N_17981,N_17833);
or U18107 (N_18107,N_17923,N_17758);
xor U18108 (N_18108,N_17765,N_17762);
or U18109 (N_18109,N_17942,N_17835);
and U18110 (N_18110,N_17777,N_17813);
and U18111 (N_18111,N_17855,N_17921);
or U18112 (N_18112,N_17800,N_17949);
nor U18113 (N_18113,N_17838,N_17778);
or U18114 (N_18114,N_17816,N_17901);
xnor U18115 (N_18115,N_17795,N_17814);
or U18116 (N_18116,N_17996,N_17793);
nand U18117 (N_18117,N_17844,N_17997);
or U18118 (N_18118,N_17963,N_17826);
and U18119 (N_18119,N_17860,N_17892);
or U18120 (N_18120,N_17881,N_17902);
or U18121 (N_18121,N_17848,N_17862);
or U18122 (N_18122,N_17972,N_17946);
nor U18123 (N_18123,N_17853,N_17955);
or U18124 (N_18124,N_17880,N_17936);
nand U18125 (N_18125,N_17964,N_17886);
nor U18126 (N_18126,N_17852,N_17938);
nor U18127 (N_18127,N_17795,N_17948);
or U18128 (N_18128,N_17975,N_17867);
xnor U18129 (N_18129,N_17813,N_17799);
nand U18130 (N_18130,N_17911,N_17757);
and U18131 (N_18131,N_17823,N_17788);
xor U18132 (N_18132,N_17891,N_17818);
and U18133 (N_18133,N_17827,N_17823);
nand U18134 (N_18134,N_17925,N_17842);
and U18135 (N_18135,N_17994,N_17933);
nand U18136 (N_18136,N_17780,N_17772);
or U18137 (N_18137,N_17882,N_17851);
nand U18138 (N_18138,N_17861,N_17761);
and U18139 (N_18139,N_17854,N_17755);
and U18140 (N_18140,N_17987,N_17955);
and U18141 (N_18141,N_17807,N_17991);
nand U18142 (N_18142,N_17817,N_17821);
xnor U18143 (N_18143,N_17844,N_17981);
nand U18144 (N_18144,N_17834,N_17847);
and U18145 (N_18145,N_17916,N_17883);
nand U18146 (N_18146,N_17923,N_17976);
or U18147 (N_18147,N_17911,N_17959);
xnor U18148 (N_18148,N_17769,N_17898);
and U18149 (N_18149,N_17789,N_17803);
or U18150 (N_18150,N_17960,N_17768);
nor U18151 (N_18151,N_17758,N_17836);
nand U18152 (N_18152,N_17928,N_17912);
nor U18153 (N_18153,N_17915,N_17765);
xnor U18154 (N_18154,N_17914,N_17934);
and U18155 (N_18155,N_17956,N_17949);
nor U18156 (N_18156,N_17897,N_17966);
nand U18157 (N_18157,N_17906,N_17878);
nor U18158 (N_18158,N_17831,N_17965);
xor U18159 (N_18159,N_17910,N_17794);
or U18160 (N_18160,N_17775,N_17965);
nand U18161 (N_18161,N_17865,N_17866);
nand U18162 (N_18162,N_17968,N_17788);
nand U18163 (N_18163,N_17941,N_17787);
nor U18164 (N_18164,N_17782,N_17751);
nand U18165 (N_18165,N_17843,N_17782);
nand U18166 (N_18166,N_17800,N_17822);
and U18167 (N_18167,N_17755,N_17895);
nor U18168 (N_18168,N_17893,N_17770);
nor U18169 (N_18169,N_17912,N_17828);
nor U18170 (N_18170,N_17826,N_17773);
xor U18171 (N_18171,N_17918,N_17984);
xnor U18172 (N_18172,N_17766,N_17935);
xor U18173 (N_18173,N_17977,N_17842);
nor U18174 (N_18174,N_17765,N_17773);
and U18175 (N_18175,N_17878,N_17955);
xor U18176 (N_18176,N_17911,N_17993);
and U18177 (N_18177,N_17873,N_17852);
and U18178 (N_18178,N_17770,N_17798);
xor U18179 (N_18179,N_17935,N_17810);
or U18180 (N_18180,N_17954,N_17980);
or U18181 (N_18181,N_17958,N_17852);
and U18182 (N_18182,N_17887,N_17824);
xor U18183 (N_18183,N_17843,N_17960);
or U18184 (N_18184,N_17809,N_17774);
xnor U18185 (N_18185,N_17873,N_17997);
nor U18186 (N_18186,N_17880,N_17857);
or U18187 (N_18187,N_17784,N_17793);
nand U18188 (N_18188,N_17787,N_17813);
xor U18189 (N_18189,N_17983,N_17950);
nor U18190 (N_18190,N_17896,N_17777);
nor U18191 (N_18191,N_17791,N_17901);
nor U18192 (N_18192,N_17960,N_17817);
nand U18193 (N_18193,N_17802,N_17775);
or U18194 (N_18194,N_17817,N_17772);
nor U18195 (N_18195,N_17868,N_17896);
xnor U18196 (N_18196,N_17811,N_17865);
nor U18197 (N_18197,N_17994,N_17993);
xor U18198 (N_18198,N_17978,N_17774);
nor U18199 (N_18199,N_17970,N_17979);
xnor U18200 (N_18200,N_17955,N_17810);
xnor U18201 (N_18201,N_17860,N_17937);
xnor U18202 (N_18202,N_17936,N_17902);
or U18203 (N_18203,N_17785,N_17974);
nor U18204 (N_18204,N_17751,N_17971);
nor U18205 (N_18205,N_17844,N_17861);
or U18206 (N_18206,N_17809,N_17812);
xor U18207 (N_18207,N_17995,N_17752);
nor U18208 (N_18208,N_17826,N_17847);
nand U18209 (N_18209,N_17832,N_17761);
nand U18210 (N_18210,N_17916,N_17964);
xnor U18211 (N_18211,N_17798,N_17987);
nand U18212 (N_18212,N_17759,N_17838);
xor U18213 (N_18213,N_17792,N_17906);
nand U18214 (N_18214,N_17909,N_17946);
xnor U18215 (N_18215,N_17919,N_17982);
or U18216 (N_18216,N_17977,N_17807);
nand U18217 (N_18217,N_17825,N_17883);
xor U18218 (N_18218,N_17935,N_17755);
and U18219 (N_18219,N_17883,N_17896);
or U18220 (N_18220,N_17885,N_17912);
nor U18221 (N_18221,N_17787,N_17959);
or U18222 (N_18222,N_17879,N_17837);
xor U18223 (N_18223,N_17803,N_17912);
or U18224 (N_18224,N_17901,N_17979);
nor U18225 (N_18225,N_17857,N_17948);
xor U18226 (N_18226,N_17922,N_17999);
and U18227 (N_18227,N_17842,N_17995);
and U18228 (N_18228,N_17877,N_17783);
nand U18229 (N_18229,N_17882,N_17767);
and U18230 (N_18230,N_17865,N_17968);
xnor U18231 (N_18231,N_17928,N_17902);
xnor U18232 (N_18232,N_17872,N_17779);
nand U18233 (N_18233,N_17890,N_17781);
nor U18234 (N_18234,N_17903,N_17868);
and U18235 (N_18235,N_17833,N_17993);
or U18236 (N_18236,N_17914,N_17971);
or U18237 (N_18237,N_17886,N_17959);
xnor U18238 (N_18238,N_17982,N_17811);
nor U18239 (N_18239,N_17913,N_17970);
or U18240 (N_18240,N_17978,N_17926);
nand U18241 (N_18241,N_17823,N_17765);
nor U18242 (N_18242,N_17977,N_17838);
nor U18243 (N_18243,N_17936,N_17916);
or U18244 (N_18244,N_17901,N_17863);
and U18245 (N_18245,N_17832,N_17843);
xor U18246 (N_18246,N_17827,N_17846);
and U18247 (N_18247,N_17978,N_17872);
nor U18248 (N_18248,N_17861,N_17967);
or U18249 (N_18249,N_17830,N_17980);
and U18250 (N_18250,N_18004,N_18104);
or U18251 (N_18251,N_18095,N_18006);
nand U18252 (N_18252,N_18149,N_18045);
nor U18253 (N_18253,N_18061,N_18221);
nand U18254 (N_18254,N_18066,N_18226);
xnor U18255 (N_18255,N_18236,N_18084);
nor U18256 (N_18256,N_18165,N_18164);
nand U18257 (N_18257,N_18182,N_18198);
xor U18258 (N_18258,N_18213,N_18009);
nor U18259 (N_18259,N_18239,N_18142);
and U18260 (N_18260,N_18148,N_18057);
nand U18261 (N_18261,N_18167,N_18209);
nor U18262 (N_18262,N_18185,N_18144);
xnor U18263 (N_18263,N_18150,N_18079);
and U18264 (N_18264,N_18056,N_18014);
nor U18265 (N_18265,N_18211,N_18080);
xor U18266 (N_18266,N_18063,N_18127);
or U18267 (N_18267,N_18133,N_18120);
nor U18268 (N_18268,N_18029,N_18065);
or U18269 (N_18269,N_18160,N_18215);
nor U18270 (N_18270,N_18169,N_18070);
nor U18271 (N_18271,N_18173,N_18137);
and U18272 (N_18272,N_18038,N_18162);
xnor U18273 (N_18273,N_18249,N_18017);
or U18274 (N_18274,N_18243,N_18074);
nor U18275 (N_18275,N_18163,N_18217);
or U18276 (N_18276,N_18122,N_18049);
nand U18277 (N_18277,N_18116,N_18112);
xnor U18278 (N_18278,N_18039,N_18033);
nor U18279 (N_18279,N_18242,N_18203);
and U18280 (N_18280,N_18090,N_18007);
nor U18281 (N_18281,N_18199,N_18062);
nand U18282 (N_18282,N_18011,N_18015);
xnor U18283 (N_18283,N_18107,N_18000);
nor U18284 (N_18284,N_18176,N_18059);
nand U18285 (N_18285,N_18114,N_18178);
nor U18286 (N_18286,N_18246,N_18105);
or U18287 (N_18287,N_18244,N_18170);
nor U18288 (N_18288,N_18096,N_18231);
nor U18289 (N_18289,N_18190,N_18050);
nor U18290 (N_18290,N_18241,N_18075);
xnor U18291 (N_18291,N_18110,N_18094);
and U18292 (N_18292,N_18027,N_18024);
and U18293 (N_18293,N_18206,N_18073);
and U18294 (N_18294,N_18078,N_18194);
nor U18295 (N_18295,N_18181,N_18135);
or U18296 (N_18296,N_18210,N_18019);
nand U18297 (N_18297,N_18184,N_18003);
and U18298 (N_18298,N_18082,N_18143);
xor U18299 (N_18299,N_18016,N_18117);
nor U18300 (N_18300,N_18060,N_18076);
nor U18301 (N_18301,N_18141,N_18155);
nor U18302 (N_18302,N_18026,N_18159);
nor U18303 (N_18303,N_18102,N_18113);
nand U18304 (N_18304,N_18175,N_18108);
xor U18305 (N_18305,N_18247,N_18161);
nor U18306 (N_18306,N_18168,N_18054);
nor U18307 (N_18307,N_18109,N_18131);
or U18308 (N_18308,N_18052,N_18077);
and U18309 (N_18309,N_18202,N_18232);
xnor U18310 (N_18310,N_18086,N_18042);
or U18311 (N_18311,N_18187,N_18130);
nor U18312 (N_18312,N_18097,N_18153);
and U18313 (N_18313,N_18058,N_18166);
nor U18314 (N_18314,N_18069,N_18180);
or U18315 (N_18315,N_18028,N_18118);
nand U18316 (N_18316,N_18010,N_18089);
xor U18317 (N_18317,N_18132,N_18124);
nor U18318 (N_18318,N_18218,N_18088);
or U18319 (N_18319,N_18068,N_18225);
or U18320 (N_18320,N_18193,N_18136);
or U18321 (N_18321,N_18195,N_18005);
or U18322 (N_18322,N_18044,N_18071);
or U18323 (N_18323,N_18126,N_18036);
nor U18324 (N_18324,N_18087,N_18013);
nand U18325 (N_18325,N_18191,N_18030);
nand U18326 (N_18326,N_18021,N_18081);
xnor U18327 (N_18327,N_18008,N_18208);
and U18328 (N_18328,N_18098,N_18222);
nand U18329 (N_18329,N_18085,N_18197);
and U18330 (N_18330,N_18158,N_18205);
or U18331 (N_18331,N_18129,N_18214);
and U18332 (N_18332,N_18034,N_18200);
nand U18333 (N_18333,N_18020,N_18228);
nand U18334 (N_18334,N_18220,N_18140);
nor U18335 (N_18335,N_18240,N_18224);
nand U18336 (N_18336,N_18235,N_18183);
and U18337 (N_18337,N_18025,N_18032);
and U18338 (N_18338,N_18207,N_18121);
nand U18339 (N_18339,N_18099,N_18152);
or U18340 (N_18340,N_18154,N_18157);
xnor U18341 (N_18341,N_18002,N_18031);
or U18342 (N_18342,N_18092,N_18023);
xnor U18343 (N_18343,N_18041,N_18156);
nor U18344 (N_18344,N_18022,N_18103);
xor U18345 (N_18345,N_18201,N_18233);
and U18346 (N_18346,N_18125,N_18227);
nor U18347 (N_18347,N_18151,N_18245);
and U18348 (N_18348,N_18192,N_18093);
nor U18349 (N_18349,N_18047,N_18186);
xnor U18350 (N_18350,N_18018,N_18229);
or U18351 (N_18351,N_18051,N_18012);
or U18352 (N_18352,N_18147,N_18046);
or U18353 (N_18353,N_18179,N_18067);
nand U18354 (N_18354,N_18040,N_18138);
and U18355 (N_18355,N_18234,N_18048);
nor U18356 (N_18356,N_18216,N_18055);
nand U18357 (N_18357,N_18146,N_18064);
and U18358 (N_18358,N_18196,N_18223);
xor U18359 (N_18359,N_18101,N_18072);
and U18360 (N_18360,N_18037,N_18111);
nand U18361 (N_18361,N_18188,N_18212);
nand U18362 (N_18362,N_18134,N_18035);
xnor U18363 (N_18363,N_18174,N_18230);
xnor U18364 (N_18364,N_18083,N_18128);
and U18365 (N_18365,N_18219,N_18119);
and U18366 (N_18366,N_18115,N_18091);
xnor U18367 (N_18367,N_18172,N_18100);
and U18368 (N_18368,N_18139,N_18053);
xnor U18369 (N_18369,N_18171,N_18177);
and U18370 (N_18370,N_18123,N_18043);
nor U18371 (N_18371,N_18204,N_18106);
xnor U18372 (N_18372,N_18145,N_18001);
nand U18373 (N_18373,N_18189,N_18238);
or U18374 (N_18374,N_18248,N_18237);
and U18375 (N_18375,N_18207,N_18137);
xnor U18376 (N_18376,N_18215,N_18141);
xor U18377 (N_18377,N_18163,N_18136);
or U18378 (N_18378,N_18149,N_18216);
xor U18379 (N_18379,N_18127,N_18015);
xnor U18380 (N_18380,N_18247,N_18097);
and U18381 (N_18381,N_18021,N_18209);
nor U18382 (N_18382,N_18025,N_18045);
nor U18383 (N_18383,N_18065,N_18173);
xnor U18384 (N_18384,N_18149,N_18201);
and U18385 (N_18385,N_18013,N_18110);
nor U18386 (N_18386,N_18197,N_18096);
or U18387 (N_18387,N_18245,N_18087);
xnor U18388 (N_18388,N_18059,N_18118);
xnor U18389 (N_18389,N_18059,N_18135);
nor U18390 (N_18390,N_18176,N_18025);
nand U18391 (N_18391,N_18095,N_18130);
or U18392 (N_18392,N_18095,N_18021);
and U18393 (N_18393,N_18004,N_18017);
nand U18394 (N_18394,N_18136,N_18114);
nor U18395 (N_18395,N_18127,N_18139);
nand U18396 (N_18396,N_18105,N_18078);
and U18397 (N_18397,N_18067,N_18182);
or U18398 (N_18398,N_18177,N_18215);
nand U18399 (N_18399,N_18103,N_18088);
and U18400 (N_18400,N_18247,N_18203);
nor U18401 (N_18401,N_18083,N_18226);
nor U18402 (N_18402,N_18026,N_18248);
xor U18403 (N_18403,N_18140,N_18187);
xor U18404 (N_18404,N_18160,N_18126);
nand U18405 (N_18405,N_18236,N_18024);
or U18406 (N_18406,N_18081,N_18229);
nor U18407 (N_18407,N_18176,N_18033);
nand U18408 (N_18408,N_18021,N_18016);
nand U18409 (N_18409,N_18246,N_18056);
nor U18410 (N_18410,N_18216,N_18182);
xor U18411 (N_18411,N_18073,N_18150);
xor U18412 (N_18412,N_18073,N_18207);
nand U18413 (N_18413,N_18106,N_18123);
nand U18414 (N_18414,N_18190,N_18087);
xor U18415 (N_18415,N_18091,N_18192);
and U18416 (N_18416,N_18182,N_18021);
nand U18417 (N_18417,N_18186,N_18142);
and U18418 (N_18418,N_18000,N_18021);
or U18419 (N_18419,N_18153,N_18152);
xor U18420 (N_18420,N_18245,N_18130);
nor U18421 (N_18421,N_18168,N_18159);
or U18422 (N_18422,N_18165,N_18107);
nand U18423 (N_18423,N_18160,N_18060);
nor U18424 (N_18424,N_18019,N_18154);
nand U18425 (N_18425,N_18096,N_18069);
nor U18426 (N_18426,N_18096,N_18223);
xnor U18427 (N_18427,N_18202,N_18089);
xnor U18428 (N_18428,N_18094,N_18231);
xor U18429 (N_18429,N_18083,N_18241);
xor U18430 (N_18430,N_18077,N_18203);
or U18431 (N_18431,N_18074,N_18209);
and U18432 (N_18432,N_18052,N_18043);
xor U18433 (N_18433,N_18092,N_18226);
and U18434 (N_18434,N_18197,N_18003);
xor U18435 (N_18435,N_18021,N_18012);
or U18436 (N_18436,N_18047,N_18042);
nand U18437 (N_18437,N_18003,N_18109);
nand U18438 (N_18438,N_18157,N_18124);
nor U18439 (N_18439,N_18044,N_18040);
or U18440 (N_18440,N_18053,N_18108);
or U18441 (N_18441,N_18162,N_18201);
nor U18442 (N_18442,N_18187,N_18117);
nand U18443 (N_18443,N_18035,N_18083);
and U18444 (N_18444,N_18162,N_18145);
or U18445 (N_18445,N_18024,N_18116);
nand U18446 (N_18446,N_18000,N_18003);
nor U18447 (N_18447,N_18031,N_18172);
xnor U18448 (N_18448,N_18021,N_18110);
xor U18449 (N_18449,N_18139,N_18217);
xor U18450 (N_18450,N_18247,N_18010);
and U18451 (N_18451,N_18188,N_18205);
or U18452 (N_18452,N_18194,N_18167);
and U18453 (N_18453,N_18164,N_18052);
or U18454 (N_18454,N_18189,N_18166);
nor U18455 (N_18455,N_18039,N_18030);
or U18456 (N_18456,N_18083,N_18205);
nor U18457 (N_18457,N_18190,N_18234);
and U18458 (N_18458,N_18020,N_18135);
nor U18459 (N_18459,N_18209,N_18117);
xor U18460 (N_18460,N_18235,N_18140);
or U18461 (N_18461,N_18144,N_18084);
xnor U18462 (N_18462,N_18096,N_18021);
or U18463 (N_18463,N_18066,N_18169);
nor U18464 (N_18464,N_18094,N_18184);
xor U18465 (N_18465,N_18212,N_18020);
and U18466 (N_18466,N_18209,N_18203);
or U18467 (N_18467,N_18181,N_18049);
xnor U18468 (N_18468,N_18181,N_18239);
and U18469 (N_18469,N_18143,N_18219);
and U18470 (N_18470,N_18141,N_18147);
and U18471 (N_18471,N_18022,N_18155);
nor U18472 (N_18472,N_18028,N_18224);
and U18473 (N_18473,N_18147,N_18041);
nand U18474 (N_18474,N_18214,N_18031);
or U18475 (N_18475,N_18110,N_18145);
or U18476 (N_18476,N_18141,N_18088);
or U18477 (N_18477,N_18079,N_18108);
nor U18478 (N_18478,N_18217,N_18075);
and U18479 (N_18479,N_18102,N_18157);
nand U18480 (N_18480,N_18243,N_18229);
and U18481 (N_18481,N_18095,N_18124);
nand U18482 (N_18482,N_18003,N_18058);
nand U18483 (N_18483,N_18111,N_18101);
nor U18484 (N_18484,N_18107,N_18049);
and U18485 (N_18485,N_18160,N_18004);
xnor U18486 (N_18486,N_18092,N_18028);
nand U18487 (N_18487,N_18068,N_18019);
nand U18488 (N_18488,N_18156,N_18229);
and U18489 (N_18489,N_18095,N_18070);
and U18490 (N_18490,N_18043,N_18051);
and U18491 (N_18491,N_18040,N_18172);
nor U18492 (N_18492,N_18113,N_18149);
nor U18493 (N_18493,N_18105,N_18069);
or U18494 (N_18494,N_18073,N_18009);
nand U18495 (N_18495,N_18212,N_18028);
xnor U18496 (N_18496,N_18212,N_18177);
and U18497 (N_18497,N_18038,N_18173);
xor U18498 (N_18498,N_18159,N_18142);
and U18499 (N_18499,N_18121,N_18246);
nor U18500 (N_18500,N_18301,N_18250);
nand U18501 (N_18501,N_18499,N_18324);
nor U18502 (N_18502,N_18497,N_18406);
and U18503 (N_18503,N_18318,N_18412);
and U18504 (N_18504,N_18458,N_18260);
and U18505 (N_18505,N_18253,N_18321);
or U18506 (N_18506,N_18465,N_18363);
and U18507 (N_18507,N_18446,N_18405);
or U18508 (N_18508,N_18258,N_18400);
and U18509 (N_18509,N_18390,N_18366);
nor U18510 (N_18510,N_18474,N_18372);
nor U18511 (N_18511,N_18352,N_18408);
and U18512 (N_18512,N_18349,N_18492);
nand U18513 (N_18513,N_18344,N_18259);
xor U18514 (N_18514,N_18384,N_18308);
xnor U18515 (N_18515,N_18304,N_18418);
nor U18516 (N_18516,N_18317,N_18359);
xor U18517 (N_18517,N_18299,N_18307);
and U18518 (N_18518,N_18353,N_18411);
nor U18519 (N_18519,N_18498,N_18319);
nor U18520 (N_18520,N_18450,N_18455);
or U18521 (N_18521,N_18402,N_18448);
nand U18522 (N_18522,N_18479,N_18496);
nor U18523 (N_18523,N_18378,N_18251);
nand U18524 (N_18524,N_18495,N_18486);
and U18525 (N_18525,N_18334,N_18470);
nor U18526 (N_18526,N_18261,N_18434);
nor U18527 (N_18527,N_18296,N_18272);
nor U18528 (N_18528,N_18427,N_18429);
nand U18529 (N_18529,N_18303,N_18395);
xor U18530 (N_18530,N_18289,N_18300);
xnor U18531 (N_18531,N_18329,N_18396);
and U18532 (N_18532,N_18462,N_18494);
nor U18533 (N_18533,N_18285,N_18331);
nor U18534 (N_18534,N_18435,N_18466);
nor U18535 (N_18535,N_18432,N_18481);
nor U18536 (N_18536,N_18404,N_18274);
and U18537 (N_18537,N_18282,N_18381);
nor U18538 (N_18538,N_18428,N_18439);
or U18539 (N_18539,N_18413,N_18312);
nand U18540 (N_18540,N_18467,N_18419);
and U18541 (N_18541,N_18364,N_18277);
nor U18542 (N_18542,N_18417,N_18382);
or U18543 (N_18543,N_18314,N_18255);
or U18544 (N_18544,N_18460,N_18355);
and U18545 (N_18545,N_18431,N_18362);
nand U18546 (N_18546,N_18383,N_18473);
or U18547 (N_18547,N_18371,N_18468);
nor U18548 (N_18548,N_18367,N_18335);
nand U18549 (N_18549,N_18409,N_18280);
xnor U18550 (N_18550,N_18488,N_18295);
or U18551 (N_18551,N_18451,N_18283);
and U18552 (N_18552,N_18420,N_18323);
xnor U18553 (N_18553,N_18273,N_18341);
nor U18554 (N_18554,N_18291,N_18373);
or U18555 (N_18555,N_18487,N_18471);
nand U18556 (N_18556,N_18370,N_18430);
nor U18557 (N_18557,N_18410,N_18310);
or U18558 (N_18558,N_18385,N_18423);
and U18559 (N_18559,N_18313,N_18340);
nand U18560 (N_18560,N_18374,N_18476);
xor U18561 (N_18561,N_18437,N_18493);
nor U18562 (N_18562,N_18337,N_18397);
xnor U18563 (N_18563,N_18266,N_18325);
and U18564 (N_18564,N_18414,N_18424);
or U18565 (N_18565,N_18482,N_18284);
xor U18566 (N_18566,N_18483,N_18354);
or U18567 (N_18567,N_18415,N_18315);
nand U18568 (N_18568,N_18421,N_18328);
xnor U18569 (N_18569,N_18464,N_18403);
nor U18570 (N_18570,N_18452,N_18268);
or U18571 (N_18571,N_18262,N_18254);
nor U18572 (N_18572,N_18379,N_18338);
nand U18573 (N_18573,N_18269,N_18438);
or U18574 (N_18574,N_18368,N_18456);
nor U18575 (N_18575,N_18477,N_18387);
or U18576 (N_18576,N_18288,N_18394);
and U18577 (N_18577,N_18270,N_18389);
xnor U18578 (N_18578,N_18440,N_18339);
nor U18579 (N_18579,N_18267,N_18290);
and U18580 (N_18580,N_18399,N_18447);
xnor U18581 (N_18581,N_18357,N_18422);
nand U18582 (N_18582,N_18436,N_18441);
nand U18583 (N_18583,N_18398,N_18469);
xnor U18584 (N_18584,N_18263,N_18459);
nand U18585 (N_18585,N_18375,N_18305);
xnor U18586 (N_18586,N_18391,N_18453);
and U18587 (N_18587,N_18484,N_18252);
xor U18588 (N_18588,N_18311,N_18297);
or U18589 (N_18589,N_18490,N_18345);
xnor U18590 (N_18590,N_18278,N_18365);
nand U18591 (N_18591,N_18347,N_18376);
nor U18592 (N_18592,N_18480,N_18326);
nor U18593 (N_18593,N_18377,N_18392);
and U18594 (N_18594,N_18265,N_18433);
nor U18595 (N_18595,N_18360,N_18287);
xnor U18596 (N_18596,N_18457,N_18401);
or U18597 (N_18597,N_18271,N_18358);
nor U18598 (N_18598,N_18425,N_18346);
nor U18599 (N_18599,N_18380,N_18361);
or U18600 (N_18600,N_18463,N_18416);
nor U18601 (N_18601,N_18336,N_18461);
and U18602 (N_18602,N_18333,N_18454);
or U18603 (N_18603,N_18472,N_18276);
and U18604 (N_18604,N_18327,N_18351);
nand U18605 (N_18605,N_18306,N_18275);
nor U18606 (N_18606,N_18302,N_18407);
or U18607 (N_18607,N_18475,N_18292);
xnor U18608 (N_18608,N_18264,N_18426);
and U18609 (N_18609,N_18309,N_18443);
nor U18610 (N_18610,N_18316,N_18279);
nor U18611 (N_18611,N_18485,N_18332);
xnor U18612 (N_18612,N_18489,N_18442);
or U18613 (N_18613,N_18256,N_18386);
xnor U18614 (N_18614,N_18342,N_18393);
xnor U18615 (N_18615,N_18293,N_18320);
xnor U18616 (N_18616,N_18388,N_18491);
xnor U18617 (N_18617,N_18281,N_18445);
nand U18618 (N_18618,N_18356,N_18348);
nor U18619 (N_18619,N_18257,N_18286);
nand U18620 (N_18620,N_18350,N_18330);
xor U18621 (N_18621,N_18298,N_18369);
xnor U18622 (N_18622,N_18294,N_18322);
xnor U18623 (N_18623,N_18444,N_18478);
and U18624 (N_18624,N_18449,N_18343);
nand U18625 (N_18625,N_18264,N_18479);
and U18626 (N_18626,N_18368,N_18455);
nor U18627 (N_18627,N_18427,N_18350);
and U18628 (N_18628,N_18465,N_18336);
xor U18629 (N_18629,N_18473,N_18326);
xnor U18630 (N_18630,N_18357,N_18276);
nand U18631 (N_18631,N_18285,N_18375);
and U18632 (N_18632,N_18448,N_18264);
or U18633 (N_18633,N_18374,N_18470);
xnor U18634 (N_18634,N_18405,N_18425);
xnor U18635 (N_18635,N_18451,N_18461);
xor U18636 (N_18636,N_18381,N_18439);
xor U18637 (N_18637,N_18317,N_18428);
or U18638 (N_18638,N_18320,N_18449);
nor U18639 (N_18639,N_18250,N_18489);
nand U18640 (N_18640,N_18385,N_18298);
xor U18641 (N_18641,N_18375,N_18411);
nor U18642 (N_18642,N_18377,N_18345);
and U18643 (N_18643,N_18319,N_18384);
nand U18644 (N_18644,N_18310,N_18460);
and U18645 (N_18645,N_18404,N_18475);
nor U18646 (N_18646,N_18266,N_18406);
or U18647 (N_18647,N_18274,N_18435);
and U18648 (N_18648,N_18284,N_18414);
nand U18649 (N_18649,N_18394,N_18341);
xor U18650 (N_18650,N_18415,N_18309);
xor U18651 (N_18651,N_18335,N_18481);
xor U18652 (N_18652,N_18257,N_18267);
nor U18653 (N_18653,N_18390,N_18274);
nand U18654 (N_18654,N_18398,N_18478);
and U18655 (N_18655,N_18417,N_18479);
and U18656 (N_18656,N_18489,N_18325);
nor U18657 (N_18657,N_18301,N_18370);
or U18658 (N_18658,N_18415,N_18422);
and U18659 (N_18659,N_18400,N_18430);
nor U18660 (N_18660,N_18410,N_18277);
xor U18661 (N_18661,N_18301,N_18403);
xnor U18662 (N_18662,N_18490,N_18467);
nand U18663 (N_18663,N_18301,N_18458);
and U18664 (N_18664,N_18263,N_18352);
and U18665 (N_18665,N_18487,N_18373);
xnor U18666 (N_18666,N_18366,N_18409);
nand U18667 (N_18667,N_18356,N_18423);
or U18668 (N_18668,N_18466,N_18426);
nand U18669 (N_18669,N_18416,N_18473);
nand U18670 (N_18670,N_18348,N_18274);
xor U18671 (N_18671,N_18399,N_18277);
xor U18672 (N_18672,N_18358,N_18260);
nand U18673 (N_18673,N_18451,N_18475);
xnor U18674 (N_18674,N_18393,N_18323);
or U18675 (N_18675,N_18267,N_18438);
or U18676 (N_18676,N_18414,N_18397);
nand U18677 (N_18677,N_18464,N_18336);
nor U18678 (N_18678,N_18376,N_18423);
xnor U18679 (N_18679,N_18433,N_18282);
nand U18680 (N_18680,N_18354,N_18437);
nand U18681 (N_18681,N_18297,N_18458);
or U18682 (N_18682,N_18343,N_18403);
and U18683 (N_18683,N_18334,N_18300);
nand U18684 (N_18684,N_18317,N_18430);
nor U18685 (N_18685,N_18473,N_18470);
or U18686 (N_18686,N_18372,N_18441);
and U18687 (N_18687,N_18400,N_18294);
xnor U18688 (N_18688,N_18358,N_18361);
and U18689 (N_18689,N_18382,N_18366);
and U18690 (N_18690,N_18424,N_18323);
xor U18691 (N_18691,N_18353,N_18459);
nor U18692 (N_18692,N_18363,N_18299);
xnor U18693 (N_18693,N_18347,N_18323);
xor U18694 (N_18694,N_18252,N_18496);
nand U18695 (N_18695,N_18447,N_18349);
nor U18696 (N_18696,N_18467,N_18445);
xnor U18697 (N_18697,N_18417,N_18409);
nand U18698 (N_18698,N_18408,N_18266);
xor U18699 (N_18699,N_18349,N_18439);
nand U18700 (N_18700,N_18333,N_18498);
nand U18701 (N_18701,N_18320,N_18403);
nor U18702 (N_18702,N_18323,N_18466);
or U18703 (N_18703,N_18489,N_18404);
nand U18704 (N_18704,N_18328,N_18279);
and U18705 (N_18705,N_18256,N_18280);
or U18706 (N_18706,N_18261,N_18279);
or U18707 (N_18707,N_18481,N_18332);
and U18708 (N_18708,N_18377,N_18268);
xor U18709 (N_18709,N_18384,N_18314);
xor U18710 (N_18710,N_18438,N_18412);
xor U18711 (N_18711,N_18270,N_18348);
and U18712 (N_18712,N_18344,N_18359);
or U18713 (N_18713,N_18452,N_18254);
or U18714 (N_18714,N_18321,N_18487);
or U18715 (N_18715,N_18365,N_18300);
nor U18716 (N_18716,N_18342,N_18450);
or U18717 (N_18717,N_18499,N_18455);
or U18718 (N_18718,N_18338,N_18485);
and U18719 (N_18719,N_18297,N_18333);
nor U18720 (N_18720,N_18312,N_18363);
nand U18721 (N_18721,N_18254,N_18371);
nor U18722 (N_18722,N_18319,N_18489);
nand U18723 (N_18723,N_18358,N_18424);
nand U18724 (N_18724,N_18308,N_18333);
xor U18725 (N_18725,N_18444,N_18347);
nor U18726 (N_18726,N_18453,N_18379);
xnor U18727 (N_18727,N_18252,N_18490);
nor U18728 (N_18728,N_18485,N_18437);
and U18729 (N_18729,N_18477,N_18264);
nor U18730 (N_18730,N_18359,N_18275);
nand U18731 (N_18731,N_18280,N_18450);
and U18732 (N_18732,N_18354,N_18456);
and U18733 (N_18733,N_18381,N_18335);
and U18734 (N_18734,N_18338,N_18307);
and U18735 (N_18735,N_18414,N_18364);
nor U18736 (N_18736,N_18340,N_18394);
xor U18737 (N_18737,N_18309,N_18465);
nand U18738 (N_18738,N_18387,N_18285);
and U18739 (N_18739,N_18483,N_18457);
nand U18740 (N_18740,N_18398,N_18425);
xor U18741 (N_18741,N_18290,N_18319);
and U18742 (N_18742,N_18494,N_18273);
xor U18743 (N_18743,N_18390,N_18427);
xor U18744 (N_18744,N_18434,N_18376);
xnor U18745 (N_18745,N_18333,N_18450);
nor U18746 (N_18746,N_18404,N_18277);
xor U18747 (N_18747,N_18326,N_18310);
or U18748 (N_18748,N_18387,N_18281);
and U18749 (N_18749,N_18386,N_18454);
xor U18750 (N_18750,N_18541,N_18613);
nand U18751 (N_18751,N_18586,N_18723);
and U18752 (N_18752,N_18601,N_18661);
or U18753 (N_18753,N_18637,N_18608);
nand U18754 (N_18754,N_18571,N_18547);
xnor U18755 (N_18755,N_18669,N_18719);
nor U18756 (N_18756,N_18698,N_18500);
or U18757 (N_18757,N_18663,N_18730);
nand U18758 (N_18758,N_18643,N_18622);
nand U18759 (N_18759,N_18697,N_18551);
nor U18760 (N_18760,N_18685,N_18548);
xor U18761 (N_18761,N_18693,N_18745);
and U18762 (N_18762,N_18516,N_18529);
nand U18763 (N_18763,N_18673,N_18714);
and U18764 (N_18764,N_18641,N_18596);
xor U18765 (N_18765,N_18528,N_18536);
xor U18766 (N_18766,N_18720,N_18672);
nand U18767 (N_18767,N_18599,N_18653);
and U18768 (N_18768,N_18503,N_18743);
or U18769 (N_18769,N_18704,N_18515);
and U18770 (N_18770,N_18690,N_18565);
and U18771 (N_18771,N_18522,N_18718);
or U18772 (N_18772,N_18629,N_18615);
or U18773 (N_18773,N_18568,N_18686);
nor U18774 (N_18774,N_18501,N_18559);
xor U18775 (N_18775,N_18736,N_18646);
and U18776 (N_18776,N_18741,N_18594);
or U18777 (N_18777,N_18550,N_18620);
xor U18778 (N_18778,N_18530,N_18569);
nand U18779 (N_18779,N_18724,N_18737);
xnor U18780 (N_18780,N_18694,N_18538);
nor U18781 (N_18781,N_18510,N_18614);
nor U18782 (N_18782,N_18593,N_18512);
nand U18783 (N_18783,N_18540,N_18519);
xor U18784 (N_18784,N_18664,N_18578);
nor U18785 (N_18785,N_18731,N_18649);
nor U18786 (N_18786,N_18572,N_18732);
or U18787 (N_18787,N_18554,N_18675);
or U18788 (N_18788,N_18577,N_18710);
nand U18789 (N_18789,N_18639,N_18648);
xor U18790 (N_18790,N_18729,N_18716);
xor U18791 (N_18791,N_18584,N_18744);
xor U18792 (N_18792,N_18630,N_18651);
nand U18793 (N_18793,N_18527,N_18705);
nand U18794 (N_18794,N_18631,N_18676);
and U18795 (N_18795,N_18655,N_18604);
nand U18796 (N_18796,N_18722,N_18588);
or U18797 (N_18797,N_18592,N_18699);
or U18798 (N_18798,N_18532,N_18702);
nor U18799 (N_18799,N_18612,N_18727);
and U18800 (N_18800,N_18553,N_18746);
and U18801 (N_18801,N_18533,N_18667);
and U18802 (N_18802,N_18566,N_18678);
nand U18803 (N_18803,N_18508,N_18658);
or U18804 (N_18804,N_18682,N_18721);
xnor U18805 (N_18805,N_18597,N_18634);
nor U18806 (N_18806,N_18602,N_18543);
nand U18807 (N_18807,N_18591,N_18660);
nand U18808 (N_18808,N_18711,N_18657);
or U18809 (N_18809,N_18726,N_18681);
and U18810 (N_18810,N_18645,N_18638);
and U18811 (N_18811,N_18507,N_18647);
nor U18812 (N_18812,N_18671,N_18742);
nand U18813 (N_18813,N_18740,N_18707);
or U18814 (N_18814,N_18625,N_18627);
xor U18815 (N_18815,N_18689,N_18546);
and U18816 (N_18816,N_18582,N_18712);
nor U18817 (N_18817,N_18650,N_18609);
xnor U18818 (N_18818,N_18652,N_18713);
nor U18819 (N_18819,N_18636,N_18688);
xnor U18820 (N_18820,N_18526,N_18715);
nor U18821 (N_18821,N_18623,N_18610);
xor U18822 (N_18822,N_18668,N_18537);
or U18823 (N_18823,N_18545,N_18574);
or U18824 (N_18824,N_18735,N_18656);
nand U18825 (N_18825,N_18747,N_18703);
and U18826 (N_18826,N_18573,N_18587);
xor U18827 (N_18827,N_18595,N_18562);
or U18828 (N_18828,N_18684,N_18534);
nor U18829 (N_18829,N_18692,N_18738);
nor U18830 (N_18830,N_18695,N_18517);
nor U18831 (N_18831,N_18556,N_18670);
nand U18832 (N_18832,N_18701,N_18600);
or U18833 (N_18833,N_18539,N_18628);
xnor U18834 (N_18834,N_18520,N_18581);
nor U18835 (N_18835,N_18531,N_18644);
and U18836 (N_18836,N_18576,N_18624);
nor U18837 (N_18837,N_18560,N_18514);
nor U18838 (N_18838,N_18666,N_18677);
or U18839 (N_18839,N_18525,N_18640);
and U18840 (N_18840,N_18563,N_18606);
or U18841 (N_18841,N_18605,N_18617);
xnor U18842 (N_18842,N_18632,N_18567);
nor U18843 (N_18843,N_18509,N_18709);
nand U18844 (N_18844,N_18748,N_18683);
xnor U18845 (N_18845,N_18662,N_18580);
and U18846 (N_18846,N_18626,N_18749);
xor U18847 (N_18847,N_18570,N_18619);
or U18848 (N_18848,N_18679,N_18603);
and U18849 (N_18849,N_18579,N_18523);
xor U18850 (N_18850,N_18505,N_18558);
nor U18851 (N_18851,N_18621,N_18552);
nand U18852 (N_18852,N_18585,N_18542);
nor U18853 (N_18853,N_18524,N_18589);
xor U18854 (N_18854,N_18511,N_18502);
nand U18855 (N_18855,N_18717,N_18708);
xnor U18856 (N_18856,N_18590,N_18564);
and U18857 (N_18857,N_18607,N_18544);
or U18858 (N_18858,N_18555,N_18506);
nor U18859 (N_18859,N_18700,N_18518);
and U18860 (N_18860,N_18642,N_18674);
nor U18861 (N_18861,N_18535,N_18504);
or U18862 (N_18862,N_18654,N_18734);
or U18863 (N_18863,N_18549,N_18557);
or U18864 (N_18864,N_18728,N_18659);
or U18865 (N_18865,N_18706,N_18635);
nand U18866 (N_18866,N_18583,N_18575);
or U18867 (N_18867,N_18513,N_18665);
and U18868 (N_18868,N_18739,N_18691);
and U18869 (N_18869,N_18611,N_18733);
xor U18870 (N_18870,N_18521,N_18687);
xor U18871 (N_18871,N_18725,N_18680);
xnor U18872 (N_18872,N_18618,N_18598);
nor U18873 (N_18873,N_18561,N_18696);
nor U18874 (N_18874,N_18616,N_18633);
xnor U18875 (N_18875,N_18543,N_18542);
xor U18876 (N_18876,N_18625,N_18676);
nand U18877 (N_18877,N_18748,N_18653);
nand U18878 (N_18878,N_18589,N_18731);
and U18879 (N_18879,N_18613,N_18637);
nor U18880 (N_18880,N_18736,N_18692);
xnor U18881 (N_18881,N_18501,N_18723);
or U18882 (N_18882,N_18701,N_18560);
and U18883 (N_18883,N_18568,N_18593);
nand U18884 (N_18884,N_18590,N_18542);
nor U18885 (N_18885,N_18692,N_18530);
or U18886 (N_18886,N_18700,N_18573);
nor U18887 (N_18887,N_18628,N_18589);
xnor U18888 (N_18888,N_18529,N_18517);
nand U18889 (N_18889,N_18598,N_18540);
or U18890 (N_18890,N_18568,N_18612);
nor U18891 (N_18891,N_18709,N_18686);
xor U18892 (N_18892,N_18719,N_18716);
nor U18893 (N_18893,N_18724,N_18708);
xor U18894 (N_18894,N_18561,N_18569);
nor U18895 (N_18895,N_18547,N_18505);
nor U18896 (N_18896,N_18597,N_18594);
xor U18897 (N_18897,N_18604,N_18682);
xor U18898 (N_18898,N_18710,N_18592);
or U18899 (N_18899,N_18592,N_18674);
nor U18900 (N_18900,N_18502,N_18562);
xor U18901 (N_18901,N_18659,N_18748);
or U18902 (N_18902,N_18646,N_18511);
and U18903 (N_18903,N_18706,N_18731);
and U18904 (N_18904,N_18691,N_18669);
nand U18905 (N_18905,N_18595,N_18552);
xor U18906 (N_18906,N_18560,N_18691);
nand U18907 (N_18907,N_18543,N_18501);
xnor U18908 (N_18908,N_18702,N_18553);
and U18909 (N_18909,N_18701,N_18577);
or U18910 (N_18910,N_18697,N_18602);
or U18911 (N_18911,N_18660,N_18512);
nand U18912 (N_18912,N_18617,N_18567);
or U18913 (N_18913,N_18694,N_18640);
nor U18914 (N_18914,N_18547,N_18564);
nor U18915 (N_18915,N_18668,N_18702);
nor U18916 (N_18916,N_18588,N_18542);
nand U18917 (N_18917,N_18712,N_18692);
xor U18918 (N_18918,N_18706,N_18701);
nand U18919 (N_18919,N_18666,N_18735);
and U18920 (N_18920,N_18501,N_18632);
xor U18921 (N_18921,N_18539,N_18715);
or U18922 (N_18922,N_18598,N_18505);
and U18923 (N_18923,N_18626,N_18515);
nand U18924 (N_18924,N_18710,N_18679);
xor U18925 (N_18925,N_18709,N_18623);
xor U18926 (N_18926,N_18622,N_18586);
nand U18927 (N_18927,N_18733,N_18720);
and U18928 (N_18928,N_18597,N_18599);
and U18929 (N_18929,N_18712,N_18739);
nor U18930 (N_18930,N_18676,N_18717);
xnor U18931 (N_18931,N_18613,N_18536);
nand U18932 (N_18932,N_18507,N_18581);
and U18933 (N_18933,N_18639,N_18739);
nor U18934 (N_18934,N_18517,N_18645);
nand U18935 (N_18935,N_18523,N_18577);
nor U18936 (N_18936,N_18688,N_18523);
or U18937 (N_18937,N_18571,N_18529);
or U18938 (N_18938,N_18520,N_18647);
nor U18939 (N_18939,N_18528,N_18560);
and U18940 (N_18940,N_18722,N_18744);
nor U18941 (N_18941,N_18650,N_18503);
xor U18942 (N_18942,N_18613,N_18696);
xnor U18943 (N_18943,N_18577,N_18638);
and U18944 (N_18944,N_18563,N_18695);
and U18945 (N_18945,N_18728,N_18612);
and U18946 (N_18946,N_18724,N_18710);
xnor U18947 (N_18947,N_18610,N_18622);
nand U18948 (N_18948,N_18526,N_18632);
and U18949 (N_18949,N_18505,N_18513);
xnor U18950 (N_18950,N_18708,N_18561);
nor U18951 (N_18951,N_18513,N_18504);
nor U18952 (N_18952,N_18729,N_18600);
and U18953 (N_18953,N_18545,N_18725);
nand U18954 (N_18954,N_18603,N_18558);
xor U18955 (N_18955,N_18531,N_18563);
or U18956 (N_18956,N_18670,N_18601);
nand U18957 (N_18957,N_18585,N_18558);
and U18958 (N_18958,N_18662,N_18639);
nor U18959 (N_18959,N_18573,N_18704);
and U18960 (N_18960,N_18535,N_18660);
nor U18961 (N_18961,N_18567,N_18719);
xnor U18962 (N_18962,N_18586,N_18652);
or U18963 (N_18963,N_18538,N_18614);
nand U18964 (N_18964,N_18527,N_18600);
xor U18965 (N_18965,N_18742,N_18682);
nor U18966 (N_18966,N_18659,N_18532);
and U18967 (N_18967,N_18508,N_18554);
and U18968 (N_18968,N_18554,N_18542);
and U18969 (N_18969,N_18635,N_18584);
and U18970 (N_18970,N_18737,N_18555);
and U18971 (N_18971,N_18528,N_18621);
nor U18972 (N_18972,N_18539,N_18710);
nor U18973 (N_18973,N_18692,N_18634);
nand U18974 (N_18974,N_18631,N_18719);
and U18975 (N_18975,N_18704,N_18598);
and U18976 (N_18976,N_18664,N_18681);
or U18977 (N_18977,N_18565,N_18738);
nor U18978 (N_18978,N_18557,N_18544);
and U18979 (N_18979,N_18511,N_18677);
nand U18980 (N_18980,N_18697,N_18501);
xor U18981 (N_18981,N_18688,N_18639);
nand U18982 (N_18982,N_18575,N_18678);
nand U18983 (N_18983,N_18554,N_18532);
or U18984 (N_18984,N_18572,N_18561);
or U18985 (N_18985,N_18527,N_18590);
or U18986 (N_18986,N_18547,N_18577);
or U18987 (N_18987,N_18552,N_18669);
nand U18988 (N_18988,N_18655,N_18714);
or U18989 (N_18989,N_18564,N_18563);
xnor U18990 (N_18990,N_18532,N_18602);
and U18991 (N_18991,N_18736,N_18650);
or U18992 (N_18992,N_18744,N_18563);
and U18993 (N_18993,N_18648,N_18594);
and U18994 (N_18994,N_18652,N_18690);
or U18995 (N_18995,N_18715,N_18533);
nor U18996 (N_18996,N_18593,N_18723);
and U18997 (N_18997,N_18594,N_18513);
and U18998 (N_18998,N_18738,N_18647);
nand U18999 (N_18999,N_18714,N_18666);
and U19000 (N_19000,N_18969,N_18924);
and U19001 (N_19001,N_18794,N_18814);
nor U19002 (N_19002,N_18930,N_18764);
nand U19003 (N_19003,N_18988,N_18864);
nand U19004 (N_19004,N_18928,N_18855);
or U19005 (N_19005,N_18879,N_18753);
nor U19006 (N_19006,N_18972,N_18990);
or U19007 (N_19007,N_18922,N_18867);
nand U19008 (N_19008,N_18888,N_18929);
nand U19009 (N_19009,N_18925,N_18936);
and U19010 (N_19010,N_18992,N_18887);
or U19011 (N_19011,N_18996,N_18792);
and U19012 (N_19012,N_18954,N_18848);
nand U19013 (N_19013,N_18883,N_18907);
xnor U19014 (N_19014,N_18785,N_18806);
or U19015 (N_19015,N_18901,N_18881);
or U19016 (N_19016,N_18761,N_18896);
xnor U19017 (N_19017,N_18933,N_18800);
or U19018 (N_19018,N_18821,N_18766);
xnor U19019 (N_19019,N_18776,N_18885);
and U19020 (N_19020,N_18935,N_18754);
nor U19021 (N_19021,N_18921,N_18895);
xnor U19022 (N_19022,N_18805,N_18947);
and U19023 (N_19023,N_18750,N_18993);
and U19024 (N_19024,N_18917,N_18900);
nor U19025 (N_19025,N_18854,N_18859);
xnor U19026 (N_19026,N_18934,N_18875);
or U19027 (N_19027,N_18852,N_18932);
nor U19028 (N_19028,N_18845,N_18948);
xor U19029 (N_19029,N_18765,N_18967);
and U19030 (N_19030,N_18816,N_18989);
nand U19031 (N_19031,N_18832,N_18795);
or U19032 (N_19032,N_18828,N_18987);
or U19033 (N_19033,N_18944,N_18787);
xor U19034 (N_19034,N_18836,N_18973);
nand U19035 (N_19035,N_18910,N_18851);
nand U19036 (N_19036,N_18965,N_18906);
and U19037 (N_19037,N_18923,N_18760);
nand U19038 (N_19038,N_18798,N_18868);
xor U19039 (N_19039,N_18861,N_18818);
nand U19040 (N_19040,N_18916,N_18788);
nand U19041 (N_19041,N_18873,N_18931);
nor U19042 (N_19042,N_18860,N_18857);
and U19043 (N_19043,N_18941,N_18886);
nor U19044 (N_19044,N_18751,N_18943);
nand U19045 (N_19045,N_18770,N_18790);
nor U19046 (N_19046,N_18889,N_18915);
or U19047 (N_19047,N_18809,N_18983);
and U19048 (N_19048,N_18774,N_18909);
nand U19049 (N_19049,N_18768,N_18862);
nand U19050 (N_19050,N_18837,N_18802);
nor U19051 (N_19051,N_18866,N_18882);
and U19052 (N_19052,N_18956,N_18918);
xor U19053 (N_19053,N_18835,N_18884);
nor U19054 (N_19054,N_18926,N_18897);
and U19055 (N_19055,N_18796,N_18758);
nor U19056 (N_19056,N_18780,N_18949);
xnor U19057 (N_19057,N_18920,N_18913);
xor U19058 (N_19058,N_18998,N_18968);
or U19059 (N_19059,N_18976,N_18823);
nand U19060 (N_19060,N_18853,N_18964);
nor U19061 (N_19061,N_18871,N_18985);
nand U19062 (N_19062,N_18804,N_18986);
and U19063 (N_19063,N_18911,N_18946);
or U19064 (N_19064,N_18892,N_18902);
or U19065 (N_19065,N_18824,N_18789);
nor U19066 (N_19066,N_18812,N_18893);
nand U19067 (N_19067,N_18844,N_18908);
nand U19068 (N_19068,N_18995,N_18994);
nor U19069 (N_19069,N_18927,N_18865);
nand U19070 (N_19070,N_18957,N_18815);
nor U19071 (N_19071,N_18919,N_18863);
or U19072 (N_19072,N_18759,N_18830);
nand U19073 (N_19073,N_18803,N_18833);
xor U19074 (N_19074,N_18813,N_18834);
nand U19075 (N_19075,N_18962,N_18979);
xor U19076 (N_19076,N_18890,N_18783);
and U19077 (N_19077,N_18829,N_18793);
xor U19078 (N_19078,N_18756,N_18846);
xor U19079 (N_19079,N_18856,N_18869);
or U19080 (N_19080,N_18784,N_18843);
nand U19081 (N_19081,N_18963,N_18763);
nand U19082 (N_19082,N_18778,N_18914);
and U19083 (N_19083,N_18755,N_18945);
nand U19084 (N_19084,N_18905,N_18953);
nor U19085 (N_19085,N_18772,N_18959);
nor U19086 (N_19086,N_18781,N_18771);
xor U19087 (N_19087,N_18840,N_18773);
and U19088 (N_19088,N_18940,N_18971);
nand U19089 (N_19089,N_18899,N_18825);
or U19090 (N_19090,N_18894,N_18938);
nor U19091 (N_19091,N_18797,N_18842);
and U19092 (N_19092,N_18958,N_18975);
nand U19093 (N_19093,N_18966,N_18762);
xor U19094 (N_19094,N_18822,N_18999);
nor U19095 (N_19095,N_18937,N_18880);
nand U19096 (N_19096,N_18847,N_18752);
nand U19097 (N_19097,N_18810,N_18838);
and U19098 (N_19098,N_18876,N_18912);
or U19099 (N_19099,N_18974,N_18970);
xor U19100 (N_19100,N_18939,N_18826);
and U19101 (N_19101,N_18977,N_18978);
nor U19102 (N_19102,N_18841,N_18782);
and U19103 (N_19103,N_18819,N_18850);
or U19104 (N_19104,N_18801,N_18791);
xor U19105 (N_19105,N_18878,N_18942);
or U19106 (N_19106,N_18903,N_18769);
nor U19107 (N_19107,N_18799,N_18877);
or U19108 (N_19108,N_18997,N_18767);
nand U19109 (N_19109,N_18991,N_18980);
and U19110 (N_19110,N_18950,N_18898);
nor U19111 (N_19111,N_18858,N_18960);
and U19112 (N_19112,N_18904,N_18891);
xnor U19113 (N_19113,N_18811,N_18952);
xnor U19114 (N_19114,N_18870,N_18872);
xnor U19115 (N_19115,N_18839,N_18827);
nor U19116 (N_19116,N_18757,N_18786);
xnor U19117 (N_19117,N_18820,N_18951);
or U19118 (N_19118,N_18808,N_18982);
nor U19119 (N_19119,N_18984,N_18849);
xnor U19120 (N_19120,N_18779,N_18955);
xor U19121 (N_19121,N_18981,N_18961);
nor U19122 (N_19122,N_18775,N_18807);
nand U19123 (N_19123,N_18817,N_18777);
nor U19124 (N_19124,N_18831,N_18874);
and U19125 (N_19125,N_18986,N_18806);
or U19126 (N_19126,N_18944,N_18936);
xnor U19127 (N_19127,N_18838,N_18890);
xnor U19128 (N_19128,N_18913,N_18778);
nor U19129 (N_19129,N_18876,N_18867);
nand U19130 (N_19130,N_18867,N_18751);
or U19131 (N_19131,N_18882,N_18930);
and U19132 (N_19132,N_18784,N_18903);
nand U19133 (N_19133,N_18977,N_18903);
or U19134 (N_19134,N_18928,N_18838);
nand U19135 (N_19135,N_18794,N_18953);
nand U19136 (N_19136,N_18784,N_18799);
and U19137 (N_19137,N_18821,N_18819);
and U19138 (N_19138,N_18824,N_18870);
xnor U19139 (N_19139,N_18911,N_18966);
and U19140 (N_19140,N_18997,N_18906);
nor U19141 (N_19141,N_18914,N_18988);
nand U19142 (N_19142,N_18841,N_18839);
xnor U19143 (N_19143,N_18780,N_18891);
xor U19144 (N_19144,N_18807,N_18819);
and U19145 (N_19145,N_18818,N_18803);
or U19146 (N_19146,N_18930,N_18761);
nand U19147 (N_19147,N_18864,N_18977);
or U19148 (N_19148,N_18879,N_18964);
nand U19149 (N_19149,N_18983,N_18853);
xnor U19150 (N_19150,N_18935,N_18828);
xor U19151 (N_19151,N_18785,N_18877);
and U19152 (N_19152,N_18945,N_18852);
nand U19153 (N_19153,N_18785,N_18853);
or U19154 (N_19154,N_18936,N_18813);
nor U19155 (N_19155,N_18792,N_18991);
nand U19156 (N_19156,N_18981,N_18945);
nor U19157 (N_19157,N_18953,N_18884);
nand U19158 (N_19158,N_18887,N_18902);
xor U19159 (N_19159,N_18938,N_18973);
nand U19160 (N_19160,N_18782,N_18905);
nand U19161 (N_19161,N_18989,N_18987);
and U19162 (N_19162,N_18919,N_18819);
nor U19163 (N_19163,N_18782,N_18929);
nand U19164 (N_19164,N_18929,N_18897);
or U19165 (N_19165,N_18867,N_18857);
and U19166 (N_19166,N_18793,N_18862);
xor U19167 (N_19167,N_18884,N_18988);
nor U19168 (N_19168,N_18815,N_18961);
nand U19169 (N_19169,N_18776,N_18838);
xor U19170 (N_19170,N_18844,N_18776);
or U19171 (N_19171,N_18957,N_18980);
xor U19172 (N_19172,N_18911,N_18783);
nand U19173 (N_19173,N_18790,N_18859);
nand U19174 (N_19174,N_18915,N_18963);
nor U19175 (N_19175,N_18863,N_18940);
or U19176 (N_19176,N_18787,N_18964);
and U19177 (N_19177,N_18827,N_18852);
nand U19178 (N_19178,N_18956,N_18838);
or U19179 (N_19179,N_18957,N_18995);
and U19180 (N_19180,N_18991,N_18795);
or U19181 (N_19181,N_18830,N_18768);
nor U19182 (N_19182,N_18844,N_18943);
or U19183 (N_19183,N_18926,N_18918);
nand U19184 (N_19184,N_18987,N_18770);
nand U19185 (N_19185,N_18960,N_18784);
xor U19186 (N_19186,N_18815,N_18765);
nand U19187 (N_19187,N_18988,N_18977);
nand U19188 (N_19188,N_18762,N_18782);
nor U19189 (N_19189,N_18945,N_18966);
and U19190 (N_19190,N_18964,N_18980);
or U19191 (N_19191,N_18893,N_18995);
and U19192 (N_19192,N_18918,N_18987);
nor U19193 (N_19193,N_18993,N_18990);
nand U19194 (N_19194,N_18816,N_18936);
or U19195 (N_19195,N_18941,N_18905);
or U19196 (N_19196,N_18827,N_18846);
nor U19197 (N_19197,N_18752,N_18967);
xor U19198 (N_19198,N_18781,N_18773);
xnor U19199 (N_19199,N_18896,N_18877);
and U19200 (N_19200,N_18774,N_18902);
nand U19201 (N_19201,N_18943,N_18929);
nand U19202 (N_19202,N_18846,N_18944);
nand U19203 (N_19203,N_18973,N_18833);
or U19204 (N_19204,N_18849,N_18804);
nor U19205 (N_19205,N_18988,N_18836);
nand U19206 (N_19206,N_18800,N_18971);
or U19207 (N_19207,N_18823,N_18795);
nand U19208 (N_19208,N_18859,N_18934);
nor U19209 (N_19209,N_18810,N_18946);
or U19210 (N_19210,N_18784,N_18760);
or U19211 (N_19211,N_18816,N_18887);
nand U19212 (N_19212,N_18802,N_18942);
nor U19213 (N_19213,N_18877,N_18762);
and U19214 (N_19214,N_18807,N_18889);
or U19215 (N_19215,N_18774,N_18787);
and U19216 (N_19216,N_18941,N_18965);
or U19217 (N_19217,N_18874,N_18788);
or U19218 (N_19218,N_18873,N_18865);
or U19219 (N_19219,N_18975,N_18972);
nand U19220 (N_19220,N_18919,N_18838);
or U19221 (N_19221,N_18767,N_18931);
nand U19222 (N_19222,N_18851,N_18809);
and U19223 (N_19223,N_18807,N_18756);
nor U19224 (N_19224,N_18751,N_18760);
or U19225 (N_19225,N_18754,N_18911);
xor U19226 (N_19226,N_18881,N_18961);
and U19227 (N_19227,N_18898,N_18831);
nor U19228 (N_19228,N_18904,N_18994);
and U19229 (N_19229,N_18804,N_18891);
nor U19230 (N_19230,N_18841,N_18820);
and U19231 (N_19231,N_18947,N_18951);
nor U19232 (N_19232,N_18862,N_18997);
and U19233 (N_19233,N_18751,N_18827);
nor U19234 (N_19234,N_18796,N_18906);
nor U19235 (N_19235,N_18958,N_18918);
xnor U19236 (N_19236,N_18994,N_18777);
nand U19237 (N_19237,N_18960,N_18850);
or U19238 (N_19238,N_18984,N_18831);
nand U19239 (N_19239,N_18903,N_18783);
xnor U19240 (N_19240,N_18871,N_18997);
or U19241 (N_19241,N_18904,N_18875);
xnor U19242 (N_19242,N_18877,N_18842);
or U19243 (N_19243,N_18838,N_18998);
and U19244 (N_19244,N_18795,N_18974);
xnor U19245 (N_19245,N_18980,N_18906);
nand U19246 (N_19246,N_18840,N_18871);
and U19247 (N_19247,N_18882,N_18946);
and U19248 (N_19248,N_18874,N_18790);
or U19249 (N_19249,N_18844,N_18876);
nand U19250 (N_19250,N_19086,N_19158);
nor U19251 (N_19251,N_19203,N_19091);
nand U19252 (N_19252,N_19126,N_19141);
nand U19253 (N_19253,N_19016,N_19041);
and U19254 (N_19254,N_19169,N_19094);
nor U19255 (N_19255,N_19178,N_19156);
and U19256 (N_19256,N_19185,N_19002);
or U19257 (N_19257,N_19088,N_19052);
or U19258 (N_19258,N_19183,N_19146);
or U19259 (N_19259,N_19054,N_19192);
nand U19260 (N_19260,N_19234,N_19006);
nor U19261 (N_19261,N_19076,N_19139);
nor U19262 (N_19262,N_19096,N_19123);
and U19263 (N_19263,N_19108,N_19160);
and U19264 (N_19264,N_19167,N_19188);
nor U19265 (N_19265,N_19067,N_19189);
and U19266 (N_19266,N_19101,N_19200);
or U19267 (N_19267,N_19119,N_19171);
and U19268 (N_19268,N_19191,N_19173);
xor U19269 (N_19269,N_19049,N_19177);
and U19270 (N_19270,N_19075,N_19204);
or U19271 (N_19271,N_19085,N_19175);
and U19272 (N_19272,N_19045,N_19174);
or U19273 (N_19273,N_19140,N_19034);
and U19274 (N_19274,N_19064,N_19065);
or U19275 (N_19275,N_19196,N_19113);
nand U19276 (N_19276,N_19093,N_19226);
nor U19277 (N_19277,N_19068,N_19100);
or U19278 (N_19278,N_19147,N_19181);
nand U19279 (N_19279,N_19029,N_19249);
nor U19280 (N_19280,N_19214,N_19179);
or U19281 (N_19281,N_19240,N_19103);
nand U19282 (N_19282,N_19025,N_19166);
xnor U19283 (N_19283,N_19057,N_19237);
nor U19284 (N_19284,N_19242,N_19236);
nand U19285 (N_19285,N_19230,N_19001);
nor U19286 (N_19286,N_19000,N_19221);
nor U19287 (N_19287,N_19161,N_19210);
xnor U19288 (N_19288,N_19186,N_19205);
nor U19289 (N_19289,N_19247,N_19013);
nand U19290 (N_19290,N_19144,N_19190);
or U19291 (N_19291,N_19035,N_19028);
and U19292 (N_19292,N_19066,N_19157);
and U19293 (N_19293,N_19056,N_19246);
nor U19294 (N_19294,N_19199,N_19176);
or U19295 (N_19295,N_19198,N_19079);
nor U19296 (N_19296,N_19211,N_19128);
nor U19297 (N_19297,N_19032,N_19219);
or U19298 (N_19298,N_19172,N_19239);
and U19299 (N_19299,N_19021,N_19072);
nand U19300 (N_19300,N_19248,N_19238);
and U19301 (N_19301,N_19009,N_19043);
nor U19302 (N_19302,N_19137,N_19020);
or U19303 (N_19303,N_19011,N_19154);
nand U19304 (N_19304,N_19110,N_19130);
or U19305 (N_19305,N_19074,N_19058);
and U19306 (N_19306,N_19047,N_19050);
nand U19307 (N_19307,N_19111,N_19129);
and U19308 (N_19308,N_19023,N_19195);
nand U19309 (N_19309,N_19228,N_19115);
xnor U19310 (N_19310,N_19084,N_19132);
nor U19311 (N_19311,N_19187,N_19117);
nor U19312 (N_19312,N_19015,N_19180);
nand U19313 (N_19313,N_19134,N_19155);
nand U19314 (N_19314,N_19099,N_19225);
nor U19315 (N_19315,N_19209,N_19212);
nand U19316 (N_19316,N_19046,N_19201);
and U19317 (N_19317,N_19112,N_19217);
nand U19318 (N_19318,N_19215,N_19102);
and U19319 (N_19319,N_19004,N_19048);
or U19320 (N_19320,N_19005,N_19193);
or U19321 (N_19321,N_19202,N_19243);
xnor U19322 (N_19322,N_19208,N_19151);
and U19323 (N_19323,N_19039,N_19107);
xnor U19324 (N_19324,N_19007,N_19061);
nand U19325 (N_19325,N_19159,N_19116);
and U19326 (N_19326,N_19133,N_19232);
and U19327 (N_19327,N_19038,N_19003);
or U19328 (N_19328,N_19019,N_19222);
and U19329 (N_19329,N_19098,N_19010);
and U19330 (N_19330,N_19145,N_19142);
nand U19331 (N_19331,N_19182,N_19168);
and U19332 (N_19332,N_19073,N_19104);
or U19333 (N_19333,N_19136,N_19149);
nand U19334 (N_19334,N_19062,N_19077);
nand U19335 (N_19335,N_19184,N_19030);
nor U19336 (N_19336,N_19031,N_19241);
nand U19337 (N_19337,N_19233,N_19163);
nor U19338 (N_19338,N_19053,N_19224);
nand U19339 (N_19339,N_19090,N_19109);
or U19340 (N_19340,N_19078,N_19033);
nor U19341 (N_19341,N_19106,N_19118);
nor U19342 (N_19342,N_19153,N_19127);
nand U19343 (N_19343,N_19089,N_19017);
and U19344 (N_19344,N_19170,N_19071);
and U19345 (N_19345,N_19024,N_19083);
or U19346 (N_19346,N_19218,N_19120);
xnor U19347 (N_19347,N_19223,N_19042);
nor U19348 (N_19348,N_19121,N_19135);
xor U19349 (N_19349,N_19213,N_19044);
nand U19350 (N_19350,N_19164,N_19070);
or U19351 (N_19351,N_19092,N_19125);
nand U19352 (N_19352,N_19040,N_19036);
nor U19353 (N_19353,N_19095,N_19082);
nor U19354 (N_19354,N_19097,N_19229);
and U19355 (N_19355,N_19069,N_19162);
nand U19356 (N_19356,N_19027,N_19197);
xor U19357 (N_19357,N_19194,N_19014);
nand U19358 (N_19358,N_19055,N_19105);
nor U19359 (N_19359,N_19051,N_19063);
or U19360 (N_19360,N_19138,N_19206);
nor U19361 (N_19361,N_19022,N_19245);
nand U19362 (N_19362,N_19235,N_19037);
and U19363 (N_19363,N_19150,N_19148);
and U19364 (N_19364,N_19143,N_19081);
xnor U19365 (N_19365,N_19122,N_19026);
nor U19366 (N_19366,N_19207,N_19018);
or U19367 (N_19367,N_19124,N_19152);
and U19368 (N_19368,N_19114,N_19059);
nand U19369 (N_19369,N_19080,N_19131);
and U19370 (N_19370,N_19165,N_19227);
xnor U19371 (N_19371,N_19087,N_19244);
nor U19372 (N_19372,N_19008,N_19216);
and U19373 (N_19373,N_19220,N_19012);
nand U19374 (N_19374,N_19060,N_19231);
nor U19375 (N_19375,N_19195,N_19147);
nand U19376 (N_19376,N_19171,N_19109);
and U19377 (N_19377,N_19084,N_19172);
xnor U19378 (N_19378,N_19199,N_19162);
and U19379 (N_19379,N_19094,N_19044);
nand U19380 (N_19380,N_19028,N_19020);
nor U19381 (N_19381,N_19196,N_19090);
nor U19382 (N_19382,N_19162,N_19156);
xnor U19383 (N_19383,N_19072,N_19095);
xor U19384 (N_19384,N_19118,N_19171);
nand U19385 (N_19385,N_19147,N_19150);
or U19386 (N_19386,N_19014,N_19198);
xnor U19387 (N_19387,N_19194,N_19157);
xor U19388 (N_19388,N_19248,N_19077);
and U19389 (N_19389,N_19171,N_19196);
nand U19390 (N_19390,N_19031,N_19049);
nor U19391 (N_19391,N_19097,N_19102);
and U19392 (N_19392,N_19207,N_19081);
and U19393 (N_19393,N_19211,N_19038);
nor U19394 (N_19394,N_19109,N_19080);
or U19395 (N_19395,N_19073,N_19021);
and U19396 (N_19396,N_19212,N_19141);
xnor U19397 (N_19397,N_19041,N_19101);
nor U19398 (N_19398,N_19000,N_19092);
nor U19399 (N_19399,N_19134,N_19131);
nand U19400 (N_19400,N_19002,N_19107);
nor U19401 (N_19401,N_19035,N_19122);
nand U19402 (N_19402,N_19198,N_19076);
xnor U19403 (N_19403,N_19080,N_19048);
or U19404 (N_19404,N_19103,N_19143);
and U19405 (N_19405,N_19129,N_19140);
and U19406 (N_19406,N_19136,N_19094);
and U19407 (N_19407,N_19052,N_19211);
nor U19408 (N_19408,N_19157,N_19161);
xnor U19409 (N_19409,N_19133,N_19121);
and U19410 (N_19410,N_19061,N_19010);
or U19411 (N_19411,N_19101,N_19155);
nor U19412 (N_19412,N_19035,N_19217);
xor U19413 (N_19413,N_19017,N_19006);
xnor U19414 (N_19414,N_19095,N_19040);
and U19415 (N_19415,N_19031,N_19148);
or U19416 (N_19416,N_19006,N_19038);
xor U19417 (N_19417,N_19067,N_19208);
nand U19418 (N_19418,N_19214,N_19104);
xor U19419 (N_19419,N_19170,N_19104);
nand U19420 (N_19420,N_19100,N_19074);
or U19421 (N_19421,N_19040,N_19177);
xnor U19422 (N_19422,N_19234,N_19062);
and U19423 (N_19423,N_19220,N_19010);
or U19424 (N_19424,N_19216,N_19218);
or U19425 (N_19425,N_19108,N_19154);
or U19426 (N_19426,N_19196,N_19222);
nand U19427 (N_19427,N_19020,N_19121);
nand U19428 (N_19428,N_19050,N_19145);
nor U19429 (N_19429,N_19121,N_19151);
nand U19430 (N_19430,N_19219,N_19226);
xnor U19431 (N_19431,N_19115,N_19016);
and U19432 (N_19432,N_19239,N_19205);
or U19433 (N_19433,N_19027,N_19224);
and U19434 (N_19434,N_19150,N_19225);
or U19435 (N_19435,N_19240,N_19033);
or U19436 (N_19436,N_19009,N_19121);
or U19437 (N_19437,N_19062,N_19213);
xor U19438 (N_19438,N_19179,N_19193);
xnor U19439 (N_19439,N_19176,N_19248);
xnor U19440 (N_19440,N_19177,N_19083);
or U19441 (N_19441,N_19138,N_19203);
nor U19442 (N_19442,N_19093,N_19157);
xnor U19443 (N_19443,N_19089,N_19008);
or U19444 (N_19444,N_19074,N_19040);
xnor U19445 (N_19445,N_19198,N_19054);
nor U19446 (N_19446,N_19211,N_19096);
nor U19447 (N_19447,N_19184,N_19069);
nor U19448 (N_19448,N_19231,N_19213);
or U19449 (N_19449,N_19235,N_19061);
xor U19450 (N_19450,N_19117,N_19176);
nor U19451 (N_19451,N_19076,N_19181);
or U19452 (N_19452,N_19248,N_19221);
or U19453 (N_19453,N_19038,N_19015);
nand U19454 (N_19454,N_19162,N_19153);
and U19455 (N_19455,N_19113,N_19077);
nor U19456 (N_19456,N_19077,N_19178);
and U19457 (N_19457,N_19153,N_19142);
or U19458 (N_19458,N_19218,N_19143);
and U19459 (N_19459,N_19122,N_19242);
and U19460 (N_19460,N_19015,N_19177);
nor U19461 (N_19461,N_19198,N_19157);
xnor U19462 (N_19462,N_19014,N_19239);
xor U19463 (N_19463,N_19155,N_19110);
xor U19464 (N_19464,N_19196,N_19207);
nand U19465 (N_19465,N_19060,N_19133);
and U19466 (N_19466,N_19240,N_19173);
xor U19467 (N_19467,N_19235,N_19000);
and U19468 (N_19468,N_19092,N_19110);
or U19469 (N_19469,N_19234,N_19101);
or U19470 (N_19470,N_19053,N_19163);
nand U19471 (N_19471,N_19029,N_19112);
nor U19472 (N_19472,N_19162,N_19229);
nand U19473 (N_19473,N_19070,N_19243);
and U19474 (N_19474,N_19137,N_19179);
xor U19475 (N_19475,N_19057,N_19202);
xnor U19476 (N_19476,N_19049,N_19111);
or U19477 (N_19477,N_19141,N_19132);
xor U19478 (N_19478,N_19036,N_19210);
and U19479 (N_19479,N_19104,N_19206);
or U19480 (N_19480,N_19161,N_19011);
nand U19481 (N_19481,N_19068,N_19169);
xnor U19482 (N_19482,N_19080,N_19218);
or U19483 (N_19483,N_19239,N_19046);
xnor U19484 (N_19484,N_19118,N_19020);
or U19485 (N_19485,N_19196,N_19110);
or U19486 (N_19486,N_19215,N_19198);
and U19487 (N_19487,N_19206,N_19038);
or U19488 (N_19488,N_19053,N_19040);
and U19489 (N_19489,N_19142,N_19208);
or U19490 (N_19490,N_19186,N_19136);
nor U19491 (N_19491,N_19085,N_19073);
or U19492 (N_19492,N_19192,N_19133);
or U19493 (N_19493,N_19000,N_19098);
xor U19494 (N_19494,N_19168,N_19029);
nor U19495 (N_19495,N_19042,N_19104);
xnor U19496 (N_19496,N_19128,N_19072);
nor U19497 (N_19497,N_19159,N_19164);
nor U19498 (N_19498,N_19220,N_19151);
or U19499 (N_19499,N_19007,N_19178);
nor U19500 (N_19500,N_19315,N_19355);
xnor U19501 (N_19501,N_19428,N_19345);
nor U19502 (N_19502,N_19285,N_19442);
nand U19503 (N_19503,N_19256,N_19347);
and U19504 (N_19504,N_19254,N_19307);
nand U19505 (N_19505,N_19297,N_19263);
nor U19506 (N_19506,N_19420,N_19333);
and U19507 (N_19507,N_19473,N_19374);
xnor U19508 (N_19508,N_19482,N_19349);
and U19509 (N_19509,N_19399,N_19364);
xnor U19510 (N_19510,N_19381,N_19351);
and U19511 (N_19511,N_19441,N_19425);
or U19512 (N_19512,N_19472,N_19252);
or U19513 (N_19513,N_19492,N_19393);
nand U19514 (N_19514,N_19447,N_19436);
and U19515 (N_19515,N_19375,N_19474);
nor U19516 (N_19516,N_19324,N_19417);
or U19517 (N_19517,N_19402,N_19437);
nand U19518 (N_19518,N_19450,N_19498);
nand U19519 (N_19519,N_19448,N_19406);
or U19520 (N_19520,N_19267,N_19359);
nor U19521 (N_19521,N_19433,N_19301);
xor U19522 (N_19522,N_19395,N_19319);
nand U19523 (N_19523,N_19386,N_19497);
and U19524 (N_19524,N_19342,N_19443);
and U19525 (N_19525,N_19274,N_19449);
xnor U19526 (N_19526,N_19348,N_19264);
nor U19527 (N_19527,N_19275,N_19266);
xnor U19528 (N_19528,N_19286,N_19404);
nand U19529 (N_19529,N_19346,N_19467);
and U19530 (N_19530,N_19369,N_19427);
nand U19531 (N_19531,N_19257,N_19332);
and U19532 (N_19532,N_19278,N_19444);
nor U19533 (N_19533,N_19268,N_19320);
nor U19534 (N_19534,N_19304,N_19314);
nor U19535 (N_19535,N_19353,N_19476);
xor U19536 (N_19536,N_19488,N_19271);
nand U19537 (N_19537,N_19489,N_19480);
xnor U19538 (N_19538,N_19251,N_19258);
xor U19539 (N_19539,N_19317,N_19331);
or U19540 (N_19540,N_19398,N_19387);
xor U19541 (N_19541,N_19466,N_19388);
or U19542 (N_19542,N_19358,N_19438);
xor U19543 (N_19543,N_19414,N_19439);
or U19544 (N_19544,N_19487,N_19394);
or U19545 (N_19545,N_19362,N_19255);
or U19546 (N_19546,N_19470,N_19343);
nand U19547 (N_19547,N_19460,N_19405);
and U19548 (N_19548,N_19323,N_19260);
and U19549 (N_19549,N_19431,N_19261);
or U19550 (N_19550,N_19360,N_19253);
and U19551 (N_19551,N_19352,N_19366);
nor U19552 (N_19552,N_19457,N_19298);
nor U19553 (N_19553,N_19306,N_19471);
xnor U19554 (N_19554,N_19400,N_19336);
nand U19555 (N_19555,N_19451,N_19294);
or U19556 (N_19556,N_19269,N_19344);
or U19557 (N_19557,N_19270,N_19340);
nor U19558 (N_19558,N_19328,N_19485);
xnor U19559 (N_19559,N_19373,N_19335);
or U19560 (N_19560,N_19290,N_19376);
xnor U19561 (N_19561,N_19415,N_19367);
xnor U19562 (N_19562,N_19280,N_19459);
nor U19563 (N_19563,N_19452,N_19377);
or U19564 (N_19564,N_19273,N_19490);
nor U19565 (N_19565,N_19327,N_19461);
or U19566 (N_19566,N_19350,N_19391);
xnor U19567 (N_19567,N_19426,N_19419);
or U19568 (N_19568,N_19311,N_19262);
xnor U19569 (N_19569,N_19334,N_19302);
nor U19570 (N_19570,N_19435,N_19378);
or U19571 (N_19571,N_19308,N_19422);
nor U19572 (N_19572,N_19318,N_19322);
or U19573 (N_19573,N_19478,N_19372);
nand U19574 (N_19574,N_19495,N_19403);
nand U19575 (N_19575,N_19293,N_19465);
xnor U19576 (N_19576,N_19287,N_19413);
nand U19577 (N_19577,N_19390,N_19316);
or U19578 (N_19578,N_19458,N_19259);
xnor U19579 (N_19579,N_19283,N_19463);
or U19580 (N_19580,N_19412,N_19289);
and U19581 (N_19581,N_19416,N_19300);
nor U19582 (N_19582,N_19385,N_19313);
or U19583 (N_19583,N_19496,N_19409);
nand U19584 (N_19584,N_19380,N_19341);
xnor U19585 (N_19585,N_19424,N_19371);
nand U19586 (N_19586,N_19408,N_19368);
nand U19587 (N_19587,N_19454,N_19410);
or U19588 (N_19588,N_19484,N_19384);
nor U19589 (N_19589,N_19464,N_19357);
and U19590 (N_19590,N_19337,N_19407);
nand U19591 (N_19591,N_19491,N_19421);
or U19592 (N_19592,N_19475,N_19279);
and U19593 (N_19593,N_19363,N_19430);
nor U19594 (N_19594,N_19493,N_19432);
and U19595 (N_19595,N_19303,N_19296);
or U19596 (N_19596,N_19312,N_19440);
nor U19597 (N_19597,N_19276,N_19329);
xor U19598 (N_19598,N_19284,N_19265);
nand U19599 (N_19599,N_19277,N_19292);
and U19600 (N_19600,N_19356,N_19309);
xor U19601 (N_19601,N_19446,N_19272);
nor U19602 (N_19602,N_19382,N_19379);
nor U19603 (N_19603,N_19383,N_19310);
xor U19604 (N_19604,N_19288,N_19305);
nand U19605 (N_19605,N_19299,N_19494);
nor U19606 (N_19606,N_19468,N_19295);
or U19607 (N_19607,N_19325,N_19429);
xnor U19608 (N_19608,N_19453,N_19321);
nand U19609 (N_19609,N_19411,N_19462);
nand U19610 (N_19610,N_19456,N_19483);
and U19611 (N_19611,N_19469,N_19434);
xor U19612 (N_19612,N_19396,N_19477);
nand U19613 (N_19613,N_19397,N_19486);
xnor U19614 (N_19614,N_19445,N_19282);
and U19615 (N_19615,N_19250,N_19401);
nor U19616 (N_19616,N_19281,N_19481);
nand U19617 (N_19617,N_19365,N_19455);
and U19618 (N_19618,N_19499,N_19370);
nand U19619 (N_19619,N_19479,N_19423);
xnor U19620 (N_19620,N_19389,N_19330);
nor U19621 (N_19621,N_19291,N_19392);
xnor U19622 (N_19622,N_19326,N_19338);
xor U19623 (N_19623,N_19361,N_19354);
or U19624 (N_19624,N_19339,N_19418);
nand U19625 (N_19625,N_19411,N_19429);
nor U19626 (N_19626,N_19367,N_19440);
nand U19627 (N_19627,N_19482,N_19376);
nand U19628 (N_19628,N_19353,N_19293);
xnor U19629 (N_19629,N_19360,N_19440);
and U19630 (N_19630,N_19499,N_19439);
nand U19631 (N_19631,N_19460,N_19338);
xor U19632 (N_19632,N_19265,N_19335);
or U19633 (N_19633,N_19314,N_19474);
nand U19634 (N_19634,N_19426,N_19421);
xor U19635 (N_19635,N_19253,N_19263);
and U19636 (N_19636,N_19255,N_19325);
nand U19637 (N_19637,N_19401,N_19281);
nand U19638 (N_19638,N_19265,N_19300);
nand U19639 (N_19639,N_19395,N_19308);
nand U19640 (N_19640,N_19420,N_19387);
nand U19641 (N_19641,N_19426,N_19397);
xor U19642 (N_19642,N_19424,N_19418);
or U19643 (N_19643,N_19427,N_19280);
nand U19644 (N_19644,N_19437,N_19430);
and U19645 (N_19645,N_19259,N_19417);
xnor U19646 (N_19646,N_19401,N_19440);
or U19647 (N_19647,N_19265,N_19309);
and U19648 (N_19648,N_19401,N_19411);
or U19649 (N_19649,N_19316,N_19317);
nor U19650 (N_19650,N_19408,N_19499);
nand U19651 (N_19651,N_19376,N_19338);
nor U19652 (N_19652,N_19327,N_19298);
and U19653 (N_19653,N_19312,N_19398);
or U19654 (N_19654,N_19409,N_19291);
nand U19655 (N_19655,N_19426,N_19485);
xnor U19656 (N_19656,N_19292,N_19488);
and U19657 (N_19657,N_19484,N_19291);
nand U19658 (N_19658,N_19398,N_19396);
xor U19659 (N_19659,N_19261,N_19494);
nor U19660 (N_19660,N_19279,N_19256);
and U19661 (N_19661,N_19283,N_19262);
or U19662 (N_19662,N_19331,N_19373);
nor U19663 (N_19663,N_19411,N_19263);
and U19664 (N_19664,N_19488,N_19348);
nor U19665 (N_19665,N_19403,N_19275);
or U19666 (N_19666,N_19380,N_19437);
nand U19667 (N_19667,N_19479,N_19359);
nor U19668 (N_19668,N_19483,N_19286);
nand U19669 (N_19669,N_19381,N_19379);
or U19670 (N_19670,N_19491,N_19398);
nand U19671 (N_19671,N_19291,N_19390);
xor U19672 (N_19672,N_19479,N_19310);
nand U19673 (N_19673,N_19477,N_19344);
and U19674 (N_19674,N_19376,N_19495);
or U19675 (N_19675,N_19385,N_19266);
and U19676 (N_19676,N_19432,N_19292);
nor U19677 (N_19677,N_19334,N_19451);
xnor U19678 (N_19678,N_19373,N_19323);
xnor U19679 (N_19679,N_19465,N_19281);
nand U19680 (N_19680,N_19455,N_19323);
or U19681 (N_19681,N_19272,N_19492);
and U19682 (N_19682,N_19252,N_19334);
nor U19683 (N_19683,N_19306,N_19401);
or U19684 (N_19684,N_19328,N_19338);
and U19685 (N_19685,N_19337,N_19488);
nand U19686 (N_19686,N_19308,N_19450);
and U19687 (N_19687,N_19496,N_19489);
xnor U19688 (N_19688,N_19467,N_19254);
nor U19689 (N_19689,N_19338,N_19418);
nand U19690 (N_19690,N_19433,N_19331);
or U19691 (N_19691,N_19480,N_19352);
and U19692 (N_19692,N_19269,N_19444);
and U19693 (N_19693,N_19478,N_19400);
or U19694 (N_19694,N_19487,N_19323);
nand U19695 (N_19695,N_19276,N_19296);
nor U19696 (N_19696,N_19465,N_19338);
xnor U19697 (N_19697,N_19411,N_19292);
xnor U19698 (N_19698,N_19353,N_19318);
and U19699 (N_19699,N_19491,N_19319);
xor U19700 (N_19700,N_19399,N_19370);
xor U19701 (N_19701,N_19443,N_19451);
nand U19702 (N_19702,N_19314,N_19255);
xnor U19703 (N_19703,N_19322,N_19368);
nor U19704 (N_19704,N_19388,N_19445);
and U19705 (N_19705,N_19376,N_19364);
nand U19706 (N_19706,N_19340,N_19470);
or U19707 (N_19707,N_19295,N_19403);
xnor U19708 (N_19708,N_19292,N_19449);
nand U19709 (N_19709,N_19372,N_19381);
nand U19710 (N_19710,N_19418,N_19386);
xor U19711 (N_19711,N_19295,N_19413);
and U19712 (N_19712,N_19401,N_19407);
nand U19713 (N_19713,N_19465,N_19330);
and U19714 (N_19714,N_19464,N_19395);
nor U19715 (N_19715,N_19267,N_19481);
or U19716 (N_19716,N_19422,N_19442);
nand U19717 (N_19717,N_19497,N_19442);
or U19718 (N_19718,N_19491,N_19433);
xor U19719 (N_19719,N_19385,N_19277);
xor U19720 (N_19720,N_19255,N_19484);
and U19721 (N_19721,N_19362,N_19420);
or U19722 (N_19722,N_19385,N_19307);
xnor U19723 (N_19723,N_19315,N_19386);
xor U19724 (N_19724,N_19401,N_19384);
and U19725 (N_19725,N_19478,N_19289);
or U19726 (N_19726,N_19326,N_19426);
and U19727 (N_19727,N_19352,N_19410);
nand U19728 (N_19728,N_19357,N_19436);
nor U19729 (N_19729,N_19301,N_19486);
nand U19730 (N_19730,N_19283,N_19411);
nand U19731 (N_19731,N_19479,N_19254);
nand U19732 (N_19732,N_19463,N_19361);
or U19733 (N_19733,N_19470,N_19260);
xnor U19734 (N_19734,N_19482,N_19450);
or U19735 (N_19735,N_19487,N_19468);
or U19736 (N_19736,N_19479,N_19420);
nand U19737 (N_19737,N_19445,N_19389);
and U19738 (N_19738,N_19402,N_19323);
nor U19739 (N_19739,N_19253,N_19432);
nand U19740 (N_19740,N_19402,N_19288);
and U19741 (N_19741,N_19482,N_19451);
or U19742 (N_19742,N_19300,N_19305);
and U19743 (N_19743,N_19450,N_19436);
xnor U19744 (N_19744,N_19472,N_19444);
nor U19745 (N_19745,N_19434,N_19350);
or U19746 (N_19746,N_19479,N_19333);
nor U19747 (N_19747,N_19370,N_19362);
and U19748 (N_19748,N_19447,N_19364);
nor U19749 (N_19749,N_19357,N_19266);
nor U19750 (N_19750,N_19578,N_19545);
or U19751 (N_19751,N_19615,N_19543);
nor U19752 (N_19752,N_19624,N_19731);
nor U19753 (N_19753,N_19567,N_19640);
or U19754 (N_19754,N_19715,N_19572);
nand U19755 (N_19755,N_19627,N_19724);
and U19756 (N_19756,N_19502,N_19618);
nand U19757 (N_19757,N_19535,N_19652);
nand U19758 (N_19758,N_19717,N_19603);
nand U19759 (N_19759,N_19656,N_19577);
and U19760 (N_19760,N_19554,N_19642);
or U19761 (N_19761,N_19564,N_19587);
or U19762 (N_19762,N_19550,N_19541);
nand U19763 (N_19763,N_19583,N_19637);
or U19764 (N_19764,N_19666,N_19730);
nor U19765 (N_19765,N_19621,N_19557);
and U19766 (N_19766,N_19584,N_19631);
or U19767 (N_19767,N_19505,N_19503);
and U19768 (N_19768,N_19542,N_19648);
nand U19769 (N_19769,N_19530,N_19510);
or U19770 (N_19770,N_19518,N_19555);
nand U19771 (N_19771,N_19500,N_19628);
or U19772 (N_19772,N_19527,N_19723);
nor U19773 (N_19773,N_19600,N_19629);
nor U19774 (N_19774,N_19690,N_19574);
nand U19775 (N_19775,N_19531,N_19607);
nand U19776 (N_19776,N_19726,N_19745);
xor U19777 (N_19777,N_19695,N_19722);
and U19778 (N_19778,N_19645,N_19619);
xor U19779 (N_19779,N_19719,N_19704);
and U19780 (N_19780,N_19683,N_19508);
nand U19781 (N_19781,N_19632,N_19720);
or U19782 (N_19782,N_19573,N_19571);
or U19783 (N_19783,N_19528,N_19699);
and U19784 (N_19784,N_19538,N_19570);
xor U19785 (N_19785,N_19625,N_19565);
nand U19786 (N_19786,N_19552,N_19714);
nor U19787 (N_19787,N_19639,N_19634);
or U19788 (N_19788,N_19622,N_19513);
nor U19789 (N_19789,N_19727,N_19739);
and U19790 (N_19790,N_19721,N_19534);
nand U19791 (N_19791,N_19654,N_19585);
or U19792 (N_19792,N_19716,N_19591);
nor U19793 (N_19793,N_19653,N_19589);
nor U19794 (N_19794,N_19507,N_19660);
nor U19795 (N_19795,N_19697,N_19743);
xnor U19796 (N_19796,N_19641,N_19678);
and U19797 (N_19797,N_19673,N_19698);
xor U19798 (N_19798,N_19630,N_19602);
or U19799 (N_19799,N_19665,N_19566);
or U19800 (N_19800,N_19604,N_19582);
xor U19801 (N_19801,N_19520,N_19676);
nor U19802 (N_19802,N_19668,N_19606);
nand U19803 (N_19803,N_19711,N_19680);
or U19804 (N_19804,N_19512,N_19701);
nor U19805 (N_19805,N_19620,N_19533);
or U19806 (N_19806,N_19563,N_19735);
and U19807 (N_19807,N_19601,N_19594);
or U19808 (N_19808,N_19738,N_19633);
nand U19809 (N_19809,N_19539,N_19526);
and U19810 (N_19810,N_19700,N_19517);
and U19811 (N_19811,N_19702,N_19609);
nor U19812 (N_19812,N_19576,N_19688);
nand U19813 (N_19813,N_19643,N_19506);
xor U19814 (N_19814,N_19655,N_19646);
nand U19815 (N_19815,N_19537,N_19669);
nand U19816 (N_19816,N_19547,N_19514);
nand U19817 (N_19817,N_19707,N_19667);
nand U19818 (N_19818,N_19741,N_19703);
or U19819 (N_19819,N_19605,N_19744);
nor U19820 (N_19820,N_19536,N_19725);
xor U19821 (N_19821,N_19663,N_19681);
nor U19822 (N_19822,N_19675,N_19623);
or U19823 (N_19823,N_19529,N_19685);
nor U19824 (N_19824,N_19511,N_19661);
and U19825 (N_19825,N_19532,N_19580);
nor U19826 (N_19826,N_19590,N_19662);
or U19827 (N_19827,N_19599,N_19558);
xor U19828 (N_19828,N_19610,N_19729);
nor U19829 (N_19829,N_19736,N_19617);
nor U19830 (N_19830,N_19689,N_19556);
and U19831 (N_19831,N_19608,N_19709);
nand U19832 (N_19832,N_19553,N_19521);
xor U19833 (N_19833,N_19677,N_19592);
or U19834 (N_19834,N_19638,N_19519);
nor U19835 (N_19835,N_19742,N_19644);
and U19836 (N_19836,N_19649,N_19692);
nand U19837 (N_19837,N_19515,N_19734);
and U19838 (N_19838,N_19706,N_19737);
xor U19839 (N_19839,N_19746,N_19635);
xor U19840 (N_19840,N_19613,N_19581);
nor U19841 (N_19841,N_19670,N_19686);
or U19842 (N_19842,N_19597,N_19616);
nand U19843 (N_19843,N_19712,N_19560);
nand U19844 (N_19844,N_19626,N_19748);
nand U19845 (N_19845,N_19569,N_19732);
nor U19846 (N_19846,N_19691,N_19728);
nor U19847 (N_19847,N_19586,N_19540);
xnor U19848 (N_19848,N_19544,N_19611);
nor U19849 (N_19849,N_19740,N_19694);
nand U19850 (N_19850,N_19525,N_19598);
xnor U19851 (N_19851,N_19693,N_19682);
xor U19852 (N_19852,N_19559,N_19708);
or U19853 (N_19853,N_19671,N_19687);
and U19854 (N_19854,N_19595,N_19658);
xor U19855 (N_19855,N_19546,N_19548);
xnor U19856 (N_19856,N_19579,N_19516);
nand U19857 (N_19857,N_19575,N_19747);
xor U19858 (N_19858,N_19523,N_19659);
nand U19859 (N_19859,N_19561,N_19524);
nor U19860 (N_19860,N_19549,N_19674);
and U19861 (N_19861,N_19733,N_19593);
xor U19862 (N_19862,N_19501,N_19696);
xor U19863 (N_19863,N_19562,N_19713);
nand U19864 (N_19864,N_19672,N_19657);
or U19865 (N_19865,N_19647,N_19664);
and U19866 (N_19866,N_19636,N_19679);
xnor U19867 (N_19867,N_19684,N_19588);
nand U19868 (N_19868,N_19568,N_19612);
nor U19869 (N_19869,N_19614,N_19509);
xnor U19870 (N_19870,N_19650,N_19651);
nand U19871 (N_19871,N_19749,N_19504);
and U19872 (N_19872,N_19551,N_19718);
nand U19873 (N_19873,N_19710,N_19522);
nor U19874 (N_19874,N_19596,N_19705);
nor U19875 (N_19875,N_19720,N_19539);
nor U19876 (N_19876,N_19564,N_19715);
or U19877 (N_19877,N_19718,N_19562);
and U19878 (N_19878,N_19538,N_19507);
nand U19879 (N_19879,N_19746,N_19601);
xor U19880 (N_19880,N_19523,N_19643);
and U19881 (N_19881,N_19716,N_19525);
or U19882 (N_19882,N_19707,N_19636);
nand U19883 (N_19883,N_19557,N_19646);
nand U19884 (N_19884,N_19503,N_19714);
nor U19885 (N_19885,N_19522,N_19601);
xnor U19886 (N_19886,N_19548,N_19591);
xnor U19887 (N_19887,N_19545,N_19687);
nand U19888 (N_19888,N_19607,N_19557);
nand U19889 (N_19889,N_19522,N_19549);
or U19890 (N_19890,N_19631,N_19715);
nor U19891 (N_19891,N_19565,N_19511);
nor U19892 (N_19892,N_19526,N_19705);
or U19893 (N_19893,N_19676,N_19670);
xnor U19894 (N_19894,N_19582,N_19576);
nand U19895 (N_19895,N_19717,N_19693);
nor U19896 (N_19896,N_19526,N_19597);
xnor U19897 (N_19897,N_19740,N_19690);
nor U19898 (N_19898,N_19701,N_19514);
and U19899 (N_19899,N_19585,N_19675);
nand U19900 (N_19900,N_19658,N_19570);
xor U19901 (N_19901,N_19719,N_19608);
nor U19902 (N_19902,N_19571,N_19612);
and U19903 (N_19903,N_19589,N_19699);
xnor U19904 (N_19904,N_19559,N_19511);
or U19905 (N_19905,N_19634,N_19536);
nand U19906 (N_19906,N_19543,N_19731);
xnor U19907 (N_19907,N_19684,N_19728);
xor U19908 (N_19908,N_19511,N_19568);
nor U19909 (N_19909,N_19685,N_19614);
nor U19910 (N_19910,N_19555,N_19528);
nor U19911 (N_19911,N_19573,N_19731);
nand U19912 (N_19912,N_19522,N_19722);
nand U19913 (N_19913,N_19743,N_19711);
and U19914 (N_19914,N_19734,N_19671);
nand U19915 (N_19915,N_19704,N_19706);
and U19916 (N_19916,N_19693,N_19712);
nor U19917 (N_19917,N_19677,N_19547);
and U19918 (N_19918,N_19614,N_19697);
and U19919 (N_19919,N_19736,N_19664);
xor U19920 (N_19920,N_19632,N_19719);
nor U19921 (N_19921,N_19748,N_19701);
and U19922 (N_19922,N_19627,N_19728);
xor U19923 (N_19923,N_19638,N_19606);
and U19924 (N_19924,N_19661,N_19512);
or U19925 (N_19925,N_19508,N_19515);
and U19926 (N_19926,N_19633,N_19657);
nand U19927 (N_19927,N_19630,N_19608);
and U19928 (N_19928,N_19627,N_19703);
xor U19929 (N_19929,N_19707,N_19595);
xnor U19930 (N_19930,N_19746,N_19531);
nor U19931 (N_19931,N_19701,N_19501);
nor U19932 (N_19932,N_19565,N_19510);
or U19933 (N_19933,N_19745,N_19681);
xnor U19934 (N_19934,N_19608,N_19517);
xnor U19935 (N_19935,N_19685,N_19741);
nor U19936 (N_19936,N_19729,N_19642);
nand U19937 (N_19937,N_19681,N_19641);
nor U19938 (N_19938,N_19614,N_19690);
nor U19939 (N_19939,N_19656,N_19624);
nor U19940 (N_19940,N_19529,N_19722);
xnor U19941 (N_19941,N_19617,N_19675);
and U19942 (N_19942,N_19724,N_19699);
or U19943 (N_19943,N_19648,N_19658);
nor U19944 (N_19944,N_19709,N_19596);
and U19945 (N_19945,N_19561,N_19670);
nand U19946 (N_19946,N_19549,N_19655);
or U19947 (N_19947,N_19501,N_19568);
or U19948 (N_19948,N_19698,N_19519);
nor U19949 (N_19949,N_19659,N_19509);
and U19950 (N_19950,N_19564,N_19645);
nor U19951 (N_19951,N_19605,N_19521);
nor U19952 (N_19952,N_19649,N_19712);
nand U19953 (N_19953,N_19604,N_19639);
and U19954 (N_19954,N_19670,N_19514);
and U19955 (N_19955,N_19741,N_19681);
and U19956 (N_19956,N_19506,N_19527);
nand U19957 (N_19957,N_19747,N_19516);
nor U19958 (N_19958,N_19713,N_19535);
nor U19959 (N_19959,N_19690,N_19558);
nand U19960 (N_19960,N_19641,N_19704);
and U19961 (N_19961,N_19610,N_19614);
nand U19962 (N_19962,N_19501,N_19745);
nor U19963 (N_19963,N_19624,N_19523);
or U19964 (N_19964,N_19532,N_19583);
and U19965 (N_19965,N_19687,N_19656);
or U19966 (N_19966,N_19699,N_19609);
xor U19967 (N_19967,N_19549,N_19562);
nor U19968 (N_19968,N_19538,N_19693);
nor U19969 (N_19969,N_19699,N_19667);
and U19970 (N_19970,N_19588,N_19584);
nor U19971 (N_19971,N_19689,N_19604);
xnor U19972 (N_19972,N_19522,N_19714);
nor U19973 (N_19973,N_19591,N_19529);
or U19974 (N_19974,N_19660,N_19558);
or U19975 (N_19975,N_19571,N_19659);
xnor U19976 (N_19976,N_19660,N_19571);
nor U19977 (N_19977,N_19641,N_19682);
nor U19978 (N_19978,N_19525,N_19563);
nand U19979 (N_19979,N_19735,N_19719);
nor U19980 (N_19980,N_19711,N_19535);
and U19981 (N_19981,N_19639,N_19653);
nand U19982 (N_19982,N_19598,N_19563);
xnor U19983 (N_19983,N_19633,N_19577);
nand U19984 (N_19984,N_19592,N_19596);
nand U19985 (N_19985,N_19655,N_19565);
and U19986 (N_19986,N_19532,N_19723);
nor U19987 (N_19987,N_19697,N_19674);
nor U19988 (N_19988,N_19570,N_19634);
and U19989 (N_19989,N_19548,N_19677);
xnor U19990 (N_19990,N_19742,N_19529);
and U19991 (N_19991,N_19505,N_19620);
xnor U19992 (N_19992,N_19683,N_19687);
nand U19993 (N_19993,N_19707,N_19739);
nand U19994 (N_19994,N_19607,N_19550);
nand U19995 (N_19995,N_19571,N_19724);
or U19996 (N_19996,N_19620,N_19545);
xor U19997 (N_19997,N_19638,N_19562);
xnor U19998 (N_19998,N_19731,N_19664);
nor U19999 (N_19999,N_19532,N_19663);
xnor UO_0 (O_0,N_19938,N_19900);
nor UO_1 (O_1,N_19873,N_19955);
and UO_2 (O_2,N_19830,N_19817);
xor UO_3 (O_3,N_19901,N_19983);
nor UO_4 (O_4,N_19928,N_19790);
nand UO_5 (O_5,N_19882,N_19871);
and UO_6 (O_6,N_19945,N_19785);
nand UO_7 (O_7,N_19761,N_19805);
xor UO_8 (O_8,N_19909,N_19925);
nand UO_9 (O_9,N_19821,N_19993);
or UO_10 (O_10,N_19895,N_19844);
xnor UO_11 (O_11,N_19890,N_19934);
xor UO_12 (O_12,N_19996,N_19984);
and UO_13 (O_13,N_19835,N_19974);
nand UO_14 (O_14,N_19898,N_19847);
nor UO_15 (O_15,N_19773,N_19939);
xor UO_16 (O_16,N_19961,N_19988);
nor UO_17 (O_17,N_19875,N_19903);
nor UO_18 (O_18,N_19798,N_19858);
nor UO_19 (O_19,N_19776,N_19941);
xor UO_20 (O_20,N_19839,N_19828);
or UO_21 (O_21,N_19850,N_19853);
nand UO_22 (O_22,N_19932,N_19896);
and UO_23 (O_23,N_19855,N_19891);
and UO_24 (O_24,N_19750,N_19775);
nor UO_25 (O_25,N_19977,N_19979);
or UO_26 (O_26,N_19788,N_19885);
nand UO_27 (O_27,N_19981,N_19926);
nand UO_28 (O_28,N_19881,N_19792);
nand UO_29 (O_29,N_19888,N_19889);
xnor UO_30 (O_30,N_19857,N_19860);
nor UO_31 (O_31,N_19783,N_19840);
and UO_32 (O_32,N_19978,N_19864);
xnor UO_33 (O_33,N_19849,N_19943);
and UO_34 (O_34,N_19794,N_19915);
and UO_35 (O_35,N_19751,N_19876);
nor UO_36 (O_36,N_19806,N_19942);
xor UO_37 (O_37,N_19877,N_19852);
nor UO_38 (O_38,N_19789,N_19770);
nor UO_39 (O_39,N_19766,N_19910);
and UO_40 (O_40,N_19762,N_19973);
nor UO_41 (O_41,N_19802,N_19989);
nand UO_42 (O_42,N_19797,N_19769);
or UO_43 (O_43,N_19758,N_19795);
and UO_44 (O_44,N_19969,N_19874);
nand UO_45 (O_45,N_19778,N_19812);
nor UO_46 (O_46,N_19980,N_19755);
nand UO_47 (O_47,N_19967,N_19917);
xor UO_48 (O_48,N_19800,N_19948);
xor UO_49 (O_49,N_19951,N_19902);
nor UO_50 (O_50,N_19958,N_19803);
and UO_51 (O_51,N_19784,N_19796);
xnor UO_52 (O_52,N_19911,N_19897);
and UO_53 (O_53,N_19827,N_19957);
xor UO_54 (O_54,N_19807,N_19968);
or UO_55 (O_55,N_19777,N_19809);
or UO_56 (O_56,N_19815,N_19754);
or UO_57 (O_57,N_19865,N_19845);
or UO_58 (O_58,N_19774,N_19834);
or UO_59 (O_59,N_19893,N_19914);
and UO_60 (O_60,N_19997,N_19818);
nand UO_61 (O_61,N_19907,N_19952);
or UO_62 (O_62,N_19819,N_19972);
nand UO_63 (O_63,N_19924,N_19870);
xnor UO_64 (O_64,N_19786,N_19994);
nand UO_65 (O_65,N_19810,N_19991);
or UO_66 (O_66,N_19808,N_19861);
nor UO_67 (O_67,N_19944,N_19990);
and UO_68 (O_68,N_19935,N_19930);
nor UO_69 (O_69,N_19933,N_19856);
or UO_70 (O_70,N_19752,N_19920);
xnor UO_71 (O_71,N_19878,N_19899);
and UO_72 (O_72,N_19886,N_19779);
nor UO_73 (O_73,N_19908,N_19929);
nor UO_74 (O_74,N_19879,N_19859);
and UO_75 (O_75,N_19867,N_19992);
nand UO_76 (O_76,N_19959,N_19999);
and UO_77 (O_77,N_19913,N_19905);
xnor UO_78 (O_78,N_19832,N_19854);
and UO_79 (O_79,N_19995,N_19804);
nor UO_80 (O_80,N_19843,N_19880);
or UO_81 (O_81,N_19962,N_19918);
or UO_82 (O_82,N_19764,N_19862);
or UO_83 (O_83,N_19842,N_19894);
nor UO_84 (O_84,N_19816,N_19987);
and UO_85 (O_85,N_19919,N_19970);
or UO_86 (O_86,N_19964,N_19963);
or UO_87 (O_87,N_19765,N_19950);
or UO_88 (O_88,N_19801,N_19823);
nor UO_89 (O_89,N_19927,N_19838);
or UO_90 (O_90,N_19863,N_19904);
nor UO_91 (O_91,N_19936,N_19824);
xnor UO_92 (O_92,N_19848,N_19940);
and UO_93 (O_93,N_19998,N_19956);
xor UO_94 (O_94,N_19966,N_19829);
xor UO_95 (O_95,N_19768,N_19960);
nor UO_96 (O_96,N_19772,N_19826);
xor UO_97 (O_97,N_19949,N_19954);
xor UO_98 (O_98,N_19837,N_19872);
and UO_99 (O_99,N_19820,N_19923);
or UO_100 (O_100,N_19912,N_19822);
or UO_101 (O_101,N_19976,N_19965);
nor UO_102 (O_102,N_19841,N_19780);
and UO_103 (O_103,N_19868,N_19799);
or UO_104 (O_104,N_19836,N_19916);
nand UO_105 (O_105,N_19759,N_19975);
or UO_106 (O_106,N_19793,N_19756);
nor UO_107 (O_107,N_19771,N_19811);
nor UO_108 (O_108,N_19906,N_19931);
and UO_109 (O_109,N_19833,N_19946);
xnor UO_110 (O_110,N_19947,N_19884);
or UO_111 (O_111,N_19757,N_19922);
nand UO_112 (O_112,N_19767,N_19985);
nand UO_113 (O_113,N_19887,N_19971);
nand UO_114 (O_114,N_19814,N_19753);
xor UO_115 (O_115,N_19869,N_19851);
and UO_116 (O_116,N_19846,N_19982);
nor UO_117 (O_117,N_19953,N_19787);
and UO_118 (O_118,N_19883,N_19763);
xor UO_119 (O_119,N_19791,N_19813);
xnor UO_120 (O_120,N_19825,N_19986);
nor UO_121 (O_121,N_19831,N_19760);
nand UO_122 (O_122,N_19866,N_19892);
and UO_123 (O_123,N_19782,N_19921);
nand UO_124 (O_124,N_19937,N_19781);
nor UO_125 (O_125,N_19787,N_19771);
nand UO_126 (O_126,N_19957,N_19952);
nor UO_127 (O_127,N_19842,N_19764);
nand UO_128 (O_128,N_19780,N_19928);
and UO_129 (O_129,N_19996,N_19822);
nand UO_130 (O_130,N_19941,N_19979);
nand UO_131 (O_131,N_19952,N_19795);
or UO_132 (O_132,N_19975,N_19779);
nor UO_133 (O_133,N_19778,N_19844);
nor UO_134 (O_134,N_19883,N_19801);
nand UO_135 (O_135,N_19842,N_19972);
and UO_136 (O_136,N_19931,N_19984);
or UO_137 (O_137,N_19930,N_19970);
and UO_138 (O_138,N_19839,N_19975);
nor UO_139 (O_139,N_19996,N_19876);
nor UO_140 (O_140,N_19979,N_19955);
xnor UO_141 (O_141,N_19984,N_19945);
xnor UO_142 (O_142,N_19868,N_19978);
nand UO_143 (O_143,N_19877,N_19933);
or UO_144 (O_144,N_19816,N_19793);
xor UO_145 (O_145,N_19968,N_19760);
and UO_146 (O_146,N_19777,N_19837);
or UO_147 (O_147,N_19785,N_19923);
nand UO_148 (O_148,N_19928,N_19961);
and UO_149 (O_149,N_19822,N_19975);
nor UO_150 (O_150,N_19981,N_19773);
nor UO_151 (O_151,N_19965,N_19789);
xnor UO_152 (O_152,N_19992,N_19866);
and UO_153 (O_153,N_19948,N_19926);
or UO_154 (O_154,N_19954,N_19922);
xor UO_155 (O_155,N_19848,N_19857);
nor UO_156 (O_156,N_19758,N_19909);
nand UO_157 (O_157,N_19883,N_19805);
xor UO_158 (O_158,N_19931,N_19752);
xnor UO_159 (O_159,N_19950,N_19794);
nor UO_160 (O_160,N_19928,N_19829);
or UO_161 (O_161,N_19822,N_19893);
or UO_162 (O_162,N_19800,N_19851);
nand UO_163 (O_163,N_19770,N_19802);
nor UO_164 (O_164,N_19833,N_19881);
nor UO_165 (O_165,N_19919,N_19787);
nand UO_166 (O_166,N_19984,N_19799);
xor UO_167 (O_167,N_19832,N_19790);
xor UO_168 (O_168,N_19947,N_19927);
and UO_169 (O_169,N_19805,N_19937);
xor UO_170 (O_170,N_19996,N_19932);
xor UO_171 (O_171,N_19993,N_19973);
or UO_172 (O_172,N_19805,N_19919);
nand UO_173 (O_173,N_19786,N_19789);
xnor UO_174 (O_174,N_19819,N_19796);
or UO_175 (O_175,N_19813,N_19980);
nand UO_176 (O_176,N_19877,N_19927);
xnor UO_177 (O_177,N_19839,N_19781);
or UO_178 (O_178,N_19982,N_19817);
and UO_179 (O_179,N_19783,N_19864);
nor UO_180 (O_180,N_19944,N_19929);
or UO_181 (O_181,N_19946,N_19973);
xnor UO_182 (O_182,N_19937,N_19836);
xnor UO_183 (O_183,N_19784,N_19868);
or UO_184 (O_184,N_19890,N_19802);
xor UO_185 (O_185,N_19990,N_19938);
nand UO_186 (O_186,N_19824,N_19898);
or UO_187 (O_187,N_19811,N_19984);
nor UO_188 (O_188,N_19842,N_19871);
xnor UO_189 (O_189,N_19924,N_19827);
nor UO_190 (O_190,N_19817,N_19767);
xnor UO_191 (O_191,N_19931,N_19975);
and UO_192 (O_192,N_19835,N_19909);
or UO_193 (O_193,N_19836,N_19751);
nand UO_194 (O_194,N_19786,N_19807);
or UO_195 (O_195,N_19885,N_19919);
and UO_196 (O_196,N_19858,N_19785);
and UO_197 (O_197,N_19823,N_19945);
nor UO_198 (O_198,N_19906,N_19922);
nor UO_199 (O_199,N_19999,N_19886);
nand UO_200 (O_200,N_19977,N_19954);
xor UO_201 (O_201,N_19964,N_19842);
nand UO_202 (O_202,N_19979,N_19839);
nor UO_203 (O_203,N_19795,N_19812);
nor UO_204 (O_204,N_19999,N_19945);
or UO_205 (O_205,N_19902,N_19822);
and UO_206 (O_206,N_19970,N_19939);
or UO_207 (O_207,N_19984,N_19804);
or UO_208 (O_208,N_19778,N_19997);
and UO_209 (O_209,N_19935,N_19900);
nor UO_210 (O_210,N_19880,N_19986);
and UO_211 (O_211,N_19763,N_19771);
or UO_212 (O_212,N_19982,N_19892);
or UO_213 (O_213,N_19900,N_19916);
xnor UO_214 (O_214,N_19974,N_19933);
xnor UO_215 (O_215,N_19823,N_19936);
or UO_216 (O_216,N_19760,N_19860);
and UO_217 (O_217,N_19992,N_19759);
nand UO_218 (O_218,N_19779,N_19762);
and UO_219 (O_219,N_19760,N_19798);
xor UO_220 (O_220,N_19859,N_19809);
or UO_221 (O_221,N_19756,N_19833);
or UO_222 (O_222,N_19857,N_19919);
and UO_223 (O_223,N_19989,N_19826);
or UO_224 (O_224,N_19992,N_19876);
and UO_225 (O_225,N_19997,N_19958);
nand UO_226 (O_226,N_19827,N_19932);
nor UO_227 (O_227,N_19947,N_19963);
or UO_228 (O_228,N_19839,N_19868);
nor UO_229 (O_229,N_19829,N_19838);
nand UO_230 (O_230,N_19757,N_19881);
nand UO_231 (O_231,N_19987,N_19935);
and UO_232 (O_232,N_19947,N_19751);
nand UO_233 (O_233,N_19947,N_19959);
nand UO_234 (O_234,N_19807,N_19826);
nor UO_235 (O_235,N_19789,N_19936);
xnor UO_236 (O_236,N_19899,N_19752);
nand UO_237 (O_237,N_19776,N_19974);
and UO_238 (O_238,N_19768,N_19946);
nand UO_239 (O_239,N_19754,N_19765);
xor UO_240 (O_240,N_19982,N_19893);
and UO_241 (O_241,N_19904,N_19783);
xor UO_242 (O_242,N_19992,N_19977);
nor UO_243 (O_243,N_19983,N_19922);
xnor UO_244 (O_244,N_19832,N_19782);
nand UO_245 (O_245,N_19935,N_19863);
or UO_246 (O_246,N_19830,N_19823);
or UO_247 (O_247,N_19834,N_19868);
or UO_248 (O_248,N_19997,N_19873);
and UO_249 (O_249,N_19781,N_19865);
nor UO_250 (O_250,N_19890,N_19760);
xnor UO_251 (O_251,N_19810,N_19927);
xor UO_252 (O_252,N_19995,N_19887);
nand UO_253 (O_253,N_19856,N_19868);
and UO_254 (O_254,N_19875,N_19956);
xnor UO_255 (O_255,N_19781,N_19950);
nand UO_256 (O_256,N_19947,N_19948);
nor UO_257 (O_257,N_19870,N_19829);
and UO_258 (O_258,N_19998,N_19806);
nand UO_259 (O_259,N_19965,N_19982);
nor UO_260 (O_260,N_19868,N_19976);
nand UO_261 (O_261,N_19992,N_19845);
nand UO_262 (O_262,N_19874,N_19952);
nand UO_263 (O_263,N_19787,N_19963);
or UO_264 (O_264,N_19765,N_19941);
nor UO_265 (O_265,N_19786,N_19976);
nor UO_266 (O_266,N_19867,N_19839);
nand UO_267 (O_267,N_19834,N_19867);
and UO_268 (O_268,N_19952,N_19834);
xnor UO_269 (O_269,N_19849,N_19879);
xor UO_270 (O_270,N_19986,N_19975);
or UO_271 (O_271,N_19908,N_19835);
nand UO_272 (O_272,N_19774,N_19846);
and UO_273 (O_273,N_19887,N_19871);
nand UO_274 (O_274,N_19904,N_19822);
xnor UO_275 (O_275,N_19857,N_19973);
nor UO_276 (O_276,N_19785,N_19780);
and UO_277 (O_277,N_19955,N_19899);
or UO_278 (O_278,N_19930,N_19773);
and UO_279 (O_279,N_19954,N_19869);
nor UO_280 (O_280,N_19918,N_19827);
xor UO_281 (O_281,N_19931,N_19933);
and UO_282 (O_282,N_19914,N_19889);
or UO_283 (O_283,N_19923,N_19879);
nor UO_284 (O_284,N_19823,N_19784);
or UO_285 (O_285,N_19958,N_19872);
and UO_286 (O_286,N_19772,N_19933);
nor UO_287 (O_287,N_19832,N_19861);
xnor UO_288 (O_288,N_19961,N_19932);
nand UO_289 (O_289,N_19804,N_19858);
or UO_290 (O_290,N_19863,N_19948);
nor UO_291 (O_291,N_19997,N_19866);
nor UO_292 (O_292,N_19979,N_19994);
and UO_293 (O_293,N_19954,N_19910);
nand UO_294 (O_294,N_19880,N_19827);
xor UO_295 (O_295,N_19926,N_19769);
nand UO_296 (O_296,N_19922,N_19927);
and UO_297 (O_297,N_19873,N_19789);
and UO_298 (O_298,N_19795,N_19843);
nor UO_299 (O_299,N_19750,N_19796);
nand UO_300 (O_300,N_19805,N_19864);
xnor UO_301 (O_301,N_19925,N_19837);
nor UO_302 (O_302,N_19958,N_19789);
nand UO_303 (O_303,N_19757,N_19944);
nor UO_304 (O_304,N_19852,N_19892);
or UO_305 (O_305,N_19913,N_19870);
nand UO_306 (O_306,N_19969,N_19799);
nand UO_307 (O_307,N_19947,N_19768);
xor UO_308 (O_308,N_19778,N_19791);
and UO_309 (O_309,N_19923,N_19855);
xnor UO_310 (O_310,N_19918,N_19848);
or UO_311 (O_311,N_19768,N_19938);
or UO_312 (O_312,N_19891,N_19978);
nand UO_313 (O_313,N_19821,N_19839);
nor UO_314 (O_314,N_19956,N_19879);
nor UO_315 (O_315,N_19888,N_19816);
xor UO_316 (O_316,N_19793,N_19845);
nor UO_317 (O_317,N_19941,N_19987);
and UO_318 (O_318,N_19934,N_19940);
nand UO_319 (O_319,N_19809,N_19769);
and UO_320 (O_320,N_19962,N_19883);
xor UO_321 (O_321,N_19883,N_19765);
and UO_322 (O_322,N_19886,N_19978);
and UO_323 (O_323,N_19912,N_19775);
or UO_324 (O_324,N_19856,N_19779);
xnor UO_325 (O_325,N_19770,N_19755);
or UO_326 (O_326,N_19930,N_19907);
and UO_327 (O_327,N_19847,N_19929);
xor UO_328 (O_328,N_19967,N_19907);
or UO_329 (O_329,N_19931,N_19760);
or UO_330 (O_330,N_19879,N_19872);
or UO_331 (O_331,N_19948,N_19931);
or UO_332 (O_332,N_19820,N_19873);
nand UO_333 (O_333,N_19792,N_19755);
nand UO_334 (O_334,N_19777,N_19858);
or UO_335 (O_335,N_19980,N_19785);
nor UO_336 (O_336,N_19845,N_19889);
or UO_337 (O_337,N_19805,N_19845);
nand UO_338 (O_338,N_19792,N_19874);
xnor UO_339 (O_339,N_19921,N_19858);
or UO_340 (O_340,N_19819,N_19978);
nor UO_341 (O_341,N_19753,N_19884);
and UO_342 (O_342,N_19762,N_19895);
nand UO_343 (O_343,N_19869,N_19992);
or UO_344 (O_344,N_19897,N_19912);
nand UO_345 (O_345,N_19863,N_19756);
nand UO_346 (O_346,N_19813,N_19899);
nor UO_347 (O_347,N_19812,N_19750);
nand UO_348 (O_348,N_19927,N_19813);
nand UO_349 (O_349,N_19856,N_19959);
nor UO_350 (O_350,N_19759,N_19808);
xor UO_351 (O_351,N_19802,N_19769);
or UO_352 (O_352,N_19772,N_19885);
nand UO_353 (O_353,N_19845,N_19953);
or UO_354 (O_354,N_19856,N_19925);
or UO_355 (O_355,N_19759,N_19959);
xnor UO_356 (O_356,N_19980,N_19825);
nor UO_357 (O_357,N_19992,N_19792);
nand UO_358 (O_358,N_19771,N_19789);
xor UO_359 (O_359,N_19990,N_19997);
xnor UO_360 (O_360,N_19880,N_19946);
and UO_361 (O_361,N_19877,N_19967);
or UO_362 (O_362,N_19771,N_19794);
nor UO_363 (O_363,N_19978,N_19956);
and UO_364 (O_364,N_19965,N_19832);
or UO_365 (O_365,N_19912,N_19870);
and UO_366 (O_366,N_19788,N_19806);
nor UO_367 (O_367,N_19848,N_19925);
and UO_368 (O_368,N_19908,N_19967);
or UO_369 (O_369,N_19932,N_19913);
nor UO_370 (O_370,N_19951,N_19818);
nand UO_371 (O_371,N_19854,N_19965);
xnor UO_372 (O_372,N_19991,N_19962);
nor UO_373 (O_373,N_19939,N_19957);
nand UO_374 (O_374,N_19769,N_19805);
and UO_375 (O_375,N_19787,N_19975);
and UO_376 (O_376,N_19797,N_19766);
or UO_377 (O_377,N_19800,N_19754);
nand UO_378 (O_378,N_19967,N_19977);
and UO_379 (O_379,N_19753,N_19996);
nand UO_380 (O_380,N_19800,N_19891);
xnor UO_381 (O_381,N_19896,N_19986);
and UO_382 (O_382,N_19954,N_19848);
or UO_383 (O_383,N_19857,N_19907);
nand UO_384 (O_384,N_19790,N_19880);
nor UO_385 (O_385,N_19844,N_19947);
nand UO_386 (O_386,N_19984,N_19857);
or UO_387 (O_387,N_19994,N_19766);
and UO_388 (O_388,N_19839,N_19799);
or UO_389 (O_389,N_19830,N_19880);
nor UO_390 (O_390,N_19929,N_19983);
nand UO_391 (O_391,N_19787,N_19985);
xor UO_392 (O_392,N_19827,N_19771);
or UO_393 (O_393,N_19979,N_19883);
xnor UO_394 (O_394,N_19830,N_19793);
nand UO_395 (O_395,N_19897,N_19938);
or UO_396 (O_396,N_19884,N_19804);
or UO_397 (O_397,N_19940,N_19835);
nor UO_398 (O_398,N_19921,N_19756);
or UO_399 (O_399,N_19878,N_19986);
nor UO_400 (O_400,N_19932,N_19917);
xnor UO_401 (O_401,N_19842,N_19883);
or UO_402 (O_402,N_19928,N_19974);
or UO_403 (O_403,N_19983,N_19768);
and UO_404 (O_404,N_19933,N_19932);
or UO_405 (O_405,N_19926,N_19771);
and UO_406 (O_406,N_19915,N_19823);
nor UO_407 (O_407,N_19971,N_19960);
or UO_408 (O_408,N_19958,N_19879);
nand UO_409 (O_409,N_19879,N_19782);
xnor UO_410 (O_410,N_19979,N_19949);
nor UO_411 (O_411,N_19897,N_19833);
or UO_412 (O_412,N_19815,N_19938);
nor UO_413 (O_413,N_19992,N_19789);
xor UO_414 (O_414,N_19944,N_19814);
or UO_415 (O_415,N_19857,N_19822);
or UO_416 (O_416,N_19864,N_19904);
or UO_417 (O_417,N_19839,N_19993);
nand UO_418 (O_418,N_19876,N_19845);
and UO_419 (O_419,N_19984,N_19866);
xor UO_420 (O_420,N_19930,N_19792);
or UO_421 (O_421,N_19837,N_19928);
or UO_422 (O_422,N_19908,N_19800);
nand UO_423 (O_423,N_19845,N_19762);
or UO_424 (O_424,N_19869,N_19772);
or UO_425 (O_425,N_19755,N_19983);
nor UO_426 (O_426,N_19950,N_19811);
xor UO_427 (O_427,N_19849,N_19966);
nand UO_428 (O_428,N_19885,N_19755);
nand UO_429 (O_429,N_19902,N_19787);
or UO_430 (O_430,N_19764,N_19810);
nor UO_431 (O_431,N_19848,N_19937);
or UO_432 (O_432,N_19775,N_19898);
nand UO_433 (O_433,N_19806,N_19809);
and UO_434 (O_434,N_19913,N_19752);
nor UO_435 (O_435,N_19950,N_19940);
nor UO_436 (O_436,N_19787,N_19842);
xnor UO_437 (O_437,N_19891,N_19877);
xnor UO_438 (O_438,N_19928,N_19959);
and UO_439 (O_439,N_19864,N_19961);
and UO_440 (O_440,N_19996,N_19916);
or UO_441 (O_441,N_19885,N_19892);
nor UO_442 (O_442,N_19859,N_19949);
or UO_443 (O_443,N_19786,N_19871);
and UO_444 (O_444,N_19873,N_19961);
and UO_445 (O_445,N_19858,N_19912);
xor UO_446 (O_446,N_19900,N_19764);
xor UO_447 (O_447,N_19861,N_19879);
and UO_448 (O_448,N_19831,N_19770);
and UO_449 (O_449,N_19832,N_19916);
and UO_450 (O_450,N_19840,N_19835);
nor UO_451 (O_451,N_19762,N_19999);
or UO_452 (O_452,N_19914,N_19811);
and UO_453 (O_453,N_19790,N_19907);
or UO_454 (O_454,N_19927,N_19995);
xor UO_455 (O_455,N_19810,N_19913);
nor UO_456 (O_456,N_19781,N_19959);
nand UO_457 (O_457,N_19912,N_19758);
nor UO_458 (O_458,N_19889,N_19987);
nor UO_459 (O_459,N_19861,N_19889);
and UO_460 (O_460,N_19870,N_19775);
nand UO_461 (O_461,N_19871,N_19970);
xor UO_462 (O_462,N_19941,N_19931);
nand UO_463 (O_463,N_19946,N_19759);
or UO_464 (O_464,N_19810,N_19957);
xnor UO_465 (O_465,N_19925,N_19842);
and UO_466 (O_466,N_19762,N_19905);
or UO_467 (O_467,N_19790,N_19820);
nand UO_468 (O_468,N_19943,N_19982);
xnor UO_469 (O_469,N_19851,N_19877);
or UO_470 (O_470,N_19755,N_19782);
and UO_471 (O_471,N_19930,N_19779);
or UO_472 (O_472,N_19900,N_19870);
nand UO_473 (O_473,N_19853,N_19933);
nor UO_474 (O_474,N_19779,N_19836);
or UO_475 (O_475,N_19925,N_19912);
xnor UO_476 (O_476,N_19796,N_19984);
nor UO_477 (O_477,N_19767,N_19997);
nor UO_478 (O_478,N_19944,N_19979);
and UO_479 (O_479,N_19778,N_19848);
nand UO_480 (O_480,N_19943,N_19967);
xor UO_481 (O_481,N_19949,N_19960);
nand UO_482 (O_482,N_19978,N_19838);
nor UO_483 (O_483,N_19892,N_19887);
and UO_484 (O_484,N_19892,N_19855);
or UO_485 (O_485,N_19832,N_19980);
or UO_486 (O_486,N_19976,N_19915);
nor UO_487 (O_487,N_19924,N_19857);
and UO_488 (O_488,N_19872,N_19933);
and UO_489 (O_489,N_19752,N_19793);
nor UO_490 (O_490,N_19902,N_19890);
or UO_491 (O_491,N_19922,N_19913);
nand UO_492 (O_492,N_19818,N_19930);
nand UO_493 (O_493,N_19846,N_19837);
and UO_494 (O_494,N_19786,N_19922);
nand UO_495 (O_495,N_19942,N_19763);
and UO_496 (O_496,N_19801,N_19856);
or UO_497 (O_497,N_19864,N_19856);
and UO_498 (O_498,N_19907,N_19973);
nand UO_499 (O_499,N_19875,N_19872);
and UO_500 (O_500,N_19982,N_19793);
or UO_501 (O_501,N_19952,N_19899);
nor UO_502 (O_502,N_19964,N_19828);
or UO_503 (O_503,N_19944,N_19787);
or UO_504 (O_504,N_19791,N_19783);
and UO_505 (O_505,N_19750,N_19799);
nor UO_506 (O_506,N_19939,N_19879);
nand UO_507 (O_507,N_19847,N_19969);
and UO_508 (O_508,N_19829,N_19900);
and UO_509 (O_509,N_19750,N_19883);
and UO_510 (O_510,N_19861,N_19758);
or UO_511 (O_511,N_19802,N_19819);
xor UO_512 (O_512,N_19853,N_19863);
nor UO_513 (O_513,N_19946,N_19963);
or UO_514 (O_514,N_19878,N_19985);
nor UO_515 (O_515,N_19921,N_19763);
nor UO_516 (O_516,N_19952,N_19835);
nand UO_517 (O_517,N_19914,N_19973);
or UO_518 (O_518,N_19925,N_19855);
nand UO_519 (O_519,N_19837,N_19939);
nor UO_520 (O_520,N_19980,N_19938);
nor UO_521 (O_521,N_19786,N_19852);
or UO_522 (O_522,N_19815,N_19973);
nand UO_523 (O_523,N_19828,N_19818);
and UO_524 (O_524,N_19788,N_19836);
and UO_525 (O_525,N_19788,N_19774);
nor UO_526 (O_526,N_19771,N_19938);
or UO_527 (O_527,N_19790,N_19855);
nor UO_528 (O_528,N_19787,N_19878);
xor UO_529 (O_529,N_19826,N_19811);
or UO_530 (O_530,N_19997,N_19799);
and UO_531 (O_531,N_19996,N_19806);
or UO_532 (O_532,N_19791,N_19968);
or UO_533 (O_533,N_19877,N_19864);
xnor UO_534 (O_534,N_19773,N_19945);
xnor UO_535 (O_535,N_19970,N_19897);
xor UO_536 (O_536,N_19830,N_19922);
or UO_537 (O_537,N_19958,N_19924);
and UO_538 (O_538,N_19950,N_19841);
nor UO_539 (O_539,N_19981,N_19902);
and UO_540 (O_540,N_19923,N_19824);
or UO_541 (O_541,N_19769,N_19851);
nand UO_542 (O_542,N_19983,N_19926);
nand UO_543 (O_543,N_19805,N_19921);
nor UO_544 (O_544,N_19943,N_19994);
nand UO_545 (O_545,N_19841,N_19818);
nor UO_546 (O_546,N_19942,N_19787);
xor UO_547 (O_547,N_19991,N_19856);
or UO_548 (O_548,N_19846,N_19804);
and UO_549 (O_549,N_19975,N_19935);
nor UO_550 (O_550,N_19960,N_19858);
or UO_551 (O_551,N_19938,N_19907);
nand UO_552 (O_552,N_19965,N_19784);
nand UO_553 (O_553,N_19837,N_19827);
nor UO_554 (O_554,N_19922,N_19965);
or UO_555 (O_555,N_19935,N_19791);
xor UO_556 (O_556,N_19975,N_19780);
and UO_557 (O_557,N_19951,N_19752);
nor UO_558 (O_558,N_19909,N_19990);
or UO_559 (O_559,N_19942,N_19777);
xor UO_560 (O_560,N_19961,N_19845);
and UO_561 (O_561,N_19775,N_19790);
or UO_562 (O_562,N_19975,N_19990);
and UO_563 (O_563,N_19849,N_19927);
nor UO_564 (O_564,N_19900,N_19833);
xor UO_565 (O_565,N_19908,N_19859);
and UO_566 (O_566,N_19938,N_19796);
and UO_567 (O_567,N_19759,N_19960);
xor UO_568 (O_568,N_19985,N_19897);
and UO_569 (O_569,N_19819,N_19866);
xnor UO_570 (O_570,N_19897,N_19887);
and UO_571 (O_571,N_19937,N_19827);
xor UO_572 (O_572,N_19866,N_19803);
nor UO_573 (O_573,N_19866,N_19929);
nand UO_574 (O_574,N_19990,N_19815);
and UO_575 (O_575,N_19913,N_19841);
and UO_576 (O_576,N_19944,N_19844);
nand UO_577 (O_577,N_19751,N_19828);
nand UO_578 (O_578,N_19899,N_19918);
nor UO_579 (O_579,N_19841,N_19755);
or UO_580 (O_580,N_19922,N_19862);
xor UO_581 (O_581,N_19931,N_19813);
nand UO_582 (O_582,N_19977,N_19792);
nand UO_583 (O_583,N_19918,N_19852);
xnor UO_584 (O_584,N_19971,N_19844);
xnor UO_585 (O_585,N_19796,N_19925);
nand UO_586 (O_586,N_19894,N_19767);
or UO_587 (O_587,N_19865,N_19912);
nand UO_588 (O_588,N_19925,N_19826);
xor UO_589 (O_589,N_19956,N_19868);
or UO_590 (O_590,N_19922,N_19979);
nor UO_591 (O_591,N_19912,N_19814);
xnor UO_592 (O_592,N_19802,N_19777);
nand UO_593 (O_593,N_19817,N_19883);
xor UO_594 (O_594,N_19941,N_19946);
nand UO_595 (O_595,N_19924,N_19917);
nor UO_596 (O_596,N_19944,N_19833);
xor UO_597 (O_597,N_19800,N_19922);
xnor UO_598 (O_598,N_19844,N_19836);
xor UO_599 (O_599,N_19947,N_19770);
nor UO_600 (O_600,N_19872,N_19871);
xor UO_601 (O_601,N_19988,N_19898);
or UO_602 (O_602,N_19762,N_19873);
or UO_603 (O_603,N_19783,N_19835);
or UO_604 (O_604,N_19797,N_19862);
and UO_605 (O_605,N_19802,N_19851);
and UO_606 (O_606,N_19881,N_19775);
nand UO_607 (O_607,N_19844,N_19980);
xor UO_608 (O_608,N_19867,N_19889);
nand UO_609 (O_609,N_19980,N_19771);
xor UO_610 (O_610,N_19821,N_19794);
and UO_611 (O_611,N_19999,N_19835);
xor UO_612 (O_612,N_19769,N_19751);
xor UO_613 (O_613,N_19760,N_19841);
and UO_614 (O_614,N_19938,N_19813);
or UO_615 (O_615,N_19831,N_19825);
nand UO_616 (O_616,N_19850,N_19985);
nor UO_617 (O_617,N_19836,N_19830);
nor UO_618 (O_618,N_19827,N_19968);
nand UO_619 (O_619,N_19909,N_19974);
nor UO_620 (O_620,N_19903,N_19778);
nand UO_621 (O_621,N_19844,N_19770);
and UO_622 (O_622,N_19869,N_19974);
or UO_623 (O_623,N_19768,N_19827);
and UO_624 (O_624,N_19992,N_19885);
xnor UO_625 (O_625,N_19912,N_19857);
nor UO_626 (O_626,N_19867,N_19949);
and UO_627 (O_627,N_19940,N_19759);
nand UO_628 (O_628,N_19779,N_19791);
nand UO_629 (O_629,N_19944,N_19772);
and UO_630 (O_630,N_19978,N_19791);
and UO_631 (O_631,N_19824,N_19895);
and UO_632 (O_632,N_19839,N_19855);
or UO_633 (O_633,N_19811,N_19869);
or UO_634 (O_634,N_19915,N_19754);
nand UO_635 (O_635,N_19783,N_19907);
nand UO_636 (O_636,N_19986,N_19861);
nor UO_637 (O_637,N_19841,N_19897);
nand UO_638 (O_638,N_19759,N_19854);
xnor UO_639 (O_639,N_19924,N_19869);
nor UO_640 (O_640,N_19971,N_19773);
xor UO_641 (O_641,N_19950,N_19776);
and UO_642 (O_642,N_19768,N_19837);
and UO_643 (O_643,N_19827,N_19821);
or UO_644 (O_644,N_19886,N_19804);
and UO_645 (O_645,N_19752,N_19902);
or UO_646 (O_646,N_19916,N_19887);
and UO_647 (O_647,N_19940,N_19898);
xnor UO_648 (O_648,N_19994,N_19933);
nor UO_649 (O_649,N_19851,N_19821);
nand UO_650 (O_650,N_19839,N_19767);
nor UO_651 (O_651,N_19750,N_19952);
and UO_652 (O_652,N_19767,N_19783);
or UO_653 (O_653,N_19994,N_19931);
nor UO_654 (O_654,N_19765,N_19872);
xor UO_655 (O_655,N_19812,N_19882);
or UO_656 (O_656,N_19863,N_19809);
nor UO_657 (O_657,N_19981,N_19887);
xor UO_658 (O_658,N_19894,N_19818);
nor UO_659 (O_659,N_19750,N_19761);
nor UO_660 (O_660,N_19991,N_19751);
nand UO_661 (O_661,N_19993,N_19849);
xor UO_662 (O_662,N_19854,N_19904);
and UO_663 (O_663,N_19924,N_19848);
xnor UO_664 (O_664,N_19884,N_19817);
and UO_665 (O_665,N_19891,N_19820);
or UO_666 (O_666,N_19972,N_19994);
or UO_667 (O_667,N_19868,N_19891);
nand UO_668 (O_668,N_19992,N_19857);
nor UO_669 (O_669,N_19840,N_19893);
nand UO_670 (O_670,N_19814,N_19988);
xor UO_671 (O_671,N_19793,N_19813);
xor UO_672 (O_672,N_19964,N_19809);
and UO_673 (O_673,N_19939,N_19807);
xnor UO_674 (O_674,N_19783,N_19804);
nand UO_675 (O_675,N_19935,N_19973);
nand UO_676 (O_676,N_19971,N_19914);
nand UO_677 (O_677,N_19952,N_19833);
nand UO_678 (O_678,N_19980,N_19936);
xnor UO_679 (O_679,N_19956,N_19950);
or UO_680 (O_680,N_19891,N_19795);
nand UO_681 (O_681,N_19808,N_19885);
xnor UO_682 (O_682,N_19963,N_19979);
nand UO_683 (O_683,N_19992,N_19802);
or UO_684 (O_684,N_19828,N_19927);
nand UO_685 (O_685,N_19901,N_19806);
or UO_686 (O_686,N_19895,N_19823);
xnor UO_687 (O_687,N_19875,N_19950);
and UO_688 (O_688,N_19907,N_19892);
and UO_689 (O_689,N_19913,N_19852);
or UO_690 (O_690,N_19959,N_19753);
nor UO_691 (O_691,N_19961,N_19828);
or UO_692 (O_692,N_19965,N_19753);
or UO_693 (O_693,N_19879,N_19877);
and UO_694 (O_694,N_19932,N_19906);
nand UO_695 (O_695,N_19802,N_19785);
nand UO_696 (O_696,N_19881,N_19823);
and UO_697 (O_697,N_19778,N_19995);
nor UO_698 (O_698,N_19762,N_19925);
and UO_699 (O_699,N_19994,N_19824);
nand UO_700 (O_700,N_19940,N_19827);
nor UO_701 (O_701,N_19790,N_19896);
nor UO_702 (O_702,N_19927,N_19951);
nand UO_703 (O_703,N_19997,N_19882);
or UO_704 (O_704,N_19815,N_19955);
and UO_705 (O_705,N_19901,N_19953);
xnor UO_706 (O_706,N_19857,N_19961);
and UO_707 (O_707,N_19830,N_19959);
or UO_708 (O_708,N_19802,N_19774);
and UO_709 (O_709,N_19906,N_19828);
nor UO_710 (O_710,N_19758,N_19989);
and UO_711 (O_711,N_19862,N_19859);
xor UO_712 (O_712,N_19754,N_19775);
and UO_713 (O_713,N_19902,N_19810);
or UO_714 (O_714,N_19897,N_19977);
and UO_715 (O_715,N_19891,N_19776);
nor UO_716 (O_716,N_19866,N_19770);
and UO_717 (O_717,N_19770,N_19876);
nor UO_718 (O_718,N_19930,N_19781);
or UO_719 (O_719,N_19829,N_19805);
and UO_720 (O_720,N_19842,N_19832);
xnor UO_721 (O_721,N_19911,N_19784);
nor UO_722 (O_722,N_19981,N_19928);
xnor UO_723 (O_723,N_19928,N_19969);
nand UO_724 (O_724,N_19997,N_19869);
nand UO_725 (O_725,N_19795,N_19837);
xor UO_726 (O_726,N_19921,N_19930);
nor UO_727 (O_727,N_19961,N_19901);
xnor UO_728 (O_728,N_19757,N_19947);
or UO_729 (O_729,N_19952,N_19970);
xnor UO_730 (O_730,N_19841,N_19919);
nor UO_731 (O_731,N_19950,N_19849);
xnor UO_732 (O_732,N_19794,N_19826);
or UO_733 (O_733,N_19906,N_19959);
and UO_734 (O_734,N_19863,N_19845);
nor UO_735 (O_735,N_19900,N_19797);
nor UO_736 (O_736,N_19915,N_19815);
nor UO_737 (O_737,N_19889,N_19895);
and UO_738 (O_738,N_19859,N_19988);
nor UO_739 (O_739,N_19823,N_19814);
xnor UO_740 (O_740,N_19966,N_19841);
or UO_741 (O_741,N_19953,N_19941);
xor UO_742 (O_742,N_19855,N_19982);
or UO_743 (O_743,N_19861,N_19823);
nor UO_744 (O_744,N_19875,N_19889);
xor UO_745 (O_745,N_19860,N_19885);
or UO_746 (O_746,N_19931,N_19946);
or UO_747 (O_747,N_19797,N_19909);
or UO_748 (O_748,N_19879,N_19834);
or UO_749 (O_749,N_19831,N_19934);
or UO_750 (O_750,N_19982,N_19812);
or UO_751 (O_751,N_19840,N_19764);
xor UO_752 (O_752,N_19913,N_19815);
nor UO_753 (O_753,N_19946,N_19996);
and UO_754 (O_754,N_19832,N_19778);
xnor UO_755 (O_755,N_19943,N_19986);
nand UO_756 (O_756,N_19923,N_19781);
nand UO_757 (O_757,N_19894,N_19927);
nand UO_758 (O_758,N_19863,N_19897);
nor UO_759 (O_759,N_19809,N_19932);
or UO_760 (O_760,N_19762,N_19940);
and UO_761 (O_761,N_19909,N_19826);
nand UO_762 (O_762,N_19812,N_19846);
and UO_763 (O_763,N_19910,N_19867);
xnor UO_764 (O_764,N_19943,N_19883);
xnor UO_765 (O_765,N_19834,N_19842);
or UO_766 (O_766,N_19836,N_19784);
and UO_767 (O_767,N_19791,N_19887);
and UO_768 (O_768,N_19821,N_19788);
and UO_769 (O_769,N_19870,N_19909);
nor UO_770 (O_770,N_19880,N_19811);
nor UO_771 (O_771,N_19955,N_19759);
and UO_772 (O_772,N_19837,N_19852);
nor UO_773 (O_773,N_19982,N_19824);
or UO_774 (O_774,N_19828,N_19907);
nor UO_775 (O_775,N_19775,N_19906);
nand UO_776 (O_776,N_19766,N_19805);
xnor UO_777 (O_777,N_19866,N_19811);
xor UO_778 (O_778,N_19954,N_19875);
nor UO_779 (O_779,N_19759,N_19761);
and UO_780 (O_780,N_19936,N_19788);
or UO_781 (O_781,N_19915,N_19854);
and UO_782 (O_782,N_19789,N_19893);
nor UO_783 (O_783,N_19750,N_19882);
nor UO_784 (O_784,N_19781,N_19778);
and UO_785 (O_785,N_19795,N_19933);
nand UO_786 (O_786,N_19908,N_19758);
nand UO_787 (O_787,N_19882,N_19918);
nor UO_788 (O_788,N_19872,N_19776);
or UO_789 (O_789,N_19859,N_19836);
xnor UO_790 (O_790,N_19968,N_19759);
or UO_791 (O_791,N_19815,N_19898);
xor UO_792 (O_792,N_19984,N_19915);
nand UO_793 (O_793,N_19750,N_19801);
and UO_794 (O_794,N_19775,N_19806);
or UO_795 (O_795,N_19884,N_19890);
nor UO_796 (O_796,N_19773,N_19751);
and UO_797 (O_797,N_19972,N_19760);
nor UO_798 (O_798,N_19768,N_19996);
nand UO_799 (O_799,N_19996,N_19887);
nand UO_800 (O_800,N_19931,N_19861);
nand UO_801 (O_801,N_19909,N_19809);
or UO_802 (O_802,N_19914,N_19775);
xor UO_803 (O_803,N_19785,N_19876);
nor UO_804 (O_804,N_19766,N_19967);
xnor UO_805 (O_805,N_19896,N_19921);
nor UO_806 (O_806,N_19819,N_19753);
nor UO_807 (O_807,N_19779,N_19969);
and UO_808 (O_808,N_19850,N_19828);
xnor UO_809 (O_809,N_19927,N_19788);
nand UO_810 (O_810,N_19893,N_19805);
and UO_811 (O_811,N_19958,N_19793);
xnor UO_812 (O_812,N_19937,N_19759);
nor UO_813 (O_813,N_19752,N_19816);
nor UO_814 (O_814,N_19932,N_19943);
or UO_815 (O_815,N_19839,N_19780);
or UO_816 (O_816,N_19759,N_19990);
nor UO_817 (O_817,N_19977,N_19843);
xor UO_818 (O_818,N_19784,N_19809);
xor UO_819 (O_819,N_19949,N_19932);
and UO_820 (O_820,N_19793,N_19912);
xnor UO_821 (O_821,N_19751,N_19914);
and UO_822 (O_822,N_19833,N_19795);
or UO_823 (O_823,N_19870,N_19750);
and UO_824 (O_824,N_19904,N_19914);
or UO_825 (O_825,N_19773,N_19834);
nand UO_826 (O_826,N_19975,N_19951);
or UO_827 (O_827,N_19907,N_19819);
and UO_828 (O_828,N_19823,N_19963);
or UO_829 (O_829,N_19941,N_19750);
or UO_830 (O_830,N_19804,N_19906);
nor UO_831 (O_831,N_19922,N_19823);
nand UO_832 (O_832,N_19843,N_19756);
or UO_833 (O_833,N_19995,N_19756);
and UO_834 (O_834,N_19765,N_19820);
or UO_835 (O_835,N_19847,N_19901);
nand UO_836 (O_836,N_19906,N_19972);
or UO_837 (O_837,N_19975,N_19925);
xor UO_838 (O_838,N_19826,N_19790);
or UO_839 (O_839,N_19941,N_19998);
nand UO_840 (O_840,N_19908,N_19815);
and UO_841 (O_841,N_19792,N_19785);
nand UO_842 (O_842,N_19819,N_19919);
nand UO_843 (O_843,N_19979,N_19986);
xor UO_844 (O_844,N_19973,N_19812);
nand UO_845 (O_845,N_19860,N_19985);
or UO_846 (O_846,N_19899,N_19849);
or UO_847 (O_847,N_19754,N_19967);
nand UO_848 (O_848,N_19844,N_19936);
or UO_849 (O_849,N_19920,N_19788);
and UO_850 (O_850,N_19834,N_19766);
nor UO_851 (O_851,N_19811,N_19887);
or UO_852 (O_852,N_19814,N_19865);
or UO_853 (O_853,N_19805,N_19857);
and UO_854 (O_854,N_19890,N_19862);
or UO_855 (O_855,N_19783,N_19917);
or UO_856 (O_856,N_19792,N_19891);
nor UO_857 (O_857,N_19861,N_19961);
nand UO_858 (O_858,N_19782,N_19913);
and UO_859 (O_859,N_19987,N_19825);
xnor UO_860 (O_860,N_19832,N_19879);
nand UO_861 (O_861,N_19805,N_19832);
nand UO_862 (O_862,N_19869,N_19922);
xnor UO_863 (O_863,N_19971,N_19891);
nor UO_864 (O_864,N_19860,N_19991);
xor UO_865 (O_865,N_19940,N_19754);
nand UO_866 (O_866,N_19831,N_19916);
nand UO_867 (O_867,N_19910,N_19779);
xor UO_868 (O_868,N_19910,N_19911);
or UO_869 (O_869,N_19873,N_19819);
nand UO_870 (O_870,N_19934,N_19901);
and UO_871 (O_871,N_19898,N_19821);
nor UO_872 (O_872,N_19911,N_19869);
or UO_873 (O_873,N_19905,N_19765);
or UO_874 (O_874,N_19765,N_19809);
and UO_875 (O_875,N_19777,N_19964);
nor UO_876 (O_876,N_19953,N_19956);
nor UO_877 (O_877,N_19967,N_19858);
and UO_878 (O_878,N_19952,N_19860);
or UO_879 (O_879,N_19827,N_19807);
or UO_880 (O_880,N_19882,N_19751);
nand UO_881 (O_881,N_19952,N_19785);
or UO_882 (O_882,N_19778,N_19792);
or UO_883 (O_883,N_19988,N_19904);
nand UO_884 (O_884,N_19861,N_19768);
xnor UO_885 (O_885,N_19760,N_19806);
nand UO_886 (O_886,N_19981,N_19912);
nand UO_887 (O_887,N_19954,N_19827);
or UO_888 (O_888,N_19988,N_19834);
xor UO_889 (O_889,N_19895,N_19959);
nor UO_890 (O_890,N_19860,N_19862);
xnor UO_891 (O_891,N_19785,N_19795);
nor UO_892 (O_892,N_19764,N_19939);
xor UO_893 (O_893,N_19871,N_19770);
or UO_894 (O_894,N_19934,N_19955);
xnor UO_895 (O_895,N_19864,N_19923);
or UO_896 (O_896,N_19808,N_19967);
or UO_897 (O_897,N_19863,N_19769);
or UO_898 (O_898,N_19787,N_19870);
nand UO_899 (O_899,N_19757,N_19774);
and UO_900 (O_900,N_19859,N_19961);
or UO_901 (O_901,N_19935,N_19869);
and UO_902 (O_902,N_19789,N_19777);
and UO_903 (O_903,N_19830,N_19858);
or UO_904 (O_904,N_19942,N_19940);
and UO_905 (O_905,N_19967,N_19809);
or UO_906 (O_906,N_19999,N_19877);
xnor UO_907 (O_907,N_19850,N_19769);
and UO_908 (O_908,N_19857,N_19948);
xor UO_909 (O_909,N_19834,N_19916);
nor UO_910 (O_910,N_19961,N_19800);
nor UO_911 (O_911,N_19874,N_19866);
or UO_912 (O_912,N_19921,N_19959);
xor UO_913 (O_913,N_19773,N_19901);
or UO_914 (O_914,N_19882,N_19768);
or UO_915 (O_915,N_19998,N_19837);
or UO_916 (O_916,N_19783,N_19854);
and UO_917 (O_917,N_19770,N_19783);
nand UO_918 (O_918,N_19993,N_19877);
xor UO_919 (O_919,N_19996,N_19878);
and UO_920 (O_920,N_19886,N_19752);
nor UO_921 (O_921,N_19934,N_19873);
and UO_922 (O_922,N_19929,N_19822);
or UO_923 (O_923,N_19875,N_19920);
nor UO_924 (O_924,N_19822,N_19923);
xor UO_925 (O_925,N_19843,N_19771);
and UO_926 (O_926,N_19963,N_19761);
xor UO_927 (O_927,N_19882,N_19963);
and UO_928 (O_928,N_19778,N_19875);
or UO_929 (O_929,N_19819,N_19824);
nor UO_930 (O_930,N_19754,N_19809);
nand UO_931 (O_931,N_19975,N_19877);
xnor UO_932 (O_932,N_19861,N_19992);
nand UO_933 (O_933,N_19989,N_19797);
or UO_934 (O_934,N_19759,N_19842);
nand UO_935 (O_935,N_19821,N_19860);
nand UO_936 (O_936,N_19992,N_19754);
nor UO_937 (O_937,N_19807,N_19879);
nand UO_938 (O_938,N_19788,N_19993);
xnor UO_939 (O_939,N_19751,N_19846);
xnor UO_940 (O_940,N_19813,N_19897);
nand UO_941 (O_941,N_19814,N_19844);
or UO_942 (O_942,N_19864,N_19947);
and UO_943 (O_943,N_19938,N_19947);
or UO_944 (O_944,N_19871,N_19766);
and UO_945 (O_945,N_19926,N_19995);
nand UO_946 (O_946,N_19864,N_19953);
and UO_947 (O_947,N_19955,N_19782);
or UO_948 (O_948,N_19896,N_19845);
xnor UO_949 (O_949,N_19870,N_19986);
xor UO_950 (O_950,N_19861,N_19983);
and UO_951 (O_951,N_19959,N_19792);
nor UO_952 (O_952,N_19974,N_19760);
and UO_953 (O_953,N_19900,N_19800);
or UO_954 (O_954,N_19819,N_19812);
xnor UO_955 (O_955,N_19778,N_19884);
nor UO_956 (O_956,N_19966,N_19809);
or UO_957 (O_957,N_19866,N_19862);
and UO_958 (O_958,N_19796,N_19980);
nor UO_959 (O_959,N_19973,N_19898);
nand UO_960 (O_960,N_19813,N_19923);
nand UO_961 (O_961,N_19905,N_19829);
xnor UO_962 (O_962,N_19936,N_19773);
nand UO_963 (O_963,N_19822,N_19940);
xor UO_964 (O_964,N_19834,N_19783);
nor UO_965 (O_965,N_19881,N_19826);
and UO_966 (O_966,N_19858,N_19890);
or UO_967 (O_967,N_19809,N_19910);
nand UO_968 (O_968,N_19970,N_19942);
nand UO_969 (O_969,N_19823,N_19827);
and UO_970 (O_970,N_19897,N_19998);
and UO_971 (O_971,N_19817,N_19790);
nor UO_972 (O_972,N_19881,N_19809);
nand UO_973 (O_973,N_19955,N_19804);
nor UO_974 (O_974,N_19943,N_19981);
and UO_975 (O_975,N_19763,N_19754);
xnor UO_976 (O_976,N_19955,N_19950);
or UO_977 (O_977,N_19799,N_19938);
and UO_978 (O_978,N_19753,N_19772);
or UO_979 (O_979,N_19923,N_19900);
xor UO_980 (O_980,N_19967,N_19821);
nor UO_981 (O_981,N_19797,N_19954);
xnor UO_982 (O_982,N_19946,N_19784);
nor UO_983 (O_983,N_19937,N_19936);
nor UO_984 (O_984,N_19760,N_19981);
and UO_985 (O_985,N_19871,N_19760);
and UO_986 (O_986,N_19789,N_19844);
and UO_987 (O_987,N_19921,N_19823);
and UO_988 (O_988,N_19761,N_19985);
nor UO_989 (O_989,N_19945,N_19927);
xnor UO_990 (O_990,N_19865,N_19889);
nand UO_991 (O_991,N_19758,N_19869);
nor UO_992 (O_992,N_19838,N_19968);
or UO_993 (O_993,N_19957,N_19779);
nor UO_994 (O_994,N_19929,N_19845);
nand UO_995 (O_995,N_19889,N_19911);
and UO_996 (O_996,N_19974,N_19891);
nor UO_997 (O_997,N_19975,N_19852);
xor UO_998 (O_998,N_19924,N_19933);
or UO_999 (O_999,N_19812,N_19976);
or UO_1000 (O_1000,N_19967,N_19776);
nor UO_1001 (O_1001,N_19802,N_19834);
nor UO_1002 (O_1002,N_19989,N_19829);
nor UO_1003 (O_1003,N_19935,N_19954);
nand UO_1004 (O_1004,N_19971,N_19915);
nor UO_1005 (O_1005,N_19883,N_19852);
and UO_1006 (O_1006,N_19820,N_19892);
xor UO_1007 (O_1007,N_19883,N_19849);
nand UO_1008 (O_1008,N_19822,N_19914);
xnor UO_1009 (O_1009,N_19947,N_19923);
or UO_1010 (O_1010,N_19792,N_19823);
xor UO_1011 (O_1011,N_19875,N_19791);
xor UO_1012 (O_1012,N_19980,N_19967);
and UO_1013 (O_1013,N_19975,N_19979);
nor UO_1014 (O_1014,N_19790,N_19988);
xnor UO_1015 (O_1015,N_19875,N_19892);
xnor UO_1016 (O_1016,N_19858,N_19988);
nand UO_1017 (O_1017,N_19795,N_19907);
and UO_1018 (O_1018,N_19884,N_19880);
xor UO_1019 (O_1019,N_19840,N_19849);
nand UO_1020 (O_1020,N_19914,N_19842);
nor UO_1021 (O_1021,N_19832,N_19826);
xor UO_1022 (O_1022,N_19973,N_19896);
nor UO_1023 (O_1023,N_19887,N_19842);
nand UO_1024 (O_1024,N_19789,N_19829);
nand UO_1025 (O_1025,N_19768,N_19761);
nor UO_1026 (O_1026,N_19980,N_19852);
nor UO_1027 (O_1027,N_19992,N_19819);
or UO_1028 (O_1028,N_19952,N_19915);
nand UO_1029 (O_1029,N_19803,N_19852);
xnor UO_1030 (O_1030,N_19842,N_19775);
or UO_1031 (O_1031,N_19962,N_19780);
or UO_1032 (O_1032,N_19759,N_19998);
xnor UO_1033 (O_1033,N_19959,N_19890);
nand UO_1034 (O_1034,N_19936,N_19808);
xnor UO_1035 (O_1035,N_19901,N_19954);
or UO_1036 (O_1036,N_19890,N_19783);
xnor UO_1037 (O_1037,N_19766,N_19791);
and UO_1038 (O_1038,N_19787,N_19956);
xor UO_1039 (O_1039,N_19799,N_19924);
and UO_1040 (O_1040,N_19976,N_19861);
nand UO_1041 (O_1041,N_19843,N_19925);
or UO_1042 (O_1042,N_19988,N_19850);
xor UO_1043 (O_1043,N_19776,N_19982);
xor UO_1044 (O_1044,N_19966,N_19978);
nor UO_1045 (O_1045,N_19929,N_19776);
nor UO_1046 (O_1046,N_19762,N_19829);
or UO_1047 (O_1047,N_19882,N_19890);
nand UO_1048 (O_1048,N_19835,N_19868);
nor UO_1049 (O_1049,N_19781,N_19915);
or UO_1050 (O_1050,N_19895,N_19904);
xnor UO_1051 (O_1051,N_19824,N_19826);
xor UO_1052 (O_1052,N_19786,N_19756);
xnor UO_1053 (O_1053,N_19929,N_19834);
nor UO_1054 (O_1054,N_19816,N_19773);
or UO_1055 (O_1055,N_19869,N_19827);
xnor UO_1056 (O_1056,N_19799,N_19814);
and UO_1057 (O_1057,N_19978,N_19756);
xor UO_1058 (O_1058,N_19849,N_19907);
nand UO_1059 (O_1059,N_19900,N_19869);
nand UO_1060 (O_1060,N_19771,N_19912);
and UO_1061 (O_1061,N_19979,N_19797);
xor UO_1062 (O_1062,N_19818,N_19833);
nand UO_1063 (O_1063,N_19883,N_19895);
xnor UO_1064 (O_1064,N_19832,N_19897);
xor UO_1065 (O_1065,N_19951,N_19948);
or UO_1066 (O_1066,N_19973,N_19869);
nor UO_1067 (O_1067,N_19884,N_19807);
nor UO_1068 (O_1068,N_19985,N_19981);
xnor UO_1069 (O_1069,N_19771,N_19952);
or UO_1070 (O_1070,N_19830,N_19826);
and UO_1071 (O_1071,N_19907,N_19886);
xor UO_1072 (O_1072,N_19901,N_19986);
and UO_1073 (O_1073,N_19990,N_19890);
and UO_1074 (O_1074,N_19758,N_19819);
or UO_1075 (O_1075,N_19752,N_19779);
and UO_1076 (O_1076,N_19839,N_19960);
or UO_1077 (O_1077,N_19993,N_19853);
or UO_1078 (O_1078,N_19904,N_19928);
nor UO_1079 (O_1079,N_19814,N_19819);
xnor UO_1080 (O_1080,N_19945,N_19995);
nand UO_1081 (O_1081,N_19885,N_19848);
nand UO_1082 (O_1082,N_19895,N_19914);
and UO_1083 (O_1083,N_19888,N_19928);
xnor UO_1084 (O_1084,N_19983,N_19807);
nand UO_1085 (O_1085,N_19825,N_19939);
or UO_1086 (O_1086,N_19768,N_19842);
nor UO_1087 (O_1087,N_19958,N_19906);
or UO_1088 (O_1088,N_19847,N_19985);
nor UO_1089 (O_1089,N_19800,N_19824);
or UO_1090 (O_1090,N_19768,N_19989);
nand UO_1091 (O_1091,N_19952,N_19887);
nand UO_1092 (O_1092,N_19863,N_19832);
nor UO_1093 (O_1093,N_19795,N_19950);
and UO_1094 (O_1094,N_19997,N_19936);
or UO_1095 (O_1095,N_19915,N_19776);
xor UO_1096 (O_1096,N_19991,N_19926);
nor UO_1097 (O_1097,N_19990,N_19923);
or UO_1098 (O_1098,N_19783,N_19998);
or UO_1099 (O_1099,N_19999,N_19853);
xnor UO_1100 (O_1100,N_19969,N_19919);
or UO_1101 (O_1101,N_19762,N_19868);
and UO_1102 (O_1102,N_19819,N_19800);
nor UO_1103 (O_1103,N_19766,N_19855);
nand UO_1104 (O_1104,N_19774,N_19929);
xnor UO_1105 (O_1105,N_19775,N_19872);
xor UO_1106 (O_1106,N_19850,N_19840);
and UO_1107 (O_1107,N_19971,N_19921);
and UO_1108 (O_1108,N_19855,N_19849);
and UO_1109 (O_1109,N_19771,N_19814);
and UO_1110 (O_1110,N_19842,N_19772);
and UO_1111 (O_1111,N_19791,N_19802);
nor UO_1112 (O_1112,N_19843,N_19904);
xor UO_1113 (O_1113,N_19958,N_19776);
and UO_1114 (O_1114,N_19896,N_19864);
xor UO_1115 (O_1115,N_19809,N_19826);
and UO_1116 (O_1116,N_19850,N_19979);
and UO_1117 (O_1117,N_19769,N_19895);
nand UO_1118 (O_1118,N_19911,N_19945);
nand UO_1119 (O_1119,N_19949,N_19887);
or UO_1120 (O_1120,N_19860,N_19923);
nor UO_1121 (O_1121,N_19871,N_19831);
or UO_1122 (O_1122,N_19901,N_19768);
or UO_1123 (O_1123,N_19902,N_19796);
and UO_1124 (O_1124,N_19994,N_19892);
xnor UO_1125 (O_1125,N_19796,N_19820);
nor UO_1126 (O_1126,N_19963,N_19754);
or UO_1127 (O_1127,N_19829,N_19957);
or UO_1128 (O_1128,N_19843,N_19803);
nor UO_1129 (O_1129,N_19850,N_19903);
nor UO_1130 (O_1130,N_19968,N_19859);
and UO_1131 (O_1131,N_19897,N_19769);
nor UO_1132 (O_1132,N_19800,N_19822);
nand UO_1133 (O_1133,N_19954,N_19782);
or UO_1134 (O_1134,N_19790,N_19892);
nand UO_1135 (O_1135,N_19860,N_19820);
and UO_1136 (O_1136,N_19918,N_19943);
or UO_1137 (O_1137,N_19780,N_19832);
nand UO_1138 (O_1138,N_19770,N_19781);
and UO_1139 (O_1139,N_19988,N_19794);
or UO_1140 (O_1140,N_19915,N_19945);
and UO_1141 (O_1141,N_19778,N_19758);
or UO_1142 (O_1142,N_19951,N_19999);
and UO_1143 (O_1143,N_19909,N_19985);
xnor UO_1144 (O_1144,N_19852,N_19791);
nor UO_1145 (O_1145,N_19797,N_19962);
or UO_1146 (O_1146,N_19965,N_19809);
and UO_1147 (O_1147,N_19803,N_19849);
and UO_1148 (O_1148,N_19878,N_19809);
nor UO_1149 (O_1149,N_19988,N_19887);
nor UO_1150 (O_1150,N_19769,N_19784);
nor UO_1151 (O_1151,N_19819,N_19847);
and UO_1152 (O_1152,N_19835,N_19955);
nand UO_1153 (O_1153,N_19788,N_19982);
xnor UO_1154 (O_1154,N_19917,N_19834);
and UO_1155 (O_1155,N_19764,N_19938);
nor UO_1156 (O_1156,N_19971,N_19783);
xnor UO_1157 (O_1157,N_19806,N_19977);
nor UO_1158 (O_1158,N_19924,N_19920);
and UO_1159 (O_1159,N_19984,N_19777);
xor UO_1160 (O_1160,N_19757,N_19780);
nor UO_1161 (O_1161,N_19844,N_19831);
nor UO_1162 (O_1162,N_19752,N_19950);
or UO_1163 (O_1163,N_19989,N_19939);
xnor UO_1164 (O_1164,N_19797,N_19802);
and UO_1165 (O_1165,N_19849,N_19957);
or UO_1166 (O_1166,N_19829,N_19982);
nand UO_1167 (O_1167,N_19761,N_19869);
xor UO_1168 (O_1168,N_19997,N_19976);
nor UO_1169 (O_1169,N_19889,N_19923);
nand UO_1170 (O_1170,N_19802,N_19762);
or UO_1171 (O_1171,N_19897,N_19825);
nand UO_1172 (O_1172,N_19818,N_19864);
and UO_1173 (O_1173,N_19985,N_19882);
xor UO_1174 (O_1174,N_19796,N_19956);
nand UO_1175 (O_1175,N_19894,N_19792);
or UO_1176 (O_1176,N_19803,N_19862);
nor UO_1177 (O_1177,N_19906,N_19766);
nor UO_1178 (O_1178,N_19821,N_19847);
or UO_1179 (O_1179,N_19893,N_19879);
nor UO_1180 (O_1180,N_19839,N_19823);
xor UO_1181 (O_1181,N_19805,N_19976);
or UO_1182 (O_1182,N_19972,N_19995);
xnor UO_1183 (O_1183,N_19846,N_19893);
nand UO_1184 (O_1184,N_19875,N_19781);
xor UO_1185 (O_1185,N_19840,N_19852);
or UO_1186 (O_1186,N_19969,N_19778);
nand UO_1187 (O_1187,N_19950,N_19905);
xnor UO_1188 (O_1188,N_19923,N_19794);
or UO_1189 (O_1189,N_19941,N_19893);
nor UO_1190 (O_1190,N_19839,N_19805);
and UO_1191 (O_1191,N_19967,N_19830);
and UO_1192 (O_1192,N_19906,N_19863);
and UO_1193 (O_1193,N_19774,N_19880);
nor UO_1194 (O_1194,N_19885,N_19952);
nand UO_1195 (O_1195,N_19908,N_19874);
and UO_1196 (O_1196,N_19786,N_19934);
nand UO_1197 (O_1197,N_19935,N_19889);
xnor UO_1198 (O_1198,N_19946,N_19900);
nor UO_1199 (O_1199,N_19988,N_19847);
or UO_1200 (O_1200,N_19828,N_19893);
or UO_1201 (O_1201,N_19796,N_19973);
xor UO_1202 (O_1202,N_19841,N_19867);
nand UO_1203 (O_1203,N_19872,N_19972);
nor UO_1204 (O_1204,N_19993,N_19884);
nand UO_1205 (O_1205,N_19895,N_19812);
or UO_1206 (O_1206,N_19887,N_19977);
nor UO_1207 (O_1207,N_19807,N_19880);
or UO_1208 (O_1208,N_19941,N_19753);
xnor UO_1209 (O_1209,N_19875,N_19790);
or UO_1210 (O_1210,N_19866,N_19896);
and UO_1211 (O_1211,N_19870,N_19824);
or UO_1212 (O_1212,N_19752,N_19914);
nor UO_1213 (O_1213,N_19815,N_19914);
nor UO_1214 (O_1214,N_19955,N_19865);
xor UO_1215 (O_1215,N_19815,N_19950);
and UO_1216 (O_1216,N_19947,N_19780);
xnor UO_1217 (O_1217,N_19826,N_19911);
and UO_1218 (O_1218,N_19914,N_19987);
xor UO_1219 (O_1219,N_19811,N_19898);
nor UO_1220 (O_1220,N_19920,N_19906);
or UO_1221 (O_1221,N_19994,N_19992);
xor UO_1222 (O_1222,N_19908,N_19882);
or UO_1223 (O_1223,N_19822,N_19757);
and UO_1224 (O_1224,N_19791,N_19940);
or UO_1225 (O_1225,N_19816,N_19964);
xor UO_1226 (O_1226,N_19884,N_19772);
xor UO_1227 (O_1227,N_19914,N_19950);
or UO_1228 (O_1228,N_19894,N_19860);
xnor UO_1229 (O_1229,N_19836,N_19850);
nor UO_1230 (O_1230,N_19831,N_19922);
xnor UO_1231 (O_1231,N_19860,N_19994);
nor UO_1232 (O_1232,N_19881,N_19908);
xnor UO_1233 (O_1233,N_19833,N_19985);
xor UO_1234 (O_1234,N_19798,N_19994);
or UO_1235 (O_1235,N_19868,N_19750);
nand UO_1236 (O_1236,N_19864,N_19948);
xnor UO_1237 (O_1237,N_19835,N_19765);
and UO_1238 (O_1238,N_19919,N_19962);
and UO_1239 (O_1239,N_19949,N_19766);
and UO_1240 (O_1240,N_19904,N_19791);
or UO_1241 (O_1241,N_19970,N_19982);
nor UO_1242 (O_1242,N_19880,N_19974);
and UO_1243 (O_1243,N_19755,N_19926);
and UO_1244 (O_1244,N_19900,N_19768);
and UO_1245 (O_1245,N_19810,N_19812);
xor UO_1246 (O_1246,N_19823,N_19869);
or UO_1247 (O_1247,N_19996,N_19969);
or UO_1248 (O_1248,N_19898,N_19765);
nand UO_1249 (O_1249,N_19866,N_19848);
and UO_1250 (O_1250,N_19780,N_19990);
or UO_1251 (O_1251,N_19956,N_19822);
xnor UO_1252 (O_1252,N_19963,N_19999);
nand UO_1253 (O_1253,N_19983,N_19930);
and UO_1254 (O_1254,N_19828,N_19773);
or UO_1255 (O_1255,N_19890,N_19910);
nor UO_1256 (O_1256,N_19786,N_19803);
nor UO_1257 (O_1257,N_19962,N_19959);
xor UO_1258 (O_1258,N_19930,N_19949);
or UO_1259 (O_1259,N_19798,N_19847);
and UO_1260 (O_1260,N_19887,N_19756);
and UO_1261 (O_1261,N_19975,N_19926);
nand UO_1262 (O_1262,N_19761,N_19861);
and UO_1263 (O_1263,N_19877,N_19948);
xnor UO_1264 (O_1264,N_19816,N_19898);
nand UO_1265 (O_1265,N_19916,N_19767);
nor UO_1266 (O_1266,N_19897,N_19932);
nand UO_1267 (O_1267,N_19882,N_19977);
nand UO_1268 (O_1268,N_19802,N_19841);
nor UO_1269 (O_1269,N_19750,N_19918);
and UO_1270 (O_1270,N_19810,N_19954);
xnor UO_1271 (O_1271,N_19801,N_19852);
or UO_1272 (O_1272,N_19953,N_19975);
nand UO_1273 (O_1273,N_19953,N_19905);
xnor UO_1274 (O_1274,N_19943,N_19911);
nand UO_1275 (O_1275,N_19882,N_19854);
xor UO_1276 (O_1276,N_19803,N_19973);
and UO_1277 (O_1277,N_19753,N_19982);
nor UO_1278 (O_1278,N_19928,N_19915);
and UO_1279 (O_1279,N_19958,N_19918);
xnor UO_1280 (O_1280,N_19765,N_19929);
nor UO_1281 (O_1281,N_19853,N_19770);
xnor UO_1282 (O_1282,N_19762,N_19857);
nand UO_1283 (O_1283,N_19821,N_19755);
xor UO_1284 (O_1284,N_19989,N_19985);
xnor UO_1285 (O_1285,N_19975,N_19754);
and UO_1286 (O_1286,N_19862,N_19877);
and UO_1287 (O_1287,N_19943,N_19968);
or UO_1288 (O_1288,N_19802,N_19895);
nor UO_1289 (O_1289,N_19884,N_19800);
and UO_1290 (O_1290,N_19769,N_19979);
xor UO_1291 (O_1291,N_19955,N_19859);
nor UO_1292 (O_1292,N_19969,N_19771);
nand UO_1293 (O_1293,N_19877,N_19969);
nor UO_1294 (O_1294,N_19923,N_19913);
and UO_1295 (O_1295,N_19823,N_19754);
and UO_1296 (O_1296,N_19826,N_19838);
nor UO_1297 (O_1297,N_19935,N_19797);
xnor UO_1298 (O_1298,N_19925,N_19774);
nand UO_1299 (O_1299,N_19960,N_19937);
and UO_1300 (O_1300,N_19809,N_19957);
and UO_1301 (O_1301,N_19786,N_19950);
or UO_1302 (O_1302,N_19967,N_19881);
and UO_1303 (O_1303,N_19924,N_19972);
and UO_1304 (O_1304,N_19784,N_19766);
or UO_1305 (O_1305,N_19819,N_19903);
nand UO_1306 (O_1306,N_19927,N_19926);
nand UO_1307 (O_1307,N_19936,N_19879);
and UO_1308 (O_1308,N_19950,N_19939);
xor UO_1309 (O_1309,N_19840,N_19941);
nand UO_1310 (O_1310,N_19887,N_19912);
xnor UO_1311 (O_1311,N_19847,N_19845);
xor UO_1312 (O_1312,N_19959,N_19835);
xnor UO_1313 (O_1313,N_19917,N_19977);
and UO_1314 (O_1314,N_19908,N_19795);
and UO_1315 (O_1315,N_19802,N_19795);
and UO_1316 (O_1316,N_19802,N_19871);
nand UO_1317 (O_1317,N_19953,N_19972);
nand UO_1318 (O_1318,N_19886,N_19986);
nor UO_1319 (O_1319,N_19864,N_19884);
xor UO_1320 (O_1320,N_19814,N_19990);
and UO_1321 (O_1321,N_19767,N_19974);
xnor UO_1322 (O_1322,N_19900,N_19912);
nor UO_1323 (O_1323,N_19821,N_19937);
xor UO_1324 (O_1324,N_19791,N_19934);
xor UO_1325 (O_1325,N_19982,N_19880);
nand UO_1326 (O_1326,N_19959,N_19833);
xor UO_1327 (O_1327,N_19976,N_19882);
nor UO_1328 (O_1328,N_19975,N_19804);
or UO_1329 (O_1329,N_19982,N_19787);
nor UO_1330 (O_1330,N_19880,N_19992);
xnor UO_1331 (O_1331,N_19762,N_19981);
nand UO_1332 (O_1332,N_19813,N_19812);
xnor UO_1333 (O_1333,N_19756,N_19766);
nor UO_1334 (O_1334,N_19886,N_19864);
xnor UO_1335 (O_1335,N_19906,N_19970);
xnor UO_1336 (O_1336,N_19963,N_19922);
and UO_1337 (O_1337,N_19909,N_19829);
or UO_1338 (O_1338,N_19879,N_19999);
nor UO_1339 (O_1339,N_19840,N_19866);
nor UO_1340 (O_1340,N_19945,N_19772);
xnor UO_1341 (O_1341,N_19861,N_19891);
xor UO_1342 (O_1342,N_19986,N_19822);
xor UO_1343 (O_1343,N_19911,N_19768);
or UO_1344 (O_1344,N_19922,N_19904);
nand UO_1345 (O_1345,N_19755,N_19808);
and UO_1346 (O_1346,N_19926,N_19920);
nand UO_1347 (O_1347,N_19991,N_19753);
xnor UO_1348 (O_1348,N_19951,N_19840);
nand UO_1349 (O_1349,N_19916,N_19905);
or UO_1350 (O_1350,N_19786,N_19797);
and UO_1351 (O_1351,N_19818,N_19897);
nand UO_1352 (O_1352,N_19765,N_19922);
or UO_1353 (O_1353,N_19790,N_19841);
nand UO_1354 (O_1354,N_19756,N_19758);
nand UO_1355 (O_1355,N_19872,N_19893);
and UO_1356 (O_1356,N_19775,N_19795);
xor UO_1357 (O_1357,N_19761,N_19833);
and UO_1358 (O_1358,N_19835,N_19779);
nand UO_1359 (O_1359,N_19773,N_19932);
nand UO_1360 (O_1360,N_19917,N_19959);
and UO_1361 (O_1361,N_19847,N_19854);
xnor UO_1362 (O_1362,N_19886,N_19959);
xor UO_1363 (O_1363,N_19763,N_19759);
xnor UO_1364 (O_1364,N_19874,N_19880);
xor UO_1365 (O_1365,N_19862,N_19788);
nand UO_1366 (O_1366,N_19867,N_19950);
and UO_1367 (O_1367,N_19817,N_19797);
and UO_1368 (O_1368,N_19963,N_19957);
xnor UO_1369 (O_1369,N_19782,N_19756);
xor UO_1370 (O_1370,N_19953,N_19981);
xnor UO_1371 (O_1371,N_19875,N_19897);
xor UO_1372 (O_1372,N_19938,N_19981);
or UO_1373 (O_1373,N_19909,N_19980);
or UO_1374 (O_1374,N_19817,N_19937);
and UO_1375 (O_1375,N_19922,N_19843);
nand UO_1376 (O_1376,N_19970,N_19928);
and UO_1377 (O_1377,N_19976,N_19912);
nand UO_1378 (O_1378,N_19795,N_19963);
or UO_1379 (O_1379,N_19958,N_19876);
or UO_1380 (O_1380,N_19984,N_19949);
xnor UO_1381 (O_1381,N_19990,N_19808);
xor UO_1382 (O_1382,N_19988,N_19976);
nand UO_1383 (O_1383,N_19932,N_19830);
nor UO_1384 (O_1384,N_19983,N_19799);
nand UO_1385 (O_1385,N_19755,N_19769);
nand UO_1386 (O_1386,N_19916,N_19878);
nor UO_1387 (O_1387,N_19875,N_19910);
nand UO_1388 (O_1388,N_19754,N_19911);
nand UO_1389 (O_1389,N_19890,N_19992);
xnor UO_1390 (O_1390,N_19844,N_19915);
or UO_1391 (O_1391,N_19934,N_19754);
xnor UO_1392 (O_1392,N_19838,N_19820);
xor UO_1393 (O_1393,N_19923,N_19890);
or UO_1394 (O_1394,N_19799,N_19956);
and UO_1395 (O_1395,N_19762,N_19909);
nand UO_1396 (O_1396,N_19835,N_19808);
nand UO_1397 (O_1397,N_19823,N_19804);
nor UO_1398 (O_1398,N_19762,N_19799);
nor UO_1399 (O_1399,N_19853,N_19892);
nand UO_1400 (O_1400,N_19854,N_19943);
and UO_1401 (O_1401,N_19835,N_19791);
and UO_1402 (O_1402,N_19998,N_19949);
nand UO_1403 (O_1403,N_19969,N_19956);
xor UO_1404 (O_1404,N_19946,N_19925);
and UO_1405 (O_1405,N_19842,N_19959);
nand UO_1406 (O_1406,N_19923,N_19978);
nand UO_1407 (O_1407,N_19978,N_19878);
nand UO_1408 (O_1408,N_19790,N_19901);
and UO_1409 (O_1409,N_19932,N_19776);
and UO_1410 (O_1410,N_19839,N_19920);
and UO_1411 (O_1411,N_19876,N_19762);
or UO_1412 (O_1412,N_19809,N_19886);
nand UO_1413 (O_1413,N_19889,N_19807);
and UO_1414 (O_1414,N_19958,N_19968);
or UO_1415 (O_1415,N_19985,N_19812);
or UO_1416 (O_1416,N_19796,N_19900);
nor UO_1417 (O_1417,N_19945,N_19969);
xor UO_1418 (O_1418,N_19975,N_19776);
nand UO_1419 (O_1419,N_19788,N_19847);
xor UO_1420 (O_1420,N_19763,N_19938);
nor UO_1421 (O_1421,N_19946,N_19828);
nor UO_1422 (O_1422,N_19804,N_19929);
nor UO_1423 (O_1423,N_19872,N_19922);
or UO_1424 (O_1424,N_19800,N_19777);
nand UO_1425 (O_1425,N_19964,N_19820);
or UO_1426 (O_1426,N_19866,N_19762);
nor UO_1427 (O_1427,N_19973,N_19752);
and UO_1428 (O_1428,N_19819,N_19973);
or UO_1429 (O_1429,N_19850,N_19782);
xor UO_1430 (O_1430,N_19990,N_19868);
or UO_1431 (O_1431,N_19967,N_19835);
or UO_1432 (O_1432,N_19795,N_19990);
nand UO_1433 (O_1433,N_19848,N_19943);
nand UO_1434 (O_1434,N_19857,N_19877);
nand UO_1435 (O_1435,N_19804,N_19993);
nor UO_1436 (O_1436,N_19960,N_19871);
nand UO_1437 (O_1437,N_19829,N_19884);
and UO_1438 (O_1438,N_19759,N_19755);
xnor UO_1439 (O_1439,N_19830,N_19815);
xnor UO_1440 (O_1440,N_19904,N_19930);
and UO_1441 (O_1441,N_19753,N_19897);
nor UO_1442 (O_1442,N_19950,N_19947);
or UO_1443 (O_1443,N_19768,N_19950);
nor UO_1444 (O_1444,N_19786,N_19770);
nor UO_1445 (O_1445,N_19844,N_19849);
xor UO_1446 (O_1446,N_19928,N_19779);
xnor UO_1447 (O_1447,N_19851,N_19881);
nor UO_1448 (O_1448,N_19917,N_19941);
xnor UO_1449 (O_1449,N_19975,N_19932);
and UO_1450 (O_1450,N_19889,N_19838);
or UO_1451 (O_1451,N_19757,N_19937);
and UO_1452 (O_1452,N_19777,N_19793);
nand UO_1453 (O_1453,N_19871,N_19841);
nor UO_1454 (O_1454,N_19918,N_19889);
and UO_1455 (O_1455,N_19826,N_19914);
xnor UO_1456 (O_1456,N_19981,N_19759);
or UO_1457 (O_1457,N_19887,N_19828);
nand UO_1458 (O_1458,N_19896,N_19870);
nor UO_1459 (O_1459,N_19918,N_19878);
or UO_1460 (O_1460,N_19865,N_19852);
and UO_1461 (O_1461,N_19875,N_19978);
nand UO_1462 (O_1462,N_19811,N_19933);
and UO_1463 (O_1463,N_19847,N_19761);
nor UO_1464 (O_1464,N_19757,N_19869);
nor UO_1465 (O_1465,N_19902,N_19765);
xor UO_1466 (O_1466,N_19853,N_19872);
xor UO_1467 (O_1467,N_19762,N_19958);
xor UO_1468 (O_1468,N_19943,N_19853);
or UO_1469 (O_1469,N_19803,N_19798);
nand UO_1470 (O_1470,N_19831,N_19876);
xnor UO_1471 (O_1471,N_19805,N_19762);
and UO_1472 (O_1472,N_19846,N_19888);
nand UO_1473 (O_1473,N_19890,N_19834);
and UO_1474 (O_1474,N_19815,N_19887);
nor UO_1475 (O_1475,N_19794,N_19792);
or UO_1476 (O_1476,N_19842,N_19811);
nand UO_1477 (O_1477,N_19871,N_19948);
nor UO_1478 (O_1478,N_19757,N_19966);
nor UO_1479 (O_1479,N_19783,N_19773);
xnor UO_1480 (O_1480,N_19938,N_19784);
xor UO_1481 (O_1481,N_19952,N_19849);
and UO_1482 (O_1482,N_19890,N_19997);
and UO_1483 (O_1483,N_19977,N_19916);
nand UO_1484 (O_1484,N_19994,N_19761);
or UO_1485 (O_1485,N_19919,N_19898);
or UO_1486 (O_1486,N_19796,N_19895);
xnor UO_1487 (O_1487,N_19908,N_19992);
xnor UO_1488 (O_1488,N_19979,N_19906);
nand UO_1489 (O_1489,N_19867,N_19770);
and UO_1490 (O_1490,N_19989,N_19995);
or UO_1491 (O_1491,N_19889,N_19942);
or UO_1492 (O_1492,N_19873,N_19870);
nand UO_1493 (O_1493,N_19884,N_19798);
or UO_1494 (O_1494,N_19888,N_19907);
nor UO_1495 (O_1495,N_19883,N_19912);
nor UO_1496 (O_1496,N_19923,N_19854);
nor UO_1497 (O_1497,N_19905,N_19941);
xnor UO_1498 (O_1498,N_19970,N_19802);
nand UO_1499 (O_1499,N_19953,N_19838);
nor UO_1500 (O_1500,N_19815,N_19820);
or UO_1501 (O_1501,N_19971,N_19825);
and UO_1502 (O_1502,N_19854,N_19833);
nand UO_1503 (O_1503,N_19896,N_19764);
nand UO_1504 (O_1504,N_19987,N_19811);
and UO_1505 (O_1505,N_19959,N_19831);
xnor UO_1506 (O_1506,N_19828,N_19782);
and UO_1507 (O_1507,N_19800,N_19993);
nor UO_1508 (O_1508,N_19818,N_19884);
nand UO_1509 (O_1509,N_19935,N_19953);
and UO_1510 (O_1510,N_19837,N_19971);
xor UO_1511 (O_1511,N_19827,N_19842);
nor UO_1512 (O_1512,N_19874,N_19808);
nor UO_1513 (O_1513,N_19925,N_19798);
nor UO_1514 (O_1514,N_19913,N_19834);
and UO_1515 (O_1515,N_19992,N_19909);
or UO_1516 (O_1516,N_19874,N_19849);
and UO_1517 (O_1517,N_19923,N_19831);
nor UO_1518 (O_1518,N_19974,N_19879);
and UO_1519 (O_1519,N_19814,N_19974);
xnor UO_1520 (O_1520,N_19771,N_19985);
nand UO_1521 (O_1521,N_19884,N_19792);
or UO_1522 (O_1522,N_19918,N_19764);
xnor UO_1523 (O_1523,N_19908,N_19933);
nand UO_1524 (O_1524,N_19826,N_19988);
nand UO_1525 (O_1525,N_19915,N_19783);
xnor UO_1526 (O_1526,N_19955,N_19852);
nor UO_1527 (O_1527,N_19797,N_19754);
xor UO_1528 (O_1528,N_19916,N_19952);
nand UO_1529 (O_1529,N_19900,N_19920);
or UO_1530 (O_1530,N_19892,N_19810);
xnor UO_1531 (O_1531,N_19895,N_19930);
nand UO_1532 (O_1532,N_19943,N_19772);
xor UO_1533 (O_1533,N_19942,N_19852);
nor UO_1534 (O_1534,N_19877,N_19870);
and UO_1535 (O_1535,N_19769,N_19790);
xor UO_1536 (O_1536,N_19881,N_19771);
nand UO_1537 (O_1537,N_19998,N_19878);
and UO_1538 (O_1538,N_19996,N_19777);
xor UO_1539 (O_1539,N_19981,N_19862);
xor UO_1540 (O_1540,N_19795,N_19780);
or UO_1541 (O_1541,N_19794,N_19964);
nand UO_1542 (O_1542,N_19869,N_19805);
xor UO_1543 (O_1543,N_19941,N_19871);
nand UO_1544 (O_1544,N_19969,N_19830);
and UO_1545 (O_1545,N_19756,N_19776);
or UO_1546 (O_1546,N_19883,N_19977);
or UO_1547 (O_1547,N_19910,N_19814);
nand UO_1548 (O_1548,N_19937,N_19847);
nand UO_1549 (O_1549,N_19816,N_19971);
nor UO_1550 (O_1550,N_19867,N_19969);
or UO_1551 (O_1551,N_19759,N_19891);
nand UO_1552 (O_1552,N_19865,N_19786);
nand UO_1553 (O_1553,N_19907,N_19826);
and UO_1554 (O_1554,N_19785,N_19771);
nor UO_1555 (O_1555,N_19896,N_19997);
xor UO_1556 (O_1556,N_19875,N_19938);
nand UO_1557 (O_1557,N_19802,N_19753);
xor UO_1558 (O_1558,N_19815,N_19785);
or UO_1559 (O_1559,N_19774,N_19786);
or UO_1560 (O_1560,N_19865,N_19862);
or UO_1561 (O_1561,N_19905,N_19903);
and UO_1562 (O_1562,N_19817,N_19927);
xnor UO_1563 (O_1563,N_19959,N_19978);
nand UO_1564 (O_1564,N_19786,N_19775);
xnor UO_1565 (O_1565,N_19919,N_19905);
nor UO_1566 (O_1566,N_19845,N_19959);
nand UO_1567 (O_1567,N_19754,N_19826);
nor UO_1568 (O_1568,N_19809,N_19816);
and UO_1569 (O_1569,N_19887,N_19999);
nand UO_1570 (O_1570,N_19826,N_19798);
nor UO_1571 (O_1571,N_19894,N_19752);
xor UO_1572 (O_1572,N_19906,N_19969);
xor UO_1573 (O_1573,N_19831,N_19821);
and UO_1574 (O_1574,N_19790,N_19975);
nor UO_1575 (O_1575,N_19920,N_19798);
nand UO_1576 (O_1576,N_19927,N_19842);
or UO_1577 (O_1577,N_19833,N_19945);
xor UO_1578 (O_1578,N_19814,N_19778);
nand UO_1579 (O_1579,N_19937,N_19963);
nand UO_1580 (O_1580,N_19861,N_19834);
xnor UO_1581 (O_1581,N_19946,N_19998);
xnor UO_1582 (O_1582,N_19802,N_19761);
nand UO_1583 (O_1583,N_19807,N_19765);
xnor UO_1584 (O_1584,N_19789,N_19772);
xnor UO_1585 (O_1585,N_19824,N_19860);
nand UO_1586 (O_1586,N_19795,N_19810);
nor UO_1587 (O_1587,N_19902,N_19824);
nor UO_1588 (O_1588,N_19946,N_19950);
and UO_1589 (O_1589,N_19853,N_19786);
xor UO_1590 (O_1590,N_19990,N_19879);
xnor UO_1591 (O_1591,N_19836,N_19879);
or UO_1592 (O_1592,N_19876,N_19766);
xnor UO_1593 (O_1593,N_19826,N_19931);
or UO_1594 (O_1594,N_19890,N_19859);
or UO_1595 (O_1595,N_19992,N_19859);
xor UO_1596 (O_1596,N_19992,N_19872);
xor UO_1597 (O_1597,N_19812,N_19958);
nor UO_1598 (O_1598,N_19871,N_19891);
xnor UO_1599 (O_1599,N_19785,N_19793);
xor UO_1600 (O_1600,N_19789,N_19867);
nor UO_1601 (O_1601,N_19859,N_19986);
nand UO_1602 (O_1602,N_19776,N_19907);
or UO_1603 (O_1603,N_19890,N_19894);
or UO_1604 (O_1604,N_19758,N_19970);
or UO_1605 (O_1605,N_19955,N_19958);
xnor UO_1606 (O_1606,N_19792,N_19843);
nor UO_1607 (O_1607,N_19989,N_19857);
and UO_1608 (O_1608,N_19859,N_19911);
and UO_1609 (O_1609,N_19771,N_19828);
or UO_1610 (O_1610,N_19850,N_19818);
xnor UO_1611 (O_1611,N_19871,N_19931);
nor UO_1612 (O_1612,N_19894,N_19928);
and UO_1613 (O_1613,N_19884,N_19853);
and UO_1614 (O_1614,N_19831,N_19970);
xor UO_1615 (O_1615,N_19803,N_19767);
xor UO_1616 (O_1616,N_19922,N_19780);
xnor UO_1617 (O_1617,N_19934,N_19937);
xor UO_1618 (O_1618,N_19923,N_19909);
nand UO_1619 (O_1619,N_19871,N_19852);
and UO_1620 (O_1620,N_19771,N_19949);
xor UO_1621 (O_1621,N_19967,N_19993);
nand UO_1622 (O_1622,N_19996,N_19971);
xor UO_1623 (O_1623,N_19957,N_19764);
xor UO_1624 (O_1624,N_19815,N_19771);
nand UO_1625 (O_1625,N_19779,N_19948);
or UO_1626 (O_1626,N_19891,N_19981);
nand UO_1627 (O_1627,N_19794,N_19832);
and UO_1628 (O_1628,N_19756,N_19940);
and UO_1629 (O_1629,N_19918,N_19879);
and UO_1630 (O_1630,N_19831,N_19956);
nand UO_1631 (O_1631,N_19910,N_19876);
nand UO_1632 (O_1632,N_19973,N_19840);
and UO_1633 (O_1633,N_19996,N_19829);
or UO_1634 (O_1634,N_19891,N_19804);
xor UO_1635 (O_1635,N_19942,N_19781);
and UO_1636 (O_1636,N_19813,N_19973);
nor UO_1637 (O_1637,N_19946,N_19878);
xnor UO_1638 (O_1638,N_19779,N_19833);
nand UO_1639 (O_1639,N_19899,N_19769);
nor UO_1640 (O_1640,N_19750,N_19956);
or UO_1641 (O_1641,N_19787,N_19997);
xor UO_1642 (O_1642,N_19822,N_19988);
or UO_1643 (O_1643,N_19808,N_19752);
and UO_1644 (O_1644,N_19981,N_19849);
nand UO_1645 (O_1645,N_19923,N_19895);
or UO_1646 (O_1646,N_19761,N_19978);
nand UO_1647 (O_1647,N_19791,N_19981);
or UO_1648 (O_1648,N_19787,N_19977);
nor UO_1649 (O_1649,N_19928,N_19858);
nor UO_1650 (O_1650,N_19930,N_19950);
and UO_1651 (O_1651,N_19817,N_19834);
nor UO_1652 (O_1652,N_19772,N_19818);
and UO_1653 (O_1653,N_19861,N_19811);
nor UO_1654 (O_1654,N_19965,N_19919);
xor UO_1655 (O_1655,N_19900,N_19968);
and UO_1656 (O_1656,N_19872,N_19956);
nor UO_1657 (O_1657,N_19853,N_19891);
or UO_1658 (O_1658,N_19823,N_19948);
xnor UO_1659 (O_1659,N_19904,N_19877);
nand UO_1660 (O_1660,N_19804,N_19928);
xnor UO_1661 (O_1661,N_19776,N_19968);
or UO_1662 (O_1662,N_19765,N_19920);
or UO_1663 (O_1663,N_19954,N_19852);
or UO_1664 (O_1664,N_19960,N_19750);
or UO_1665 (O_1665,N_19834,N_19979);
nand UO_1666 (O_1666,N_19889,N_19851);
xor UO_1667 (O_1667,N_19785,N_19796);
or UO_1668 (O_1668,N_19767,N_19872);
or UO_1669 (O_1669,N_19851,N_19942);
or UO_1670 (O_1670,N_19892,N_19977);
or UO_1671 (O_1671,N_19976,N_19801);
nand UO_1672 (O_1672,N_19955,N_19933);
xor UO_1673 (O_1673,N_19888,N_19911);
nor UO_1674 (O_1674,N_19762,N_19869);
nor UO_1675 (O_1675,N_19970,N_19765);
or UO_1676 (O_1676,N_19865,N_19944);
xor UO_1677 (O_1677,N_19765,N_19975);
nand UO_1678 (O_1678,N_19856,N_19782);
xor UO_1679 (O_1679,N_19945,N_19872);
nand UO_1680 (O_1680,N_19778,N_19920);
nor UO_1681 (O_1681,N_19867,N_19952);
xnor UO_1682 (O_1682,N_19832,N_19905);
and UO_1683 (O_1683,N_19965,N_19988);
nor UO_1684 (O_1684,N_19859,N_19806);
and UO_1685 (O_1685,N_19842,N_19805);
nor UO_1686 (O_1686,N_19913,N_19888);
nand UO_1687 (O_1687,N_19833,N_19934);
nand UO_1688 (O_1688,N_19779,N_19795);
or UO_1689 (O_1689,N_19947,N_19951);
nor UO_1690 (O_1690,N_19809,N_19947);
or UO_1691 (O_1691,N_19859,N_19761);
and UO_1692 (O_1692,N_19844,N_19941);
nand UO_1693 (O_1693,N_19989,N_19978);
xnor UO_1694 (O_1694,N_19817,N_19886);
nand UO_1695 (O_1695,N_19827,N_19943);
nor UO_1696 (O_1696,N_19860,N_19792);
nand UO_1697 (O_1697,N_19835,N_19932);
or UO_1698 (O_1698,N_19923,N_19815);
or UO_1699 (O_1699,N_19752,N_19895);
xor UO_1700 (O_1700,N_19859,N_19861);
xor UO_1701 (O_1701,N_19980,N_19791);
and UO_1702 (O_1702,N_19772,N_19841);
nor UO_1703 (O_1703,N_19827,N_19955);
nor UO_1704 (O_1704,N_19943,N_19779);
and UO_1705 (O_1705,N_19926,N_19794);
and UO_1706 (O_1706,N_19767,N_19971);
nand UO_1707 (O_1707,N_19863,N_19763);
and UO_1708 (O_1708,N_19775,N_19850);
xor UO_1709 (O_1709,N_19906,N_19901);
nand UO_1710 (O_1710,N_19837,N_19877);
nor UO_1711 (O_1711,N_19808,N_19809);
nand UO_1712 (O_1712,N_19885,N_19784);
nor UO_1713 (O_1713,N_19924,N_19922);
or UO_1714 (O_1714,N_19900,N_19951);
nand UO_1715 (O_1715,N_19805,N_19780);
nand UO_1716 (O_1716,N_19800,N_19876);
nor UO_1717 (O_1717,N_19873,N_19779);
nand UO_1718 (O_1718,N_19942,N_19983);
xor UO_1719 (O_1719,N_19958,N_19985);
xnor UO_1720 (O_1720,N_19879,N_19839);
xnor UO_1721 (O_1721,N_19820,N_19996);
nor UO_1722 (O_1722,N_19893,N_19957);
or UO_1723 (O_1723,N_19904,N_19857);
nand UO_1724 (O_1724,N_19968,N_19970);
nand UO_1725 (O_1725,N_19972,N_19829);
nand UO_1726 (O_1726,N_19885,N_19752);
xnor UO_1727 (O_1727,N_19998,N_19770);
nand UO_1728 (O_1728,N_19812,N_19966);
nor UO_1729 (O_1729,N_19845,N_19858);
or UO_1730 (O_1730,N_19961,N_19789);
nor UO_1731 (O_1731,N_19847,N_19793);
xor UO_1732 (O_1732,N_19944,N_19853);
xor UO_1733 (O_1733,N_19783,N_19911);
nor UO_1734 (O_1734,N_19755,N_19819);
and UO_1735 (O_1735,N_19929,N_19942);
or UO_1736 (O_1736,N_19999,N_19947);
and UO_1737 (O_1737,N_19793,N_19998);
or UO_1738 (O_1738,N_19904,N_19992);
nor UO_1739 (O_1739,N_19779,N_19971);
or UO_1740 (O_1740,N_19903,N_19790);
or UO_1741 (O_1741,N_19885,N_19764);
nand UO_1742 (O_1742,N_19942,N_19967);
nor UO_1743 (O_1743,N_19926,N_19852);
or UO_1744 (O_1744,N_19993,N_19773);
nand UO_1745 (O_1745,N_19934,N_19836);
and UO_1746 (O_1746,N_19960,N_19886);
nor UO_1747 (O_1747,N_19865,N_19855);
nand UO_1748 (O_1748,N_19922,N_19998);
nand UO_1749 (O_1749,N_19907,N_19839);
and UO_1750 (O_1750,N_19852,N_19885);
and UO_1751 (O_1751,N_19929,N_19855);
nand UO_1752 (O_1752,N_19931,N_19877);
or UO_1753 (O_1753,N_19856,N_19940);
and UO_1754 (O_1754,N_19800,N_19796);
and UO_1755 (O_1755,N_19969,N_19964);
or UO_1756 (O_1756,N_19937,N_19927);
nand UO_1757 (O_1757,N_19903,N_19794);
and UO_1758 (O_1758,N_19990,N_19971);
xor UO_1759 (O_1759,N_19785,N_19782);
nand UO_1760 (O_1760,N_19907,N_19793);
xor UO_1761 (O_1761,N_19832,N_19934);
nor UO_1762 (O_1762,N_19789,N_19890);
and UO_1763 (O_1763,N_19896,N_19799);
and UO_1764 (O_1764,N_19978,N_19943);
xor UO_1765 (O_1765,N_19805,N_19890);
xor UO_1766 (O_1766,N_19752,N_19955);
and UO_1767 (O_1767,N_19784,N_19840);
or UO_1768 (O_1768,N_19990,N_19996);
or UO_1769 (O_1769,N_19850,N_19958);
nor UO_1770 (O_1770,N_19859,N_19870);
and UO_1771 (O_1771,N_19760,N_19811);
and UO_1772 (O_1772,N_19965,N_19920);
xor UO_1773 (O_1773,N_19881,N_19992);
or UO_1774 (O_1774,N_19841,N_19924);
or UO_1775 (O_1775,N_19984,N_19808);
xnor UO_1776 (O_1776,N_19886,N_19869);
xor UO_1777 (O_1777,N_19778,N_19856);
nand UO_1778 (O_1778,N_19856,N_19762);
and UO_1779 (O_1779,N_19952,N_19769);
and UO_1780 (O_1780,N_19925,N_19827);
nand UO_1781 (O_1781,N_19934,N_19977);
or UO_1782 (O_1782,N_19991,N_19917);
nand UO_1783 (O_1783,N_19758,N_19893);
nand UO_1784 (O_1784,N_19858,N_19907);
nor UO_1785 (O_1785,N_19796,N_19920);
nor UO_1786 (O_1786,N_19944,N_19835);
and UO_1787 (O_1787,N_19932,N_19784);
nand UO_1788 (O_1788,N_19802,N_19904);
or UO_1789 (O_1789,N_19973,N_19781);
or UO_1790 (O_1790,N_19783,N_19955);
xor UO_1791 (O_1791,N_19815,N_19910);
or UO_1792 (O_1792,N_19780,N_19873);
nor UO_1793 (O_1793,N_19893,N_19836);
nand UO_1794 (O_1794,N_19979,N_19989);
or UO_1795 (O_1795,N_19954,N_19961);
nor UO_1796 (O_1796,N_19950,N_19982);
xor UO_1797 (O_1797,N_19767,N_19878);
nor UO_1798 (O_1798,N_19939,N_19803);
or UO_1799 (O_1799,N_19886,N_19785);
nand UO_1800 (O_1800,N_19931,N_19811);
nor UO_1801 (O_1801,N_19881,N_19883);
and UO_1802 (O_1802,N_19800,N_19862);
nand UO_1803 (O_1803,N_19764,N_19944);
xnor UO_1804 (O_1804,N_19779,N_19789);
nor UO_1805 (O_1805,N_19874,N_19781);
or UO_1806 (O_1806,N_19843,N_19991);
nor UO_1807 (O_1807,N_19900,N_19931);
nand UO_1808 (O_1808,N_19911,N_19770);
and UO_1809 (O_1809,N_19920,N_19833);
and UO_1810 (O_1810,N_19791,N_19883);
nand UO_1811 (O_1811,N_19942,N_19959);
xnor UO_1812 (O_1812,N_19834,N_19880);
xor UO_1813 (O_1813,N_19940,N_19895);
and UO_1814 (O_1814,N_19856,N_19826);
nand UO_1815 (O_1815,N_19979,N_19786);
xor UO_1816 (O_1816,N_19940,N_19760);
xor UO_1817 (O_1817,N_19881,N_19781);
nor UO_1818 (O_1818,N_19753,N_19789);
and UO_1819 (O_1819,N_19897,N_19980);
xor UO_1820 (O_1820,N_19793,N_19758);
nand UO_1821 (O_1821,N_19974,N_19823);
or UO_1822 (O_1822,N_19908,N_19948);
or UO_1823 (O_1823,N_19767,N_19951);
xor UO_1824 (O_1824,N_19946,N_19872);
nand UO_1825 (O_1825,N_19790,N_19808);
nand UO_1826 (O_1826,N_19864,N_19888);
nand UO_1827 (O_1827,N_19934,N_19882);
or UO_1828 (O_1828,N_19869,N_19793);
nand UO_1829 (O_1829,N_19994,N_19768);
nand UO_1830 (O_1830,N_19804,N_19972);
or UO_1831 (O_1831,N_19766,N_19799);
or UO_1832 (O_1832,N_19855,N_19763);
xnor UO_1833 (O_1833,N_19836,N_19888);
nand UO_1834 (O_1834,N_19861,N_19800);
nor UO_1835 (O_1835,N_19775,N_19983);
and UO_1836 (O_1836,N_19989,N_19828);
nor UO_1837 (O_1837,N_19857,N_19993);
and UO_1838 (O_1838,N_19973,N_19936);
nand UO_1839 (O_1839,N_19935,N_19916);
nand UO_1840 (O_1840,N_19937,N_19760);
nor UO_1841 (O_1841,N_19819,N_19959);
nor UO_1842 (O_1842,N_19964,N_19834);
nor UO_1843 (O_1843,N_19799,N_19953);
nor UO_1844 (O_1844,N_19868,N_19849);
nand UO_1845 (O_1845,N_19991,N_19778);
xor UO_1846 (O_1846,N_19898,N_19851);
and UO_1847 (O_1847,N_19994,N_19918);
or UO_1848 (O_1848,N_19819,N_19881);
nor UO_1849 (O_1849,N_19807,N_19817);
and UO_1850 (O_1850,N_19802,N_19991);
and UO_1851 (O_1851,N_19909,N_19946);
nand UO_1852 (O_1852,N_19899,N_19894);
xnor UO_1853 (O_1853,N_19815,N_19924);
or UO_1854 (O_1854,N_19780,N_19906);
and UO_1855 (O_1855,N_19999,N_19905);
nand UO_1856 (O_1856,N_19837,N_19874);
or UO_1857 (O_1857,N_19830,N_19825);
and UO_1858 (O_1858,N_19956,N_19843);
or UO_1859 (O_1859,N_19796,N_19836);
nor UO_1860 (O_1860,N_19935,N_19773);
and UO_1861 (O_1861,N_19862,N_19876);
or UO_1862 (O_1862,N_19910,N_19831);
and UO_1863 (O_1863,N_19990,N_19873);
or UO_1864 (O_1864,N_19767,N_19759);
xnor UO_1865 (O_1865,N_19938,N_19919);
xnor UO_1866 (O_1866,N_19778,N_19912);
nand UO_1867 (O_1867,N_19863,N_19998);
nand UO_1868 (O_1868,N_19843,N_19782);
nor UO_1869 (O_1869,N_19946,N_19786);
xor UO_1870 (O_1870,N_19940,N_19951);
and UO_1871 (O_1871,N_19996,N_19907);
nor UO_1872 (O_1872,N_19901,N_19881);
or UO_1873 (O_1873,N_19983,N_19884);
nor UO_1874 (O_1874,N_19849,N_19998);
or UO_1875 (O_1875,N_19892,N_19927);
nor UO_1876 (O_1876,N_19983,N_19981);
xnor UO_1877 (O_1877,N_19856,N_19841);
xor UO_1878 (O_1878,N_19911,N_19872);
xnor UO_1879 (O_1879,N_19930,N_19911);
or UO_1880 (O_1880,N_19980,N_19809);
nand UO_1881 (O_1881,N_19863,N_19847);
and UO_1882 (O_1882,N_19943,N_19923);
nand UO_1883 (O_1883,N_19852,N_19941);
and UO_1884 (O_1884,N_19932,N_19984);
nand UO_1885 (O_1885,N_19814,N_19784);
and UO_1886 (O_1886,N_19777,N_19871);
and UO_1887 (O_1887,N_19833,N_19994);
or UO_1888 (O_1888,N_19894,N_19900);
nor UO_1889 (O_1889,N_19924,N_19918);
or UO_1890 (O_1890,N_19773,N_19926);
xor UO_1891 (O_1891,N_19873,N_19775);
nor UO_1892 (O_1892,N_19816,N_19930);
and UO_1893 (O_1893,N_19793,N_19773);
nor UO_1894 (O_1894,N_19999,N_19982);
xnor UO_1895 (O_1895,N_19964,N_19992);
nand UO_1896 (O_1896,N_19880,N_19906);
xor UO_1897 (O_1897,N_19826,N_19934);
and UO_1898 (O_1898,N_19820,N_19883);
and UO_1899 (O_1899,N_19907,N_19823);
nor UO_1900 (O_1900,N_19927,N_19941);
xor UO_1901 (O_1901,N_19836,N_19758);
nor UO_1902 (O_1902,N_19931,N_19982);
or UO_1903 (O_1903,N_19975,N_19755);
nor UO_1904 (O_1904,N_19951,N_19803);
xnor UO_1905 (O_1905,N_19835,N_19904);
nor UO_1906 (O_1906,N_19872,N_19884);
nand UO_1907 (O_1907,N_19756,N_19860);
or UO_1908 (O_1908,N_19823,N_19893);
or UO_1909 (O_1909,N_19984,N_19868);
and UO_1910 (O_1910,N_19826,N_19780);
nand UO_1911 (O_1911,N_19918,N_19797);
xnor UO_1912 (O_1912,N_19768,N_19891);
or UO_1913 (O_1913,N_19866,N_19959);
and UO_1914 (O_1914,N_19965,N_19876);
or UO_1915 (O_1915,N_19870,N_19951);
and UO_1916 (O_1916,N_19965,N_19900);
nor UO_1917 (O_1917,N_19822,N_19879);
and UO_1918 (O_1918,N_19908,N_19807);
xnor UO_1919 (O_1919,N_19910,N_19857);
nand UO_1920 (O_1920,N_19949,N_19989);
nand UO_1921 (O_1921,N_19894,N_19789);
and UO_1922 (O_1922,N_19839,N_19949);
nand UO_1923 (O_1923,N_19912,N_19872);
or UO_1924 (O_1924,N_19768,N_19955);
xnor UO_1925 (O_1925,N_19916,N_19985);
xnor UO_1926 (O_1926,N_19916,N_19889);
xor UO_1927 (O_1927,N_19809,N_19851);
nor UO_1928 (O_1928,N_19750,N_19992);
or UO_1929 (O_1929,N_19898,N_19758);
or UO_1930 (O_1930,N_19847,N_19995);
nor UO_1931 (O_1931,N_19988,N_19953);
nor UO_1932 (O_1932,N_19834,N_19887);
or UO_1933 (O_1933,N_19810,N_19904);
nand UO_1934 (O_1934,N_19833,N_19953);
nand UO_1935 (O_1935,N_19863,N_19860);
nand UO_1936 (O_1936,N_19795,N_19943);
or UO_1937 (O_1937,N_19754,N_19867);
and UO_1938 (O_1938,N_19914,N_19991);
nor UO_1939 (O_1939,N_19975,N_19778);
nor UO_1940 (O_1940,N_19901,N_19923);
xnor UO_1941 (O_1941,N_19879,N_19900);
nand UO_1942 (O_1942,N_19919,N_19829);
xor UO_1943 (O_1943,N_19869,N_19751);
nand UO_1944 (O_1944,N_19879,N_19830);
nand UO_1945 (O_1945,N_19912,N_19796);
xor UO_1946 (O_1946,N_19951,N_19857);
or UO_1947 (O_1947,N_19979,N_19829);
nand UO_1948 (O_1948,N_19751,N_19756);
or UO_1949 (O_1949,N_19985,N_19815);
and UO_1950 (O_1950,N_19954,N_19816);
nand UO_1951 (O_1951,N_19794,N_19999);
or UO_1952 (O_1952,N_19764,N_19952);
xnor UO_1953 (O_1953,N_19757,N_19980);
nor UO_1954 (O_1954,N_19752,N_19875);
xor UO_1955 (O_1955,N_19782,N_19950);
xor UO_1956 (O_1956,N_19907,N_19912);
and UO_1957 (O_1957,N_19885,N_19820);
nor UO_1958 (O_1958,N_19838,N_19823);
and UO_1959 (O_1959,N_19977,N_19929);
nand UO_1960 (O_1960,N_19960,N_19832);
xor UO_1961 (O_1961,N_19963,N_19960);
nand UO_1962 (O_1962,N_19970,N_19789);
nand UO_1963 (O_1963,N_19921,N_19887);
xor UO_1964 (O_1964,N_19918,N_19921);
xor UO_1965 (O_1965,N_19923,N_19921);
and UO_1966 (O_1966,N_19840,N_19997);
and UO_1967 (O_1967,N_19844,N_19761);
xnor UO_1968 (O_1968,N_19917,N_19911);
xor UO_1969 (O_1969,N_19798,N_19888);
nor UO_1970 (O_1970,N_19757,N_19938);
xnor UO_1971 (O_1971,N_19985,N_19994);
nor UO_1972 (O_1972,N_19782,N_19889);
or UO_1973 (O_1973,N_19787,N_19852);
nand UO_1974 (O_1974,N_19852,N_19855);
xnor UO_1975 (O_1975,N_19854,N_19830);
nand UO_1976 (O_1976,N_19872,N_19903);
nand UO_1977 (O_1977,N_19794,N_19872);
xor UO_1978 (O_1978,N_19923,N_19841);
xor UO_1979 (O_1979,N_19942,N_19857);
and UO_1980 (O_1980,N_19831,N_19881);
xnor UO_1981 (O_1981,N_19898,N_19756);
and UO_1982 (O_1982,N_19998,N_19892);
nor UO_1983 (O_1983,N_19757,N_19801);
or UO_1984 (O_1984,N_19800,N_19839);
and UO_1985 (O_1985,N_19797,N_19770);
nand UO_1986 (O_1986,N_19875,N_19868);
xor UO_1987 (O_1987,N_19771,N_19772);
nor UO_1988 (O_1988,N_19892,N_19772);
nand UO_1989 (O_1989,N_19752,N_19785);
nor UO_1990 (O_1990,N_19988,N_19820);
xor UO_1991 (O_1991,N_19812,N_19938);
and UO_1992 (O_1992,N_19771,N_19800);
nor UO_1993 (O_1993,N_19764,N_19979);
or UO_1994 (O_1994,N_19960,N_19880);
xnor UO_1995 (O_1995,N_19906,N_19803);
or UO_1996 (O_1996,N_19779,N_19776);
nand UO_1997 (O_1997,N_19959,N_19988);
nor UO_1998 (O_1998,N_19810,N_19975);
xnor UO_1999 (O_1999,N_19966,N_19900);
nand UO_2000 (O_2000,N_19959,N_19780);
xor UO_2001 (O_2001,N_19804,N_19857);
and UO_2002 (O_2002,N_19799,N_19918);
or UO_2003 (O_2003,N_19853,N_19860);
and UO_2004 (O_2004,N_19979,N_19840);
or UO_2005 (O_2005,N_19992,N_19781);
and UO_2006 (O_2006,N_19966,N_19871);
nand UO_2007 (O_2007,N_19881,N_19988);
or UO_2008 (O_2008,N_19853,N_19899);
nor UO_2009 (O_2009,N_19874,N_19897);
and UO_2010 (O_2010,N_19972,N_19940);
nor UO_2011 (O_2011,N_19887,N_19780);
and UO_2012 (O_2012,N_19750,N_19804);
xor UO_2013 (O_2013,N_19775,N_19942);
xor UO_2014 (O_2014,N_19959,N_19765);
nor UO_2015 (O_2015,N_19900,N_19756);
nand UO_2016 (O_2016,N_19832,N_19808);
or UO_2017 (O_2017,N_19805,N_19816);
xnor UO_2018 (O_2018,N_19917,N_19994);
nand UO_2019 (O_2019,N_19879,N_19794);
nor UO_2020 (O_2020,N_19786,N_19932);
and UO_2021 (O_2021,N_19961,N_19787);
and UO_2022 (O_2022,N_19948,N_19769);
nand UO_2023 (O_2023,N_19999,N_19934);
nor UO_2024 (O_2024,N_19853,N_19962);
or UO_2025 (O_2025,N_19773,N_19839);
xnor UO_2026 (O_2026,N_19992,N_19831);
nand UO_2027 (O_2027,N_19816,N_19850);
nor UO_2028 (O_2028,N_19989,N_19873);
nor UO_2029 (O_2029,N_19851,N_19793);
or UO_2030 (O_2030,N_19821,N_19858);
or UO_2031 (O_2031,N_19982,N_19956);
xor UO_2032 (O_2032,N_19837,N_19766);
xnor UO_2033 (O_2033,N_19807,N_19902);
or UO_2034 (O_2034,N_19851,N_19882);
nand UO_2035 (O_2035,N_19853,N_19910);
or UO_2036 (O_2036,N_19975,N_19934);
xnor UO_2037 (O_2037,N_19853,N_19930);
and UO_2038 (O_2038,N_19838,N_19976);
or UO_2039 (O_2039,N_19832,N_19869);
nor UO_2040 (O_2040,N_19869,N_19798);
or UO_2041 (O_2041,N_19874,N_19759);
xnor UO_2042 (O_2042,N_19771,N_19915);
or UO_2043 (O_2043,N_19783,N_19762);
nand UO_2044 (O_2044,N_19854,N_19980);
and UO_2045 (O_2045,N_19761,N_19881);
and UO_2046 (O_2046,N_19883,N_19788);
nor UO_2047 (O_2047,N_19856,N_19968);
xor UO_2048 (O_2048,N_19773,N_19983);
and UO_2049 (O_2049,N_19961,N_19895);
nand UO_2050 (O_2050,N_19866,N_19941);
xnor UO_2051 (O_2051,N_19915,N_19979);
xor UO_2052 (O_2052,N_19776,N_19954);
and UO_2053 (O_2053,N_19905,N_19978);
nor UO_2054 (O_2054,N_19972,N_19789);
nand UO_2055 (O_2055,N_19982,N_19954);
xor UO_2056 (O_2056,N_19795,N_19924);
or UO_2057 (O_2057,N_19856,N_19977);
nor UO_2058 (O_2058,N_19882,N_19796);
xor UO_2059 (O_2059,N_19988,N_19753);
nor UO_2060 (O_2060,N_19933,N_19921);
nand UO_2061 (O_2061,N_19778,N_19782);
xor UO_2062 (O_2062,N_19814,N_19858);
nand UO_2063 (O_2063,N_19811,N_19763);
nand UO_2064 (O_2064,N_19847,N_19888);
and UO_2065 (O_2065,N_19819,N_19955);
and UO_2066 (O_2066,N_19942,N_19945);
nand UO_2067 (O_2067,N_19982,N_19978);
xor UO_2068 (O_2068,N_19777,N_19779);
and UO_2069 (O_2069,N_19901,N_19951);
nor UO_2070 (O_2070,N_19789,N_19902);
or UO_2071 (O_2071,N_19974,N_19946);
nand UO_2072 (O_2072,N_19880,N_19852);
nand UO_2073 (O_2073,N_19977,N_19757);
xor UO_2074 (O_2074,N_19846,N_19986);
and UO_2075 (O_2075,N_19959,N_19920);
nand UO_2076 (O_2076,N_19930,N_19958);
and UO_2077 (O_2077,N_19772,N_19786);
and UO_2078 (O_2078,N_19971,N_19807);
and UO_2079 (O_2079,N_19859,N_19778);
and UO_2080 (O_2080,N_19914,N_19859);
and UO_2081 (O_2081,N_19855,N_19996);
or UO_2082 (O_2082,N_19828,N_19960);
and UO_2083 (O_2083,N_19896,N_19818);
xnor UO_2084 (O_2084,N_19777,N_19768);
or UO_2085 (O_2085,N_19827,N_19915);
nand UO_2086 (O_2086,N_19945,N_19935);
nor UO_2087 (O_2087,N_19908,N_19999);
nand UO_2088 (O_2088,N_19955,N_19843);
and UO_2089 (O_2089,N_19999,N_19874);
or UO_2090 (O_2090,N_19977,N_19877);
nand UO_2091 (O_2091,N_19819,N_19938);
or UO_2092 (O_2092,N_19940,N_19763);
and UO_2093 (O_2093,N_19953,N_19837);
xnor UO_2094 (O_2094,N_19854,N_19937);
nand UO_2095 (O_2095,N_19758,N_19754);
nand UO_2096 (O_2096,N_19967,N_19953);
nor UO_2097 (O_2097,N_19803,N_19765);
nor UO_2098 (O_2098,N_19875,N_19800);
nand UO_2099 (O_2099,N_19832,N_19983);
or UO_2100 (O_2100,N_19877,N_19953);
or UO_2101 (O_2101,N_19759,N_19784);
nor UO_2102 (O_2102,N_19856,N_19753);
xnor UO_2103 (O_2103,N_19895,N_19928);
xnor UO_2104 (O_2104,N_19756,N_19862);
xnor UO_2105 (O_2105,N_19972,N_19878);
and UO_2106 (O_2106,N_19977,N_19807);
xnor UO_2107 (O_2107,N_19892,N_19893);
nor UO_2108 (O_2108,N_19882,N_19920);
xnor UO_2109 (O_2109,N_19789,N_19759);
and UO_2110 (O_2110,N_19943,N_19814);
xnor UO_2111 (O_2111,N_19894,N_19848);
or UO_2112 (O_2112,N_19989,N_19946);
and UO_2113 (O_2113,N_19869,N_19939);
or UO_2114 (O_2114,N_19895,N_19861);
nor UO_2115 (O_2115,N_19940,N_19906);
nor UO_2116 (O_2116,N_19830,N_19798);
or UO_2117 (O_2117,N_19937,N_19986);
nor UO_2118 (O_2118,N_19896,N_19804);
and UO_2119 (O_2119,N_19881,N_19783);
nor UO_2120 (O_2120,N_19895,N_19938);
xor UO_2121 (O_2121,N_19757,N_19895);
or UO_2122 (O_2122,N_19853,N_19913);
and UO_2123 (O_2123,N_19899,N_19890);
or UO_2124 (O_2124,N_19889,N_19818);
and UO_2125 (O_2125,N_19767,N_19873);
xor UO_2126 (O_2126,N_19810,N_19832);
or UO_2127 (O_2127,N_19964,N_19971);
nand UO_2128 (O_2128,N_19914,N_19978);
or UO_2129 (O_2129,N_19985,N_19759);
nand UO_2130 (O_2130,N_19923,N_19893);
and UO_2131 (O_2131,N_19877,N_19943);
nor UO_2132 (O_2132,N_19887,N_19790);
or UO_2133 (O_2133,N_19900,N_19889);
xnor UO_2134 (O_2134,N_19914,N_19990);
xor UO_2135 (O_2135,N_19797,N_19805);
or UO_2136 (O_2136,N_19930,N_19791);
xnor UO_2137 (O_2137,N_19961,N_19903);
xor UO_2138 (O_2138,N_19855,N_19769);
or UO_2139 (O_2139,N_19917,N_19968);
nor UO_2140 (O_2140,N_19763,N_19972);
nor UO_2141 (O_2141,N_19850,N_19891);
or UO_2142 (O_2142,N_19967,N_19761);
nor UO_2143 (O_2143,N_19784,N_19970);
nand UO_2144 (O_2144,N_19937,N_19873);
or UO_2145 (O_2145,N_19974,N_19753);
nand UO_2146 (O_2146,N_19958,N_19833);
or UO_2147 (O_2147,N_19776,N_19952);
nand UO_2148 (O_2148,N_19838,N_19770);
xnor UO_2149 (O_2149,N_19971,N_19810);
xor UO_2150 (O_2150,N_19840,N_19900);
or UO_2151 (O_2151,N_19879,N_19770);
nand UO_2152 (O_2152,N_19751,N_19778);
xnor UO_2153 (O_2153,N_19922,N_19817);
and UO_2154 (O_2154,N_19906,N_19900);
nor UO_2155 (O_2155,N_19781,N_19876);
and UO_2156 (O_2156,N_19919,N_19800);
and UO_2157 (O_2157,N_19923,N_19835);
and UO_2158 (O_2158,N_19828,N_19880);
or UO_2159 (O_2159,N_19945,N_19905);
nand UO_2160 (O_2160,N_19839,N_19923);
or UO_2161 (O_2161,N_19885,N_19824);
nand UO_2162 (O_2162,N_19857,N_19863);
and UO_2163 (O_2163,N_19820,N_19901);
nor UO_2164 (O_2164,N_19939,N_19757);
or UO_2165 (O_2165,N_19793,N_19932);
nor UO_2166 (O_2166,N_19962,N_19821);
or UO_2167 (O_2167,N_19801,N_19950);
and UO_2168 (O_2168,N_19911,N_19955);
nand UO_2169 (O_2169,N_19992,N_19927);
and UO_2170 (O_2170,N_19761,N_19991);
xnor UO_2171 (O_2171,N_19916,N_19808);
nand UO_2172 (O_2172,N_19905,N_19926);
xor UO_2173 (O_2173,N_19826,N_19968);
nand UO_2174 (O_2174,N_19876,N_19975);
or UO_2175 (O_2175,N_19988,N_19930);
and UO_2176 (O_2176,N_19873,N_19998);
and UO_2177 (O_2177,N_19843,N_19858);
nand UO_2178 (O_2178,N_19772,N_19782);
xor UO_2179 (O_2179,N_19888,N_19963);
nor UO_2180 (O_2180,N_19997,N_19757);
xor UO_2181 (O_2181,N_19902,N_19779);
xor UO_2182 (O_2182,N_19881,N_19984);
nand UO_2183 (O_2183,N_19833,N_19753);
nand UO_2184 (O_2184,N_19975,N_19937);
nand UO_2185 (O_2185,N_19906,N_19963);
or UO_2186 (O_2186,N_19891,N_19785);
nand UO_2187 (O_2187,N_19916,N_19802);
or UO_2188 (O_2188,N_19905,N_19895);
and UO_2189 (O_2189,N_19975,N_19996);
or UO_2190 (O_2190,N_19872,N_19918);
nor UO_2191 (O_2191,N_19843,N_19974);
xnor UO_2192 (O_2192,N_19967,N_19789);
and UO_2193 (O_2193,N_19996,N_19889);
nand UO_2194 (O_2194,N_19803,N_19815);
and UO_2195 (O_2195,N_19871,N_19848);
and UO_2196 (O_2196,N_19966,N_19840);
xor UO_2197 (O_2197,N_19854,N_19897);
xnor UO_2198 (O_2198,N_19807,N_19838);
nand UO_2199 (O_2199,N_19918,N_19792);
nand UO_2200 (O_2200,N_19826,N_19954);
nor UO_2201 (O_2201,N_19861,N_19988);
nand UO_2202 (O_2202,N_19945,N_19760);
and UO_2203 (O_2203,N_19868,N_19905);
and UO_2204 (O_2204,N_19963,N_19886);
nor UO_2205 (O_2205,N_19758,N_19792);
and UO_2206 (O_2206,N_19824,N_19893);
and UO_2207 (O_2207,N_19865,N_19900);
nand UO_2208 (O_2208,N_19852,N_19767);
or UO_2209 (O_2209,N_19894,N_19910);
and UO_2210 (O_2210,N_19813,N_19867);
xnor UO_2211 (O_2211,N_19882,N_19990);
and UO_2212 (O_2212,N_19867,N_19993);
or UO_2213 (O_2213,N_19958,N_19986);
and UO_2214 (O_2214,N_19967,N_19930);
nor UO_2215 (O_2215,N_19930,N_19813);
nor UO_2216 (O_2216,N_19945,N_19761);
nor UO_2217 (O_2217,N_19802,N_19926);
nor UO_2218 (O_2218,N_19948,N_19913);
or UO_2219 (O_2219,N_19769,N_19873);
or UO_2220 (O_2220,N_19923,N_19840);
nand UO_2221 (O_2221,N_19817,N_19887);
and UO_2222 (O_2222,N_19879,N_19844);
and UO_2223 (O_2223,N_19836,N_19806);
nand UO_2224 (O_2224,N_19797,N_19942);
and UO_2225 (O_2225,N_19798,N_19867);
and UO_2226 (O_2226,N_19843,N_19933);
nor UO_2227 (O_2227,N_19957,N_19822);
xor UO_2228 (O_2228,N_19987,N_19885);
and UO_2229 (O_2229,N_19775,N_19892);
xnor UO_2230 (O_2230,N_19852,N_19909);
xor UO_2231 (O_2231,N_19789,N_19963);
xor UO_2232 (O_2232,N_19991,N_19882);
nor UO_2233 (O_2233,N_19833,N_19984);
or UO_2234 (O_2234,N_19797,N_19751);
xor UO_2235 (O_2235,N_19877,N_19781);
and UO_2236 (O_2236,N_19780,N_19837);
or UO_2237 (O_2237,N_19883,N_19785);
or UO_2238 (O_2238,N_19786,N_19867);
nor UO_2239 (O_2239,N_19834,N_19761);
nor UO_2240 (O_2240,N_19884,N_19848);
nor UO_2241 (O_2241,N_19790,N_19828);
or UO_2242 (O_2242,N_19877,N_19846);
nand UO_2243 (O_2243,N_19973,N_19940);
nor UO_2244 (O_2244,N_19993,N_19889);
and UO_2245 (O_2245,N_19792,N_19955);
xor UO_2246 (O_2246,N_19846,N_19861);
and UO_2247 (O_2247,N_19802,N_19894);
xor UO_2248 (O_2248,N_19865,N_19782);
or UO_2249 (O_2249,N_19777,N_19921);
nor UO_2250 (O_2250,N_19893,N_19954);
nor UO_2251 (O_2251,N_19906,N_19987);
and UO_2252 (O_2252,N_19997,N_19975);
and UO_2253 (O_2253,N_19923,N_19851);
nand UO_2254 (O_2254,N_19885,N_19939);
nand UO_2255 (O_2255,N_19914,N_19982);
nor UO_2256 (O_2256,N_19995,N_19883);
and UO_2257 (O_2257,N_19824,N_19927);
nor UO_2258 (O_2258,N_19775,N_19966);
nand UO_2259 (O_2259,N_19807,N_19852);
nand UO_2260 (O_2260,N_19848,N_19758);
nor UO_2261 (O_2261,N_19846,N_19931);
nand UO_2262 (O_2262,N_19950,N_19894);
nand UO_2263 (O_2263,N_19983,N_19770);
xnor UO_2264 (O_2264,N_19757,N_19851);
nor UO_2265 (O_2265,N_19848,N_19831);
nor UO_2266 (O_2266,N_19818,N_19753);
xnor UO_2267 (O_2267,N_19833,N_19820);
xor UO_2268 (O_2268,N_19960,N_19827);
nand UO_2269 (O_2269,N_19824,N_19803);
nor UO_2270 (O_2270,N_19996,N_19921);
or UO_2271 (O_2271,N_19929,N_19973);
or UO_2272 (O_2272,N_19928,N_19921);
nor UO_2273 (O_2273,N_19833,N_19773);
or UO_2274 (O_2274,N_19855,N_19751);
nand UO_2275 (O_2275,N_19912,N_19768);
and UO_2276 (O_2276,N_19968,N_19870);
or UO_2277 (O_2277,N_19863,N_19866);
nand UO_2278 (O_2278,N_19915,N_19759);
nand UO_2279 (O_2279,N_19828,N_19834);
nor UO_2280 (O_2280,N_19795,N_19822);
or UO_2281 (O_2281,N_19940,N_19800);
nor UO_2282 (O_2282,N_19873,N_19833);
xnor UO_2283 (O_2283,N_19984,N_19936);
nand UO_2284 (O_2284,N_19802,N_19856);
nand UO_2285 (O_2285,N_19870,N_19993);
nor UO_2286 (O_2286,N_19902,N_19960);
nor UO_2287 (O_2287,N_19929,N_19826);
or UO_2288 (O_2288,N_19940,N_19928);
nand UO_2289 (O_2289,N_19781,N_19991);
nand UO_2290 (O_2290,N_19916,N_19972);
nor UO_2291 (O_2291,N_19948,N_19995);
nor UO_2292 (O_2292,N_19973,N_19992);
xor UO_2293 (O_2293,N_19862,N_19760);
xnor UO_2294 (O_2294,N_19766,N_19883);
or UO_2295 (O_2295,N_19868,N_19884);
nand UO_2296 (O_2296,N_19794,N_19842);
and UO_2297 (O_2297,N_19762,N_19826);
or UO_2298 (O_2298,N_19806,N_19890);
xnor UO_2299 (O_2299,N_19849,N_19819);
and UO_2300 (O_2300,N_19985,N_19851);
or UO_2301 (O_2301,N_19973,N_19923);
nand UO_2302 (O_2302,N_19868,N_19972);
xnor UO_2303 (O_2303,N_19954,N_19966);
nor UO_2304 (O_2304,N_19973,N_19757);
nand UO_2305 (O_2305,N_19752,N_19764);
or UO_2306 (O_2306,N_19882,N_19914);
and UO_2307 (O_2307,N_19837,N_19853);
nand UO_2308 (O_2308,N_19862,N_19880);
and UO_2309 (O_2309,N_19815,N_19909);
or UO_2310 (O_2310,N_19757,N_19880);
or UO_2311 (O_2311,N_19853,N_19964);
or UO_2312 (O_2312,N_19919,N_19798);
and UO_2313 (O_2313,N_19996,N_19869);
nand UO_2314 (O_2314,N_19985,N_19874);
or UO_2315 (O_2315,N_19791,N_19960);
nor UO_2316 (O_2316,N_19798,N_19859);
nor UO_2317 (O_2317,N_19959,N_19834);
nor UO_2318 (O_2318,N_19928,N_19987);
xor UO_2319 (O_2319,N_19751,N_19885);
or UO_2320 (O_2320,N_19841,N_19898);
xor UO_2321 (O_2321,N_19921,N_19900);
nor UO_2322 (O_2322,N_19932,N_19775);
or UO_2323 (O_2323,N_19754,N_19891);
and UO_2324 (O_2324,N_19893,N_19755);
and UO_2325 (O_2325,N_19900,N_19864);
nand UO_2326 (O_2326,N_19842,N_19758);
nor UO_2327 (O_2327,N_19970,N_19795);
or UO_2328 (O_2328,N_19985,N_19845);
nor UO_2329 (O_2329,N_19835,N_19993);
and UO_2330 (O_2330,N_19818,N_19856);
xor UO_2331 (O_2331,N_19894,N_19823);
or UO_2332 (O_2332,N_19781,N_19795);
nor UO_2333 (O_2333,N_19924,N_19786);
nor UO_2334 (O_2334,N_19890,N_19781);
nand UO_2335 (O_2335,N_19851,N_19814);
and UO_2336 (O_2336,N_19933,N_19782);
nor UO_2337 (O_2337,N_19806,N_19866);
and UO_2338 (O_2338,N_19917,N_19795);
or UO_2339 (O_2339,N_19759,N_19932);
nand UO_2340 (O_2340,N_19857,N_19759);
or UO_2341 (O_2341,N_19759,N_19790);
nand UO_2342 (O_2342,N_19951,N_19775);
and UO_2343 (O_2343,N_19767,N_19990);
nor UO_2344 (O_2344,N_19868,N_19885);
or UO_2345 (O_2345,N_19783,N_19948);
or UO_2346 (O_2346,N_19880,N_19819);
or UO_2347 (O_2347,N_19836,N_19854);
nor UO_2348 (O_2348,N_19776,N_19788);
or UO_2349 (O_2349,N_19804,N_19999);
xor UO_2350 (O_2350,N_19897,N_19765);
or UO_2351 (O_2351,N_19752,N_19901);
or UO_2352 (O_2352,N_19960,N_19770);
nand UO_2353 (O_2353,N_19779,N_19826);
nor UO_2354 (O_2354,N_19755,N_19753);
nand UO_2355 (O_2355,N_19874,N_19994);
nor UO_2356 (O_2356,N_19768,N_19922);
xnor UO_2357 (O_2357,N_19932,N_19870);
and UO_2358 (O_2358,N_19759,N_19868);
nand UO_2359 (O_2359,N_19937,N_19875);
nand UO_2360 (O_2360,N_19838,N_19756);
or UO_2361 (O_2361,N_19919,N_19917);
nor UO_2362 (O_2362,N_19857,N_19900);
nor UO_2363 (O_2363,N_19804,N_19867);
or UO_2364 (O_2364,N_19914,N_19829);
and UO_2365 (O_2365,N_19959,N_19794);
and UO_2366 (O_2366,N_19917,N_19790);
nand UO_2367 (O_2367,N_19969,N_19782);
or UO_2368 (O_2368,N_19891,N_19859);
nand UO_2369 (O_2369,N_19917,N_19892);
or UO_2370 (O_2370,N_19838,N_19923);
and UO_2371 (O_2371,N_19912,N_19924);
or UO_2372 (O_2372,N_19966,N_19942);
nor UO_2373 (O_2373,N_19863,N_19850);
xor UO_2374 (O_2374,N_19956,N_19937);
nor UO_2375 (O_2375,N_19798,N_19885);
nor UO_2376 (O_2376,N_19773,N_19896);
nand UO_2377 (O_2377,N_19944,N_19782);
xor UO_2378 (O_2378,N_19878,N_19852);
and UO_2379 (O_2379,N_19891,N_19813);
xnor UO_2380 (O_2380,N_19854,N_19917);
nand UO_2381 (O_2381,N_19778,N_19827);
and UO_2382 (O_2382,N_19757,N_19811);
nand UO_2383 (O_2383,N_19803,N_19808);
nor UO_2384 (O_2384,N_19921,N_19939);
nand UO_2385 (O_2385,N_19796,N_19881);
and UO_2386 (O_2386,N_19773,N_19849);
nor UO_2387 (O_2387,N_19950,N_19787);
nor UO_2388 (O_2388,N_19797,N_19967);
or UO_2389 (O_2389,N_19771,N_19943);
xor UO_2390 (O_2390,N_19805,N_19985);
nand UO_2391 (O_2391,N_19907,N_19917);
or UO_2392 (O_2392,N_19945,N_19893);
and UO_2393 (O_2393,N_19803,N_19842);
nand UO_2394 (O_2394,N_19886,N_19764);
nor UO_2395 (O_2395,N_19961,N_19753);
or UO_2396 (O_2396,N_19918,N_19821);
nor UO_2397 (O_2397,N_19929,N_19899);
xnor UO_2398 (O_2398,N_19934,N_19908);
xnor UO_2399 (O_2399,N_19780,N_19880);
or UO_2400 (O_2400,N_19928,N_19881);
nor UO_2401 (O_2401,N_19905,N_19812);
and UO_2402 (O_2402,N_19953,N_19891);
and UO_2403 (O_2403,N_19937,N_19897);
and UO_2404 (O_2404,N_19884,N_19799);
xor UO_2405 (O_2405,N_19890,N_19840);
nor UO_2406 (O_2406,N_19920,N_19795);
or UO_2407 (O_2407,N_19768,N_19966);
or UO_2408 (O_2408,N_19780,N_19814);
nand UO_2409 (O_2409,N_19873,N_19967);
and UO_2410 (O_2410,N_19838,N_19933);
xnor UO_2411 (O_2411,N_19873,N_19844);
and UO_2412 (O_2412,N_19816,N_19783);
xor UO_2413 (O_2413,N_19833,N_19808);
xnor UO_2414 (O_2414,N_19923,N_19964);
and UO_2415 (O_2415,N_19981,N_19832);
or UO_2416 (O_2416,N_19807,N_19851);
nor UO_2417 (O_2417,N_19834,N_19902);
xor UO_2418 (O_2418,N_19924,N_19953);
nand UO_2419 (O_2419,N_19991,N_19888);
and UO_2420 (O_2420,N_19827,N_19811);
xor UO_2421 (O_2421,N_19992,N_19858);
and UO_2422 (O_2422,N_19846,N_19945);
or UO_2423 (O_2423,N_19828,N_19963);
and UO_2424 (O_2424,N_19785,N_19965);
nand UO_2425 (O_2425,N_19791,N_19763);
xor UO_2426 (O_2426,N_19791,N_19901);
and UO_2427 (O_2427,N_19978,N_19870);
and UO_2428 (O_2428,N_19762,N_19989);
nand UO_2429 (O_2429,N_19860,N_19998);
nor UO_2430 (O_2430,N_19754,N_19996);
nand UO_2431 (O_2431,N_19757,N_19889);
and UO_2432 (O_2432,N_19877,N_19922);
xor UO_2433 (O_2433,N_19979,N_19841);
xnor UO_2434 (O_2434,N_19916,N_19841);
nor UO_2435 (O_2435,N_19822,N_19807);
xnor UO_2436 (O_2436,N_19854,N_19776);
xnor UO_2437 (O_2437,N_19968,N_19840);
or UO_2438 (O_2438,N_19953,N_19982);
or UO_2439 (O_2439,N_19841,N_19761);
xor UO_2440 (O_2440,N_19821,N_19875);
nand UO_2441 (O_2441,N_19904,N_19945);
and UO_2442 (O_2442,N_19756,N_19939);
nand UO_2443 (O_2443,N_19832,N_19939);
nand UO_2444 (O_2444,N_19870,N_19868);
xnor UO_2445 (O_2445,N_19765,N_19750);
nand UO_2446 (O_2446,N_19844,N_19812);
or UO_2447 (O_2447,N_19947,N_19794);
nand UO_2448 (O_2448,N_19901,N_19990);
and UO_2449 (O_2449,N_19942,N_19864);
xor UO_2450 (O_2450,N_19977,N_19960);
and UO_2451 (O_2451,N_19992,N_19976);
nand UO_2452 (O_2452,N_19971,N_19836);
or UO_2453 (O_2453,N_19863,N_19921);
nand UO_2454 (O_2454,N_19935,N_19938);
or UO_2455 (O_2455,N_19888,N_19990);
nand UO_2456 (O_2456,N_19827,N_19840);
or UO_2457 (O_2457,N_19829,N_19927);
or UO_2458 (O_2458,N_19934,N_19756);
xnor UO_2459 (O_2459,N_19973,N_19894);
nand UO_2460 (O_2460,N_19889,N_19849);
or UO_2461 (O_2461,N_19962,N_19835);
nor UO_2462 (O_2462,N_19907,N_19871);
or UO_2463 (O_2463,N_19996,N_19862);
and UO_2464 (O_2464,N_19976,N_19938);
and UO_2465 (O_2465,N_19999,N_19923);
nor UO_2466 (O_2466,N_19757,N_19862);
xnor UO_2467 (O_2467,N_19883,N_19907);
and UO_2468 (O_2468,N_19794,N_19913);
nand UO_2469 (O_2469,N_19876,N_19852);
xnor UO_2470 (O_2470,N_19760,N_19821);
or UO_2471 (O_2471,N_19758,N_19984);
and UO_2472 (O_2472,N_19998,N_19829);
or UO_2473 (O_2473,N_19751,N_19776);
or UO_2474 (O_2474,N_19818,N_19848);
nand UO_2475 (O_2475,N_19867,N_19933);
nor UO_2476 (O_2476,N_19961,N_19889);
and UO_2477 (O_2477,N_19921,N_19808);
xor UO_2478 (O_2478,N_19795,N_19824);
and UO_2479 (O_2479,N_19757,N_19783);
xnor UO_2480 (O_2480,N_19969,N_19761);
and UO_2481 (O_2481,N_19792,N_19759);
or UO_2482 (O_2482,N_19861,N_19981);
nand UO_2483 (O_2483,N_19780,N_19952);
and UO_2484 (O_2484,N_19845,N_19844);
or UO_2485 (O_2485,N_19986,N_19946);
or UO_2486 (O_2486,N_19948,N_19924);
nand UO_2487 (O_2487,N_19912,N_19903);
nand UO_2488 (O_2488,N_19878,N_19893);
xor UO_2489 (O_2489,N_19897,N_19959);
xnor UO_2490 (O_2490,N_19816,N_19957);
or UO_2491 (O_2491,N_19945,N_19962);
and UO_2492 (O_2492,N_19953,N_19970);
xor UO_2493 (O_2493,N_19785,N_19777);
nor UO_2494 (O_2494,N_19965,N_19877);
nor UO_2495 (O_2495,N_19950,N_19763);
or UO_2496 (O_2496,N_19864,N_19808);
and UO_2497 (O_2497,N_19849,N_19759);
nor UO_2498 (O_2498,N_19998,N_19943);
and UO_2499 (O_2499,N_19938,N_19912);
endmodule